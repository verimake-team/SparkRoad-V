// Verilog netlist created by TD v4.5.12562
// Mon Sep 30 17:08:49 2019

`timescale 1ns / 1ps
module M0demo  // ../RTL/M0demo.v(4)
  (
  NRST,
  SWCLKTCK,
  TDI,
  XTAL1,
  nTRST,
  uart0_rxd,
  P0,
  TDO,
  XTAL2,
  uart0_txd,
  uart0_txen,
  SWDIOTMS,
  b_pad_gpio_porta
  );

  input NRST;  // ../RTL/M0demo.v(7)
  input SWCLKTCK;  // ../RTL/M0demo.v(15)
  input TDI;  // ../RTL/M0demo.v(12)
  input XTAL1;  // ../RTL/M0demo.v(5)
  input nTRST;  // ../RTL/M0demo.v(11)
  input uart0_rxd;  // ../RTL/M0demo.v(19)
  output [15:0] P0;  // ../RTL/M0demo.v(8)
  output TDO;  // ../RTL/M0demo.v(13)
  output XTAL2;  // ../RTL/M0demo.v(6)
  output uart0_txd;  // ../RTL/M0demo.v(20)
  output uart0_txen;  // ../RTL/M0demo.v(21)
  inout SWDIOTMS;  // ../RTL/M0demo.v(14)
  inout [7:0] b_pad_gpio_porta;  // ../RTL/M0demo.v(17)

  parameter BE = 0;
  parameter BKPT = 4;
  parameter DBG = 1;
  parameter NUMIRQ = 32;
  parameter SMUL = 0;
  parameter SYST = 1;
  parameter WIC = 1;
  parameter WICLINES = 34;
  parameter WPT = 2;
  wire [7:0] b_pad_gpio_porta_pad;  // ../RTL/M0demo.v(17)
  wire [13:0] n0;
  wire [13:0] n1;
  wire [31:0] \u_cmsdk_mcu/HADDR ;  // ../RTL/cmsdk_mcu.v(103)
  wire [2:0] \u_cmsdk_mcu/HSIZE ;  // ../RTL/cmsdk_mcu.v(105)
  wire [1:0] \u_cmsdk_mcu/HTRANS ;  // ../RTL/cmsdk_mcu.v(104)
  wire [31:0] \u_cmsdk_mcu/HWDATA ;  // ../RTL/cmsdk_mcu.v(107)
  wire [31:0] \u_cmsdk_mcu/flash_hrdata ;  // ../RTL/cmsdk_mcu.v(113)
  wire [15:0] \u_cmsdk_mcu/p0_altfunc ;  // ../RTL/cmsdk_mcu.v(140)
  wire [15:0] \u_cmsdk_mcu/p0_out ;  // ../RTL/cmsdk_mcu.v(138)
  wire [15:0] \u_cmsdk_mcu/p0_outen ;  // ../RTL/cmsdk_mcu.v(139)
  wire [15:0] \u_cmsdk_mcu/p1_altfunc ;  // ../RTL/cmsdk_mcu.v(145)
  wire [15:0] \u_cmsdk_mcu/p1_in ;  // ../RTL/cmsdk_mcu.v(142)
  wire [15:0] \u_cmsdk_mcu/p1_out ;  // ../RTL/cmsdk_mcu.v(143)
  wire [15:0] \u_cmsdk_mcu/p1_outen ;  // ../RTL/cmsdk_mcu.v(144)
  wire [31:0] \u_cmsdk_mcu/sram_hrdata ;  // ../RTL/cmsdk_mcu.v(119)
  wire [31:0] \u_cmsdk_mcu/u_ahb_ram/buf_hwaddr ;  // ../RTL/AHB2MEM.v(30)
  wire [31:0] \u_cmsdk_mcu/u_ahb_ram/hwdata_mask ;  // ../RTL/AHB2MEM.v(28)
  wire [31:0] \u_cmsdk_mcu/u_ahb_ram/n13 ;
  wire [31:0] \u_cmsdk_mcu/u_ahb_ram/n5 ;
  wire [31:0] \u_cmsdk_mcu/u_ahb_rom/n13 ;
  wire [2:0] \u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/reset_sync_reg ;  // ../RTL/cmsdk_mcu_clkctrl.v(62)
  wire [31:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/apbsubsys_interrupt ;  // ../RTL/cmsdk_mcu_system.v(307)
  wire [15:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr ;  // ../RTL/cmsdk_mcu_system.v(304)
  wire [11:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR ;  // ../RTL/cmsdk_ahb_gpio.v(76)
  wire [1:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOSIZE ;  // ../RTL/cmsdk_ahb_gpio.v(78)
  wire [31:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n13 ;
  wire [15:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/new_masked_int ;  // ../RTL/cmsdk_iop_gpio.v(517)
  wire [15:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/nxt_dout_padded ;  // ../RTL/cmsdk_iop_gpio.v(263)
  wire [15:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_altfuncset ;  // ../RTL/cmsdk_iop_gpio.v(361)
  wire [15:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_doutenset ;  // ../RTL/cmsdk_iop_gpio.v(322)
  wire [15:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inten_padded ;  // ../RTL/cmsdk_iop_gpio.v(397)
  wire [15:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intenset ;  // ../RTL/cmsdk_iop_gpio.v(399)
  wire [15:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpol_padded ;  // ../RTL/cmsdk_iop_gpio.v(474)
  wire [15:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpolset ;  // ../RTL/cmsdk_iop_gpio.v(476)
  wire [15:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttype_padded ;  // ../RTL/cmsdk_iop_gpio.v(435)
  wire [15:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttypeset ;  // ../RTL/cmsdk_iop_gpio.v(437)
  wire  \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/mux0_b0/B1_0 ;
  wire  \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/mux0_b1/B1_0 ;
  wire  \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/mux0_b10/B1_0 ;
  wire  \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/mux0_b11/B1_0 ;
  wire  \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/mux0_b12/B1_0 ;
  wire  \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/mux0_b13/B1_0 ;
  wire  \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/mux0_b14/B1_0 ;
  wire  \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/mux0_b15/B1_0 ;
  wire  \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/mux0_b2/B1_0 ;
  wire  \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/mux0_b3/B1_0 ;
  wire  \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/mux0_b4/B1_0 ;
  wire  \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/mux0_b5/B1_0 ;
  wire  \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/mux0_b6/B1_0 ;
  wire  \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/mux0_b7/B1_0 ;
  wire  \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/mux0_b8/B1_0 ;
  wire  \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/mux0_b9/B1_0 ;
  wire [15:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_masked_int ;  // ../RTL/cmsdk_iop_gpio.v(517)
  wire [15:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_raw_int ;  // ../RTL/cmsdk_iop_gpio.v(129)
  wire [15:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/nxt_dout_padded ;  // ../RTL/cmsdk_iop_gpio.v(263)
  wire [15:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_altfuncset ;  // ../RTL/cmsdk_iop_gpio.v(361)
  wire [15:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_doutenset ;  // ../RTL/cmsdk_iop_gpio.v(322)
  wire [15:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync1 ;  // ../RTL/cmsdk_iop_gpio.v(238)
  wire [15:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 ;  // ../RTL/cmsdk_iop_gpio.v(239)
  wire [15:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inten_padded ;  // ../RTL/cmsdk_iop_gpio.v(397)
  wire [15:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intenset ;  // ../RTL/cmsdk_iop_gpio.v(399)
  wire [15:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpol_padded ;  // ../RTL/cmsdk_iop_gpio.v(474)
  wire [15:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpolset ;  // ../RTL/cmsdk_iop_gpio.v(476)
  wire [15:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded ;  // ../RTL/cmsdk_iop_gpio.v(435)
  wire [15:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttypeset ;  // ../RTL/cmsdk_iop_gpio.v(437)
  wire [15:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_last_datain ;  // ../RTL/cmsdk_iop_gpio.v(549)
  wire [31:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n31 ;
  wire [31:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n33 ;
  wire [31:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n35 ;
  wire [31:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n37 ;
  wire [9:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel ;  // ../RTL/cmsdk_ahb_slave_mux.v(95)
  wire [7:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_int_polarity ;  // ../RTL/gpio.v(60)
  wire [7:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inten ;  // ../RTL/gpio.v(61)
  wire [7:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_intmask ;  // ../RTL/gpio.v(62)
  wire [7:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inttype_level ;  // ../RTL/gpio.v(67)
  wire [7:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_raw_intstatus ;  // ../RTL/gpio.v(73)
  wire [7:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_ddr ;  // ../RTL/gpio.v(75)
  wire [7:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_dr ;  // ../RTL/gpio.v(76)
  wire [31:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/int_gpio_ls_sync ;  // ../RTL/gpio_apbif.v(98)
  wire [31:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n81 ;
  wire  \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/sel0_b0/B1_0 ;
  wire  \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/sel0_b1/B1_0 ;
  wire  \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/sel0_b2/B1_0 ;
  wire  \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/sel0_b3/B1_0 ;
  wire  \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/sel0_b4/B1_0 ;
  wire  \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/sel0_b5/B1_0 ;
  wire  \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/sel0_b6/B1_0 ;
  wire  \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/sel0_b7/B1_0 ;
  wire [7:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/ed_int_d1 ;  // ../RTL/gpio_ctrl.v(70)
  wire [7:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/gpio_ext_porta_int ;  // ../RTL/gpio_ctrl.v(72)
  wire [7:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/gpio_intr_ed_pm ;  // ../RTL/gpio_ctrl.v(74)
  wire [7:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/int_pre_in ;  // ../RTL/gpio_ctrl.v(79)
  wire [7:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/int_s1 ;  // ../RTL/gpio_ctrl.v(80)
  wire [7:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/ls_int_in ;  // ../RTL/gpio_ctrl.v(83)
  wire [1:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/intr_stat_set ;  // ../RTL/cmsdk_apb_uart.v(147)
  wire  \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/mux3_b4/B1_0 ;
  wire  \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/mux3_b5/B1_0 ;
  wire  \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/mux3_b6/B1_0 ;
  wire [3:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n102 ;
  wire [7:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n26 ;
  wire [7:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n28 ;
  wire [15:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n37 ;
  wire [3:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n43 ;
  wire [3:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n55 ;
  wire [3:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n67 ;
  wire [3:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n92 ;
  wire [3:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_baud_cntr_f ;  // ../RTL/cmsdk_apb_uart.v(125)
  wire [15:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_baud_cntr_i ;  // ../RTL/cmsdk_apb_uart.v(123)
  wire [4:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_rx_state ;  // ../RTL/cmsdk_apb_uart.v(176)
  wire [4:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_rx_tick_cnt ;  // ../RTL/cmsdk_apb_uart.v(179)
  wire [7:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_tx_shift_buf ;  // ../RTL/cmsdk_apb_uart.v(158)
  wire [4:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_tx_state ;  // ../RTL/cmsdk_apb_uart.v(152)
  wire [4:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_tx_tick_cnt ;  // ../RTL/cmsdk_apb_uart.v(156)
  wire [7:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/read_mux_byte0 ;  // ../RTL/cmsdk_apb_uart.v(109)
  wire [7:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/read_mux_byte0_reg ;  // ../RTL/cmsdk_apb_uart.v(110)
  wire [3:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_f ;  // ../RTL/cmsdk_apb_uart.v(124)
  wire [15:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_i ;  // ../RTL/cmsdk_apb_uart.v(122)
  wire [19:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div ;  // ../RTL/cmsdk_apb_uart.v(118)
  wire [6:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_ctrl ;  // ../RTL/cmsdk_apb_uart.v(115)
  wire [7:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_rx_buf ;  // ../RTL/cmsdk_apb_uart.v(117)
  wire [7:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_tx_buf ;  // ../RTL/cmsdk_apb_uart.v(116)
  wire [6:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_shift_buf ;  // ../RTL/cmsdk_apb_uart.v(182)
  wire [3:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_state ;  // ../RTL/cmsdk_apb_uart.v(175)
  wire [3:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_tick_cnt ;  // ../RTL/cmsdk_apb_uart.v(178)
  wire [2:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rxd_lpf ;  // ../RTL/cmsdk_apb_uart.v(170)
  wire [7:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_shift_buf ;  // ../RTL/cmsdk_apb_uart.v(157)
  wire [3:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_state ;  // ../RTL/cmsdk_apb_uart.v(151)
  wire [3:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_tick_cnt ;  // ../RTL/cmsdk_apb_uart.v(155)
  wire [31:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gpio0_prdata ;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(185)
  wire [15:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/i_paddr ;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(170)
  wire [2:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/next_state ;  // ../RTL/cmsdk_ahb_to_apb.v(89)
  wire [31:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/rwdata_reg ;  // ../RTL/cmsdk_ahb_to_apb.v(90)
  wire [2:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/state_reg ;  // ../RTL/cmsdk_ahb_to_apb.v(80)
  wire [31:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_apb_slave_mux/n117 ;
  wire [31:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_apb_slave_mux/n118 ;
  wire  \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/mux3_b0/B1_0 ;
  wire [31:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/n19 ;
  wire [2:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/n38 ;
  wire [3:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/nxt_byte_strobe ;  // ../RTL/cmsdk_mcu_sysctrl.v(119)
  wire [2:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/nxt_resetinfo ;  // ../RTL/cmsdk_mcu_sysctrl.v(302)
  wire [11:2] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr ;  // ../RTL/cmsdk_mcu_sysctrl.v(123)
  wire [3:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_byte_strobe ;  // ../RTL/cmsdk_mcu_sysctrl.v(120)
  wire [2:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_resetinfo ;  // ../RTL/cmsdk_mcu_sysctrl.v(109)
  wire [31:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 ;  // ../RTL/cortexm0ds_logic.v(1528)
  wire [23:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6gpw6 ;  // ../RTL/cortexm0ds_logic.v(1545)
  wire [31:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mifpw6 ;  // ../RTL/cortexm0ds_logic.v(1531)
  wire [30:2] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 ;  // ../RTL/cortexm0ds_logic.v(1523)
  wire [31:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ntkbx6 ;  // ../RTL/cortexm0ds_logic.v(1719)
  wire [31:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nvkbx6 ;  // ../RTL/cortexm0ds_logic.v(1720)
  wire [33:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 ;  // ../RTL/cortexm0ds_logic.v(1721)
  wire [1:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pkhpw6 ;  // ../RTL/cortexm0ds_logic.v(1577)
  wire [30:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 ;  // ../RTL/cortexm0ds_logic.v(1527)
  wire [31:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgfpw6 ;  // ../RTL/cortexm0ds_logic.v(1530)
  wire [7:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vnfpw6 ;  // ../RTL/cortexm0ds_logic.v(1534)
  wire [33:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vrkbx6 ;  // ../RTL/cortexm0ds_logic.v(1718)
  wire [8:1] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xlfpw6 ;  // ../RTL/cortexm0ds_logic.v(1533)
  wire [6:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zehpw6 ;  // ../RTL/cortexm0ds_logic.v(1573)
  wire [30:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 ;  // ../RTL/cortexm0ds_logic.v(1537)
  wire [9:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/haddr_reg ;  // ../RTL/cmsdk_ahb_cs_rom_table.v(118)
  wire NRST_pad;  // ../RTL/M0demo.v(7)
  wire SWCLKTCK_pad;  // ../RTL/M0demo.v(15)
  wire XTAL1_pad;  // ../RTL/M0demo.v(5)
  wire XTAL1_wire;  // ../RTL/M0demo.v(25)
  wire XTAL2_pad;  // ../RTL/M0demo.v(6)
  wire _al_u1000_o;
  wire _al_u1001_o;
  wire _al_u1002_o;
  wire _al_u1003_o;
  wire _al_u1004_o;
  wire _al_u1006_o;
  wire _al_u1008_o;
  wire _al_u1010_o;
  wire _al_u1011_o;
  wire _al_u1012_o;
  wire _al_u1013_o;
  wire _al_u1015_o;
  wire _al_u1016_o;
  wire _al_u1017_o;
  wire _al_u1018_o;
  wire _al_u1020_o;
  wire _al_u1023_o;
  wire _al_u1024_o;
  wire _al_u1025_o;
  wire _al_u1026_o;
  wire _al_u1027_o;
  wire _al_u1028_o;
  wire _al_u1030_o;
  wire _al_u1032_o;
  wire _al_u1033_o;
  wire _al_u1034_o;
  wire _al_u1035_o;
  wire _al_u1039_o;
  wire _al_u1040_o;
  wire _al_u1048_o;
  wire _al_u1055_o;
  wire _al_u1058_o;
  wire _al_u1061_o;
  wire _al_u1064_o;
  wire _al_u1065_o;
  wire _al_u1066_o;
  wire _al_u1070_o;
  wire _al_u1071_o;
  wire _al_u1073_o;
  wire _al_u1076_o;
  wire _al_u1077_o;
  wire _al_u1078_o;
  wire _al_u1079_o;
  wire _al_u1082_o;
  wire _al_u1083_o;
  wire _al_u1085_o;
  wire _al_u1088_o;
  wire _al_u1089_o;
  wire _al_u1090_o;
  wire _al_u1091_o;
  wire _al_u1094_o;
  wire _al_u1095_o;
  wire _al_u1096_o;
  wire _al_u1097_o;
  wire _al_u1100_o;
  wire _al_u1101_o;
  wire _al_u1102_o;
  wire _al_u1103_o;
  wire _al_u1106_o;
  wire _al_u1107_o;
  wire _al_u1109_o;
  wire _al_u1112_o;
  wire _al_u1113_o;
  wire _al_u1114_o;
  wire _al_u1115_o;
  wire _al_u1118_o;
  wire _al_u1119_o;
  wire _al_u1121_o;
  wire _al_u1124_o;
  wire _al_u1125_o;
  wire _al_u1126_o;
  wire _al_u1131_o;
  wire _al_u1132_o;
  wire _al_u1133_o;
  wire _al_u1137_o;
  wire _al_u1138_o;
  wire _al_u1139_o;
  wire _al_u1142_o;
  wire _al_u1143_o;
  wire _al_u1144_o;
  wire _al_u1145_o;
  wire _al_u1148_o;
  wire _al_u1149_o;
  wire _al_u1150_o;
  wire _al_u1151_o;
  wire _al_u1154_o;
  wire _al_u1155_o;
  wire _al_u1156_o;
  wire _al_u1157_o;
  wire _al_u1160_o;
  wire _al_u1161_o;
  wire _al_u1162_o;
  wire _al_u1163_o;
  wire _al_u1166_o;
  wire _al_u1167_o;
  wire _al_u1168_o;
  wire _al_u1169_o;
  wire _al_u1173_o;
  wire _al_u1174_o;
  wire _al_u1175_o;
  wire _al_u1178_o;
  wire _al_u1179_o;
  wire _al_u1181_o;
  wire _al_u1184_o;
  wire _al_u1185_o;
  wire _al_u1186_o;
  wire _al_u1187_o;
  wire _al_u1190_o;
  wire _al_u1193_o;
  wire _al_u1196_o;
  wire _al_u1197_o;
  wire _al_u1198_o;
  wire _al_u1202_o;
  wire _al_u1203_o;
  wire _al_u1204_o;
  wire _al_u1208_o;
  wire _al_u1209_o;
  wire _al_u1210_o;
  wire _al_u1211_o;
  wire _al_u1215_o;
  wire _al_u1216_o;
  wire _al_u1217_o;
  wire _al_u1220_o;
  wire _al_u1221_o;
  wire _al_u1223_o;
  wire _al_u1226_o;
  wire _al_u1227_o;
  wire _al_u1228_o;
  wire _al_u1229_o;
  wire _al_u1232_o;
  wire _al_u1233_o;
  wire _al_u1234_o;
  wire _al_u1235_o;
  wire _al_u1238_o;
  wire _al_u1239_o;
  wire _al_u1240_o;
  wire _al_u1241_o;
  wire _al_u1244_o;
  wire _al_u1245_o;
  wire _al_u1246_o;
  wire _al_u1247_o;
  wire _al_u1250_o;
  wire _al_u1251_o;
  wire _al_u1253_o;
  wire _al_u1255_o;
  wire _al_u1257_o;
  wire _al_u1264_o;
  wire _al_u1266_o;
  wire _al_u1268_o;
  wire _al_u1269_o;
  wire _al_u1270_o;
  wire _al_u1271_o;
  wire _al_u1273_o;
  wire _al_u1276_o;
  wire _al_u1281_o;
  wire _al_u1282_o;
  wire _al_u1285_o;
  wire _al_u1286_o;
  wire _al_u1288_o;
  wire _al_u1289_o;
  wire _al_u1290_o;
  wire _al_u1291_o;
  wire _al_u1292_o;
  wire _al_u1293_o;
  wire _al_u1294_o;
  wire _al_u1296_o;
  wire _al_u1297_o;
  wire _al_u1299_o;
  wire _al_u1301_o;
  wire _al_u1304_o;
  wire _al_u1305_o;
  wire _al_u1307_o;
  wire _al_u1308_o;
  wire _al_u1309_o;
  wire _al_u1310_o;
  wire _al_u1311_o;
  wire _al_u1316_o;
  wire _al_u1319_o;
  wire _al_u1323_o;
  wire _al_u1327_o;
  wire _al_u1328_o;
  wire _al_u1329_o;
  wire _al_u1331_o;
  wire _al_u1332_o;
  wire _al_u1333_o;
  wire _al_u1334_o;
  wire _al_u1336_o;
  wire _al_u1337_o;
  wire _al_u1339_o;
  wire _al_u1341_o;
  wire _al_u1342_o;
  wire _al_u1343_o;
  wire _al_u1344_o;
  wire _al_u1345_o;
  wire _al_u1346_o;
  wire _al_u1347_o;
  wire _al_u1348_o;
  wire _al_u1350_o;
  wire _al_u1351_o;
  wire _al_u1354_o;
  wire _al_u1357_o;
  wire _al_u1359_o;
  wire _al_u1360_o;
  wire _al_u1363_o;
  wire _al_u1364_o;
  wire _al_u1366_o;
  wire _al_u1367_o;
  wire _al_u1370_o;
  wire _al_u1372_o;
  wire _al_u1375_o;
  wire _al_u1376_o;
  wire _al_u1379_o;
  wire _al_u1380_o;
  wire _al_u1381_o;
  wire _al_u1382_o;
  wire _al_u1383_o;
  wire _al_u1385_o;
  wire _al_u1387_o;
  wire _al_u1390_o;
  wire _al_u1391_o;
  wire _al_u1393_o;
  wire _al_u1394_o;
  wire _al_u1395_o;
  wire _al_u1396_o;
  wire _al_u1397_o;
  wire _al_u1399_o;
  wire _al_u1400_o;
  wire _al_u1401_o;
  wire _al_u1402_o;
  wire _al_u1403_o;
  wire _al_u1404_o;
  wire _al_u1405_o;
  wire _al_u1407_o;
  wire _al_u1408_o;
  wire _al_u1409_o;
  wire _al_u1410_o;
  wire _al_u1411_o;
  wire _al_u1412_o;
  wire _al_u1413_o;
  wire _al_u1415_o;
  wire _al_u1416_o;
  wire _al_u1417_o;
  wire _al_u1418_o;
  wire _al_u1419_o;
  wire _al_u1420_o;
  wire _al_u1421_o;
  wire _al_u1423_o;
  wire _al_u1424_o;
  wire _al_u1425_o;
  wire _al_u1426_o;
  wire _al_u1427_o;
  wire _al_u1428_o;
  wire _al_u1429_o;
  wire _al_u1431_o;
  wire _al_u1432_o;
  wire _al_u1433_o;
  wire _al_u1435_o;
  wire _al_u1436_o;
  wire _al_u1437_o;
  wire _al_u1439_o;
  wire _al_u1440_o;
  wire _al_u1441_o;
  wire _al_u1443_o;
  wire _al_u1444_o;
  wire _al_u1445_o;
  wire _al_u1447_o;
  wire _al_u1448_o;
  wire _al_u1449_o;
  wire _al_u1450_o;
  wire _al_u1451_o;
  wire _al_u1452_o;
  wire _al_u1453_o;
  wire _al_u1455_o;
  wire _al_u1456_o;
  wire _al_u1457_o;
  wire _al_u1458_o;
  wire _al_u1459_o;
  wire _al_u1460_o;
  wire _al_u1461_o;
  wire _al_u1463_o;
  wire _al_u1464_o;
  wire _al_u1465_o;
  wire _al_u1466_o;
  wire _al_u1467_o;
  wire _al_u1468_o;
  wire _al_u1469_o;
  wire _al_u1471_o;
  wire _al_u1472_o;
  wire _al_u1473_o;
  wire _al_u1474_o;
  wire _al_u1475_o;
  wire _al_u1476_o;
  wire _al_u1477_o;
  wire _al_u1479_o;
  wire _al_u1480_o;
  wire _al_u1481_o;
  wire _al_u1483_o;
  wire _al_u1484_o;
  wire _al_u1485_o;
  wire _al_u1487_o;
  wire _al_u1488_o;
  wire _al_u1489_o;
  wire _al_u1490_o;
  wire _al_u1491_o;
  wire _al_u1492_o;
  wire _al_u1493_o;
  wire _al_u1495_o;
  wire _al_u1496_o;
  wire _al_u1497_o;
  wire _al_u1498_o;
  wire _al_u1499_o;
  wire _al_u1500_o;
  wire _al_u1503_o;
  wire _al_u1504_o;
  wire _al_u1505_o;
  wire _al_u1506_o;
  wire _al_u1507_o;
  wire _al_u1508_o;
  wire _al_u1511_o;
  wire _al_u1512_o;
  wire _al_u1513_o;
  wire _al_u1514_o;
  wire _al_u1515_o;
  wire _al_u1516_o;
  wire _al_u1519_o;
  wire _al_u1520_o;
  wire _al_u1521_o;
  wire _al_u1522_o;
  wire _al_u1523_o;
  wire _al_u1524_o;
  wire _al_u1525_o;
  wire _al_u1527_o;
  wire _al_u1528_o;
  wire _al_u1529_o;
  wire _al_u1531_o;
  wire _al_u1532_o;
  wire _al_u1533_o;
  wire _al_u1535_o;
  wire _al_u1536_o;
  wire _al_u1537_o;
  wire _al_u1538_o;
  wire _al_u1539_o;
  wire _al_u1540_o;
  wire _al_u1541_o;
  wire _al_u1543_o;
  wire _al_u1544_o;
  wire _al_u1545_o;
  wire _al_u1546_o;
  wire _al_u1547_o;
  wire _al_u1548_o;
  wire _al_u1551_o;
  wire _al_u1552_o;
  wire _al_u1553_o;
  wire _al_u1554_o;
  wire _al_u1555_o;
  wire _al_u1556_o;
  wire _al_u1559_o;
  wire _al_u1560_o;
  wire _al_u1561_o;
  wire _al_u1562_o;
  wire _al_u1563_o;
  wire _al_u1564_o;
  wire _al_u1567_o;
  wire _al_u1568_o;
  wire _al_u1569_o;
  wire _al_u1570_o;
  wire _al_u1571_o;
  wire _al_u1572_o;
  wire _al_u1573_o;
  wire _al_u1575_o;
  wire _al_u1576_o;
  wire _al_u1577_o;
  wire _al_u1578_o;
  wire _al_u1579_o;
  wire _al_u1580_o;
  wire _al_u1581_o;
  wire _al_u1582_o;
  wire _al_u1583_o;
  wire _al_u1584_o;
  wire _al_u1586_o;
  wire _al_u1587_o;
  wire _al_u1588_o;
  wire _al_u1589_o;
  wire _al_u1590_o;
  wire _al_u1591_o;
  wire _al_u1592_o;
  wire _al_u1594_o;
  wire _al_u1595_o;
  wire _al_u1596_o;
  wire _al_u1597_o;
  wire _al_u1598_o;
  wire _al_u1599_o;
  wire _al_u1600_o;
  wire _al_u1602_o;
  wire _al_u1603_o;
  wire _al_u1604_o;
  wire _al_u1605_o;
  wire _al_u1606_o;
  wire _al_u1607_o;
  wire _al_u1608_o;
  wire _al_u1610_o;
  wire _al_u1611_o;
  wire _al_u1612_o;
  wire _al_u1613_o;
  wire _al_u1614_o;
  wire _al_u1615_o;
  wire _al_u1616_o;
  wire _al_u1618_o;
  wire _al_u1619_o;
  wire _al_u1620_o;
  wire _al_u1621_o;
  wire _al_u1622_o;
  wire _al_u1623_o;
  wire _al_u1624_o;
  wire _al_u1626_o;
  wire _al_u1627_o;
  wire _al_u1628_o;
  wire _al_u1629_o;
  wire _al_u1630_o;
  wire _al_u1631_o;
  wire _al_u1632_o;
  wire _al_u1634_o;
  wire _al_u1635_o;
  wire _al_u1636_o;
  wire _al_u1638_o;
  wire _al_u1642_o;
  wire _al_u1643_o;
  wire _al_u1644_o;
  wire _al_u1646_o;
  wire _al_u1648_o;
  wire _al_u1652_o;
  wire _al_u1654_o;
  wire _al_u1656_o;
  wire _al_u1657_o;
  wire _al_u1658_o;
  wire _al_u1659_o;
  wire _al_u1660_o;
  wire _al_u1662_o;
  wire _al_u1663_o;
  wire _al_u1664_o;
  wire _al_u1667_o;
  wire _al_u1668_o;
  wire _al_u1670_o;
  wire _al_u1675_o;
  wire _al_u1676_o;
  wire _al_u1679_o;
  wire _al_u1681_o;
  wire _al_u1683_o;
  wire _al_u1685_o;
  wire _al_u1687_o;
  wire _al_u1689_o;
  wire _al_u1690_o;
  wire _al_u1692_o;
  wire _al_u1694_o;
  wire _al_u1695_o;
  wire _al_u1697_o;
  wire _al_u1699_o;
  wire _al_u1701_o;
  wire _al_u1703_o;
  wire _al_u1704_o;
  wire _al_u1706_o;
  wire _al_u1708_o;
  wire _al_u1710_o;
  wire _al_u1712_o;
  wire _al_u1713_o;
  wire _al_u1715_o;
  wire _al_u1716_o;
  wire _al_u1718_o;
  wire _al_u1720_o;
  wire _al_u1721_o;
  wire _al_u1723_o;
  wire _al_u1724_o;
  wire _al_u1726_o;
  wire _al_u1727_o;
  wire _al_u1730_o;
  wire _al_u1733_o;
  wire _al_u1734_o;
  wire _al_u1737_o;
  wire _al_u1741_o;
  wire _al_u1743_o;
  wire _al_u1749_o;
  wire _al_u1751_o;
  wire _al_u1752_o;
  wire _al_u1753_o;
  wire _al_u1755_o;
  wire _al_u1756_o;
  wire _al_u1757_o;
  wire _al_u1758_o;
  wire _al_u1759_o;
  wire _al_u1761_o;
  wire _al_u1762_o;
  wire _al_u1763_o;
  wire _al_u1765_o;
  wire _al_u1767_o;
  wire _al_u1768_o;
  wire _al_u1769_o;
  wire _al_u1770_o;
  wire _al_u1772_o;
  wire _al_u1774_o;
  wire _al_u1775_o;
  wire _al_u1777_o;
  wire _al_u1778_o;
  wire _al_u1779_o;
  wire _al_u1781_o;
  wire _al_u1782_o;
  wire _al_u1783_o;
  wire _al_u1784_o;
  wire _al_u1785_o;
  wire _al_u1787_o;
  wire _al_u1788_o;
  wire _al_u1791_o;
  wire _al_u1793_o;
  wire _al_u1794_o;
  wire _al_u1796_o;
  wire _al_u1797_o;
  wire _al_u1799_o;
  wire _al_u1801_o;
  wire _al_u1802_o;
  wire _al_u1803_o;
  wire _al_u1804_o;
  wire _al_u1806_o;
  wire _al_u1808_o;
  wire _al_u1809_o;
  wire _al_u1810_o;
  wire _al_u1811_o;
  wire _al_u1812_o;
  wire _al_u1813_o;
  wire _al_u1815_o;
  wire _al_u1816_o;
  wire _al_u1817_o;
  wire _al_u1818_o;
  wire _al_u1819_o;
  wire _al_u1820_o;
  wire _al_u1821_o;
  wire _al_u1823_o;
  wire _al_u1824_o;
  wire _al_u1826_o;
  wire _al_u1827_o;
  wire _al_u1829_o;
  wire _al_u1830_o;
  wire _al_u1832_o;
  wire _al_u1833_o;
  wire _al_u1835_o;
  wire _al_u1836_o;
  wire _al_u1838_o;
  wire _al_u1839_o;
  wire _al_u1841_o;
  wire _al_u1843_o;
  wire _al_u1844_o;
  wire _al_u1846_o;
  wire _al_u1848_o;
  wire _al_u1850_o;
  wire _al_u1852_o;
  wire _al_u1854_o;
  wire _al_u1856_o;
  wire _al_u1858_o;
  wire _al_u1859_o;
  wire _al_u1861_o;
  wire _al_u1862_o;
  wire _al_u1864_o;
  wire _al_u1865_o;
  wire _al_u1867_o;
  wire _al_u1868_o;
  wire _al_u1875_o;
  wire _al_u1881_o;
  wire _al_u1882_o;
  wire _al_u1883_o;
  wire _al_u1885_o;
  wire _al_u1886_o;
  wire _al_u1887_o;
  wire _al_u1888_o;
  wire _al_u1891_o;
  wire _al_u1892_o;
  wire _al_u1893_o;
  wire _al_u1894_o;
  wire _al_u1895_o;
  wire _al_u1896_o;
  wire _al_u1899_o;
  wire _al_u1900_o;
  wire _al_u1902_o;
  wire _al_u1905_o;
  wire _al_u1906_o;
  wire _al_u1907_o;
  wire _al_u1910_o;
  wire _al_u1911_o;
  wire _al_u1912_o;
  wire _al_u1913_o;
  wire _al_u1915_o;
  wire _al_u1916_o;
  wire _al_u1917_o;
  wire _al_u1919_o;
  wire _al_u1920_o;
  wire _al_u1921_o;
  wire _al_u1923_o;
  wire _al_u1924_o;
  wire _al_u1925_o;
  wire _al_u1926_o;
  wire _al_u1928_o;
  wire _al_u1929_o;
  wire _al_u1930_o;
  wire _al_u1932_o;
  wire _al_u1933_o;
  wire _al_u1934_o;
  wire _al_u1935_o;
  wire _al_u1937_o;
  wire _al_u1938_o;
  wire _al_u1939_o;
  wire _al_u1941_o;
  wire _al_u1942_o;
  wire _al_u1943_o;
  wire _al_u1944_o;
  wire _al_u1946_o;
  wire _al_u1947_o;
  wire _al_u1948_o;
  wire _al_u1950_o;
  wire _al_u1951_o;
  wire _al_u1952_o;
  wire _al_u1953_o;
  wire _al_u1955_o;
  wire _al_u1956_o;
  wire _al_u1957_o;
  wire _al_u1959_o;
  wire _al_u1960_o;
  wire _al_u1961_o;
  wire _al_u1962_o;
  wire _al_u1964_o;
  wire _al_u1965_o;
  wire _al_u1966_o;
  wire _al_u1967_o;
  wire _al_u1968_o;
  wire _al_u1969_o;
  wire _al_u1971_o;
  wire _al_u1972_o;
  wire _al_u1973_o;
  wire _al_u1974_o;
  wire _al_u1975_o;
  wire _al_u1976_o;
  wire _al_u1977_o;
  wire _al_u1979_o;
  wire _al_u1982_o;
  wire _al_u1983_o;
  wire _al_u1986_o;
  wire _al_u1987_o;
  wire _al_u1988_o;
  wire _al_u1993_o;
  wire _al_u2032_o;
  wire _al_u2033_o;
  wire _al_u2034_o;
  wire _al_u2035_o;
  wire _al_u2036_o;
  wire _al_u2037_o;
  wire _al_u2038_o;
  wire _al_u2040_o;
  wire _al_u2055_o;
  wire _al_u2056_o;
  wire _al_u2057_o;
  wire _al_u2059_o;
  wire _al_u2060_o;
  wire _al_u2061_o;
  wire _al_u2062_o;
  wire _al_u2063_o;
  wire _al_u2077_o;
  wire _al_u2078_o;
  wire _al_u2079_o;
  wire _al_u2080_o;
  wire _al_u2081_o;
  wire _al_u2082_o;
  wire _al_u2083_o;
  wire _al_u2084_o;
  wire _al_u2085_o;
  wire _al_u2099_o;
  wire _al_u2100_o;
  wire _al_u2101_o;
  wire _al_u2102_o;
  wire _al_u2104_o;
  wire _al_u2105_o;
  wire _al_u2106_o;
  wire _al_u2107_o;
  wire _al_u2121_o;
  wire _al_u2122_o;
  wire _al_u2123_o;
  wire _al_u2124_o;
  wire _al_u2125_o;
  wire _al_u2126_o;
  wire _al_u2127_o;
  wire _al_u2128_o;
  wire _al_u2129_o;
  wire _al_u2143_o;
  wire _al_u2144_o;
  wire _al_u2145_o;
  wire _al_u2146_o;
  wire _al_u2148_o;
  wire _al_u2149_o;
  wire _al_u2150_o;
  wire _al_u2151_o;
  wire _al_u2165_o;
  wire _al_u2166_o;
  wire _al_u2167_o;
  wire _al_u2168_o;
  wire _al_u2170_o;
  wire _al_u2171_o;
  wire _al_u2173_o;
  wire _al_u2201_o;
  wire _al_u2202_o;
  wire _al_u2203_o;
  wire _al_u2204_o;
  wire _al_u2205_o;
  wire _al_u2207_o;
  wire _al_u2208_o;
  wire _al_u2210_o;
  wire _al_u2211_o;
  wire _al_u2212_o;
  wire _al_u2213_o;
  wire _al_u2215_o;
  wire _al_u2216_o;
  wire _al_u2217_o;
  wire _al_u2219_o;
  wire _al_u2220_o;
  wire _al_u2221_o;
  wire _al_u2223_o;
  wire _al_u2224_o;
  wire _al_u2225_o;
  wire _al_u2228_o;
  wire _al_u2229_o;
  wire _al_u2230_o;
  wire _al_u2231_o;
  wire _al_u2233_o;
  wire _al_u2234_o;
  wire _al_u2235_o;
  wire _al_u2237_o;
  wire _al_u2238_o;
  wire _al_u2239_o;
  wire _al_u2240_o;
  wire _al_u2242_o;
  wire _al_u2243_o;
  wire _al_u2244_o;
  wire _al_u2246_o;
  wire _al_u2247_o;
  wire _al_u2248_o;
  wire _al_u2250_o;
  wire _al_u2251_o;
  wire _al_u2252_o;
  wire _al_u2255_o;
  wire _al_u2256_o;
  wire _al_u2257_o;
  wire _al_u2259_o;
  wire _al_u2260_o;
  wire _al_u2261_o;
  wire _al_u2262_o;
  wire _al_u2264_o;
  wire _al_u2265_o;
  wire _al_u2266_o;
  wire _al_u2267_o;
  wire _al_u2268_o;
  wire _al_u2269_o;
  wire _al_u2270_o;
  wire _al_u2272_o;
  wire _al_u2274_o;
  wire _al_u2275_o;
  wire _al_u2276_o;
  wire _al_u2277_o;
  wire _al_u2278_o;
  wire _al_u2279_o;
  wire _al_u2280_o;
  wire _al_u2281_o;
  wire _al_u2283_o;
  wire _al_u2284_o;
  wire _al_u2285_o;
  wire _al_u2288_o;
  wire _al_u2289_o;
  wire _al_u2290_o;
  wire _al_u2292_o;
  wire _al_u2293_o;
  wire _al_u2295_o;
  wire _al_u2296_o;
  wire _al_u2297_o;
  wire _al_u2298_o;
  wire _al_u2299_o;
  wire _al_u2305_o;
  wire _al_u2306_o;
  wire _al_u2309_o;
  wire _al_u2312_o;
  wire _al_u2315_o;
  wire _al_u2317_o;
  wire _al_u2319_o;
  wire _al_u2321_o;
  wire _al_u2323_o;
  wire _al_u2325_o;
  wire _al_u2327_o;
  wire _al_u2329_o;
  wire _al_u2331_o;
  wire _al_u2333_o;
  wire _al_u2335_o;
  wire _al_u2337_o;
  wire _al_u2339_o;
  wire _al_u2341_o;
  wire _al_u2343_o;
  wire _al_u2345_o;
  wire _al_u2347_o;
  wire _al_u2349_o;
  wire _al_u2351_o;
  wire _al_u2353_o;
  wire _al_u2355_o;
  wire _al_u2357_o;
  wire _al_u2359_o;
  wire _al_u2361_o;
  wire _al_u2364_o;
  wire _al_u2365_o;
  wire _al_u2366_o;
  wire _al_u2367_o;
  wire _al_u2369_o;
  wire _al_u2370_o;
  wire _al_u2371_o;
  wire _al_u2373_o;
  wire _al_u2375_o;
  wire _al_u2376_o;
  wire _al_u2377_o;
  wire _al_u2378_o;
  wire _al_u2379_o;
  wire _al_u2380_o;
  wire _al_u2381_o;
  wire _al_u2382_o;
  wire _al_u2386_o;
  wire _al_u2387_o;
  wire _al_u2388_o;
  wire _al_u2389_o;
  wire _al_u2390_o;
  wire _al_u2392_o;
  wire _al_u2393_o;
  wire _al_u2395_o;
  wire _al_u2396_o;
  wire _al_u2397_o;
  wire _al_u2398_o;
  wire _al_u2399_o;
  wire _al_u2403_o;
  wire _al_u2404_o;
  wire _al_u2405_o;
  wire _al_u2406_o;
  wire _al_u2407_o;
  wire _al_u2409_o;
  wire _al_u2411_o;
  wire _al_u2412_o;
  wire _al_u2413_o;
  wire _al_u2414_o;
  wire _al_u2415_o;
  wire _al_u2416_o;
  wire _al_u2417_o;
  wire _al_u2418_o;
  wire _al_u2419_o;
  wire _al_u2420_o;
  wire _al_u2423_o;
  wire _al_u2424_o;
  wire _al_u2425_o;
  wire _al_u2426_o;
  wire _al_u2427_o;
  wire _al_u2428_o;
  wire _al_u2429_o;
  wire _al_u2433_o;
  wire _al_u2434_o;
  wire _al_u2435_o;
  wire _al_u2437_o;
  wire _al_u2438_o;
  wire _al_u2439_o;
  wire _al_u2441_o;
  wire _al_u2442_o;
  wire _al_u2443_o;
  wire _al_u2445_o;
  wire _al_u2446_o;
  wire _al_u2447_o;
  wire _al_u2449_o;
  wire _al_u2450_o;
  wire _al_u2451_o;
  wire _al_u2453_o;
  wire _al_u2454_o;
  wire _al_u2455_o;
  wire _al_u2458_o;
  wire _al_u2459_o;
  wire _al_u2460_o;
  wire _al_u2461_o;
  wire _al_u2463_o;
  wire _al_u2464_o;
  wire _al_u2467_o;
  wire _al_u2468_o;
  wire _al_u2469_o;
  wire _al_u2470_o;
  wire _al_u2476_o;
  wire _al_u2478_o;
  wire _al_u2480_o;
  wire _al_u2482_o;
  wire _al_u2484_o;
  wire _al_u2488_o;
  wire _al_u2490_o;
  wire _al_u2492_o;
  wire _al_u2494_o;
  wire _al_u2496_o;
  wire _al_u2500_o;
  wire _al_u2502_o;
  wire _al_u2504_o;
  wire _al_u2506_o;
  wire _al_u2508_o;
  wire _al_u2512_o;
  wire _al_u2514_o;
  wire _al_u2516_o;
  wire _al_u2518_o;
  wire _al_u2520_o;
  wire _al_u2642_o;
  wire _al_u2643_o;
  wire _al_u2644_o;
  wire _al_u2646_o;
  wire _al_u2647_o;
  wire _al_u2648_o;
  wire _al_u2649_o;
  wire _al_u2650_o;
  wire _al_u2717_o;
  wire _al_u2721_o;
  wire _al_u2724_o;
  wire _al_u2725_o;
  wire _al_u2728_o;
  wire _al_u2729_o;
  wire _al_u2733_o;
  wire _al_u2740_o;
  wire _al_u2741_o;
  wire _al_u2746_o;
  wire _al_u2747_o;
  wire _al_u2748_o;
  wire _al_u2749_o;
  wire _al_u2750_o;
  wire _al_u2751_o;
  wire _al_u2754_o;
  wire _al_u2755_o;
  wire _al_u2756_o;
  wire _al_u2758_o;
  wire _al_u2759_o;
  wire _al_u2760_o;
  wire _al_u2761_o;
  wire _al_u2763_o;
  wire _al_u2764_o;
  wire _al_u2766_o;
  wire _al_u2767_o;
  wire _al_u2770_o;
  wire _al_u2771_o;
  wire _al_u2772_o;
  wire _al_u2773_o;
  wire _al_u2774_o;
  wire _al_u2776_o;
  wire _al_u2778_o;
  wire _al_u2779_o;
  wire _al_u2782_o;
  wire _al_u2783_o;
  wire _al_u2784_o;
  wire _al_u2785_o;
  wire _al_u2786_o;
  wire _al_u2787_o;
  wire _al_u2789_o;
  wire _al_u2790_o;
  wire _al_u2791_o;
  wire _al_u2793_o;
  wire _al_u2794_o;
  wire _al_u2800_o;
  wire _al_u2802_o;
  wire _al_u2803_o;
  wire _al_u2804_o;
  wire _al_u2808_o;
  wire _al_u2809_o;
  wire _al_u2810_o;
  wire _al_u2813_o;
  wire _al_u2815_o;
  wire _al_u2816_o;
  wire _al_u2817_o;
  wire _al_u2818_o;
  wire _al_u2824_o;
  wire _al_u2825_o;
  wire _al_u2827_o;
  wire _al_u2829_o;
  wire _al_u2832_o;
  wire _al_u2834_o;
  wire _al_u2835_o;
  wire _al_u2836_o;
  wire _al_u2837_o;
  wire _al_u2839_o;
  wire _al_u2840_o;
  wire _al_u2841_o;
  wire _al_u2843_o;
  wire _al_u2845_o;
  wire _al_u2846_o;
  wire _al_u2847_o;
  wire _al_u2849_o;
  wire _al_u2855_o;
  wire _al_u2857_o;
  wire _al_u2858_o;
  wire _al_u2860_o;
  wire _al_u2861_o;
  wire _al_u2862_o;
  wire _al_u2863_o;
  wire _al_u2865_o;
  wire _al_u2866_o;
  wire _al_u2867_o;
  wire _al_u2868_o;
  wire _al_u2869_o;
  wire _al_u2870_o;
  wire _al_u2871_o;
  wire _al_u2872_o;
  wire _al_u2873_o;
  wire _al_u2875_o;
  wire _al_u2877_o;
  wire _al_u2878_o;
  wire _al_u2881_o;
  wire _al_u2882_o;
  wire _al_u2920_o;
  wire _al_u2921_o;
  wire _al_u2937_o;
  wire _al_u2953_o;
  wire _al_u2969_o;
  wire _al_u2985_o;
  wire _al_u2986_o;
  wire _al_u2988_o;
  wire _al_u2990_o;
  wire _al_u2992_o;
  wire _al_u3000_o;
  wire _al_u3002_o;
  wire _al_u3004_o;
  wire _al_u3006_o;
  wire _al_u3008_o;
  wire _al_u3010_o;
  wire _al_u3012_o;
  wire _al_u3015_o;
  wire _al_u3017_o;
  wire _al_u3020_o;
  wire _al_u3021_o;
  wire _al_u3022_o;
  wire _al_u3023_o;
  wire _al_u3024_o;
  wire _al_u3026_o;
  wire _al_u3027_o;
  wire _al_u3029_o;
  wire _al_u3030_o;
  wire _al_u3032_o;
  wire _al_u3034_o;
  wire _al_u3035_o;
  wire _al_u3040_o;
  wire _al_u3041_o;
  wire _al_u3046_o;
  wire _al_u3047_o;
  wire _al_u3052_o;
  wire _al_u3053_o;
  wire _al_u3057_o;
  wire _al_u3058_o;
  wire _al_u3062_o;
  wire _al_u3063_o;
  wire _al_u3067_o;
  wire _al_u3068_o;
  wire _al_u3072_o;
  wire _al_u3073_o;
  wire _al_u3075_o;
  wire _al_u3076_o;
  wire _al_u3078_o;
  wire _al_u3079_o;
  wire _al_u3080_o;
  wire _al_u3081_o;
  wire _al_u3082_o;
  wire _al_u3083_o;
  wire _al_u3085_o;
  wire _al_u3086_o;
  wire _al_u3087_o;
  wire _al_u3091_o;
  wire _al_u3092_o;
  wire _al_u3094_o;
  wire _al_u3096_o;
  wire _al_u3097_o;
  wire _al_u3100_o;
  wire _al_u3101_o;
  wire _al_u3102_o;
  wire _al_u3103_o;
  wire _al_u3104_o;
  wire _al_u3105_o;
  wire _al_u3106_o;
  wire _al_u3107_o;
  wire _al_u3108_o;
  wire _al_u3109_o;
  wire _al_u3110_o;
  wire _al_u3111_o;
  wire _al_u3114_o;
  wire _al_u3115_o;
  wire _al_u3117_o;
  wire _al_u3118_o;
  wire _al_u3119_o;
  wire _al_u3120_o;
  wire _al_u3121_o;
  wire _al_u3122_o;
  wire _al_u3124_o;
  wire _al_u3126_o;
  wire _al_u3127_o;
  wire _al_u3129_o;
  wire _al_u3132_o;
  wire _al_u3133_o;
  wire _al_u3148_o;
  wire _al_u3149_o;
  wire _al_u3150_o;
  wire _al_u3151_o;
  wire _al_u3152_o;
  wire _al_u3156_o;
  wire _al_u3157_o;
  wire _al_u3158_o;
  wire _al_u3159_o;
  wire _al_u3160_o;
  wire _al_u3164_o;
  wire _al_u3165_o;
  wire _al_u3166_o;
  wire _al_u3167_o;
  wire _al_u3169_o;
  wire _al_u3170_o;
  wire _al_u3173_o;
  wire _al_u3174_o;
  wire _al_u3175_o;
  wire _al_u3176_o;
  wire _al_u3179_o;
  wire _al_u3180_o;
  wire _al_u3181_o;
  wire _al_u3183_o;
  wire _al_u3184_o;
  wire _al_u3185_o;
  wire _al_u3186_o;
  wire _al_u3187_o;
  wire _al_u3189_o;
  wire _al_u3190_o;
  wire _al_u3191_o;
  wire _al_u3193_o;
  wire _al_u3196_o;
  wire _al_u3197_o;
  wire _al_u3198_o;
  wire _al_u3199_o;
  wire _al_u3201_o;
  wire _al_u3202_o;
  wire _al_u3203_o;
  wire _al_u3205_o;
  wire _al_u3206_o;
  wire _al_u3208_o;
  wire _al_u3210_o;
  wire _al_u3211_o;
  wire _al_u3214_o;
  wire _al_u3215_o;
  wire _al_u3216_o;
  wire _al_u3217_o;
  wire _al_u3218_o;
  wire _al_u3219_o;
  wire _al_u3221_o;
  wire _al_u3222_o;
  wire _al_u3223_o;
  wire _al_u3224_o;
  wire _al_u3225_o;
  wire _al_u3226_o;
  wire _al_u3227_o;
  wire _al_u3229_o;
  wire _al_u3230_o;
  wire _al_u3233_o;
  wire _al_u3234_o;
  wire _al_u3235_o;
  wire _al_u3236_o;
  wire _al_u3237_o;
  wire _al_u3238_o;
  wire _al_u3239_o;
  wire _al_u3240_o;
  wire _al_u3242_o;
  wire _al_u3243_o;
  wire _al_u3245_o;
  wire _al_u3246_o;
  wire _al_u3248_o;
  wire _al_u3249_o;
  wire _al_u3255_o;
  wire _al_u3256_o;
  wire _al_u3258_o;
  wire _al_u3259_o;
  wire _al_u3268_o;
  wire _al_u3270_o;
  wire _al_u3271_o;
  wire _al_u3274_o;
  wire _al_u3275_o;
  wire _al_u3279_o;
  wire _al_u3280_o;
  wire _al_u3281_o;
  wire _al_u3286_o;
  wire _al_u3287_o;
  wire _al_u3305_o;
  wire _al_u3306_o;
  wire _al_u3307_o;
  wire _al_u3308_o;
  wire _al_u3309_o;
  wire _al_u3312_o;
  wire _al_u3313_o;
  wire _al_u3314_o;
  wire _al_u3318_o;
  wire _al_u3319_o;
  wire _al_u3320_o;
  wire _al_u3322_o;
  wire _al_u3323_o;
  wire _al_u3324_o;
  wire _al_u3325_o;
  wire _al_u3326_o;
  wire _al_u3327_o;
  wire _al_u3328_o;
  wire _al_u3329_o;
  wire _al_u3333_o;
  wire _al_u3334_o;
  wire _al_u3335_o;
  wire _al_u3337_o;
  wire _al_u3338_o;
  wire _al_u3339_o;
  wire _al_u3342_o;
  wire _al_u3343_o;
  wire _al_u3345_o;
  wire _al_u3348_o;
  wire _al_u3350_o;
  wire _al_u3352_o;
  wire _al_u3355_o;
  wire _al_u3356_o;
  wire _al_u3357_o;
  wire _al_u3358_o;
  wire _al_u3359_o;
  wire _al_u3360_o;
  wire _al_u3361_o;
  wire _al_u3365_o;
  wire _al_u3366_o;
  wire _al_u3367_o;
  wire _al_u3368_o;
  wire _al_u3369_o;
  wire _al_u3370_o;
  wire _al_u3371_o;
  wire _al_u3372_o;
  wire _al_u3378_o;
  wire _al_u3381_o;
  wire _al_u3384_o;
  wire _al_u3385_o;
  wire _al_u3387_o;
  wire _al_u3388_o;
  wire _al_u3390_o;
  wire _al_u3391_o;
  wire _al_u3392_o;
  wire _al_u3393_o;
  wire _al_u3395_o;
  wire _al_u3396_o;
  wire _al_u3397_o;
  wire _al_u3398_o;
  wire _al_u3399_o;
  wire _al_u3400_o;
  wire _al_u3401_o;
  wire _al_u3402_o;
  wire _al_u3405_o;
  wire _al_u3410_o;
  wire _al_u3414_o;
  wire _al_u3415_o;
  wire _al_u3416_o;
  wire _al_u3419_o;
  wire _al_u3420_o;
  wire _al_u3421_o;
  wire _al_u3422_o;
  wire _al_u3423_o;
  wire _al_u3424_o;
  wire _al_u3429_o;
  wire _al_u3430_o;
  wire _al_u3431_o;
  wire _al_u3434_o;
  wire _al_u3435_o;
  wire _al_u3438_o;
  wire _al_u3439_o;
  wire _al_u3440_o;
  wire _al_u3441_o;
  wire _al_u3442_o;
  wire _al_u3443_o;
  wire _al_u3445_o;
  wire _al_u3446_o;
  wire _al_u3448_o;
  wire _al_u3449_o;
  wire _al_u3450_o;
  wire _al_u3451_o;
  wire _al_u3453_o;
  wire _al_u3454_o;
  wire _al_u3456_o;
  wire _al_u3457_o;
  wire _al_u3460_o;
  wire _al_u3461_o;
  wire _al_u3462_o;
  wire _al_u3463_o;
  wire _al_u3465_o;
  wire _al_u3466_o;
  wire _al_u3467_o;
  wire _al_u3468_o;
  wire _al_u3470_o;
  wire _al_u3471_o;
  wire _al_u3472_o;
  wire _al_u3473_o;
  wire _al_u3476_o;
  wire _al_u3477_o;
  wire _al_u3478_o;
  wire _al_u3479_o;
  wire _al_u3481_o;
  wire _al_u3482_o;
  wire _al_u3483_o;
  wire _al_u3486_o;
  wire _al_u3487_o;
  wire _al_u3488_o;
  wire _al_u3489_o;
  wire _al_u3491_o;
  wire _al_u3492_o;
  wire _al_u3493_o;
  wire _al_u3494_o;
  wire _al_u3497_o;
  wire _al_u3498_o;
  wire _al_u3499_o;
  wire _al_u3502_o;
  wire _al_u3503_o;
  wire _al_u3504_o;
  wire _al_u3507_o;
  wire _al_u3508_o;
  wire _al_u3509_o;
  wire _al_u3512_o;
  wire _al_u3513_o;
  wire _al_u3514_o;
  wire _al_u3515_o;
  wire _al_u3517_o;
  wire _al_u3518_o;
  wire _al_u3519_o;
  wire _al_u3520_o;
  wire _al_u3522_o;
  wire _al_u3523_o;
  wire _al_u3524_o;
  wire _al_u3527_o;
  wire _al_u3528_o;
  wire _al_u3529_o;
  wire _al_u3530_o;
  wire _al_u3532_o;
  wire _al_u3533_o;
  wire _al_u3534_o;
  wire _al_u3535_o;
  wire _al_u3538_o;
  wire _al_u3539_o;
  wire _al_u3540_o;
  wire _al_u3542_o;
  wire _al_u3544_o;
  wire _al_u3547_o;
  wire _al_u3549_o;
  wire _al_u3552_o;
  wire _al_u3553_o;
  wire _al_u3554_o;
  wire _al_u3555_o;
  wire _al_u3556_o;
  wire _al_u3557_o;
  wire _al_u3558_o;
  wire _al_u3559_o;
  wire _al_u355_o;
  wire _al_u3560_o;
  wire _al_u3561_o;
  wire _al_u3562_o;
  wire _al_u3563_o;
  wire _al_u3564_o;
  wire _al_u3565_o;
  wire _al_u3568_o;
  wire _al_u3569_o;
  wire _al_u3570_o;
  wire _al_u3571_o;
  wire _al_u3573_o;
  wire _al_u3574_o;
  wire _al_u3575_o;
  wire _al_u3576_o;
  wire _al_u3578_o;
  wire _al_u3579_o;
  wire _al_u357_o;
  wire _al_u3580_o;
  wire _al_u3581_o;
  wire _al_u3582_o;
  wire _al_u3583_o;
  wire _al_u3584_o;
  wire _al_u3585_o;
  wire _al_u3586_o;
  wire _al_u3587_o;
  wire _al_u3588_o;
  wire _al_u358_o;
  wire _al_u3591_o;
  wire _al_u3592_o;
  wire _al_u3593_o;
  wire _al_u3596_o;
  wire _al_u3597_o;
  wire _al_u359_o;
  wire _al_u3601_o;
  wire _al_u3603_o;
  wire _al_u3608_o;
  wire _al_u3609_o;
  wire _al_u360_o;
  wire _al_u3610_o;
  wire _al_u3611_o;
  wire _al_u3612_o;
  wire _al_u3613_o;
  wire _al_u3614_o;
  wire _al_u3615_o;
  wire _al_u3617_o;
  wire _al_u3618_o;
  wire _al_u3620_o;
  wire _al_u3621_o;
  wire _al_u3622_o;
  wire _al_u3624_o;
  wire _al_u3625_o;
  wire _al_u3626_o;
  wire _al_u3627_o;
  wire _al_u3628_o;
  wire _al_u3629_o;
  wire _al_u3630_o;
  wire _al_u3631_o;
  wire _al_u3632_o;
  wire _al_u3633_o;
  wire _al_u3634_o;
  wire _al_u3635_o;
  wire _al_u3636_o;
  wire _al_u3637_o;
  wire _al_u3638_o;
  wire _al_u3639_o;
  wire _al_u3640_o;
  wire _al_u3641_o;
  wire _al_u3643_o;
  wire _al_u3646_o;
  wire _al_u3647_o;
  wire _al_u3648_o;
  wire _al_u3649_o;
  wire _al_u364_o;
  wire _al_u3650_o;
  wire _al_u3652_o;
  wire _al_u3653_o;
  wire _al_u3654_o;
  wire _al_u3655_o;
  wire _al_u3657_o;
  wire _al_u3658_o;
  wire _al_u3659_o;
  wire _al_u3661_o;
  wire _al_u3662_o;
  wire _al_u3663_o;
  wire _al_u3664_o;
  wire _al_u3665_o;
  wire _al_u3666_o;
  wire _al_u3667_o;
  wire _al_u3669_o;
  wire _al_u3670_o;
  wire _al_u3672_o;
  wire _al_u3673_o;
  wire _al_u3674_o;
  wire _al_u3675_o;
  wire _al_u3677_o;
  wire _al_u3678_o;
  wire _al_u3679_o;
  wire _al_u367_o;
  wire _al_u3680_o;
  wire _al_u3681_o;
  wire _al_u3683_o;
  wire _al_u3684_o;
  wire _al_u3686_o;
  wire _al_u3688_o;
  wire _al_u368_o;
  wire _al_u3690_o;
  wire _al_u3691_o;
  wire _al_u3692_o;
  wire _al_u3693_o;
  wire _al_u3694_o;
  wire _al_u3695_o;
  wire _al_u3696_o;
  wire _al_u3697_o;
  wire _al_u3699_o;
  wire _al_u3700_o;
  wire _al_u3701_o;
  wire _al_u3702_o;
  wire _al_u3703_o;
  wire _al_u3704_o;
  wire _al_u3705_o;
  wire _al_u3706_o;
  wire _al_u3707_o;
  wire _al_u3708_o;
  wire _al_u3709_o;
  wire _al_u370_o;
  wire _al_u3710_o;
  wire _al_u3713_o;
  wire _al_u3715_o;
  wire _al_u3716_o;
  wire _al_u3717_o;
  wire _al_u3718_o;
  wire _al_u3719_o;
  wire _al_u3720_o;
  wire _al_u3721_o;
  wire _al_u3722_o;
  wire _al_u3724_o;
  wire _al_u3725_o;
  wire _al_u3726_o;
  wire _al_u3727_o;
  wire _al_u3728_o;
  wire _al_u3729_o;
  wire _al_u3730_o;
  wire _al_u3731_o;
  wire _al_u3732_o;
  wire _al_u3733_o;
  wire _al_u3734_o;
  wire _al_u3735_o;
  wire _al_u3736_o;
  wire _al_u3738_o;
  wire _al_u3739_o;
  wire _al_u3740_o;
  wire _al_u3741_o;
  wire _al_u3742_o;
  wire _al_u3743_o;
  wire _al_u3744_o;
  wire _al_u3745_o;
  wire _al_u3747_o;
  wire _al_u3748_o;
  wire _al_u3749_o;
  wire _al_u374_o;
  wire _al_u3750_o;
  wire _al_u3753_o;
  wire _al_u3754_o;
  wire _al_u3755_o;
  wire _al_u3758_o;
  wire _al_u3769_o;
  wire _al_u3776_o;
  wire _al_u3777_o;
  wire _al_u3779_o;
  wire _al_u3780_o;
  wire _al_u3781_o;
  wire _al_u3782_o;
  wire _al_u3783_o;
  wire _al_u3784_o;
  wire _al_u3787_o;
  wire _al_u3788_o;
  wire _al_u3789_o;
  wire _al_u3790_o;
  wire _al_u3791_o;
  wire _al_u3792_o;
  wire _al_u3793_o;
  wire _al_u3794_o;
  wire _al_u3795_o;
  wire _al_u3796_o;
  wire _al_u3797_o;
  wire _al_u3798_o;
  wire _al_u3799_o;
  wire _al_u379_o;
  wire _al_u3800_o;
  wire _al_u3801_o;
  wire _al_u3803_o;
  wire _al_u3804_o;
  wire _al_u3805_o;
  wire _al_u3806_o;
  wire _al_u3807_o;
  wire _al_u3808_o;
  wire _al_u3810_o;
  wire _al_u3811_o;
  wire _al_u3812_o;
  wire _al_u3813_o;
  wire _al_u3814_o;
  wire _al_u3815_o;
  wire _al_u3816_o;
  wire _al_u3817_o;
  wire _al_u3818_o;
  wire _al_u3819_o;
  wire _al_u3820_o;
  wire _al_u3821_o;
  wire _al_u3822_o;
  wire _al_u3823_o;
  wire _al_u3824_o;
  wire _al_u3825_o;
  wire _al_u3826_o;
  wire _al_u3827_o;
  wire _al_u3829_o;
  wire _al_u3830_o;
  wire _al_u3831_o;
  wire _al_u3832_o;
  wire _al_u3833_o;
  wire _al_u3834_o;
  wire _al_u3835_o;
  wire _al_u3836_o;
  wire _al_u3837_o;
  wire _al_u3838_o;
  wire _al_u3839_o;
  wire _al_u3840_o;
  wire _al_u3841_o;
  wire _al_u3843_o;
  wire _al_u3844_o;
  wire _al_u3845_o;
  wire _al_u3846_o;
  wire _al_u3847_o;
  wire _al_u3848_o;
  wire _al_u3849_o;
  wire _al_u3851_o;
  wire _al_u3853_o;
  wire _al_u3854_o;
  wire _al_u3855_o;
  wire _al_u3856_o;
  wire _al_u3857_o;
  wire _al_u3858_o;
  wire _al_u3859_o;
  wire _al_u3869_o;
  wire _al_u3870_o;
  wire _al_u3872_o;
  wire _al_u3874_o;
  wire _al_u3875_o;
  wire _al_u3878_o;
  wire _al_u3879_o;
  wire _al_u3880_o;
  wire _al_u3882_o;
  wire _al_u3884_o;
  wire _al_u3885_o;
  wire _al_u3887_o;
  wire _al_u3889_o;
  wire _al_u388_o;
  wire _al_u3891_o;
  wire _al_u3892_o;
  wire _al_u3893_o;
  wire _al_u3894_o;
  wire _al_u3895_o;
  wire _al_u3896_o;
  wire _al_u3897_o;
  wire _al_u3898_o;
  wire _al_u3900_o;
  wire _al_u3901_o;
  wire _al_u3902_o;
  wire _al_u3903_o;
  wire _al_u3904_o;
  wire _al_u3905_o;
  wire _al_u3906_o;
  wire _al_u3907_o;
  wire _al_u3908_o;
  wire _al_u3909_o;
  wire _al_u3910_o;
  wire _al_u3911_o;
  wire _al_u3912_o;
  wire _al_u3914_o;
  wire _al_u3915_o;
  wire _al_u3916_o;
  wire _al_u3917_o;
  wire _al_u3918_o;
  wire _al_u3919_o;
  wire _al_u3920_o;
  wire _al_u3921_o;
  wire _al_u3922_o;
  wire _al_u3924_o;
  wire _al_u3925_o;
  wire _al_u3926_o;
  wire _al_u3927_o;
  wire _al_u3929_o;
  wire _al_u3931_o;
  wire _al_u3932_o;
  wire _al_u3934_o;
  wire _al_u3935_o;
  wire _al_u3937_o;
  wire _al_u3938_o;
  wire _al_u3940_o;
  wire _al_u3941_o;
  wire _al_u3943_o;
  wire _al_u3944_o;
  wire _al_u3946_o;
  wire _al_u3947_o;
  wire _al_u3949_o;
  wire _al_u3950_o;
  wire _al_u3952_o;
  wire _al_u3953_o;
  wire _al_u3955_o;
  wire _al_u3956_o;
  wire _al_u3958_o;
  wire _al_u3959_o;
  wire _al_u3961_o;
  wire _al_u3962_o;
  wire _al_u3964_o;
  wire _al_u3966_o;
  wire _al_u3967_o;
  wire _al_u3969_o;
  wire _al_u3970_o;
  wire _al_u3972_o;
  wire _al_u3973_o;
  wire _al_u3975_o;
  wire _al_u3976_o;
  wire _al_u3978_o;
  wire _al_u3979_o;
  wire _al_u3981_o;
  wire _al_u3982_o;
  wire _al_u3984_o;
  wire _al_u3985_o;
  wire _al_u3987_o;
  wire _al_u3988_o;
  wire _al_u3990_o;
  wire _al_u3991_o;
  wire _al_u3993_o;
  wire _al_u3994_o;
  wire _al_u3995_o;
  wire _al_u3996_o;
  wire _al_u3997_o;
  wire _al_u4000_o;
  wire _al_u4001_o;
  wire _al_u4002_o;
  wire _al_u4003_o;
  wire _al_u4004_o;
  wire _al_u4007_o;
  wire _al_u4008_o;
  wire _al_u4009_o;
  wire _al_u4010_o;
  wire _al_u4011_o;
  wire _al_u4012_o;
  wire _al_u4013_o;
  wire _al_u4014_o;
  wire _al_u4015_o;
  wire _al_u4016_o;
  wire _al_u4017_o;
  wire _al_u4018_o;
  wire _al_u4019_o;
  wire _al_u4021_o;
  wire _al_u4022_o;
  wire _al_u4023_o;
  wire _al_u4025_o;
  wire _al_u4027_o;
  wire _al_u4028_o;
  wire _al_u4029_o;
  wire _al_u4030_o;
  wire _al_u4031_o;
  wire _al_u4032_o;
  wire _al_u4034_o;
  wire _al_u4035_o;
  wire _al_u4036_o;
  wire _al_u4037_o;
  wire _al_u4038_o;
  wire _al_u4039_o;
  wire _al_u4040_o;
  wire _al_u4041_o;
  wire _al_u4042_o;
  wire _al_u4043_o;
  wire _al_u4044_o;
  wire _al_u4045_o;
  wire _al_u4046_o;
  wire _al_u4048_o;
  wire _al_u4049_o;
  wire _al_u4052_o;
  wire _al_u4055_o;
  wire _al_u4056_o;
  wire _al_u4058_o;
  wire _al_u405_o;
  wire _al_u4060_o;
  wire _al_u4061_o;
  wire _al_u4063_o;
  wire _al_u4065_o;
  wire _al_u4066_o;
  wire _al_u4068_o;
  wire _al_u4070_o;
  wire _al_u4071_o;
  wire _al_u4073_o;
  wire _al_u4075_o;
  wire _al_u4076_o;
  wire _al_u4078_o;
  wire _al_u4080_o;
  wire _al_u4081_o;
  wire _al_u4083_o;
  wire _al_u4085_o;
  wire _al_u4086_o;
  wire _al_u4088_o;
  wire _al_u4090_o;
  wire _al_u4091_o;
  wire _al_u4093_o;
  wire _al_u4095_o;
  wire _al_u4096_o;
  wire _al_u4098_o;
  wire _al_u4100_o;
  wire _al_u4101_o;
  wire _al_u4103_o;
  wire _al_u4105_o;
  wire _al_u4106_o;
  wire _al_u4108_o;
  wire _al_u4110_o;
  wire _al_u4111_o;
  wire _al_u4113_o;
  wire _al_u4115_o;
  wire _al_u4116_o;
  wire _al_u4118_o;
  wire _al_u4120_o;
  wire _al_u4121_o;
  wire _al_u4123_o;
  wire _al_u4125_o;
  wire _al_u4126_o;
  wire _al_u4128_o;
  wire _al_u4130_o;
  wire _al_u4131_o;
  wire _al_u4133_o;
  wire _al_u4135_o;
  wire _al_u4136_o;
  wire _al_u4138_o;
  wire _al_u4140_o;
  wire _al_u4141_o;
  wire _al_u4143_o;
  wire _al_u4145_o;
  wire _al_u4146_o;
  wire _al_u4147_o;
  wire _al_u4148_o;
  wire _al_u4150_o;
  wire _al_u4151_o;
  wire _al_u4152_o;
  wire _al_u4153_o;
  wire _al_u4154_o;
  wire _al_u4155_o;
  wire _al_u4156_o;
  wire _al_u4157_o;
  wire _al_u4158_o;
  wire _al_u4159_o;
  wire _al_u4160_o;
  wire _al_u4161_o;
  wire _al_u4162_o;
  wire _al_u4163_o;
  wire _al_u4164_o;
  wire _al_u4165_o;
  wire _al_u4166_o;
  wire _al_u4168_o;
  wire _al_u4169_o;
  wire _al_u4170_o;
  wire _al_u4171_o;
  wire _al_u4172_o;
  wire _al_u4173_o;
  wire _al_u4175_o;
  wire _al_u4181_o;
  wire _al_u4182_o;
  wire _al_u4183_o;
  wire _al_u4184_o;
  wire _al_u4188_o;
  wire _al_u4189_o;
  wire _al_u4190_o;
  wire _al_u4191_o;
  wire _al_u4194_o;
  wire _al_u4195_o;
  wire _al_u4196_o;
  wire _al_u4197_o;
  wire _al_u4200_o;
  wire _al_u4201_o;
  wire _al_u4204_o;
  wire _al_u4205_o;
  wire _al_u4208_o;
  wire _al_u4209_o;
  wire _al_u4212_o;
  wire _al_u4213_o;
  wire _al_u4216_o;
  wire _al_u4217_o;
  wire _al_u4218_o;
  wire _al_u4219_o;
  wire _al_u4222_o;
  wire _al_u4223_o;
  wire _al_u4224_o;
  wire _al_u4225_o;
  wire _al_u4228_o;
  wire _al_u4229_o;
  wire _al_u4230_o;
  wire _al_u4231_o;
  wire _al_u4234_o;
  wire _al_u4235_o;
  wire _al_u4236_o;
  wire _al_u4237_o;
  wire _al_u4239_o;
  wire _al_u4240_o;
  wire _al_u4242_o;
  wire _al_u4243_o;
  wire _al_u4244_o;
  wire _al_u4245_o;
  wire _al_u4246_o;
  wire _al_u4247_o;
  wire _al_u4248_o;
  wire _al_u4249_o;
  wire _al_u4251_o;
  wire _al_u4252_o;
  wire _al_u4256_o;
  wire _al_u4258_o;
  wire _al_u4259_o;
  wire _al_u4260_o;
  wire _al_u4261_o;
  wire _al_u4262_o;
  wire _al_u4263_o;
  wire _al_u4266_o;
  wire _al_u4267_o;
  wire _al_u4269_o;
  wire _al_u4271_o;
  wire _al_u4272_o;
  wire _al_u4273_o;
  wire _al_u4274_o;
  wire _al_u4278_o;
  wire _al_u4280_o;
  wire _al_u4281_o;
  wire _al_u4282_o;
  wire _al_u4283_o;
  wire _al_u4284_o;
  wire _al_u4289_o;
  wire _al_u4290_o;
  wire _al_u4291_o;
  wire _al_u4292_o;
  wire _al_u4293_o;
  wire _al_u4294_o;
  wire _al_u4295_o;
  wire _al_u4297_o;
  wire _al_u4300_o;
  wire _al_u4302_o;
  wire _al_u4304_o;
  wire _al_u4305_o;
  wire _al_u4306_o;
  wire _al_u4308_o;
  wire _al_u4309_o;
  wire _al_u4310_o;
  wire _al_u4311_o;
  wire _al_u4312_o;
  wire _al_u4313_o;
  wire _al_u4314_o;
  wire _al_u4315_o;
  wire _al_u4316_o;
  wire _al_u4317_o;
  wire _al_u4318_o;
  wire _al_u4319_o;
  wire _al_u4320_o;
  wire _al_u4322_o;
  wire _al_u4323_o;
  wire _al_u4324_o;
  wire _al_u4325_o;
  wire _al_u4326_o;
  wire _al_u4327_o;
  wire _al_u4328_o;
  wire _al_u4329_o;
  wire _al_u4330_o;
  wire _al_u4331_o;
  wire _al_u4332_o;
  wire _al_u4333_o;
  wire _al_u4334_o;
  wire _al_u4336_o;
  wire _al_u4337_o;
  wire _al_u4338_o;
  wire _al_u4339_o;
  wire _al_u4340_o;
  wire _al_u4341_o;
  wire _al_u4342_o;
  wire _al_u4343_o;
  wire _al_u4344_o;
  wire _al_u4345_o;
  wire _al_u4346_o;
  wire _al_u4350_o;
  wire _al_u4351_o;
  wire _al_u4352_o;
  wire _al_u4353_o;
  wire _al_u4354_o;
  wire _al_u4355_o;
  wire _al_u4356_o;
  wire _al_u4357_o;
  wire _al_u4358_o;
  wire _al_u4359_o;
  wire _al_u4360_o;
  wire _al_u4361_o;
  wire _al_u4362_o;
  wire _al_u4363_o;
  wire _al_u4364_o;
  wire _al_u4367_o;
  wire _al_u4368_o;
  wire _al_u4371_o;
  wire _al_u4372_o;
  wire _al_u4373_o;
  wire _al_u4374_o;
  wire _al_u4375_o;
  wire _al_u4376_o;
  wire _al_u4377_o;
  wire _al_u4378_o;
  wire _al_u4379_o;
  wire _al_u4380_o;
  wire _al_u4381_o;
  wire _al_u4382_o;
  wire _al_u4383_o;
  wire _al_u4384_o;
  wire _al_u4385_o;
  wire _al_u4386_o;
  wire _al_u4387_o;
  wire _al_u4388_o;
  wire _al_u4389_o;
  wire _al_u4390_o;
  wire _al_u4391_o;
  wire _al_u4392_o;
  wire _al_u4393_o;
  wire _al_u4395_o;
  wire _al_u4396_o;
  wire _al_u4397_o;
  wire _al_u4398_o;
  wire _al_u4399_o;
  wire _al_u4400_o;
  wire _al_u4401_o;
  wire _al_u4402_o;
  wire _al_u4403_o;
  wire _al_u4404_o;
  wire _al_u4405_o;
  wire _al_u4406_o;
  wire _al_u4407_o;
  wire _al_u4408_o;
  wire _al_u4409_o;
  wire _al_u4410_o;
  wire _al_u4411_o;
  wire _al_u4412_o;
  wire _al_u4413_o;
  wire _al_u4414_o;
  wire _al_u4415_o;
  wire _al_u4416_o;
  wire _al_u4419_o;
  wire _al_u4421_o;
  wire _al_u4422_o;
  wire _al_u4423_o;
  wire _al_u4425_o;
  wire _al_u4426_o;
  wire _al_u4438_o;
  wire _al_u4450_o;
  wire _al_u4451_o;
  wire _al_u4452_o;
  wire _al_u4455_o;
  wire _al_u4456_o;
  wire _al_u4457_o;
  wire _al_u4459_o;
  wire _al_u4460_o;
  wire _al_u4461_o;
  wire _al_u4462_o;
  wire _al_u4463_o;
  wire _al_u4464_o;
  wire _al_u4465_o;
  wire _al_u4466_o;
  wire _al_u4467_o;
  wire _al_u4468_o;
  wire _al_u4470_o;
  wire _al_u4471_o;
  wire _al_u4472_o;
  wire _al_u4473_o;
  wire _al_u4474_o;
  wire _al_u4475_o;
  wire _al_u4476_o;
  wire _al_u4478_o;
  wire _al_u4480_o;
  wire _al_u4481_o;
  wire _al_u4483_o;
  wire _al_u4484_o;
  wire _al_u4485_o;
  wire _al_u4486_o;
  wire _al_u4487_o;
  wire _al_u4488_o;
  wire _al_u4490_o;
  wire _al_u4492_o;
  wire _al_u4495_o;
  wire _al_u4499_o;
  wire _al_u4500_o;
  wire _al_u4501_o;
  wire _al_u4509_o;
  wire _al_u4511_o;
  wire _al_u4512_o;
  wire _al_u4513_o;
  wire _al_u4514_o;
  wire _al_u4515_o;
  wire _al_u4516_o;
  wire _al_u4517_o;
  wire _al_u4519_o;
  wire _al_u4520_o;
  wire _al_u4521_o;
  wire _al_u4523_o;
  wire _al_u4524_o;
  wire _al_u4525_o;
  wire _al_u4526_o;
  wire _al_u4527_o;
  wire _al_u4528_o;
  wire _al_u4529_o;
  wire _al_u452_o;
  wire _al_u4530_o;
  wire _al_u4532_o;
  wire _al_u4533_o;
  wire _al_u4534_o;
  wire _al_u4535_o;
  wire _al_u4537_o;
  wire _al_u4539_o;
  wire _al_u453_o;
  wire _al_u4542_o;
  wire _al_u4544_o;
  wire _al_u4545_o;
  wire _al_u4546_o;
  wire _al_u4548_o;
  wire _al_u4549_o;
  wire _al_u4550_o;
  wire _al_u4551_o;
  wire _al_u4552_o;
  wire _al_u4553_o;
  wire _al_u4557_o;
  wire _al_u4558_o;
  wire _al_u4559_o;
  wire _al_u4560_o;
  wire _al_u4561_o;
  wire _al_u4562_o;
  wire _al_u4563_o;
  wire _al_u4564_o;
  wire _al_u4566_o;
  wire _al_u4567_o;
  wire _al_u4568_o;
  wire _al_u4569_o;
  wire _al_u456_o;
  wire _al_u4571_o;
  wire _al_u4573_o;
  wire _al_u4574_o;
  wire _al_u4575_o;
  wire _al_u4576_o;
  wire _al_u4577_o;
  wire _al_u4578_o;
  wire _al_u4580_o;
  wire _al_u4581_o;
  wire _al_u4582_o;
  wire _al_u4583_o;
  wire _al_u4584_o;
  wire _al_u4586_o;
  wire _al_u4587_o;
  wire _al_u4588_o;
  wire _al_u4589_o;
  wire _al_u4591_o;
  wire _al_u4592_o;
  wire _al_u4593_o;
  wire _al_u4594_o;
  wire _al_u4595_o;
  wire _al_u4596_o;
  wire _al_u4597_o;
  wire _al_u4598_o;
  wire _al_u4599_o;
  wire _al_u4600_o;
  wire _al_u4601_o;
  wire _al_u4602_o;
  wire _al_u4603_o;
  wire _al_u4604_o;
  wire _al_u4605_o;
  wire _al_u4607_o;
  wire _al_u4608_o;
  wire _al_u4609_o;
  wire _al_u4610_o;
  wire _al_u4611_o;
  wire _al_u4612_o;
  wire _al_u4613_o;
  wire _al_u4616_o;
  wire _al_u4617_o;
  wire _al_u4618_o;
  wire _al_u4619_o;
  wire _al_u4620_o;
  wire _al_u4621_o;
  wire _al_u4623_o;
  wire _al_u4624_o;
  wire _al_u4625_o;
  wire _al_u4626_o;
  wire _al_u4627_o;
  wire _al_u4628_o;
  wire _al_u4629_o;
  wire _al_u462_o;
  wire _al_u4631_o;
  wire _al_u4633_o;
  wire _al_u4634_o;
  wire _al_u4635_o;
  wire _al_u4636_o;
  wire _al_u4637_o;
  wire _al_u4638_o;
  wire _al_u4639_o;
  wire _al_u463_o;
  wire _al_u4642_o;
  wire _al_u4643_o;
  wire _al_u4644_o;
  wire _al_u4645_o;
  wire _al_u4646_o;
  wire _al_u4647_o;
  wire _al_u4649_o;
  wire _al_u4650_o;
  wire _al_u4651_o;
  wire _al_u4652_o;
  wire _al_u4653_o;
  wire _al_u4654_o;
  wire _al_u4655_o;
  wire _al_u4657_o;
  wire _al_u4659_o;
  wire _al_u465_o;
  wire _al_u4660_o;
  wire _al_u4661_o;
  wire _al_u4662_o;
  wire _al_u4663_o;
  wire _al_u4664_o;
  wire _al_u4665_o;
  wire _al_u4668_o;
  wire _al_u4669_o;
  wire _al_u4670_o;
  wire _al_u4671_o;
  wire _al_u4672_o;
  wire _al_u4673_o;
  wire _al_u4675_o;
  wire _al_u4676_o;
  wire _al_u4677_o;
  wire _al_u4678_o;
  wire _al_u4679_o;
  wire _al_u467_o;
  wire _al_u4680_o;
  wire _al_u4681_o;
  wire _al_u4682_o;
  wire _al_u4683_o;
  wire _al_u4684_o;
  wire _al_u4685_o;
  wire _al_u4686_o;
  wire _al_u4687_o;
  wire _al_u4688_o;
  wire _al_u4689_o;
  wire _al_u4690_o;
  wire _al_u4692_o;
  wire _al_u4693_o;
  wire _al_u4694_o;
  wire _al_u4695_o;
  wire _al_u4697_o;
  wire _al_u4698_o;
  wire _al_u4699_o;
  wire _al_u4700_o;
  wire _al_u4701_o;
  wire _al_u4702_o;
  wire _al_u4703_o;
  wire _al_u4704_o;
  wire _al_u4705_o;
  wire _al_u4706_o;
  wire _al_u4708_o;
  wire _al_u4709_o;
  wire _al_u470_o;
  wire _al_u4711_o;
  wire _al_u4712_o;
  wire _al_u4713_o;
  wire _al_u4716_o;
  wire _al_u4717_o;
  wire _al_u4718_o;
  wire _al_u4719_o;
  wire _al_u4720_o;
  wire _al_u4722_o;
  wire _al_u4723_o;
  wire _al_u4724_o;
  wire _al_u4725_o;
  wire _al_u4726_o;
  wire _al_u4727_o;
  wire _al_u4728_o;
  wire _al_u4729_o;
  wire _al_u472_o;
  wire _al_u4730_o;
  wire _al_u4731_o;
  wire _al_u4732_o;
  wire _al_u4733_o;
  wire _al_u4734_o;
  wire _al_u4735_o;
  wire _al_u4736_o;
  wire _al_u4737_o;
  wire _al_u473_o;
  wire _al_u4740_o;
  wire _al_u4741_o;
  wire _al_u4742_o;
  wire _al_u4743_o;
  wire _al_u4744_o;
  wire _al_u4746_o;
  wire _al_u4747_o;
  wire _al_u4749_o;
  wire _al_u4750_o;
  wire _al_u4751_o;
  wire _al_u4752_o;
  wire _al_u4753_o;
  wire _al_u4754_o;
  wire _al_u4755_o;
  wire _al_u4756_o;
  wire _al_u4757_o;
  wire _al_u4758_o;
  wire _al_u475_o;
  wire _al_u4760_o;
  wire _al_u4761_o;
  wire _al_u4762_o;
  wire _al_u4763_o;
  wire _al_u4764_o;
  wire _al_u4766_o;
  wire _al_u4767_o;
  wire _al_u4768_o;
  wire _al_u4769_o;
  wire _al_u4770_o;
  wire _al_u4772_o;
  wire _al_u4773_o;
  wire _al_u4774_o;
  wire _al_u4775_o;
  wire _al_u4776_o;
  wire _al_u4777_o;
  wire _al_u4780_o;
  wire _al_u4781_o;
  wire _al_u4782_o;
  wire _al_u4783_o;
  wire _al_u4784_o;
  wire _al_u4786_o;
  wire _al_u4787_o;
  wire _al_u4788_o;
  wire _al_u4789_o;
  wire _al_u478_o;
  wire _al_u4790_o;
  wire _al_u4792_o;
  wire _al_u4793_o;
  wire _al_u4794_o;
  wire _al_u4795_o;
  wire _al_u4796_o;
  wire _al_u4797_o;
  wire _al_u4801_o;
  wire _al_u4802_o;
  wire _al_u4803_o;
  wire _al_u4804_o;
  wire _al_u4805_o;
  wire _al_u4806_o;
  wire _al_u4807_o;
  wire _al_u4808_o;
  wire _al_u4809_o;
  wire _al_u480_o;
  wire _al_u4810_o;
  wire _al_u4811_o;
  wire _al_u4812_o;
  wire _al_u4814_o;
  wire _al_u4815_o;
  wire _al_u4816_o;
  wire _al_u4817_o;
  wire _al_u481_o;
  wire _al_u4820_o;
  wire _al_u4821_o;
  wire _al_u4822_o;
  wire _al_u4823_o;
  wire _al_u4824_o;
  wire _al_u4826_o;
  wire _al_u4827_o;
  wire _al_u4828_o;
  wire _al_u4829_o;
  wire _al_u482_o;
  wire _al_u4830_o;
  wire _al_u4832_o;
  wire _al_u4833_o;
  wire _al_u4834_o;
  wire _al_u4835_o;
  wire _al_u4836_o;
  wire _al_u4837_o;
  wire _al_u4838_o;
  wire _al_u483_o;
  wire _al_u4841_o;
  wire _al_u4842_o;
  wire _al_u4844_o;
  wire _al_u4845_o;
  wire _al_u4846_o;
  wire _al_u4847_o;
  wire _al_u4848_o;
  wire _al_u4849_o;
  wire _al_u4850_o;
  wire _al_u4851_o;
  wire _al_u4852_o;
  wire _al_u4853_o;
  wire _al_u4854_o;
  wire _al_u4855_o;
  wire _al_u4857_o;
  wire _al_u4858_o;
  wire _al_u4859_o;
  wire _al_u4860_o;
  wire _al_u4861_o;
  wire _al_u4862_o;
  wire _al_u4863_o;
  wire _al_u4865_o;
  wire _al_u4866_o;
  wire _al_u4867_o;
  wire _al_u486_o;
  wire _al_u4871_o;
  wire _al_u4872_o;
  wire _al_u4873_o;
  wire _al_u4874_o;
  wire _al_u4875_o;
  wire _al_u4876_o;
  wire _al_u4877_o;
  wire _al_u4878_o;
  wire _al_u4879_o;
  wire _al_u487_o;
  wire _al_u4880_o;
  wire _al_u4881_o;
  wire _al_u4882_o;
  wire _al_u4884_o;
  wire _al_u4885_o;
  wire _al_u4886_o;
  wire _al_u4887_o;
  wire _al_u488_o;
  wire _al_u4890_o;
  wire _al_u4891_o;
  wire _al_u4892_o;
  wire _al_u4893_o;
  wire _al_u4894_o;
  wire _al_u4896_o;
  wire _al_u4897_o;
  wire _al_u4898_o;
  wire _al_u489_o;
  wire _al_u4900_o;
  wire _al_u4901_o;
  wire _al_u4902_o;
  wire _al_u4903_o;
  wire _al_u4904_o;
  wire _al_u4905_o;
  wire _al_u4906_o;
  wire _al_u4908_o;
  wire _al_u4909_o;
  wire _al_u4910_o;
  wire _al_u4912_o;
  wire _al_u4914_o;
  wire _al_u4916_o;
  wire _al_u4917_o;
  wire _al_u4918_o;
  wire _al_u4919_o;
  wire _al_u491_o;
  wire _al_u4920_o;
  wire _al_u4921_o;
  wire _al_u4922_o;
  wire _al_u4923_o;
  wire _al_u4925_o;
  wire _al_u4927_o;
  wire _al_u4928_o;
  wire _al_u492_o;
  wire _al_u4930_o;
  wire _al_u4931_o;
  wire _al_u4932_o;
  wire _al_u4934_o;
  wire _al_u4935_o;
  wire _al_u4937_o;
  wire _al_u4938_o;
  wire _al_u4939_o;
  wire _al_u493_o;
  wire _al_u4940_o;
  wire _al_u4941_o;
  wire _al_u4942_o;
  wire _al_u4943_o;
  wire _al_u4944_o;
  wire _al_u4945_o;
  wire _al_u4946_o;
  wire _al_u4947_o;
  wire _al_u4948_o;
  wire _al_u4949_o;
  wire _al_u494_o;
  wire _al_u4950_o;
  wire _al_u4951_o;
  wire _al_u4953_o;
  wire _al_u4954_o;
  wire _al_u4955_o;
  wire _al_u4957_o;
  wire _al_u4959_o;
  wire _al_u4961_o;
  wire _al_u4963_o;
  wire _al_u4965_o;
  wire _al_u4967_o;
  wire _al_u4969_o;
  wire _al_u496_o;
  wire _al_u4970_o;
  wire _al_u4971_o;
  wire _al_u4973_o;
  wire _al_u4974_o;
  wire _al_u4975_o;
  wire _al_u4977_o;
  wire _al_u497_o;
  wire _al_u4981_o;
  wire _al_u4982_o;
  wire _al_u4983_o;
  wire _al_u4984_o;
  wire _al_u4985_o;
  wire _al_u4986_o;
  wire _al_u4987_o;
  wire _al_u4988_o;
  wire _al_u4989_o;
  wire _al_u498_o;
  wire _al_u4990_o;
  wire _al_u4993_o;
  wire _al_u4994_o;
  wire _al_u499_o;
  wire _al_u5000_o;
  wire _al_u5001_o;
  wire _al_u5003_o;
  wire _al_u5006_o;
  wire _al_u5009_o;
  wire _al_u5017_o;
  wire _al_u5020_o;
  wire _al_u5021_o;
  wire _al_u5023_o;
  wire _al_u5024_o;
  wire _al_u5025_o;
  wire _al_u5026_o;
  wire _al_u5028_o;
  wire _al_u5029_o;
  wire _al_u5030_o;
  wire _al_u5031_o;
  wire _al_u5032_o;
  wire _al_u5036_o;
  wire _al_u5037_o;
  wire _al_u5038_o;
  wire _al_u5039_o;
  wire _al_u5040_o;
  wire _al_u5044_o;
  wire _al_u5047_o;
  wire _al_u5048_o;
  wire _al_u5049_o;
  wire _al_u5050_o;
  wire _al_u5051_o;
  wire _al_u5052_o;
  wire _al_u5053_o;
  wire _al_u5055_o;
  wire _al_u5056_o;
  wire _al_u5057_o;
  wire _al_u5058_o;
  wire _al_u5059_o;
  wire _al_u5061_o;
  wire _al_u5062_o;
  wire _al_u5063_o;
  wire _al_u5066_o;
  wire _al_u5067_o;
  wire _al_u5069_o;
  wire _al_u5070_o;
  wire _al_u5071_o;
  wire _al_u5072_o;
  wire _al_u5073_o;
  wire _al_u5074_o;
  wire _al_u5075_o;
  wire _al_u5076_o;
  wire _al_u5078_o;
  wire _al_u5080_o;
  wire _al_u5081_o;
  wire _al_u5082_o;
  wire _al_u5083_o;
  wire _al_u5084_o;
  wire _al_u5085_o;
  wire _al_u5086_o;
  wire _al_u5087_o;
  wire _al_u5088_o;
  wire _al_u5090_o;
  wire _al_u5091_o;
  wire _al_u5092_o;
  wire _al_u5094_o;
  wire _al_u5095_o;
  wire _al_u5096_o;
  wire _al_u5097_o;
  wire _al_u5098_o;
  wire _al_u5099_o;
  wire _al_u5100_o;
  wire _al_u5101_o;
  wire _al_u5103_o;
  wire _al_u5104_o;
  wire _al_u5105_o;
  wire _al_u5107_o;
  wire _al_u5108_o;
  wire _al_u5109_o;
  wire _al_u5110_o;
  wire _al_u5111_o;
  wire _al_u5112_o;
  wire _al_u5113_o;
  wire _al_u5114_o;
  wire _al_u5116_o;
  wire _al_u5117_o;
  wire _al_u5118_o;
  wire _al_u5119_o;
  wire _al_u5120_o;
  wire _al_u5121_o;
  wire _al_u5122_o;
  wire _al_u5125_o;
  wire _al_u5126_o;
  wire _al_u5127_o;
  wire _al_u5128_o;
  wire _al_u5130_o;
  wire _al_u5131_o;
  wire _al_u5132_o;
  wire _al_u5133_o;
  wire _al_u5134_o;
  wire _al_u5135_o;
  wire _al_u5136_o;
  wire _al_u5137_o;
  wire _al_u5138_o;
  wire _al_u5139_o;
  wire _al_u5140_o;
  wire _al_u5141_o;
  wire _al_u5142_o;
  wire _al_u5143_o;
  wire _al_u5144_o;
  wire _al_u5145_o;
  wire _al_u5146_o;
  wire _al_u5147_o;
  wire _al_u5148_o;
  wire _al_u5149_o;
  wire _al_u5151_o;
  wire _al_u5152_o;
  wire _al_u5153_o;
  wire _al_u5154_o;
  wire _al_u5156_o;
  wire _al_u5157_o;
  wire _al_u5159_o;
  wire _al_u5163_o;
  wire _al_u5164_o;
  wire _al_u5165_o;
  wire _al_u5166_o;
  wire _al_u5167_o;
  wire _al_u5168_o;
  wire _al_u5169_o;
  wire _al_u5171_o;
  wire _al_u5173_o;
  wire _al_u5176_o;
  wire _al_u5177_o;
  wire _al_u5178_o;
  wire _al_u5179_o;
  wire _al_u5180_o;
  wire _al_u5181_o;
  wire _al_u5183_o;
  wire _al_u5186_o;
  wire _al_u5187_o;
  wire _al_u5188_o;
  wire _al_u5189_o;
  wire _al_u5190_o;
  wire _al_u5191_o;
  wire _al_u5192_o;
  wire _al_u5193_o;
  wire _al_u5194_o;
  wire _al_u5196_o;
  wire _al_u5197_o;
  wire _al_u5198_o;
  wire _al_u5199_o;
  wire _al_u5200_o;
  wire _al_u5201_o;
  wire _al_u5203_o;
  wire _al_u5204_o;
  wire _al_u5206_o;
  wire _al_u5207_o;
  wire _al_u5208_o;
  wire _al_u5213_o;
  wire _al_u5214_o;
  wire _al_u5215_o;
  wire _al_u5216_o;
  wire _al_u5217_o;
  wire _al_u5218_o;
  wire _al_u5219_o;
  wire _al_u5220_o;
  wire _al_u5222_o;
  wire _al_u5223_o;
  wire _al_u5224_o;
  wire _al_u5225_o;
  wire _al_u5229_o;
  wire _al_u5230_o;
  wire _al_u5231_o;
  wire _al_u5232_o;
  wire _al_u5233_o;
  wire _al_u5235_o;
  wire _al_u5236_o;
  wire _al_u5237_o;
  wire _al_u5238_o;
  wire _al_u5239_o;
  wire _al_u5240_o;
  wire _al_u5241_o;
  wire _al_u5242_o;
  wire _al_u5243_o;
  wire _al_u5245_o;
  wire _al_u5246_o;
  wire _al_u5251_o;
  wire _al_u5252_o;
  wire _al_u5253_o;
  wire _al_u5254_o;
  wire _al_u5255_o;
  wire _al_u5256_o;
  wire _al_u5257_o;
  wire _al_u5258_o;
  wire _al_u5260_o;
  wire _al_u5261_o;
  wire _al_u5262_o;
  wire _al_u5263_o;
  wire _al_u5264_o;
  wire _al_u5265_o;
  wire _al_u5266_o;
  wire _al_u5267_o;
  wire _al_u5268_o;
  wire _al_u526_o;
  wire _al_u5271_o;
  wire _al_u5274_o;
  wire _al_u5275_o;
  wire _al_u5276_o;
  wire _al_u5278_o;
  wire _al_u5280_o;
  wire _al_u5282_o;
  wire _al_u5284_o;
  wire _al_u5285_o;
  wire _al_u5286_o;
  wire _al_u5287_o;
  wire _al_u5288_o;
  wire _al_u5291_o;
  wire _al_u5292_o;
  wire _al_u5293_o;
  wire _al_u5294_o;
  wire _al_u5295_o;
  wire _al_u5296_o;
  wire _al_u5297_o;
  wire _al_u5298_o;
  wire _al_u5299_o;
  wire _al_u529_o;
  wire _al_u5300_o;
  wire _al_u5301_o;
  wire _al_u5302_o;
  wire _al_u5303_o;
  wire _al_u5304_o;
  wire _al_u5305_o;
  wire _al_u5307_o;
  wire _al_u5308_o;
  wire _al_u530_o;
  wire _al_u5310_o;
  wire _al_u5311_o;
  wire _al_u5312_o;
  wire _al_u5313_o;
  wire _al_u5315_o;
  wire _al_u5316_o;
  wire _al_u5317_o;
  wire _al_u5318_o;
  wire _al_u5319_o;
  wire _al_u5320_o;
  wire _al_u5321_o;
  wire _al_u5323_o;
  wire _al_u5324_o;
  wire _al_u5325_o;
  wire _al_u5327_o;
  wire _al_u5328_o;
  wire _al_u5329_o;
  wire _al_u5331_o;
  wire _al_u5332_o;
  wire _al_u5333_o;
  wire _al_u5334_o;
  wire _al_u5335_o;
  wire _al_u5336_o;
  wire _al_u5337_o;
  wire _al_u5338_o;
  wire _al_u5339_o;
  wire _al_u533_o;
  wire _al_u5340_o;
  wire _al_u5341_o;
  wire _al_u5344_o;
  wire _al_u5345_o;
  wire _al_u5346_o;
  wire _al_u5347_o;
  wire _al_u5348_o;
  wire _al_u5349_o;
  wire _al_u5351_o;
  wire _al_u5352_o;
  wire _al_u5353_o;
  wire _al_u5354_o;
  wire _al_u5355_o;
  wire _al_u5357_o;
  wire _al_u5358_o;
  wire _al_u5359_o;
  wire _al_u5360_o;
  wire _al_u5361_o;
  wire _al_u5362_o;
  wire _al_u5364_o;
  wire _al_u5365_o;
  wire _al_u5366_o;
  wire _al_u5369_o;
  wire _al_u5370_o;
  wire _al_u5371_o;
  wire _al_u5375_o;
  wire _al_u5376_o;
  wire _al_u5377_o;
  wire _al_u5378_o;
  wire _al_u5379_o;
  wire _al_u5380_o;
  wire _al_u5381_o;
  wire _al_u5382_o;
  wire _al_u5383_o;
  wire _al_u5384_o;
  wire _al_u5385_o;
  wire _al_u5386_o;
  wire _al_u5387_o;
  wire _al_u5389_o;
  wire _al_u5390_o;
  wire _al_u5392_o;
  wire _al_u5394_o;
  wire _al_u5395_o;
  wire _al_u5396_o;
  wire _al_u5398_o;
  wire _al_u5399_o;
  wire _al_u5400_o;
  wire _al_u5403_o;
  wire _al_u5407_o;
  wire _al_u5408_o;
  wire _al_u540_o;
  wire _al_u5411_o;
  wire _al_u5412_o;
  wire _al_u5413_o;
  wire _al_u5415_o;
  wire _al_u5416_o;
  wire _al_u5417_o;
  wire _al_u5419_o;
  wire _al_u5420_o;
  wire _al_u5421_o;
  wire _al_u5424_o;
  wire _al_u5425_o;
  wire _al_u5426_o;
  wire _al_u5428_o;
  wire _al_u5429_o;
  wire _al_u5430_o;
  wire _al_u5431_o;
  wire _al_u5433_o;
  wire _al_u5435_o;
  wire _al_u5437_o;
  wire _al_u5438_o;
  wire _al_u5439_o;
  wire _al_u543_o;
  wire _al_u5441_o;
  wire _al_u5442_o;
  wire _al_u5444_o;
  wire _al_u5445_o;
  wire _al_u5446_o;
  wire _al_u5448_o;
  wire _al_u5449_o;
  wire _al_u544_o;
  wire _al_u5451_o;
  wire _al_u5452_o;
  wire _al_u5453_o;
  wire _al_u5454_o;
  wire _al_u5455_o;
  wire _al_u5457_o;
  wire _al_u5458_o;
  wire _al_u5460_o;
  wire _al_u5462_o;
  wire _al_u5463_o;
  wire _al_u5465_o;
  wire _al_u5466_o;
  wire _al_u5467_o;
  wire _al_u5468_o;
  wire _al_u546_o;
  wire _al_u5470_o;
  wire _al_u5471_o;
  wire _al_u5473_o;
  wire _al_u5474_o;
  wire _al_u5476_o;
  wire _al_u5477_o;
  wire _al_u5478_o;
  wire _al_u5479_o;
  wire _al_u5481_o;
  wire _al_u5482_o;
  wire _al_u5484_o;
  wire _al_u5485_o;
  wire _al_u5486_o;
  wire _al_u5487_o;
  wire _al_u5488_o;
  wire _al_u5489_o;
  wire _al_u5493_o;
  wire _al_u5495_o;
  wire _al_u5497_o;
  wire _al_u5498_o;
  wire _al_u5499_o;
  wire _al_u5501_o;
  wire _al_u5504_o;
  wire _al_u5505_o;
  wire _al_u5507_o;
  wire _al_u5508_o;
  wire _al_u5510_o;
  wire _al_u5511_o;
  wire _al_u5513_o;
  wire _al_u5514_o;
  wire _al_u5515_o;
  wire _al_u5516_o;
  wire _al_u5518_o;
  wire _al_u5519_o;
  wire _al_u5520_o;
  wire _al_u5522_o;
  wire _al_u5523_o;
  wire _al_u5524_o;
  wire _al_u552_o;
  wire _al_u5531_o;
  wire _al_u5532_o;
  wire _al_u5533_o;
  wire _al_u5534_o;
  wire _al_u5536_o;
  wire _al_u5537_o;
  wire _al_u5539_o;
  wire _al_u553_o;
  wire _al_u5541_o;
  wire _al_u5542_o;
  wire _al_u5544_o;
  wire _al_u5546_o;
  wire _al_u5547_o;
  wire _al_u5549_o;
  wire _al_u554_o;
  wire _al_u5550_o;
  wire _al_u5552_o;
  wire _al_u5553_o;
  wire _al_u5554_o;
  wire _al_u5556_o;
  wire _al_u5558_o;
  wire _al_u5559_o;
  wire _al_u555_o;
  wire _al_u5561_o;
  wire _al_u5562_o;
  wire _al_u5564_o;
  wire _al_u5565_o;
  wire _al_u5567_o;
  wire _al_u5568_o;
  wire _al_u556_o;
  wire _al_u5570_o;
  wire _al_u5571_o;
  wire _al_u5573_o;
  wire _al_u5574_o;
  wire _al_u5575_o;
  wire _al_u5577_o;
  wire _al_u5578_o;
  wire _al_u557_o;
  wire _al_u5580_o;
  wire _al_u5581_o;
  wire _al_u5582_o;
  wire _al_u5583_o;
  wire _al_u5584_o;
  wire _al_u5585_o;
  wire _al_u5587_o;
  wire _al_u5588_o;
  wire _al_u5590_o;
  wire _al_u5591_o;
  wire _al_u5592_o;
  wire _al_u5593_o;
  wire _al_u5594_o;
  wire _al_u5595_o;
  wire _al_u5597_o;
  wire _al_u5598_o;
  wire _al_u5599_o;
  wire _al_u5600_o;
  wire _al_u5601_o;
  wire _al_u5603_o;
  wire _al_u5604_o;
  wire _al_u5605_o;
  wire _al_u5607_o;
  wire _al_u5608_o;
  wire _al_u5609_o;
  wire _al_u560_o;
  wire _al_u5614_o;
  wire _al_u5616_o;
  wire _al_u5618_o;
  wire _al_u5619_o;
  wire _al_u5620_o;
  wire _al_u5622_o;
  wire _al_u5623_o;
  wire _al_u5625_o;
  wire _al_u5626_o;
  wire _al_u5629_o;
  wire _al_u5632_o;
  wire _al_u5633_o;
  wire _al_u5635_o;
  wire _al_u5636_o;
  wire _al_u5637_o;
  wire _al_u5638_o;
  wire _al_u5643_o;
  wire _al_u5644_o;
  wire _al_u5647_o;
  wire _al_u5648_o;
  wire _al_u5649_o;
  wire _al_u5650_o;
  wire _al_u5651_o;
  wire _al_u5652_o;
  wire _al_u5654_o;
  wire _al_u5655_o;
  wire _al_u5656_o;
  wire _al_u5657_o;
  wire _al_u5658_o;
  wire _al_u5659_o;
  wire _al_u5660_o;
  wire _al_u5661_o;
  wire _al_u5663_o;
  wire _al_u5664_o;
  wire _al_u5665_o;
  wire _al_u5666_o;
  wire _al_u5667_o;
  wire _al_u5668_o;
  wire _al_u566_o;
  wire _al_u5670_o;
  wire _al_u5671_o;
  wire _al_u5672_o;
  wire _al_u5673_o;
  wire _al_u5674_o;
  wire _al_u5675_o;
  wire _al_u5676_o;
  wire _al_u5677_o;
  wire _al_u5678_o;
  wire _al_u5679_o;
  wire _al_u5680_o;
  wire _al_u5682_o;
  wire _al_u5683_o;
  wire _al_u5684_o;
  wire _al_u5685_o;
  wire _al_u5687_o;
  wire _al_u5688_o;
  wire _al_u5689_o;
  wire _al_u5690_o;
  wire _al_u5692_o;
  wire _al_u5693_o;
  wire _al_u5694_o;
  wire _al_u5695_o;
  wire _al_u5696_o;
  wire _al_u5697_o;
  wire _al_u5698_o;
  wire _al_u5699_o;
  wire _al_u569_o;
  wire _al_u5700_o;
  wire _al_u5701_o;
  wire _al_u5702_o;
  wire _al_u5704_o;
  wire _al_u5705_o;
  wire _al_u5706_o;
  wire _al_u5707_o;
  wire _al_u5708_o;
  wire _al_u5709_o;
  wire _al_u5710_o;
  wire _al_u5711_o;
  wire _al_u5712_o;
  wire _al_u5713_o;
  wire _al_u5714_o;
  wire _al_u5715_o;
  wire _al_u5716_o;
  wire _al_u5717_o;
  wire _al_u5718_o;
  wire _al_u5719_o;
  wire _al_u571_o;
  wire _al_u5720_o;
  wire _al_u5721_o;
  wire _al_u5722_o;
  wire _al_u5723_o;
  wire _al_u5724_o;
  wire _al_u5725_o;
  wire _al_u5726_o;
  wire _al_u5727_o;
  wire _al_u5728_o;
  wire _al_u5729_o;
  wire _al_u572_o;
  wire _al_u5730_o;
  wire _al_u5731_o;
  wire _al_u5732_o;
  wire _al_u5733_o;
  wire _al_u5734_o;
  wire _al_u5735_o;
  wire _al_u5736_o;
  wire _al_u5737_o;
  wire _al_u5738_o;
  wire _al_u5739_o;
  wire _al_u573_o;
  wire _al_u5740_o;
  wire _al_u5741_o;
  wire _al_u5742_o;
  wire _al_u5743_o;
  wire _al_u5744_o;
  wire _al_u5745_o;
  wire _al_u5746_o;
  wire _al_u5747_o;
  wire _al_u5748_o;
  wire _al_u5749_o;
  wire _al_u574_o;
  wire _al_u5750_o;
  wire _al_u5751_o;
  wire _al_u5752_o;
  wire _al_u5753_o;
  wire _al_u5754_o;
  wire _al_u5755_o;
  wire _al_u5756_o;
  wire _al_u5757_o;
  wire _al_u5758_o;
  wire _al_u5759_o;
  wire _al_u575_o;
  wire _al_u5760_o;
  wire _al_u5761_o;
  wire _al_u5762_o;
  wire _al_u5763_o;
  wire _al_u5764_o;
  wire _al_u5765_o;
  wire _al_u5766_o;
  wire _al_u5767_o;
  wire _al_u5768_o;
  wire _al_u5769_o;
  wire _al_u576_o;
  wire _al_u5770_o;
  wire _al_u5771_o;
  wire _al_u5772_o;
  wire _al_u5773_o;
  wire _al_u5774_o;
  wire _al_u5775_o;
  wire _al_u5776_o;
  wire _al_u5777_o;
  wire _al_u5778_o;
  wire _al_u5779_o;
  wire _al_u5780_o;
  wire _al_u5782_o;
  wire _al_u5783_o;
  wire _al_u5784_o;
  wire _al_u5785_o;
  wire _al_u5786_o;
  wire _al_u5787_o;
  wire _al_u5788_o;
  wire _al_u5789_o;
  wire _al_u5790_o;
  wire _al_u5791_o;
  wire _al_u5792_o;
  wire _al_u5793_o;
  wire _al_u5794_o;
  wire _al_u5795_o;
  wire _al_u5796_o;
  wire _al_u5797_o;
  wire _al_u5798_o;
  wire _al_u5799_o;
  wire _al_u5800_o;
  wire _al_u5801_o;
  wire _al_u5802_o;
  wire _al_u5803_o;
  wire _al_u5804_o;
  wire _al_u5805_o;
  wire _al_u5806_o;
  wire _al_u5807_o;
  wire _al_u5808_o;
  wire _al_u5809_o;
  wire _al_u580_o;
  wire _al_u5810_o;
  wire _al_u5812_o;
  wire _al_u5813_o;
  wire _al_u5814_o;
  wire _al_u5816_o;
  wire _al_u5818_o;
  wire _al_u581_o;
  wire _al_u5820_o;
  wire _al_u5822_o;
  wire _al_u5824_o;
  wire _al_u5826_o;
  wire _al_u5828_o;
  wire _al_u582_o;
  wire _al_u5830_o;
  wire _al_u5832_o;
  wire _al_u5834_o;
  wire _al_u5836_o;
  wire _al_u5843_o;
  wire _al_u5845_o;
  wire _al_u5848_o;
  wire _al_u584_o;
  wire _al_u5850_o;
  wire _al_u5851_o;
  wire _al_u5853_o;
  wire _al_u5854_o;
  wire _al_u5856_o;
  wire _al_u5857_o;
  wire _al_u5858_o;
  wire _al_u5859_o;
  wire _al_u585_o;
  wire _al_u5860_o;
  wire _al_u5861_o;
  wire _al_u5862_o;
  wire _al_u5864_o;
  wire _al_u5865_o;
  wire _al_u5866_o;
  wire _al_u5868_o;
  wire _al_u5869_o;
  wire _al_u5870_o;
  wire _al_u5871_o;
  wire _al_u5872_o;
  wire _al_u5873_o;
  wire _al_u5874_o;
  wire _al_u5875_o;
  wire _al_u5878_o;
  wire _al_u5879_o;
  wire _al_u587_o;
  wire _al_u5880_o;
  wire _al_u5883_o;
  wire _al_u5884_o;
  wire _al_u5885_o;
  wire _al_u5886_o;
  wire _al_u5887_o;
  wire _al_u5888_o;
  wire _al_u5889_o;
  wire _al_u588_o;
  wire _al_u5890_o;
  wire _al_u5891_o;
  wire _al_u5892_o;
  wire _al_u5893_o;
  wire _al_u5894_o;
  wire _al_u5896_o;
  wire _al_u5897_o;
  wire _al_u5899_o;
  wire _al_u5900_o;
  wire _al_u5903_o;
  wire _al_u5904_o;
  wire _al_u5905_o;
  wire _al_u5906_o;
  wire _al_u5908_o;
  wire _al_u5909_o;
  wire _al_u5910_o;
  wire _al_u5911_o;
  wire _al_u5912_o;
  wire _al_u5913_o;
  wire _al_u5915_o;
  wire _al_u5916_o;
  wire _al_u5917_o;
  wire _al_u5918_o;
  wire _al_u5919_o;
  wire _al_u591_o;
  wire _al_u5920_o;
  wire _al_u5921_o;
  wire _al_u5922_o;
  wire _al_u5924_o;
  wire _al_u5925_o;
  wire _al_u5926_o;
  wire _al_u5927_o;
  wire _al_u5929_o;
  wire _al_u5930_o;
  wire _al_u5931_o;
  wire _al_u5932_o;
  wire _al_u5933_o;
  wire _al_u5934_o;
  wire _al_u5935_o;
  wire _al_u5936_o;
  wire _al_u5937_o;
  wire _al_u5938_o;
  wire _al_u593_o;
  wire _al_u5940_o;
  wire _al_u5941_o;
  wire _al_u5942_o;
  wire _al_u5943_o;
  wire _al_u5945_o;
  wire _al_u5946_o;
  wire _al_u5947_o;
  wire _al_u5948_o;
  wire _al_u5950_o;
  wire _al_u5951_o;
  wire _al_u5952_o;
  wire _al_u5953_o;
  wire _al_u5954_o;
  wire _al_u5955_o;
  wire _al_u5956_o;
  wire _al_u5957_o;
  wire _al_u5958_o;
  wire _al_u5959_o;
  wire _al_u5960_o;
  wire _al_u5961_o;
  wire _al_u5963_o;
  wire _al_u5964_o;
  wire _al_u5966_o;
  wire _al_u5968_o;
  wire _al_u5969_o;
  wire _al_u5970_o;
  wire _al_u5971_o;
  wire _al_u5972_o;
  wire _al_u5973_o;
  wire _al_u5974_o;
  wire _al_u5977_o;
  wire _al_u5979_o;
  wire _al_u597_o;
  wire _al_u5980_o;
  wire _al_u5983_o;
  wire _al_u5984_o;
  wire _al_u5985_o;
  wire _al_u5987_o;
  wire _al_u5988_o;
  wire _al_u5990_o;
  wire _al_u5991_o;
  wire _al_u5993_o;
  wire _al_u5995_o;
  wire _al_u5998_o;
  wire _al_u6000_o;
  wire _al_u6002_o;
  wire _al_u6003_o;
  wire _al_u6004_o;
  wire _al_u6005_o;
  wire _al_u6006_o;
  wire _al_u6007_o;
  wire _al_u6008_o;
  wire _al_u6009_o;
  wire _al_u6010_o;
  wire _al_u6011_o;
  wire _al_u6013_o;
  wire _al_u6014_o;
  wire _al_u6015_o;
  wire _al_u6016_o;
  wire _al_u6017_o;
  wire _al_u6018_o;
  wire _al_u6021_o;
  wire _al_u6023_o;
  wire _al_u6024_o;
  wire _al_u6025_o;
  wire _al_u6026_o;
  wire _al_u6027_o;
  wire _al_u6028_o;
  wire _al_u6029_o;
  wire _al_u6030_o;
  wire _al_u6032_o;
  wire _al_u6033_o;
  wire _al_u6034_o;
  wire _al_u6035_o;
  wire _al_u6036_o;
  wire _al_u6037_o;
  wire _al_u6039_o;
  wire _al_u6040_o;
  wire _al_u6041_o;
  wire _al_u6042_o;
  wire _al_u6043_o;
  wire _al_u6044_o;
  wire _al_u6045_o;
  wire _al_u6046_o;
  wire _al_u6047_o;
  wire _al_u6049_o;
  wire _al_u604_o;
  wire _al_u6050_o;
  wire _al_u6052_o;
  wire _al_u6053_o;
  wire _al_u6054_o;
  wire _al_u6055_o;
  wire _al_u6056_o;
  wire _al_u6057_o;
  wire _al_u6059_o;
  wire _al_u6060_o;
  wire _al_u6061_o;
  wire _al_u6062_o;
  wire _al_u6063_o;
  wire _al_u6064_o;
  wire _al_u6065_o;
  wire _al_u6066_o;
  wire _al_u6067_o;
  wire _al_u6068_o;
  wire _al_u6069_o;
  wire _al_u606_o;
  wire _al_u6070_o;
  wire _al_u6071_o;
  wire _al_u6073_o;
  wire _al_u6074_o;
  wire _al_u6075_o;
  wire _al_u6076_o;
  wire _al_u6077_o;
  wire _al_u6078_o;
  wire _al_u6079_o;
  wire _al_u607_o;
  wire _al_u6080_o;
  wire _al_u6081_o;
  wire _al_u6082_o;
  wire _al_u6084_o;
  wire _al_u6085_o;
  wire _al_u6086_o;
  wire _al_u6087_o;
  wire _al_u6088_o;
  wire _al_u6089_o;
  wire _al_u6091_o;
  wire _al_u6092_o;
  wire _al_u6094_o;
  wire _al_u6095_o;
  wire _al_u6096_o;
  wire _al_u6099_o;
  wire _al_u609_o;
  wire _al_u6100_o;
  wire _al_u6101_o;
  wire _al_u6102_o;
  wire _al_u6103_o;
  wire _al_u6104_o;
  wire _al_u6105_o;
  wire _al_u6106_o;
  wire _al_u6108_o;
  wire _al_u6109_o;
  wire _al_u6112_o;
  wire _al_u6113_o;
  wire _al_u6115_o;
  wire _al_u6116_o;
  wire _al_u6118_o;
  wire _al_u6120_o;
  wire _al_u6121_o;
  wire _al_u6122_o;
  wire _al_u6123_o;
  wire _al_u6124_o;
  wire _al_u6125_o;
  wire _al_u6127_o;
  wire _al_u6128_o;
  wire _al_u6129_o;
  wire _al_u6130_o;
  wire _al_u6133_o;
  wire _al_u6134_o;
  wire _al_u6135_o;
  wire _al_u6137_o;
  wire _al_u6138_o;
  wire _al_u6139_o;
  wire _al_u6141_o;
  wire _al_u6142_o;
  wire _al_u6144_o;
  wire _al_u6145_o;
  wire _al_u6147_o;
  wire _al_u6149_o;
  wire _al_u6150_o;
  wire _al_u6151_o;
  wire _al_u6153_o;
  wire _al_u6154_o;
  wire _al_u6155_o;
  wire _al_u6157_o;
  wire _al_u6158_o;
  wire _al_u6159_o;
  wire _al_u6160_o;
  wire _al_u6161_o;
  wire _al_u6163_o;
  wire _al_u6164_o;
  wire _al_u6166_o;
  wire _al_u6167_o;
  wire _al_u6168_o;
  wire _al_u6169_o;
  wire _al_u6170_o;
  wire _al_u6171_o;
  wire _al_u6172_o;
  wire _al_u6173_o;
  wire _al_u6174_o;
  wire _al_u6175_o;
  wire _al_u6176_o;
  wire _al_u6177_o;
  wire _al_u6180_o;
  wire _al_u6181_o;
  wire _al_u6182_o;
  wire _al_u6183_o;
  wire _al_u6184_o;
  wire _al_u6185_o;
  wire _al_u6186_o;
  wire _al_u6187_o;
  wire _al_u6188_o;
  wire _al_u6189_o;
  wire _al_u6190_o;
  wire _al_u6191_o;
  wire _al_u6192_o;
  wire _al_u6193_o;
  wire _al_u6194_o;
  wire _al_u6196_o;
  wire _al_u6197_o;
  wire _al_u6198_o;
  wire _al_u6200_o;
  wire _al_u6201_o;
  wire _al_u6202_o;
  wire _al_u6203_o;
  wire _al_u6205_o;
  wire _al_u6206_o;
  wire _al_u6207_o;
  wire _al_u6208_o;
  wire _al_u6210_o;
  wire _al_u6211_o;
  wire _al_u6214_o;
  wire _al_u6216_o;
  wire _al_u6217_o;
  wire _al_u6218_o;
  wire _al_u6219_o;
  wire _al_u6220_o;
  wire _al_u6222_o;
  wire _al_u6225_o;
  wire _al_u6226_o;
  wire _al_u6227_o;
  wire _al_u6228_o;
  wire _al_u6229_o;
  wire _al_u6230_o;
  wire _al_u6231_o;
  wire _al_u6232_o;
  wire _al_u6233_o;
  wire _al_u6234_o;
  wire _al_u6235_o;
  wire _al_u6236_o;
  wire _al_u6237_o;
  wire _al_u6238_o;
  wire _al_u6240_o;
  wire _al_u6241_o;
  wire _al_u6242_o;
  wire _al_u6243_o;
  wire _al_u6244_o;
  wire _al_u6246_o;
  wire _al_u6248_o;
  wire _al_u6249_o;
  wire _al_u6251_o;
  wire _al_u6252_o;
  wire _al_u6253_o;
  wire _al_u6254_o;
  wire _al_u6255_o;
  wire _al_u6256_o;
  wire _al_u6257_o;
  wire _al_u6258_o;
  wire _al_u6259_o;
  wire _al_u6260_o;
  wire _al_u6261_o;
  wire _al_u6262_o;
  wire _al_u6263_o;
  wire _al_u6264_o;
  wire _al_u6265_o;
  wire _al_u6266_o;
  wire _al_u6267_o;
  wire _al_u6268_o;
  wire _al_u6269_o;
  wire _al_u6271_o;
  wire _al_u6273_o;
  wire _al_u6274_o;
  wire _al_u6275_o;
  wire _al_u6276_o;
  wire _al_u6277_o;
  wire _al_u6278_o;
  wire _al_u6279_o;
  wire _al_u6280_o;
  wire _al_u6281_o;
  wire _al_u6284_o;
  wire _al_u6285_o;
  wire _al_u6286_o;
  wire _al_u6287_o;
  wire _al_u6288_o;
  wire _al_u6289_o;
  wire _al_u6290_o;
  wire _al_u6291_o;
  wire _al_u6292_o;
  wire _al_u6293_o;
  wire _al_u6294_o;
  wire _al_u6295_o;
  wire _al_u6296_o;
  wire _al_u6298_o;
  wire _al_u6300_o;
  wire _al_u6302_o;
  wire _al_u6304_o;
  wire _al_u6306_o;
  wire _al_u6307_o;
  wire _al_u6308_o;
  wire _al_u6310_o;
  wire _al_u6311_o;
  wire _al_u6312_o;
  wire _al_u6313_o;
  wire _al_u6314_o;
  wire _al_u6315_o;
  wire _al_u6316_o;
  wire _al_u6317_o;
  wire _al_u6318_o;
  wire _al_u6319_o;
  wire _al_u6320_o;
  wire _al_u6321_o;
  wire _al_u6322_o;
  wire _al_u6323_o;
  wire _al_u6324_o;
  wire _al_u6325_o;
  wire _al_u6326_o;
  wire _al_u6327_o;
  wire _al_u6328_o;
  wire _al_u6329_o;
  wire _al_u6331_o;
  wire _al_u6332_o;
  wire _al_u6333_o;
  wire _al_u6335_o;
  wire _al_u6336_o;
  wire _al_u6337_o;
  wire _al_u6338_o;
  wire _al_u6339_o;
  wire _al_u6341_o;
  wire _al_u6342_o;
  wire _al_u6343_o;
  wire _al_u6344_o;
  wire _al_u6345_o;
  wire _al_u6347_o;
  wire _al_u6348_o;
  wire _al_u6349_o;
  wire _al_u6350_o;
  wire _al_u6351_o;
  wire _al_u6352_o;
  wire _al_u6353_o;
  wire _al_u6354_o;
  wire _al_u6355_o;
  wire _al_u6356_o;
  wire _al_u6357_o;
  wire _al_u6358_o;
  wire _al_u6360_o;
  wire _al_u6361_o;
  wire _al_u6362_o;
  wire _al_u6363_o;
  wire _al_u6364_o;
  wire _al_u6365_o;
  wire _al_u6367_o;
  wire _al_u6368_o;
  wire _al_u6369_o;
  wire _al_u6370_o;
  wire _al_u6371_o;
  wire _al_u6372_o;
  wire _al_u6373_o;
  wire _al_u637_o;
  wire _al_u6380_o;
  wire _al_u6381_o;
  wire _al_u6382_o;
  wire _al_u6383_o;
  wire _al_u6384_o;
  wire _al_u6385_o;
  wire _al_u6388_o;
  wire _al_u6389_o;
  wire _al_u6390_o;
  wire _al_u6392_o;
  wire _al_u6393_o;
  wire _al_u6394_o;
  wire _al_u6395_o;
  wire _al_u6396_o;
  wire _al_u6397_o;
  wire _al_u6398_o;
  wire _al_u6399_o;
  wire _al_u6400_o;
  wire _al_u6401_o;
  wire _al_u6402_o;
  wire _al_u6403_o;
  wire _al_u6404_o;
  wire _al_u6405_o;
  wire _al_u6406_o;
  wire _al_u6407_o;
  wire _al_u6408_o;
  wire _al_u6409_o;
  wire _al_u6410_o;
  wire _al_u6411_o;
  wire _al_u6412_o;
  wire _al_u6413_o;
  wire _al_u6416_o;
  wire _al_u6417_o;
  wire _al_u6418_o;
  wire _al_u6419_o;
  wire _al_u6420_o;
  wire _al_u6421_o;
  wire _al_u6422_o;
  wire _al_u6423_o;
  wire _al_u6431_o;
  wire _al_u6432_o;
  wire _al_u6433_o;
  wire _al_u6434_o;
  wire _al_u6435_o;
  wire _al_u6436_o;
  wire _al_u6437_o;
  wire _al_u6438_o;
  wire _al_u6439_o;
  wire _al_u6440_o;
  wire _al_u6441_o;
  wire _al_u6442_o;
  wire _al_u6443_o;
  wire _al_u6444_o;
  wire _al_u6446_o;
  wire _al_u6447_o;
  wire _al_u6448_o;
  wire _al_u6449_o;
  wire _al_u6450_o;
  wire _al_u6451_o;
  wire _al_u6452_o;
  wire _al_u6453_o;
  wire _al_u6454_o;
  wire _al_u6455_o;
  wire _al_u6457_o;
  wire _al_u6458_o;
  wire _al_u6459_o;
  wire _al_u6460_o;
  wire _al_u6461_o;
  wire _al_u6463_o;
  wire _al_u6464_o;
  wire _al_u6467_o;
  wire _al_u6468_o;
  wire _al_u6469_o;
  wire _al_u6471_o;
  wire _al_u6472_o;
  wire _al_u6473_o;
  wire _al_u6475_o;
  wire _al_u6476_o;
  wire _al_u6477_o;
  wire _al_u6478_o;
  wire _al_u6479_o;
  wire _al_u6480_o;
  wire _al_u6481_o;
  wire _al_u6482_o;
  wire _al_u6483_o;
  wire _al_u6484_o;
  wire _al_u6491_o;
  wire _al_u6492_o;
  wire _al_u6493_o;
  wire _al_u6494_o;
  wire _al_u6495_o;
  wire _al_u6497_o;
  wire _al_u6498_o;
  wire _al_u6499_o;
  wire _al_u6500_o;
  wire _al_u6501_o;
  wire _al_u6502_o;
  wire _al_u6503_o;
  wire _al_u6504_o;
  wire _al_u6505_o;
  wire _al_u6507_o;
  wire _al_u6508_o;
  wire _al_u6509_o;
  wire _al_u650_o;
  wire _al_u6510_o;
  wire _al_u6511_o;
  wire _al_u6512_o;
  wire _al_u6513_o;
  wire _al_u6515_o;
  wire _al_u6518_o;
  wire _al_u6519_o;
  wire _al_u6520_o;
  wire _al_u6521_o;
  wire _al_u6522_o;
  wire _al_u6524_o;
  wire _al_u6525_o;
  wire _al_u6526_o;
  wire _al_u6527_o;
  wire _al_u6528_o;
  wire _al_u6529_o;
  wire _al_u6530_o;
  wire _al_u6531_o;
  wire _al_u6532_o;
  wire _al_u6533_o;
  wire _al_u6534_o;
  wire _al_u6535_o;
  wire _al_u6538_o;
  wire _al_u6540_o;
  wire _al_u6541_o;
  wire _al_u6542_o;
  wire _al_u6543_o;
  wire _al_u6544_o;
  wire _al_u6545_o;
  wire _al_u6546_o;
  wire _al_u6547_o;
  wire _al_u6548_o;
  wire _al_u6549_o;
  wire _al_u6550_o;
  wire _al_u6551_o;
  wire _al_u6552_o;
  wire _al_u6553_o;
  wire _al_u6554_o;
  wire _al_u6555_o;
  wire _al_u6556_o;
  wire _al_u6557_o;
  wire _al_u6558_o;
  wire _al_u6560_o;
  wire _al_u6562_o;
  wire _al_u6563_o;
  wire _al_u6564_o;
  wire _al_u6565_o;
  wire _al_u6566_o;
  wire _al_u6567_o;
  wire _al_u6568_o;
  wire _al_u6569_o;
  wire _al_u6570_o;
  wire _al_u6571_o;
  wire _al_u6572_o;
  wire _al_u6573_o;
  wire _al_u6574_o;
  wire _al_u6575_o;
  wire _al_u6576_o;
  wire _al_u6577_o;
  wire _al_u6578_o;
  wire _al_u6579_o;
  wire _al_u6580_o;
  wire _al_u6581_o;
  wire _al_u6582_o;
  wire _al_u6583_o;
  wire _al_u6584_o;
  wire _al_u6586_o;
  wire _al_u6587_o;
  wire _al_u6588_o;
  wire _al_u6589_o;
  wire _al_u6590_o;
  wire _al_u6591_o;
  wire _al_u6592_o;
  wire _al_u6593_o;
  wire _al_u6596_o;
  wire _al_u6599_o;
  wire _al_u6600_o;
  wire _al_u6601_o;
  wire _al_u6602_o;
  wire _al_u6603_o;
  wire _al_u6604_o;
  wire _al_u6605_o;
  wire _al_u6610_o;
  wire _al_u6611_o;
  wire _al_u6612_o;
  wire _al_u6614_o;
  wire _al_u6615_o;
  wire _al_u6616_o;
  wire _al_u6617_o;
  wire _al_u6619_o;
  wire _al_u6620_o;
  wire _al_u6621_o;
  wire _al_u6624_o;
  wire _al_u6625_o;
  wire _al_u6626_o;
  wire _al_u6627_o;
  wire _al_u6628_o;
  wire _al_u6629_o;
  wire _al_u6631_o;
  wire _al_u6632_o;
  wire _al_u6633_o;
  wire _al_u6634_o;
  wire _al_u6635_o;
  wire _al_u6636_o;
  wire _al_u6637_o;
  wire _al_u6638_o;
  wire _al_u6639_o;
  wire _al_u6640_o;
  wire _al_u6641_o;
  wire _al_u6643_o;
  wire _al_u6645_o;
  wire _al_u6646_o;
  wire _al_u6647_o;
  wire _al_u6648_o;
  wire _al_u6649_o;
  wire _al_u6650_o;
  wire _al_u6651_o;
  wire _al_u6652_o;
  wire _al_u6653_o;
  wire _al_u6654_o;
  wire _al_u6655_o;
  wire _al_u6656_o;
  wire _al_u6658_o;
  wire _al_u6659_o;
  wire _al_u6660_o;
  wire _al_u6661_o;
  wire _al_u6662_o;
  wire _al_u6663_o;
  wire _al_u6664_o;
  wire _al_u6665_o;
  wire _al_u6666_o;
  wire _al_u6667_o;
  wire _al_u6668_o;
  wire _al_u6669_o;
  wire _al_u6670_o;
  wire _al_u6672_o;
  wire _al_u6673_o;
  wire _al_u6674_o;
  wire _al_u6675_o;
  wire _al_u6676_o;
  wire _al_u6677_o;
  wire _al_u6679_o;
  wire _al_u6680_o;
  wire _al_u6681_o;
  wire _al_u6682_o;
  wire _al_u6683_o;
  wire _al_u6684_o;
  wire _al_u6686_o;
  wire _al_u6687_o;
  wire _al_u6688_o;
  wire _al_u6689_o;
  wire _al_u6690_o;
  wire _al_u6691_o;
  wire _al_u6692_o;
  wire _al_u6693_o;
  wire _al_u6694_o;
  wire _al_u6695_o;
  wire _al_u6696_o;
  wire _al_u6697_o;
  wire _al_u6698_o;
  wire _al_u6699_o;
  wire _al_u6700_o;
  wire _al_u6701_o;
  wire _al_u6702_o;
  wire _al_u6703_o;
  wire _al_u6706_o;
  wire _al_u6708_o;
  wire _al_u6709_o;
  wire _al_u6710_o;
  wire _al_u6711_o;
  wire _al_u6712_o;
  wire _al_u6713_o;
  wire _al_u6714_o;
  wire _al_u6715_o;
  wire _al_u6716_o;
  wire _al_u6717_o;
  wire _al_u6718_o;
  wire _al_u6719_o;
  wire _al_u6720_o;
  wire _al_u6721_o;
  wire _al_u6722_o;
  wire _al_u6723_o;
  wire _al_u6724_o;
  wire _al_u6725_o;
  wire _al_u6727_o;
  wire _al_u6728_o;
  wire _al_u6729_o;
  wire _al_u6730_o;
  wire _al_u6731_o;
  wire _al_u6732_o;
  wire _al_u6733_o;
  wire _al_u6734_o;
  wire _al_u6735_o;
  wire _al_u6737_o;
  wire _al_u6738_o;
  wire _al_u6740_o;
  wire _al_u6741_o;
  wire _al_u6742_o;
  wire _al_u6743_o;
  wire _al_u6744_o;
  wire _al_u6745_o;
  wire _al_u6746_o;
  wire _al_u6749_o;
  wire _al_u6751_o;
  wire _al_u6752_o;
  wire _al_u6753_o;
  wire _al_u6754_o;
  wire _al_u6755_o;
  wire _al_u6756_o;
  wire _al_u6757_o;
  wire _al_u6758_o;
  wire _al_u6759_o;
  wire _al_u6760_o;
  wire _al_u6761_o;
  wire _al_u6762_o;
  wire _al_u6765_o;
  wire _al_u6767_o;
  wire _al_u6769_o;
  wire _al_u6771_o;
  wire _al_u6773_o;
  wire _al_u6775_o;
  wire _al_u6776_o;
  wire _al_u6778_o;
  wire _al_u677_o;
  wire _al_u6780_o;
  wire _al_u6782_o;
  wire _al_u6784_o;
  wire _al_u6786_o;
  wire _al_u6788_o;
  wire _al_u678_o;
  wire _al_u6790_o;
  wire _al_u6792_o;
  wire _al_u6794_o;
  wire _al_u6795_o;
  wire _al_u6796_o;
  wire _al_u6797_o;
  wire _al_u6798_o;
  wire _al_u6799_o;
  wire _al_u679_o;
  wire _al_u6800_o;
  wire _al_u6801_o;
  wire _al_u6802_o;
  wire _al_u6803_o;
  wire _al_u6805_o;
  wire _al_u6806_o;
  wire _al_u6807_o;
  wire _al_u6808_o;
  wire _al_u6809_o;
  wire _al_u680_o;
  wire _al_u6810_o;
  wire _al_u6811_o;
  wire _al_u6812_o;
  wire _al_u6814_o;
  wire _al_u6817_o;
  wire _al_u6819_o;
  wire _al_u681_o;
  wire _al_u6820_o;
  wire _al_u6821_o;
  wire _al_u6822_o;
  wire _al_u6823_o;
  wire _al_u6824_o;
  wire _al_u6825_o;
  wire _al_u6826_o;
  wire _al_u6827_o;
  wire _al_u6828_o;
  wire _al_u6829_o;
  wire _al_u682_o;
  wire _al_u6830_o;
  wire _al_u6832_o;
  wire _al_u6833_o;
  wire _al_u6836_o;
  wire _al_u6838_o;
  wire _al_u6841_o;
  wire _al_u6842_o;
  wire _al_u6844_o;
  wire _al_u6846_o;
  wire _al_u6848_o;
  wire _al_u6850_o;
  wire _al_u6852_o;
  wire _al_u6853_o;
  wire _al_u6855_o;
  wire _al_u6856_o;
  wire _al_u6857_o;
  wire _al_u6858_o;
  wire _al_u6859_o;
  wire _al_u685_o;
  wire _al_u6861_o;
  wire _al_u6866_o;
  wire _al_u6867_o;
  wire _al_u6868_o;
  wire _al_u6869_o;
  wire _al_u6870_o;
  wire _al_u6871_o;
  wire _al_u6872_o;
  wire _al_u6874_o;
  wire _al_u6875_o;
  wire _al_u6876_o;
  wire _al_u6878_o;
  wire _al_u6879_o;
  wire _al_u6881_o;
  wire _al_u6882_o;
  wire _al_u6884_o;
  wire _al_u6885_o;
  wire _al_u6887_o;
  wire _al_u6888_o;
  wire _al_u6890_o;
  wire _al_u6891_o;
  wire _al_u6892_o;
  wire _al_u6894_o;
  wire _al_u6897_o;
  wire _al_u6898_o;
  wire _al_u6900_o;
  wire _al_u6901_o;
  wire _al_u6903_o;
  wire _al_u6904_o;
  wire _al_u6907_o;
  wire _al_u6908_o;
  wire _al_u6910_o;
  wire _al_u6913_o;
  wire _al_u6914_o;
  wire _al_u6915_o;
  wire _al_u6917_o;
  wire _al_u6918_o;
  wire _al_u6920_o;
  wire _al_u6921_o;
  wire _al_u6923_o;
  wire _al_u6924_o;
  wire _al_u6925_o;
  wire _al_u6926_o;
  wire _al_u6929_o;
  wire _al_u692_o;
  wire _al_u6930_o;
  wire _al_u6931_o;
  wire _al_u6932_o;
  wire _al_u6934_o;
  wire _al_u6935_o;
  wire _al_u6937_o;
  wire _al_u6938_o;
  wire _al_u6941_o;
  wire _al_u6942_o;
  wire _al_u6945_o;
  wire _al_u6946_o;
  wire _al_u6947_o;
  wire _al_u6948_o;
  wire _al_u6949_o;
  wire _al_u6950_o;
  wire _al_u6951_o;
  wire _al_u6952_o;
  wire _al_u6953_o;
  wire _al_u6954_o;
  wire _al_u6956_o;
  wire _al_u6957_o;
  wire _al_u6958_o;
  wire _al_u695_o;
  wire _al_u6960_o;
  wire _al_u6961_o;
  wire _al_u6962_o;
  wire _al_u6964_o;
  wire _al_u6965_o;
  wire _al_u6966_o;
  wire _al_u6967_o;
  wire _al_u6968_o;
  wire _al_u6969_o;
  wire _al_u696_o;
  wire _al_u6970_o;
  wire _al_u6972_o;
  wire _al_u6975_o;
  wire _al_u6977_o;
  wire _al_u6978_o;
  wire _al_u6979_o;
  wire _al_u697_o;
  wire _al_u6980_o;
  wire _al_u6981_o;
  wire _al_u6983_o;
  wire _al_u6984_o;
  wire _al_u6985_o;
  wire _al_u6987_o;
  wire _al_u6988_o;
  wire _al_u6989_o;
  wire _al_u698_o;
  wire _al_u6992_o;
  wire _al_u6993_o;
  wire _al_u6994_o;
  wire _al_u6996_o;
  wire _al_u6997_o;
  wire _al_u6998_o;
  wire _al_u7000_o;
  wire _al_u7001_o;
  wire _al_u7002_o;
  wire _al_u7005_o;
  wire _al_u7006_o;
  wire _al_u7008_o;
  wire _al_u7009_o;
  wire _al_u700_o;
  wire _al_u7010_o;
  wire _al_u7012_o;
  wire _al_u7013_o;
  wire _al_u7014_o;
  wire _al_u7015_o;
  wire _al_u7016_o;
  wire _al_u7018_o;
  wire _al_u7020_o;
  wire _al_u7021_o;
  wire _al_u7022_o;
  wire _al_u7023_o;
  wire _al_u7024_o;
  wire _al_u7025_o;
  wire _al_u7027_o;
  wire _al_u7028_o;
  wire _al_u702_o;
  wire _al_u7030_o;
  wire _al_u7031_o;
  wire _al_u7032_o;
  wire _al_u7034_o;
  wire _al_u7035_o;
  wire _al_u7036_o;
  wire _al_u7038_o;
  wire _al_u7039_o;
  wire _al_u7040_o;
  wire _al_u7041_o;
  wire _al_u7044_o;
  wire _al_u7045_o;
  wire _al_u7047_o;
  wire _al_u7048_o;
  wire _al_u7049_o;
  wire _al_u7051_o;
  wire _al_u7052_o;
  wire _al_u7053_o;
  wire _al_u7056_o;
  wire _al_u7057_o;
  wire _al_u7059_o;
  wire _al_u705_o;
  wire _al_u7060_o;
  wire _al_u7062_o;
  wire _al_u7064_o;
  wire _al_u7065_o;
  wire _al_u7068_o;
  wire _al_u7069_o;
  wire _al_u7071_o;
  wire _al_u7072_o;
  wire _al_u7074_o;
  wire _al_u7075_o;
  wire _al_u7077_o;
  wire _al_u7078_o;
  wire _al_u7080_o;
  wire _al_u7081_o;
  wire _al_u7083_o;
  wire _al_u7084_o;
  wire _al_u7085_o;
  wire _al_u7087_o;
  wire _al_u7088_o;
  wire _al_u7090_o;
  wire _al_u7092_o;
  wire _al_u7093_o;
  wire _al_u7094_o;
  wire _al_u7096_o;
  wire _al_u7097_o;
  wire _al_u7099_o;
  wire _al_u7100_o;
  wire _al_u7101_o;
  wire _al_u7103_o;
  wire _al_u7104_o;
  wire _al_u7105_o;
  wire _al_u7108_o;
  wire _al_u7109_o;
  wire _al_u7112_o;
  wire _al_u7113_o;
  wire _al_u7116_o;
  wire _al_u7117_o;
  wire _al_u7119_o;
  wire _al_u711_o;
  wire _al_u7120_o;
  wire _al_u7121_o;
  wire _al_u7122_o;
  wire _al_u7124_o;
  wire _al_u7125_o;
  wire _al_u7126_o;
  wire _al_u7128_o;
  wire _al_u7130_o;
  wire _al_u7131_o;
  wire _al_u7133_o;
  wire _al_u7135_o;
  wire _al_u7137_o;
  wire _al_u7139_o;
  wire _al_u7141_o;
  wire _al_u7144_o;
  wire _al_u7146_o;
  wire _al_u7148_o;
  wire _al_u714_o;
  wire _al_u7151_o;
  wire _al_u7154_o;
  wire _al_u7157_o;
  wire _al_u7160_o;
  wire _al_u7163_o;
  wire _al_u7166_o;
  wire _al_u7169_o;
  wire _al_u7172_o;
  wire _al_u7175_o;
  wire _al_u7178_o;
  wire _al_u717_o;
  wire _al_u7181_o;
  wire _al_u7184_o;
  wire _al_u7187_o;
  wire _al_u718_o;
  wire _al_u7190_o;
  wire _al_u7193_o;
  wire _al_u7195_o;
  wire _al_u7198_o;
  wire _al_u719_o;
  wire _al_u7201_o;
  wire _al_u7204_o;
  wire _al_u7206_o;
  wire _al_u7207_o;
  wire _al_u7208_o;
  wire _al_u720_o;
  wire _al_u7211_o;
  wire _al_u7214_o;
  wire _al_u7217_o;
  wire _al_u7220_o;
  wire _al_u7222_o;
  wire _al_u7223_o;
  wire _al_u7224_o;
  wire _al_u7225_o;
  wire _al_u723_o;
  wire _al_u725_o;
  wire _al_u726_o;
  wire _al_u729_o;
  wire _al_u731_o;
  wire _al_u732_o;
  wire _al_u735_o;
  wire _al_u736_o;
  wire _al_u737_o;
  wire _al_u738_o;
  wire _al_u741_o;
  wire _al_u742_o;
  wire _al_u744_o;
  wire _al_u747_o;
  wire _al_u749_o;
  wire _al_u750_o;
  wire _al_u753_o;
  wire _al_u754_o;
  wire _al_u755_o;
  wire _al_u756_o;
  wire _al_u759_o;
  wire _al_u760_o;
  wire _al_u761_o;
  wire _al_u762_o;
  wire _al_u765_o;
  wire _al_u766_o;
  wire _al_u767_o;
  wire _al_u768_o;
  wire _al_u771_o;
  wire _al_u772_o;
  wire _al_u774_o;
  wire _al_u777_o;
  wire _al_u778_o;
  wire _al_u779_o;
  wire _al_u780_o;
  wire _al_u783_o;
  wire _al_u786_o;
  wire _al_u789_o;
  wire _al_u790_o;
  wire _al_u792_o;
  wire _al_u795_o;
  wire _al_u796_o;
  wire _al_u797_o;
  wire _al_u798_o;
  wire _al_u801_o;
  wire _al_u802_o;
  wire _al_u804_o;
  wire _al_u807_o;
  wire _al_u808_o;
  wire _al_u809_o;
  wire _al_u813_o;
  wire _al_u814_o;
  wire _al_u815_o;
  wire _al_u816_o;
  wire _al_u819_o;
  wire _al_u821_o;
  wire _al_u822_o;
  wire _al_u823_o;
  wire _al_u825_o;
  wire _al_u828_o;
  wire _al_u831_o;
  wire _al_u832_o;
  wire _al_u833_o;
  wire _al_u837_o;
  wire _al_u839_o;
  wire _al_u840_o;
  wire _al_u843_o;
  wire _al_u844_o;
  wire _al_u846_o;
  wire _al_u849_o;
  wire _al_u850_o;
  wire _al_u851_o;
  wire _al_u852_o;
  wire _al_u855_o;
  wire _al_u858_o;
  wire _al_u861_o;
  wire _al_u862_o;
  wire _al_u864_o;
  wire _al_u867_o;
  wire _al_u868_o;
  wire _al_u869_o;
  wire _al_u870_o;
  wire _al_u873_o;
  wire _al_u874_o;
  wire _al_u875_o;
  wire _al_u876_o;
  wire _al_u879_o;
  wire _al_u880_o;
  wire _al_u882_o;
  wire _al_u885_o;
  wire _al_u886_o;
  wire _al_u887_o;
  wire _al_u888_o;
  wire _al_u891_o;
  wire _al_u892_o;
  wire _al_u894_o;
  wire _al_u897_o;
  wire _al_u898_o;
  wire _al_u899_o;
  wire _al_u900_o;
  wire _al_u903_o;
  wire _al_u904_o;
  wire _al_u906_o;
  wire _al_u908_o;
  wire _al_u909_o;
  wire _al_u912_o;
  wire _al_u913_o;
  wire _al_u914_o;
  wire _al_u916_o;
  wire _al_u920_o;
  wire _al_u922_o;
  wire _al_u923_o;
  wire _al_u924_o;
  wire _al_u925_o;
  wire _al_u926_o;
  wire _al_u927_o;
  wire _al_u930_o;
  wire _al_u931_o;
  wire _al_u932_o;
  wire _al_u933_o;
  wire _al_u935_o;
  wire _al_u938_o;
  wire _al_u939_o;
  wire _al_u940_o;
  wire _al_u941_o;
  wire _al_u942_o;
  wire _al_u944_o;
  wire _al_u945_o;
  wire _al_u946_o;
  wire _al_u948_o;
  wire _al_u951_o;
  wire _al_u952_o;
  wire _al_u953_o;
  wire _al_u954_o;
  wire _al_u955_o;
  wire _al_u956_o;
  wire _al_u958_o;
  wire _al_u960_o;
  wire _al_u963_o;
  wire _al_u964_o;
  wire _al_u965_o;
  wire _al_u966_o;
  wire _al_u967_o;
  wire _al_u968_o;
  wire _al_u970_o;
  wire _al_u972_o;
  wire _al_u975_o;
  wire _al_u976_o;
  wire _al_u977_o;
  wire _al_u978_o;
  wire _al_u979_o;
  wire _al_u980_o;
  wire _al_u982_o;
  wire _al_u984_o;
  wire _al_u987_o;
  wire _al_u988_o;
  wire _al_u989_o;
  wire _al_u990_o;
  wire _al_u991_o;
  wire _al_u992_o;
  wire _al_u994_o;
  wire _al_u996_o;
  wire _al_u999_o;
  wire \u1/c0 ;
  wire \u1/c1 ;
  wire \u1/c10 ;
  wire \u1/c11 ;
  wire \u1/c12 ;
  wire \u1/c13 ;
  wire \u1/c2 ;
  wire \u1/c3 ;
  wire \u1/c4 ;
  wire \u1/c5 ;
  wire \u1/c6 ;
  wire \u1/c7 ;
  wire \u1/c8 ;
  wire \u1/c9 ;
  wire \u2/c0 ;
  wire \u2/c1 ;
  wire \u2/c10 ;
  wire \u2/c11 ;
  wire \u2/c12 ;
  wire \u2/c13 ;
  wire \u2/c2 ;
  wire \u2/c3 ;
  wire \u2/c4 ;
  wire \u2/c5 ;
  wire \u2/c6 ;
  wire \u2/c7 ;
  wire \u2/c8 ;
  wire \u2/c9 ;
  wire \u_M0clkpll/clk0_buf ;  // al_ip/M0clkpll.v(34)
  wire \u_cmsdk_mcu/HWRITE ;  // ../RTL/cmsdk_mcu.v(106)
  wire \u_cmsdk_mcu/LOCKUPRESET ;  // ../RTL/cmsdk_mcu.v(86)
  wire \u_cmsdk_mcu/SYSRESETREQ ;  // ../RTL/cmsdk_mcu.v(78)
  wire \u_cmsdk_mcu/dbg_swdo ;  // ../RTL/cmsdk_mcu.v(166)
  wire \u_cmsdk_mcu/dbg_swdo_en ;  // ../RTL/cmsdk_mcu.v(165)
  wire \u_cmsdk_mcu/flash_hsel ;  // ../RTL/cmsdk_mcu.v(111)
  wire \u_cmsdk_mcu/n1 ;
  wire \u_cmsdk_mcu/sram_hsel ;  // ../RTL/cmsdk_mcu.v(117)
  wire \u_cmsdk_mcu/u_ahb_ram/mux3_b0_sel_is_2_o ;
  wire \u_cmsdk_mcu/u_ahb_ram/n16 ;
  wire \u_cmsdk_mcu/u_ahb_ram/n2 ;
  wire \u_cmsdk_mcu/u_ahb_ram/we ;  // ../RTL/AHB2MEM.v(29)
  wire \u_cmsdk_mcu/u_ahb_rom/n16 ;
  wire \u_cmsdk_mcu/u_ahb_rom/n2 ;
  wire \u_cmsdk_mcu/u_ahb_rom/we ;  // ../RTL/AHB2MEM.v(29)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/dbgrst_reg ;  // ../RTL/cmsdk_mcu_clkctrl.v(66)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/nxt_hrst ;  // ../RTL/cmsdk_mcu_clkctrl.v(65)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ;  // ../RTL/cmsdk_mcu_clkctrl.v(67)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/DBGRESTARTED ;  // ../RTL/cmsdk_mcu_system.v(171)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/HADDR[27]_lutinv ;  // ../RTL/cmsdk_mcu_system.v(80)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/SLEEPHOLDACKn ;  // ../RTL/cmsdk_mcu_system.v(121)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/apbsys_hreadyout ;  // ../RTL/cmsdk_mcu_system.v(251)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/apbsys_hsel ;  // ../RTL/cmsdk_mcu_system.v(250)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/cpu0cdbgpwrupreq ;  // ../RTL/cmsdk_mcu_system.v(342)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_hsel ;  // ../RTL/cmsdk_mcu_system.v(255)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/gpio1_hsel ;  // ../RTL/cmsdk_mcu_system.v(260)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/remap_ctrl ;  // ../RTL/cmsdk_mcu_system.v(301)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/sysctrl_hsel ;  // ../RTL/cmsdk_mcu_system.v(265)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/sysrom_hsel ;  // ../RTL/cmsdk_mcu_system.v(286)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOSEL ;  // ../RTL/cmsdk_ahb_gpio.v(75)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOTRANS ;  // ../RTL/cmsdk_ahb_gpio.v(79)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOWRITE ;  // ../RTL/cmsdk_ahb_gpio.v(77)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_ahb_to_gpio/n0 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/mux4_b10_sel_is_4_o ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n101 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n103 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n105 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n107 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n109 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n111 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n113 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n115 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n117 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n119 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n121 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n123 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n125 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n127 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n129 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n12_lutinv ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n133 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n136 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n144 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n146 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n148 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n150 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n152 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n154 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n156 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n158 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n160 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n162 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n164 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n166 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n168 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n170 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n172 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n174 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n178 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n181 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n189 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n191 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n193 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n195 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n197 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n199 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n201 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n203 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n205 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n207 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n209 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n211 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n213 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n215 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n217 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n219 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n223 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n226 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n234 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n236 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n238 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n240 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n242 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n244 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n246 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n248 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n24_lutinv ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n250 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n252 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n254 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n256 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n258 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n260 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n262 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n264 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n26_lutinv ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n271 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n273 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n275 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n277 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n279 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n281 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n283 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n285 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n287 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n289 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n291 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n293 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n295 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n297 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n299 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n301 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n34 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n39 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n43 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n46 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n54 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n56 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n58 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n60 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n62 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n64 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n66 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n68 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n70 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n72 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n74 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n76 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n78 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n80 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n82 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n84 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n88 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n91 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n99 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_dout_normal_write0 ;  // ../RTL/cmsdk_iop_gpio.v(265)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_dout_normal_write1 ;  // ../RTL/cmsdk_iop_gpio.v(266)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intclr_normal_write0 ;  // ../RTL/cmsdk_iop_gpio.v(514)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intclr_normal_write1 ;  // ../RTL/cmsdk_iop_gpio.v(515)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[0] ;  // ../RTL/cmsdk_ahb_gpio.v(67)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[10] ;  // ../RTL/cmsdk_ahb_gpio.v(67)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[11] ;  // ../RTL/cmsdk_ahb_gpio.v(67)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[12] ;  // ../RTL/cmsdk_ahb_gpio.v(67)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[13] ;  // ../RTL/cmsdk_ahb_gpio.v(67)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[14] ;  // ../RTL/cmsdk_ahb_gpio.v(67)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[15] ;  // ../RTL/cmsdk_ahb_gpio.v(67)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[1] ;  // ../RTL/cmsdk_ahb_gpio.v(67)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[2] ;  // ../RTL/cmsdk_ahb_gpio.v(67)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[3] ;  // ../RTL/cmsdk_ahb_gpio.v(67)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[4] ;  // ../RTL/cmsdk_ahb_gpio.v(67)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[5] ;  // ../RTL/cmsdk_ahb_gpio.v(67)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[6] ;  // ../RTL/cmsdk_ahb_gpio.v(67)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[7] ;  // ../RTL/cmsdk_ahb_gpio.v(67)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[8] ;  // ../RTL/cmsdk_ahb_gpio.v(67)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[9] ;  // ../RTL/cmsdk_ahb_gpio.v(67)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/IOSEL ;  // ../RTL/cmsdk_ahb_gpio.v(75)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_ahb_to_gpio/n0 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n101 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n103 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n105 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n107 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n109 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n111 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n113 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n115 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n117 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n119 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n121 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n123 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n125 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n127 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n129 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n133 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n136 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n144 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n146 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n148 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n150 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n152 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n154 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n156 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n158 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n160 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n162 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n164 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n166 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n168 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n170 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n172 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n174 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n178 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n181 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n189 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n191 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n193 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n195 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n197 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n199 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n201 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n203 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n205 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n207 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n209 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n211 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n213 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n215 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n217 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n219 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n223 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n226 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n234 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n236 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n238 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n240 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n242 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n244 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n246 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n248 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n250 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n252 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n254 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n256 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n258 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n260 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n262 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n264 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n271 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n273 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n275 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n277 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n279 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n281 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n283 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n285 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n287 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n289 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n291 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n293 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n295 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n297 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n299 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n301 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n304 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n34 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n39 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n43 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n46 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n54 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n56 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n58 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n60 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n62 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n64 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n66 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n68 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n70 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n72 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n74 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n76 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n78 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n80 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n82 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n84 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n88 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n91 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n99 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_dout_normal_write0 ;  // ../RTL/cmsdk_iop_gpio.v(265)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_dout_normal_write1 ;  // ../RTL/cmsdk_iop_gpio.v(266)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intclr_normal_write0 ;  // ../RTL/cmsdk_iop_gpio.v(514)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intclr_normal_write1 ;  // ../RTL/cmsdk_iop_gpio.v(515)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n11 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n43 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[10] ;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(104)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[11] ;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(104)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] ;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(104)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] ;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(104)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[4] ;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(104)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[5] ;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(104)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[6] ;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(104)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[7] ;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(104)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[8] ;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(104)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[9] ;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(104)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PWRITE ;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(105)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_ls_sync ;  // ../RTL/gpio.v(68)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n12_lutinv ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n40 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n43 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n49 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n52 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n55 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n58 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n6 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n61 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n63 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n68 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/n28 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/n36 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/n44 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/n52 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/n60 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/n68 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/n76 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/n84 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/BAUDTICK ;  // ../RTL/cmsdk_apb_uart.v(76)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add0/c0 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add0/c1 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add0/c2 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add0/c3 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add1/c0 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add1/c1 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add1/c2 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add1/c3 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add2/c0 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add2/c1 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add2/c2 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add2/c3 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add3/c0 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add3/c1 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add3/c2 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add3/c3 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/baud_updated ;  // ../RTL/cmsdk_apb_uart.v(128)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/lt0_c0 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/lt0_c1 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/lt0_c2 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/lt0_c3 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/lt0_c4 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/lt2/o_1_lutinv ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/mux4_b6_sel_is_13_o ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/mux9_b10_sel_is_3_o ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n100 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n106 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n114 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n117 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n17 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n20 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n25_lutinv ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n27_lutinv ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n31 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n38 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n40_lutinv ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n44 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n46 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n48 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n50 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n53 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n61 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n63 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n74 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n7_lutinv ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n88_lutinv ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n9_lutinv ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_rx_buf_full ;  // ../RTL/cmsdk_apb_uart.v(185)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_rx_overrun ;  // ../RTL/cmsdk_apb_uart.v(139)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_tx_overrun ;  // ../RTL/cmsdk_apb_uart.v(140)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_txd ;  // ../RTL/cmsdk_apb_uart.v(163)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/read_enable ;  // ../RTL/cmsdk_apb_uart.v(102)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_rx_overrun ;  // ../RTL/cmsdk_apb_uart.v(135)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_tx_overrun ;  // ../RTL/cmsdk_apb_uart.v(137)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reload_i ;  // ../RTL/cmsdk_apb_uart.v(129)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_buf_full ;  // ../RTL/cmsdk_apb_uart.v(184)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_overrun ;  // ../RTL/cmsdk_apb_uart.v(136)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_shift_in ;  // ../RTL/cmsdk_apb_uart.v(172)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_state_inc ;  // ../RTL/cmsdk_apb_uart.v(181)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_state_update ;  // ../RTL/cmsdk_apb_uart.v(177)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rxbuf_sample ;  // ../RTL/cmsdk_apb_uart.v(186)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rxd_sync_1 ;  // ../RTL/cmsdk_apb_uart.v(168)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rxd_sync_2 ;  // ../RTL/cmsdk_apb_uart.v(169)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/c0 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/c1 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/c10 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/c11 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/c12 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/c13 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/c14 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/c15 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/c2 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/c3 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/c4 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/c5 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/c6 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/c7 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/c8 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/c9 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub1/c0 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub1/c1 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub1/c2 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub1/c3 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_buf_full ;  // ../RTL/cmsdk_apb_uart.v(161)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_overrun ;  // ../RTL/cmsdk_apb_uart.v(138)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_state_inc ;  // ../RTL/cmsdk_apb_uart.v(154)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_state_update ;  // ../RTL/cmsdk_apb_uart.v(153)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/update_reg_txd ;  // ../RTL/cmsdk_apb_uart.v(164)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/update_rx_tick_cnt ;  // ../RTL/cmsdk_apb_uart.v(180)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/write_enable ;  // ../RTL/cmsdk_apb_uart.v(103)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/write_enable00 ;  // ../RTL/cmsdk_apb_uart.v(104)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/write_enable08 ;  // ../RTL/cmsdk_apb_uart.v(106)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/write_enable0c ;  // ../RTL/cmsdk_apb_uart.v(107)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/write_enable10 ;  // ../RTL/cmsdk_apb_uart.v(108)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/n1 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/apb_tran_end ;  // ../RTL/cmsdk_ahb_to_apb.v(88)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_apb_slave_mux/n0 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_apb_slave_mux/n4 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/uart0_txovrint ;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(248)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/ahb_access ;  // ../RTL/cmsdk_mcu_sysctrl.v(116)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/ahb_read ;  // ../RTL/cmsdk_mcu_sysctrl.v(118)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/ahb_write ;  // ../RTL/cmsdk_mcu_sysctrl.v(117)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/mux4_b6_sel_is_13_o ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/mux6_b3_sel_is_2_o ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/n34_lutinv ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_lockupreset_write ;  // ../RTL/cmsdk_mcu_sysctrl.v(280)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_read_enable ;  // ../RTL/cmsdk_mcu_sysctrl.v(121)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_remap_write ;  // ../RTL/cmsdk_mcu_sysctrl.v(240)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_resetinfo_en ;  // ../RTL/cmsdk_mcu_sysctrl.v(309)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_resetinfo_write ;  // ../RTL/cmsdk_mcu_sysctrl.v(297)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_write_enable ;  // ../RTL/cmsdk_mcu_sysctrl.v(122)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/HALTED ;  // ../RTL/CORTEXM0INTEGRATION.v(70)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A00iu6 ;  // ../RTL/cortexm0ds_logic.v(303)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A0fow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1047)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A0mow6 ;  // ../RTL/cortexm0ds_logic.v(1141)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A1zhu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(290)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A25iu6 ;  // ../RTL/cortexm0ds_logic.v(371)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A2cpw6 ;  // ../RTL/cortexm0ds_logic.v(1489)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A2lhu6 ;  // ../RTL/cortexm0ds_logic.v(138)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A2qiu6 ;  // ../RTL/cortexm0ds_logic.v(652)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A2yhu6 ;  // ../RTL/cortexm0ds_logic.v(277)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A3biu6 ;  // ../RTL/cortexm0ds_logic.v(452)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A3iiu6 ;  // ../RTL/cortexm0ds_logic.v(545)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A3ipw6 ;  // ../RTL/cortexm0ds_logic.v(1584)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A3xhu6 ;  // ../RTL/cortexm0ds_logic.v(264)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A4phu6 ;  // ../RTL/cortexm0ds_logic.v(158)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A4pow6 ;  // ../RTL/cortexm0ds_logic.v(1182)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A59pw6 ;  // ../RTL/cortexm0ds_logic.v(1450)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A5ipw6 ;  // ../RTL/cortexm0ds_logic.v(1584)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A5vhu6 ;  // ../RTL/cortexm0ds_logic.v(238)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A6cbx6 ;  // ../RTL/cortexm0ds_logic.v(1701)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A70iu6 ;  // ../RTL/cortexm0ds_logic.v(306)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A85ju6_lutinv ;  // ../RTL/cortexm0ds_logic.v(855)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A8ihu6 ;  // ../RTL/cortexm0ds_logic.v(130)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A95iu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(374)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A9rhu6 ;  // ../RTL/cortexm0ds_logic.v(186)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A9row6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1211)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aa2bx6 ;  // ../RTL/cortexm0ds_logic.v(1683)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aaiiu6 ;  // ../RTL/cortexm0ds_logic.v(548)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ab9ax6 ;  // ../RTL/cortexm0ds_logic.v(1630)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Abphu6 ;  // ../RTL/cortexm0ds_logic.v(160)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Acebx6 ;  // ../RTL/cortexm0ds_logic.v(1705)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Acohu6 ;  // ../RTL/cortexm0ds_logic.v(147)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Acvhu6 ;  // ../RTL/cortexm0ds_logic.v(241)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ad7ax6 ;  // ../RTL/cortexm0ds_logic.v(1626)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ad8pw6 ;  // ../RTL/cortexm0ds_logic.v(1440)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Admiu6 ;  // ../RTL/cortexm0ds_logic.v(602)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aduhu6 ;  // ../RTL/cortexm0ds_logic.v(228)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(309)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae7iu6 ;  // ../RTL/cortexm0ds_logic.v(402)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Afkiu6 ;  // ../RTL/cortexm0ds_logic.v(576)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ag5iu6 ;  // ../RTL/cortexm0ds_logic.v(376)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Agjiu6 ;  // ../RTL/cortexm0ds_logic.v(563)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Agyhu6 ;  // ../RTL/cortexm0ds_logic.v(283)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahcow6 ;  // ../RTL/cortexm0ds_logic.v(1013)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahdax6 ;  // ../RTL/cortexm0ds_logic.v(1638)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahdbx6 ;  // ../RTL/cortexm0ds_logic.v(1704)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahlpw6 ;  // ../RTL/cortexm0ds_logic.v(1590)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahqow6 ;  // ../RTL/cortexm0ds_logic.v(1200)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahwiu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(738)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ai2ju6_lutinv ;  // ../RTL/cortexm0ds_logic.v(818)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aj1ju6 ;  // ../RTL/cortexm0ds_logic.v(805)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ajgiu6 ;  // ../RTL/cortexm0ds_logic.v(524)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ajohu6 ;  // ../RTL/cortexm0ds_logic.v(150)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Akuow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1255)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Alkhu6 ;  // ../RTL/cortexm0ds_logic.v(137)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Alziu6 ;  // ../RTL/cortexm0ds_logic.v(779)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Am5ju6_lutinv ;  // ../RTL/cortexm0ds_logic.v(860)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Am6iu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(392)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Am7ow6 ;  // ../RTL/cortexm0ds_logic.v(948)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Amsow6 ;  // ../RTL/cortexm0ds_logic.v(1229)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Amupw6 ;  // ../RTL/cortexm0ds_logic.v(1607)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Anciu6 ;  // ../RTL/cortexm0ds_logic.v(472)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Anrhu6 ;  // ../RTL/cortexm0ds_logic.v(192)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aoeax6 ;  // ../RTL/cortexm0ds_logic.v(1640)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Apaiu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(446)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Apcax6 ;  // ../RTL/cortexm0ds_logic.v(1636)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aphiu6 ;  // ../RTL/cortexm0ds_logic.v(540)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Apihu6 ;  // ../RTL/cortexm0ds_logic.v(132)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aq2pw6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1364)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aqgiu6 ;  // ../RTL/cortexm0ds_logic.v(527)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aqniu6 ;  // ../RTL/cortexm0ds_logic.v(621)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ar1bx6 ;  // ../RTL/cortexm0ds_logic.v(1682)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ar1iu6 ;  // ../RTL/cortexm0ds_logic.v(327)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Asupw6 ;  // ../RTL/cortexm0ds_logic.v(1607)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/At2bx6 ;  // ../RTL/cortexm0ds_logic.v(1684)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujiu6 ;  // ../RTL/cortexm0ds_logic.v(569)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 ;  // ../RTL/cortexm0ds_logic.v(1587)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Auyax6 ;  // ../RTL/cortexm0ds_logic.v(1677)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Av3ju6 ;  // ../RTL/cortexm0ds_logic.v(836)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Avwiu6 ;  // ../RTL/cortexm0ds_logic.v(743)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Avzax6 ;  // ../RTL/cortexm0ds_logic.v(1679)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aw4bx6 ;  // ../RTL/cortexm0ds_logic.v(1688)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Awwow6 ;  // ../RTL/cortexm0ds_logic.v(1286)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Axohu6 ;  // ../RTL/cortexm0ds_logic.v(155)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ay1iu6 ;  // ../RTL/cortexm0ds_logic.v(329)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ay8iu6 ;  // ../RTL/cortexm0ds_logic.v(423)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ayuhu6 ;  // ../RTL/cortexm0ds_logic.v(236)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Az3bx6 ;  // ../RTL/cortexm0ds_logic.v(1686)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Azeiu6 ;  // ../RTL/cortexm0ds_logic.v(504)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Azliu6 ;  // ../RTL/cortexm0ds_logic.v(597)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B0biu6 ;  // ../RTL/cortexm0ds_logic.v(450)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B0cow6 ;  // ../RTL/cortexm0ds_logic.v(1007)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B0iiu6 ;  // ../RTL/cortexm0ds_logic.v(544)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B1phu6 ;  // ../RTL/cortexm0ds_logic.v(157)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B29iu6 ;  // ../RTL/cortexm0ds_logic.v(424)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B2vhu6 ;  // ../RTL/cortexm0ds_logic.v(237)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B3fiu6 ;  // ../RTL/cortexm0ds_logic.v(505)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B3gbx6 ;  // ../RTL/cortexm0ds_logic.v(1708)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B40iu6 ;  // ../RTL/cortexm0ds_logic.v(305)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B4epw6 ;  // ../RTL/cortexm0ds_logic.v(1516)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B4fow6 ;  // ../RTL/cortexm0ds_logic.v(1048)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B4mow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1142)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B6dow6 ;  // ../RTL/cortexm0ds_logic.v(1022)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B74iu6 ;  // ../RTL/cortexm0ds_logic.v(359)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B79bx6 ;  // ../RTL/cortexm0ds_logic.v(1696)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B7lpw6 ;  // ../RTL/cortexm0ds_logic.v(1590)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B7xhu6 ;  // ../RTL/cortexm0ds_logic.v(266)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B8bow6 ;  // ../RTL/cortexm0ds_logic.v(996)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B8phu6 ;  // ../RTL/cortexm0ds_logic.v(159)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B91ju6 ;  // ../RTL/cortexm0ds_logic.v(801)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B9eax6 ;  // ../RTL/cortexm0ds_logic.v(1639)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B9jbx6 ;  // ../RTL/cortexm0ds_logic.v(1714)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bagow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1064)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bamiu6 ;  // ../RTL/cortexm0ds_logic.v(601)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bauhu6 ;  // ../RTL/cortexm0ds_logic.v(227)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bb0iu6 ;  // ../RTL/cortexm0ds_logic.v(307)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bbliu6 ;  // ../RTL/cortexm0ds_logic.v(588)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bc3bx6 ;  // ../RTL/cortexm0ds_logic.v(1685)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bcabx6 ;  // ../RTL/cortexm0ds_logic.v(1698)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bccax6 ;  // ../RTL/cortexm0ds_logic.v(1636)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bcdbx6 ;  // ../RTL/cortexm0ds_logic.v(1703)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bcgax6 ;  // ../RTL/cortexm0ds_logic.v(1643)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bciax6 ;  // ../RTL/cortexm0ds_logic.v(1647)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bclpw6 ;  // ../RTL/cortexm0ds_logic.v(1590)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bddow6 ;  // ../RTL/cortexm0ds_logic.v(1025)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bewiu6 ;  // ../RTL/cortexm0ds_logic.v(736)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bf3qw6 ;  // ../RTL/cortexm0ds_logic.v(1623)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bfphu6 ;  // ../RTL/cortexm0ds_logic.v(162)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bg9iu6 ;  // ../RTL/cortexm0ds_logic.v(430)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bggiu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(523)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bgohu6 ;  // ../RTL/cortexm0ds_logic.v(149)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bguiu6 ;  // ../RTL/cortexm0ds_logic.v(710)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bi0iu6 ;  // ../RTL/cortexm0ds_logic.v(310)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Biaax6 ;  // ../RTL/cortexm0ds_logic.v(1632)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bimow6 ;  // ../RTL/cortexm0ds_logic.v(1147)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bisiu6 ;  // ../RTL/cortexm0ds_logic.v(684)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bithu6 ;  // ../RTL/cortexm0ds_logic.v(216)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bk7ax6 ;  // ../RTL/cortexm0ds_logic.v(1627)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bngax6 ;  // ../RTL/cortexm0ds_logic.v(1644)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bnohu6 ;  // ../RTL/cortexm0ds_logic.v(151)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bofiu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(513)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bomiu6 ;  // ../RTL/cortexm0ds_logic.v(606)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bouhu6 ;  // ../RTL/cortexm0ds_logic.v(232)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bp2qw6 ;  // ../RTL/cortexm0ds_logic.v(1622)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bpliu6 ;  // ../RTL/cortexm0ds_logic.v(593)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bq9ax6 ;  // ../RTL/cortexm0ds_logic.v(1631)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bqzhu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(300)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bs4iu6 ;  // ../RTL/cortexm0ds_logic.v(367)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bs4pw6 ;  // ../RTL/cortexm0ds_logic.v(1392)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bsxhu6 ;  // ../RTL/cortexm0ds_logic.v(274)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bt2qw6 ;  // ../RTL/cortexm0ds_logic.v(1622)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Btbbx6 ;  // ../RTL/cortexm0ds_logic.v(1700)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Btoiu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(635)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bu2pw6 ;  // ../RTL/cortexm0ds_logic.v(1366)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bu6bx6 ;  // ../RTL/cortexm0ds_logic.v(1691)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Buabx6 ;  // ../RTL/cortexm0ds_logic.v(1699)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Buohu6 ;  // ../RTL/cortexm0ds_logic.v(154)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bvaax6 ;  // ../RTL/cortexm0ds_logic.v(1633)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bvfbx6 ;  // ../RTL/cortexm0ds_logic.v(1708)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bvuhu6 ;  // ../RTL/cortexm0ds_logic.v(235)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bwdax6 ;  // ../RTL/cortexm0ds_logic.v(1639)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bwliu6 ;  // ../RTL/cortexm0ds_logic.v(596)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bx2qw6 ;  // ../RTL/cortexm0ds_logic.v(1622)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bxbax6 ;  // ../RTL/cortexm0ds_logic.v(1635)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bxdpw6 ;  // ../RTL/cortexm0ds_logic.v(1514)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bxeow6 ;  // ../RTL/cortexm0ds_logic.v(1046)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bxzhu6 ;  // ../RTL/cortexm0ds_logic.v(302)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/By4ju6 ;  // ../RTL/cortexm0ds_logic.v(851)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bziiu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(557)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bzxhu6 ;  // ../RTL/cortexm0ds_logic.v(276)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C07bx6 ;  // ../RTL/cortexm0ds_logic.v(1692)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C0fiu6 ;  // ../RTL/cortexm0ds_logic.v(504)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C10bx6 ;  // ../RTL/cortexm0ds_logic.v(1679)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C10iu6 ;  // ../RTL/cortexm0ds_logic.v(304)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C14bx6 ;  // ../RTL/cortexm0ds_logic.v(1686)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C1epw6 ;  // ../RTL/cortexm0ds_logic.v(1515)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C1fax6 ;  // ../RTL/cortexm0ds_logic.v(1641)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C1wpw6 ;  // ../RTL/cortexm0ds_logic.v(1610)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C2ypw6 ;  // ../RTL/cortexm0ds_logic.v(1613)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C30bx6 ;  // ../RTL/cortexm0ds_logic.v(1679)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C34ju6 ;  // ../RTL/cortexm0ds_logic.v(839)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C3wpw6 ;  // ../RTL/cortexm0ds_logic.v(1610)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C3yhu6 ;  // ../RTL/cortexm0ds_logic.v(278)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C4dax6 ;  // ../RTL/cortexm0ds_logic.v(1637)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C4ihu6 ;  // ../RTL/cortexm0ds_logic.v(130)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C4iiu6 ;  // ../RTL/cortexm0ds_logic.v(546)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C50bx6 ;  // ../RTL/cortexm0ds_logic.v(1680)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C53iu6 ;  // ../RTL/cortexm0ds_logic.v(345)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C5gbx6 ;  // ../RTL/cortexm0ds_logic.v(1708)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C5phu6 ;  // ../RTL/cortexm0ds_logic.v(158)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C6vhu6 ;  // ../RTL/cortexm0ds_logic.v(239)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C72qw6 ;  // ../RTL/cortexm0ds_logic.v(1621)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C7miu6 ;  // ../RTL/cortexm0ds_logic.v(600)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C7now6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1157)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C80iu6 ;  // ../RTL/cortexm0ds_logic.v(306)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C8fow6 ;  // ../RTL/cortexm0ds_logic.v(1050)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C8liu6 ;  // ../RTL/cortexm0ds_logic.v(587)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C96pw6 ;  // ../RTL/cortexm0ds_logic.v(1411)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ca1bx6 ;  // ../RTL/cortexm0ds_logic.v(1682)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cayhu6 ;  // ../RTL/cortexm0ds_logic.v(280)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cbbiu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(455)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cc2bx6 ;  // ../RTL/cortexm0ds_logic.v(1683)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cccbx6 ;  // ../RTL/cortexm0ds_logic.v(1701)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cchiu6 ;  // ../RTL/cortexm0ds_logic.v(535)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ccphu6 ;  // ../RTL/cortexm0ds_logic.v(161)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cdohu6 ;  // ../RTL/cortexm0ds_logic.v(148)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ceabx6 ;  // ../RTL/cortexm0ds_logic.v(1698)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cemiu6 ;  // ../RTL/cortexm0ds_logic.v(603)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cenow6 ;  // ../RTL/cortexm0ds_logic.v(1159)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ceuhu6 ;  // ../RTL/cortexm0ds_logic.v(228)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cf7iu6 ;  // ../RTL/cortexm0ds_logic.v(403)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cfliu6 ;  // ../RTL/cortexm0ds_logic.v(590)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cfthu6 ;  // ../RTL/cortexm0ds_logic.v(215)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cfvpw6 ;  // ../RTL/cortexm0ds_logic.v(1609)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cfziu6 ;  // ../RTL/cortexm0ds_logic.v(777)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cg5ju6_lutinv ;  // ../RTL/cortexm0ds_logic.v(858)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cgkiu6 ;  // ../RTL/cortexm0ds_logic.v(577)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ch5iu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(377)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Chkhu6 ;  // ../RTL/cortexm0ds_logic.v(136)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Chwpw6 ;  // ../RTL/cortexm0ds_logic.v(1610)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ciqow6 ;  // ../RTL/cortexm0ds_logic.v(1201)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cjiow6 ;  // ../RTL/cortexm0ds_logic.v(1094)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cjqpw6 ;  // ../RTL/cortexm0ds_logic.v(1600)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cjwpw6 ;  // ../RTL/cortexm0ds_logic.v(1611)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ckniu6 ;  // ../RTL/cortexm0ds_logic.v(618)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ckohu6 ;  // ../RTL/cortexm0ds_logic.v(150)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cl1iu6 ;  // ../RTL/cortexm0ds_logic.v(325)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Clihu6 ;  // ../RTL/cortexm0ds_logic.v(131)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cmthu6 ;  // ../RTL/cortexm0ds_logic.v(218)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cmziu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(780)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cn7ow6 ;  // ../RTL/cortexm0ds_logic.v(949)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cncbx6 ;  // ../RTL/cortexm0ds_logic.v(1702)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cndbx6 ;  // ../RTL/cortexm0ds_logic.v(1704)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cokbx6 ;  // ../RTL/cortexm0ds_logic.v(1717)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Coupw6 ;  // ../RTL/cortexm0ds_logic.v(1607)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cpqow6 ;  // ../RTL/cortexm0ds_logic.v(1203)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cq3qw6 ;  // ../RTL/cortexm0ds_logic.v(1624)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cqoiu6 ;  // ../RTL/cortexm0ds_logic.v(634)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Crniu6 ;  // ../RTL/cortexm0ds_logic.v(621)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Crohu6 ;  // ../RTL/cortexm0ds_logic.v(153)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cs1iu6 ;  // ../RTL/cortexm0ds_logic.v(327)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cs7ju6_lutinv ;  // ../RTL/cortexm0ds_logic.v(889)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Csmiu6 ;  // ../RTL/cortexm0ds_logic.v(608)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Csnow6 ;  // ../RTL/cortexm0ds_logic.v(1164)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Csuhu6 ;  // ../RTL/cortexm0ds_logic.v(234)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ctliu6 ;  // ../RTL/cortexm0ds_logic.v(595)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ctthu6 ;  // ../RTL/cortexm0ds_logic.v(221)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cvciu6 ;  // ../RTL/cortexm0ds_logic.v(475)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cwiiu6 ;  // ../RTL/cortexm0ds_logic.v(556)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cwxhu6 ;  // ../RTL/cortexm0ds_logic.v(275)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cwyax6 ;  // ../RTL/cortexm0ds_logic.v(1677)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cxcbx6 ;  // ../RTL/cortexm0ds_logic.v(1702)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cxzax6 ;  // ../RTL/cortexm0ds_logic.v(1679)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cy4bx6 ;  // ../RTL/cortexm0ds_logic.v(1688)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cy9iu6 ;  // ../RTL/cortexm0ds_logic.v(436)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cydbx6 ;  // ../RTL/cortexm0ds_logic.v(1704)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cykhu6 ;  // ../RTL/cortexm0ds_logic.v(138)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cyohu6 ;  // ../RTL/cortexm0ds_logic.v(156)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cz7ju6 ;  // ../RTL/cortexm0ds_logic.v(891)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cz8iu6 ;  // ../RTL/cortexm0ds_logic.v(423)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Czmiu6 ;  // ../RTL/cortexm0ds_logic.v(611)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Czuhu6 ;  // ../RTL/cortexm0ds_logic.v(236)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Czzax6 ;  // ../RTL/cortexm0ds_logic.v(1679)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D0jiu6 ;  // ../RTL/cortexm0ds_logic.v(557)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D0yhu6 ;  // ../RTL/cortexm0ds_logic.v(277)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D14pw6 ;  // ../RTL/cortexm0ds_logic.v(1382)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D1aax6 ;  // ../RTL/cortexm0ds_logic.v(1631)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D2opw6 ;  // ../RTL/cortexm0ds_logic.v(1595)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D2phu6 ;  // ../RTL/cortexm0ds_logic.v(157)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D2rpw6 ;  // ../RTL/cortexm0ds_logic.v(1601)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D31ju6 ;  // ../RTL/cortexm0ds_logic.v(799)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D39iu6 ;  // ../RTL/cortexm0ds_logic.v(425)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D3vhu6 ;  // ../RTL/cortexm0ds_logic.v(238)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D43qw6 ;  // ../RTL/cortexm0ds_logic.v(1623)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D4miu6 ;  // ../RTL/cortexm0ds_logic.v(599)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D50iu6 ;  // ../RTL/cortexm0ds_logic.v(305)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D5eiu6 ;  // ../RTL/cortexm0ds_logic.v(492)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D5epw6 ;  // ../RTL/cortexm0ds_logic.v(1517)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D6kiu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(573)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D6sow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1223)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D70bx6 ;  // ../RTL/cortexm0ds_logic.v(1680)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D7gbx6 ;  // ../RTL/cortexm0ds_logic.v(1709)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D84iu6 ;  // ../RTL/cortexm0ds_logic.v(360)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D8iiu6 ;  // ../RTL/cortexm0ds_logic.v(547)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D8xhu6 ;  // ../RTL/cortexm0ds_logic.v(266)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D99ax6 ;  // ../RTL/cortexm0ds_logic.v(1630)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D9phu6 ;  // ../RTL/cortexm0ds_logic.v(160)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Daebx6 ;  // ../RTL/cortexm0ds_logic.v(1705)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dagiu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(521)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Daiax6 ;  // ../RTL/cortexm0ds_logic.v(1647)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dbmiu6 ;  // ../RTL/cortexm0ds_logic.v(602)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dbuhu6 ;  // ../RTL/cortexm0ds_logic.v(227)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dc0iu6 ;  // ../RTL/cortexm0ds_logic.v(308)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dcziu6 ;  // ../RTL/cortexm0ds_logic.v(776)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dd7ow6 ;  // ../RTL/cortexm0ds_logic.v(945)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ddkiu6 ;  // ../RTL/cortexm0ds_logic.v(576)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Df4iu6 ;  // ../RTL/cortexm0ds_logic.v(362)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dfbax6 ;  // ../RTL/cortexm0ds_logic.v(1634)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dfqow6 ;  // ../RTL/cortexm0ds_logic.v(1200)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dg2qw6 ;  // ../RTL/cortexm0ds_logic.v(1621)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dgapw6 ;  // ../RTL/cortexm0ds_logic.v(1467)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dgphu6 ;  // ../RTL/cortexm0ds_logic.v(162)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dhniu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(617)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dhohu6 ;  // ../RTL/cortexm0ds_logic.v(149)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dhvhu6 ;  // ../RTL/cortexm0ds_logic.v(243)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Di1iu6 ;  // ../RTL/cortexm0ds_logic.v(323)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Di3qw6 ;  // ../RTL/cortexm0ds_logic.v(1624)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Difiu6 ;  // ../RTL/cortexm0ds_logic.v(511)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Djthu6 ;  // ../RTL/cortexm0ds_logic.v(217)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dk6pw6 ;  // ../RTL/cortexm0ds_logic.v(1415)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dk7ow6 ;  // ../RTL/cortexm0ds_logic.v(947)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dk9bx6 ;  // ../RTL/cortexm0ds_logic.v(1696)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dkeow6 ;  // ../RTL/cortexm0ds_logic.v(1041)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dkkiu6 ;  // ../RTL/cortexm0ds_logic.v(578)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dm6bx6 ;  // ../RTL/cortexm0ds_logic.v(1691)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dmeax6 ;  // ../RTL/cortexm0ds_logic.v(1640)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dmiiu6 ;  // ../RTL/cortexm0ds_logic.v(552)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dmqhu6 ;  // ../RTL/cortexm0ds_logic.v(178)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dmqow6 ;  // ../RTL/cortexm0ds_logic.v(1202)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dncax6 ;  // ../RTL/cortexm0ds_logic.v(1636)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Doohu6 ;  // ../RTL/cortexm0ds_logic.v(152)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dooow6 ;  // ../RTL/cortexm0ds_logic.v(1176)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dpuhu6 ;  // ../RTL/cortexm0ds_logic.v(232)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dpwpw6 ;  // ../RTL/cortexm0ds_logic.v(1611)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dqfhu6 ;  // ../RTL/cortexm0ds_logic.v(125)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dqthu6 ;  // ../RTL/cortexm0ds_logic.v(219)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dr7ow6 ;  // ../RTL/cortexm0ds_logic.v(950)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Drcbx6 ;  // ../RTL/cortexm0ds_logic.v(1702)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Drhhu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(129)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Drkiu6 ;  // ../RTL/cortexm0ds_logic.v(581)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Drzow6 ;  // ../RTL/cortexm0ds_logic.v(1324)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ds4ju6_lutinv ;  // ../RTL/cortexm0ds_logic.v(849)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dsrhu6 ;  // ../RTL/cortexm0ds_logic.v(193)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dt1bx6 ;  // ../RTL/cortexm0ds_logic.v(1682)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dt4iu6 ;  // ../RTL/cortexm0ds_logic.v(368)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dtjow6 ;  // ../RTL/cortexm0ds_logic.v(1111)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dtxhu6 ;  // ../RTL/cortexm0ds_logic.v(274)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dugax6 ;  // ../RTL/cortexm0ds_logic.v(1644)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dv2bx6 ;  // ../RTL/cortexm0ds_logic.v(1684)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dv9iu6 ;  // ../RTL/cortexm0ds_logic.v(435)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dw1iu6 ;  // ../RTL/cortexm0ds_logic.v(329)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dwuhu6 ;  // ../RTL/cortexm0ds_logic.v(235)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 ;  // ../RTL/cortexm0ds_logic.v(1609)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dyeow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1046)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dyzhu6 ;  // ../RTL/cortexm0ds_logic.v(303)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dzdow6 ;  // ../RTL/cortexm0ds_logic.v(1033)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dzvpw6 ;  // ../RTL/cortexm0ds_logic.v(1610)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E05bx6 ;  // ../RTL/cortexm0ds_logic.v(1688)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E0ihu6 ;  // ../RTL/cortexm0ds_logic.v(130)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E0vhu6 ;  // ../RTL/cortexm0ds_logic.v(237)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E17ju6_lutinv ;  // ../RTL/cortexm0ds_logic.v(879)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E18iu6 ;  // ../RTL/cortexm0ds_logic.v(411)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E1fiu6 ;  // ../RTL/cortexm0ds_logic.v(504)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E1miu6 ;  // ../RTL/cortexm0ds_logic.v(598)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E20iu6 ;  // ../RTL/cortexm0ds_logic.v(304)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E2epw6 ;  // ../RTL/cortexm0ds_logic.v(1516)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E2liu6 ;  // ../RTL/cortexm0ds_logic.v(585)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E34bx6 ;  // ../RTL/cortexm0ds_logic.v(1686)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E3sow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1222)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E4yhu6 ;  // ../RTL/cortexm0ds_logic.v(278)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E4yow6 ;  // ../RTL/cortexm0ds_logic.v(1303)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E54iu6 ;  // ../RTL/cortexm0ds_logic.v(359)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E5jow6 ;  // ../RTL/cortexm0ds_logic.v(1102)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E6iax6 ;  // ../RTL/cortexm0ds_logic.v(1647)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E7vhu6 ;  // ../RTL/cortexm0ds_logic.v(239)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E8iax6 ;  // ../RTL/cortexm0ds_logic.v(1647)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E8miu6 ;  // ../RTL/cortexm0ds_logic.v(601)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E8now6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1157)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E8uow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1251)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E90bx6 ;  // ../RTL/cortexm0ds_logic.v(1680)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E90iu6 ;  // ../RTL/cortexm0ds_logic.v(307)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E97ax6 ;  // ../RTL/cortexm0ds_logic.v(1626)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E9mow6 ;  // ../RTL/cortexm0ds_logic.v(1144)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ea7ow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(944)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eafax6 ;  // ../RTL/cortexm0ds_logic.v(1641)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eagax6 ;  // ../RTL/cortexm0ds_logic.v(1643)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eariu6 ;  // ../RTL/cortexm0ds_logic.v(668)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eazow6 ;  // ../RTL/cortexm0ds_logic.v(1318)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eblhu6 ;  // ../RTL/cortexm0ds_logic.v(139)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eccow6 ;  // ../RTL/cortexm0ds_logic.v(1011)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eciiu6 ;  // ../RTL/cortexm0ds_logic.v(549)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Edapw6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1466)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Edphu6 ;  // ../RTL/cortexm0ds_logic.v(161)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ee3bx6 ;  // ../RTL/cortexm0ds_logic.v(1685)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eegiu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(523)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eeohu6 ;  // ../RTL/cortexm0ds_logic.v(148)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ef7ju6 ;  // ../RTL/cortexm0ds_logic.v(884)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ef8iu6 ;  // ../RTL/cortexm0ds_logic.v(416)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Efdax6 ;  // ../RTL/cortexm0ds_logic.v(1638)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eg7iu6 ;  // ../RTL/cortexm0ds_logic.v(403)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Egaax6 ;  // ../RTL/cortexm0ds_logic.v(1632)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Egthu6 ;  // ../RTL/cortexm0ds_logic.v(216)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Egziu6 ;  // ../RTL/cortexm0ds_logic.v(777)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ;  // ../RTL/cortexm0ds_logic.v(390)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ehqpw6 ;  // ../RTL/cortexm0ds_logic.v(1600)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eidow6 ;  // ../RTL/cortexm0ds_logic.v(1027)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eirhu6 ;  // ../RTL/cortexm0ds_logic.v(190)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ejaju6_lutinv ;  // ../RTL/cortexm0ds_logic.v(926)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ejbpw6 ;  // ../RTL/cortexm0ds_logic.v(1482)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ejcow6 ;  // ../RTL/cortexm0ds_logic.v(1014)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ekhiu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(538)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Elgax6 ;  // ../RTL/cortexm0ds_logic.v(1644)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Elnpw6 ;  // ../RTL/cortexm0ds_logic.v(1594)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Elohu6 ;  // ../RTL/cortexm0ds_logic.v(151)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Emmiu6 ;  // ../RTL/cortexm0ds_logic.v(606)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Enthu6 ;  // ../RTL/cortexm0ds_logic.v(218)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eoyiu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(767)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ep4ju6 ;  // ../RTL/cortexm0ds_logic.v(848)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Epciu6 ;  // ../RTL/cortexm0ds_logic.v(473)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Epjiu6 ;  // ../RTL/cortexm0ds_logic.v(567)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Epyhu6 ;  // ../RTL/cortexm0ds_logic.v(286)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eq4pw6 ;  // ../RTL/cortexm0ds_logic.v(1391)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eqqow6 ;  // ../RTL/cortexm0ds_logic.v(1204)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Erbbx6 ;  // ../RTL/cortexm0ds_logic.v(1700)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eriow6 ;  // ../RTL/cortexm0ds_logic.v(1097)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Esabx6 ;  // ../RTL/cortexm0ds_logic.v(1698)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Esohu6 ;  // ../RTL/cortexm0ds_logic.v(153)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Et8iu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(421)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Etfbx6 ;  // ../RTL/cortexm0ds_logic.v(1708)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Etfiu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(515)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Etmiu6 ;  // ../RTL/cortexm0ds_logic.v(608)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Etuhu6 ;  // ../RTL/cortexm0ds_logic.v(234)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eudax6 ;  // ../RTL/cortexm0ds_logic.v(1639)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eukhu6 ;  // ../RTL/cortexm0ds_logic.v(137)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Evbax6 ;  // ../RTL/cortexm0ds_logic.v(1635)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Evhpw6 ;  // ../RTL/cortexm0ds_logic.v(1584)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Evkiu6 ;  // ../RTL/cortexm0ds_logic.v(582)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Evzhu6 ;  // ../RTL/cortexm0ds_logic.v(302)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ewjiu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(569)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ewrow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1219)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Exxhu6 ;  // ../RTL/cortexm0ds_logic.v(276)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eyihu6 ;  // ../RTL/cortexm0ds_logic.v(132)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eyyax6 ;  // ../RTL/cortexm0ds_logic.v(1677)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ez1ju6 ;  // ../RTL/cortexm0ds_logic.v(811)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ezohu6 ;  // ../RTL/cortexm0ds_logic.v(156)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F0eow6 ;  // ../RTL/cortexm0ds_logic.v(1034)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F0riu6 ;  // ../RTL/cortexm0ds_logic.v(664)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F14ju6 ;  // ../RTL/cortexm0ds_logic.v(839)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F15pw6 ;  // ../RTL/cortexm0ds_logic.v(1395)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F17ax6 ;  // ../RTL/cortexm0ds_logic.v(1626)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F1jiu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(558)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F1yhu6 ;  // ../RTL/cortexm0ds_logic.v(277)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F24iu6 ;  // ../RTL/cortexm0ds_logic.v(358)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F26bx6 ;  // ../RTL/cortexm0ds_logic.v(1690)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F2dax6 ;  // ../RTL/cortexm0ds_logic.v(1637)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F2xhu6 ;  // ../RTL/cortexm0ds_logic.v(264)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F3phu6 ;  // ../RTL/cortexm0ds_logic.v(157)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F42iu6 ;  // ../RTL/cortexm0ds_logic.v(332)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F4iax6 ;  // ../RTL/cortexm0ds_logic.v(1647)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F4ibx6 ;  // ../RTL/cortexm0ds_logic.v(1712)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F4vhu6 ;  // ../RTL/cortexm0ds_logic.v(238)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F57ju6_lutinv ;  // ../RTL/cortexm0ds_logic.v(880)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F58iu6 ;  // ../RTL/cortexm0ds_logic.v(412)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F59bx6 ;  // ../RTL/cortexm0ds_logic.v(1695)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F5miu6 ;  // ../RTL/cortexm0ds_logic.v(599)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F5uow6 ;  // ../RTL/cortexm0ds_logic.v(1249)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F60iu6 ;  // ../RTL/cortexm0ds_logic.v(306)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F6dbx6 ;  // ../RTL/cortexm0ds_logic.v(1703)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F6eiu6 ;  // ../RTL/cortexm0ds_logic.v(493)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F6ziu6 ;  // ../RTL/cortexm0ds_logic.v(774)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F7eax6 ;  // ../RTL/cortexm0ds_logic.v(1639)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F7jbx6 ;  // ../RTL/cortexm0ds_logic.v(1714)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F7zhu6 ;  // ../RTL/cortexm0ds_logic.v(293)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F85iu6 ;  // ../RTL/cortexm0ds_logic.v(373)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F8cbx6 ;  // ../RTL/cortexm0ds_logic.v(1701)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F8dbx6 ;  // ../RTL/cortexm0ds_logic.v(1703)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F8row6 ;  // ../RTL/cortexm0ds_logic.v(1210)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F94iu6 ;  // ../RTL/cortexm0ds_logic.v(360)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F9gbx6 ;  // ../RTL/cortexm0ds_logic.v(1709)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F9vpw6 ;  // ../RTL/cortexm0ds_logic.v(1608)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Facax6 ;  // ../RTL/cortexm0ds_logic.v(1636)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Facbx6 ;  // ../RTL/cortexm0ds_logic.v(1701)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Faoiu6 ;  // ../RTL/cortexm0ds_logic.v(628)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Faphu6 ;  // ../RTL/cortexm0ds_logic.v(160)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fb0bx6 ;  // ../RTL/cortexm0ds_logic.v(1680)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fb1ju6 ;  // ../RTL/cortexm0ds_logic.v(802)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fbvhu6 ;  // ../RTL/cortexm0ds_logic.v(241)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fc1bx6 ;  // ../RTL/cortexm0ds_logic.v(1682)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fcuhu6 ;  // ../RTL/cortexm0ds_logic.v(228)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fd7iu6 ;  // ../RTL/cortexm0ds_logic.v(402)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fdfow6 ;  // ../RTL/cortexm0ds_logic.v(1052)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fe2bx6 ;  // ../RTL/cortexm0ds_logic.v(1683)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ffqiu6 ;  // ../RTL/cortexm0ds_logic.v(657)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ffrow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1213)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ffyhu6 ;  // ../RTL/cortexm0ds_logic.v(282)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fgpiu6 ;  // ../RTL/cortexm0ds_logic.v(644)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fgqow6 ;  // ../RTL/cortexm0ds_logic.v(1200)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fhoiu6 ;  // ../RTL/cortexm0ds_logic.v(631)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fi1ju6 ;  // ../RTL/cortexm0ds_logic.v(805)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Finiu6 ;  // ../RTL/cortexm0ds_logic.v(618)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fivhu6 ;  // ../RTL/cortexm0ds_logic.v(243)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fj1iu6 ;  // ../RTL/cortexm0ds_logic.v(324)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fj8ax6 ;  // ../RTL/cortexm0ds_logic.v(1628)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fjdbx6 ;  // ../RTL/cortexm0ds_logic.v(1704)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fkliu6 ;  // ../RTL/cortexm0ds_logic.v(592)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fkrpw6 ;  // ../RTL/cortexm0ds_logic.v(1602)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fl2qw6 ;  // ../RTL/cortexm0ds_logic.v(1622)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fldbx6 ;  // ../RTL/cortexm0ds_logic.v(1704)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fllow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1135)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Flyiu6 ;  // ../RTL/cortexm0ds_logic.v(766)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fm6ow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(935)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fm7ax6 ;  // ../RTL/cortexm0ds_logic.v(1627)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fnnpw6 ;  // ../RTL/cortexm0ds_logic.v(1594)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fnpiu6 ;  // ../RTL/cortexm0ds_logic.v(646)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fnqow6 ;  // ../RTL/cortexm0ds_logic.v(1203)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fnwiu6 ;  // ../RTL/cortexm0ds_logic.v(740)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fo9ax6 ;  // ../RTL/cortexm0ds_logic.v(1631)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fpaow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(989)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fpgiu6 ;  // ../RTL/cortexm0ds_logic.v(527)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fpnpw6 ;  // ../RTL/cortexm0ds_logic.v(1595)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fpohu6 ;  // ../RTL/cortexm0ds_logic.v(152)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fquhu6 ;  // ../RTL/cortexm0ds_logic.v(233)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Frthu6 ;  // ../RTL/cortexm0ds_logic.v(220)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Frziu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(781)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fs6iu6 ;  // ../RTL/cortexm0ds_logic.v(394)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fsdiu6 ;  // ../RTL/cortexm0ds_logic.v(488)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ftaax6 ;  // ../RTL/cortexm0ds_logic.v(1633)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fucow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1018)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fuxhu6 ;  // ../RTL/cortexm0ds_logic.v(274)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fvcbx6 ;  // ../RTL/cortexm0ds_logic.v(1702)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fviow6 ;  // ../RTL/cortexm0ds_logic.v(1099)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fwohu6 ;  // ../RTL/cortexm0ds_logic.v(155)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fx9ow6 ;  // ../RTL/cortexm0ds_logic.v(979)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fxuhu6 ;  // ../RTL/cortexm0ds_logic.v(235)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fy8ow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(966)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fyliu6 ;  // ../RTL/cortexm0ds_logic.v(597)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fzkiu6 ;  // ../RTL/cortexm0ds_logic.v(584)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fzsow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1234)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fzzhu6 ;  // ../RTL/cortexm0ds_logic.v(303)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G0phu6 ;  // ../RTL/cortexm0ds_logic.v(156)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G0pow6 ;  // ../RTL/cortexm0ds_logic.v(1181)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G0zax6 ;  // ../RTL/cortexm0ds_logic.v(1678)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G1aow6 ;  // ../RTL/cortexm0ds_logic.v(981)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G1vhu6 ;  // ../RTL/cortexm0ds_logic.v(237)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G25bx6 ;  // ../RTL/cortexm0ds_logic.v(1688)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G2fiu6 ;  // ../RTL/cortexm0ds_logic.v(505)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G2iax6 ;  // ../RTL/cortexm0ds_logic.v(1647)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G2miu6 ;  // ../RTL/cortexm0ds_logic.v(598)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G30iu6 ;  // ../RTL/cortexm0ds_logic.v(305)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G3eiu6 ;  // ../RTL/cortexm0ds_logic.v(492)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G3epw6 ;  // ../RTL/cortexm0ds_logic.v(1516)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G54bx6 ;  // ../RTL/cortexm0ds_logic.v(1686)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G64iu6 ;  // ../RTL/cortexm0ds_logic.v(359)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G6cow6 ;  // ../RTL/cortexm0ds_logic.v(1009)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G6xhu6 ;  // ../RTL/cortexm0ds_logic.v(266)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G6xow6 ;  // ../RTL/cortexm0ds_logic.v(1290)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G79ax6 ;  // ../RTL/cortexm0ds_logic.v(1630)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G7aiu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(440)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G7lhu6 ;  // ../RTL/cortexm0ds_logic.v(138)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G7phu6 ;  // ../RTL/cortexm0ds_logic.v(159)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G81ju6 ;  // ../RTL/cortexm0ds_logic.v(801)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G8ebx6 ;  // ../RTL/cortexm0ds_logic.v(1705)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G8how6 ;  // ../RTL/cortexm0ds_logic.v(1077)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G8vhu6 ;  // ../RTL/cortexm0ds_logic.v(240)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G9fiu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(507)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G9uhu6 ;  // ../RTL/cortexm0ds_logic.v(227)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G9uow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1251)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ga0iu6 ;  // ../RTL/cortexm0ds_logic.v(307)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gbvpw6 ;  // ../RTL/cortexm0ds_logic.v(1608)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gc1qw6 ;  // ../RTL/cortexm0ds_logic.v(1619)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gc6ow6 ;  // ../RTL/cortexm0ds_logic.v(931)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gcjiu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(562)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gd0bx6 ;  // ../RTL/cortexm0ds_logic.v(1680)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gd4pw6 ;  // ../RTL/cortexm0ds_logic.v(1386)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gdihu6 ;  // ../RTL/cortexm0ds_logic.v(131)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gdjow6 ;  // ../RTL/cortexm0ds_logic.v(1105)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gdqow6 ;  // ../RTL/cortexm0ds_logic.v(1199)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gebow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(999)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gephu6 ;  // ../RTL/cortexm0ds_logic.v(162)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gf1ju6 ;  // ../RTL/cortexm0ds_logic.v(804)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gfniu6 ;  // ../RTL/cortexm0ds_logic.v(617)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gfvhu6 ;  // ../RTL/cortexm0ds_logic.v(242)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ggabx6 ;  // ../RTL/cortexm0ds_logic.v(1698)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gggow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1066)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gglhu6 ;  // ../RTL/cortexm0ds_logic.v(139)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ghthu6 ;  // ../RTL/cortexm0ds_logic.v(216)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gihbx6 ;  // ../RTL/cortexm0ds_logic.v(1711)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gk3ju6_lutinv ;  // ../RTL/cortexm0ds_logic.v(832)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gk4iu6 ;  // ../RTL/cortexm0ds_logic.v(364)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gk4pw6 ;  // ../RTL/cortexm0ds_logic.v(1389)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gkcow6 ;  // ../RTL/cortexm0ds_logic.v(1014)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gkeax6 ;  // ../RTL/cortexm0ds_logic.v(1640)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gkqow6 ;  // ../RTL/cortexm0ds_logic.v(1202)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gkwiu6 ;  // ../RTL/cortexm0ds_logic.v(739)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gl1qw6 ;  // ../RTL/cortexm0ds_logic.v(1620)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Glaiu6 ;  // ../RTL/cortexm0ds_logic.v(445)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Glphu6 ;  // ../RTL/cortexm0ds_logic.v(164)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gmohu6 ;  // ../RTL/cortexm0ds_logic.v(151)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gn8iu6 ;  // ../RTL/cortexm0ds_logic.v(419)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gnqpw6 ;  // ../RTL/cortexm0ds_logic.v(1600)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gnuhu6 ;  // ../RTL/cortexm0ds_logic.v(232)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Go0iu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(312)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Golpw6 ;  // ../RTL/cortexm0ds_logic.v(1591)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gothu6 ;  // ../RTL/cortexm0ds_logic.v(219)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gpeow6 ;  // ../RTL/cortexm0ds_logic.v(1043)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gpqpw6 ;  // ../RTL/cortexm0ds_logic.v(1600)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gpsow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1230)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gpyiu6 ;  // ../RTL/cortexm0ds_logic.v(767)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gq4ju6_lutinv ;  // ../RTL/cortexm0ds_logic.v(848)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gqkhu6 ;  // ../RTL/cortexm0ds_logic.v(137)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gqrow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1217)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gr2qw6 ;  // ../RTL/cortexm0ds_logic.v(1622)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Grxhu6 ;  // ../RTL/cortexm0ds_logic.v(273)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gtohu6 ;  // ../RTL/cortexm0ds_logic.v(154)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Guihu6 ;  // ../RTL/cortexm0ds_logic.v(132)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gumiu6 ;  // ../RTL/cortexm0ds_logic.v(609)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Guuhu6 ;  // ../RTL/cortexm0ds_logic.v(234)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gv1bx6 ;  // ../RTL/cortexm0ds_logic.v(1683)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gw6bx6 ;  // ../RTL/cortexm0ds_logic.v(1691)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gwdpw6 ;  // ../RTL/cortexm0ds_logic.v(1514)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gweow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1046)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gwhhu6 ;  // ../RTL/cortexm0ds_logic.v(129)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gwkiu6 ;  // ../RTL/cortexm0ds_logic.v(583)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gwwpw6 ;  // ../RTL/cortexm0ds_logic.v(1611)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gwxpw6 ;  // ../RTL/cortexm0ds_logic.v(1613)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gwzhu6 ;  // ../RTL/cortexm0ds_logic.v(302)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gx2bx6 ;  // ../RTL/cortexm0ds_logic.v(1684)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gxrow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1220)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gy3ju6 ;  // ../RTL/cortexm0ds_logic.v(838)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gylpw6 ;  // ../RTL/cortexm0ds_logic.v(1591)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gyxhu6 ;  // ../RTL/cortexm0ds_logic.v(276)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gyxpw6 ;  // ../RTL/cortexm0ds_logic.v(1613)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gz6ax6 ;  // ../RTL/cortexm0ds_logic.v(1625)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gzeax6 ;  // ../RTL/cortexm0ds_logic.v(1641)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gzphu6 ;  // ../RTL/cortexm0ds_logic.v(169)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H00iu6 ;  // ../RTL/cortexm0ds_logic.v(303)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H00pw6 ;  // ../RTL/cortexm0ds_logic.v(1328)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H0ebx6 ;  // ../RTL/cortexm0ds_logic.v(1705)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H1shu6 ;  // ../RTL/cortexm0ds_logic.v(197)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H1zhu6 ;  // ../RTL/cortexm0ds_logic.v(290)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H25iu6 ;  // ../RTL/cortexm0ds_logic.v(371)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H2qiu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(652)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H2yhu6 ;  // ../RTL/cortexm0ds_logic.v(277)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H34iu6 ;  // ../RTL/cortexm0ds_logic.v(358)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H3bpw6 ;  // ../RTL/cortexm0ds_logic.v(1476)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H3lpw6 ;  // ../RTL/cortexm0ds_logic.v(1590)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H3xhu6 ;  // ../RTL/cortexm0ds_logic.v(264)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H43iu6 ;  // ../RTL/cortexm0ds_logic.v(345)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H4bax6 ;  // ../RTL/cortexm0ds_logic.v(1633)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H4phu6 ;  // ../RTL/cortexm0ds_logic.v(158)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H4ypw6 ;  // ../RTL/cortexm0ds_logic.v(1613)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H4zax6 ;  // ../RTL/cortexm0ds_logic.v(1678)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H5vhu6 ;  // ../RTL/cortexm0ds_logic.v(238)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H70iu6 ;  // ../RTL/cortexm0ds_logic.v(306)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H7hbx6 ;  // ../RTL/cortexm0ds_logic.v(1710)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H8gax6 ;  // ../RTL/cortexm0ds_logic.v(1643)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ha3ju6_lutinv ;  // ../RTL/cortexm0ds_logic.v(829)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ha4pw6 ;  // ../RTL/cortexm0ds_logic.v(1385)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Habiu6 ;  // ../RTL/cortexm0ds_logic.v(454)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Halax6 ;  // ../RTL/cortexm0ds_logic.v(1653)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hbbow6 ;  // ../RTL/cortexm0ds_logic.v(998)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hbgbx6 ;  // ../RTL/cortexm0ds_logic.v(1709)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hbphu6 ;  // ../RTL/cortexm0ds_logic.v(160)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hbpow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1185)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hcgiu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(522)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hcohu6 ;  // ../RTL/cortexm0ds_logic.v(147)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hcuiu6 ;  // ../RTL/cortexm0ds_logic.v(709)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hcvhu6 ;  // ../RTL/cortexm0ds_logic.v(241)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hd8iu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(415)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hdbax6 ;  // ../RTL/cortexm0ds_logic.v(1634)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hdfax6 ;  // ../RTL/cortexm0ds_logic.v(1642)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hduhu6 ;  // ../RTL/cortexm0ds_logic.v(228)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/He7iu6 ;  // ../RTL/cortexm0ds_logic.v(402)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Heaax6 ;  // ../RTL/cortexm0ds_logic.v(1632)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hemow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1146)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hf0bx6 ;  // ../RTL/cortexm0ds_logic.v(1680)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hfkiu6 ;  // ../RTL/cortexm0ds_logic.v(576)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hfshu6 ;  // ../RTL/cortexm0ds_logic.v(202)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hg3bx6 ;  // ../RTL/cortexm0ds_logic.v(1685)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hg7ax6 ;  // ../RTL/cortexm0ds_logic.v(1626)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hgrpw6 ;  // ../RTL/cortexm0ds_logic.v(1601)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hhqow6 ;  // ../RTL/cortexm0ds_logic.v(1200)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hhvpw6 ;  // ../RTL/cortexm0ds_logic.v(1609)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hi9bx6 ;  // ../RTL/cortexm0ds_logic.v(1696)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ;  // ../RTL/cortexm0ds_logic.v(1601)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hjgax6 ;  // ../RTL/cortexm0ds_logic.v(1644)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hjohu6 ;  // ../RTL/cortexm0ds_logic.v(150)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hkgow6 ;  // ../RTL/cortexm0ds_logic.v(1068)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hlcax6 ;  // ../RTL/cortexm0ds_logic.v(1636)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hlliu6 ;  // ../RTL/cortexm0ds_logic.v(592)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hlwpw6 ;  // ../RTL/cortexm0ds_logic.v(1611)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hlziu6 ;  // ../RTL/cortexm0ds_logic.v(779)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hm7ow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(948)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hmbax6 ;  // ../RTL/cortexm0ds_logic.v(1634)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hndow6 ;  // ../RTL/cortexm0ds_logic.v(1029)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hoiiu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(553)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hpbbx6 ;  // ../RTL/cortexm0ds_logic.v(1700)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hpcbx6 ;  // ../RTL/cortexm0ds_logic.v(1702)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hphiu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(540)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hqabx6 ;  // ../RTL/cortexm0ds_logic.v(1698)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hqgiu6 ;  // ../RTL/cortexm0ds_logic.v(527)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hrfbx6 ;  // ../RTL/cortexm0ds_logic.v(1708)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hruhu6 ;  // ../RTL/cortexm0ds_logic.v(233)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hs8ow6 ;  // ../RTL/cortexm0ds_logic.v(964)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hsdax6 ;  // ../RTL/cortexm0ds_logic.v(1639)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hsliu6 ;  // ../RTL/cortexm0ds_logic.v(595)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Htbax6 ;  // ../RTL/cortexm0ds_logic.v(1635)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Htmpw6 ;  // ../RTL/cortexm0ds_logic.v(1593)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Htshu6 ;  // ../RTL/cortexm0ds_logic.v(207)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Htyiu6 ;  // ../RTL/cortexm0ds_logic.v(769)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hvcow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1018)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hviiu6 ;  // ../RTL/cortexm0ds_logic.v(556)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hvqhu6 ;  // ../RTL/cortexm0ds_logic.v(181)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hw8ax6 ;  // ../RTL/cortexm0ds_logic.v(1629)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hwaiu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(449)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hwhiu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(543)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hwhpw6 ;  // ../RTL/cortexm0ds_logic.v(1584)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hxohu6 ;  // ../RTL/cortexm0ds_logic.v(155)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hy1pw6 ;  // ../RTL/cortexm0ds_logic.v(1354)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hymiu6 ;  // ../RTL/cortexm0ds_logic.v(610)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hyuhu6 ;  // ../RTL/cortexm0ds_logic.v(236)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hz0iu6 ;  // ../RTL/cortexm0ds_logic.v(316)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hz0pw6 ;  // ../RTL/cortexm0ds_logic.v(1341)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hz9ax6 ;  // ../RTL/cortexm0ds_logic.v(1631)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hzliu6 ;  // ../RTL/cortexm0ds_logic.v(597)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I0dax6 ;  // ../RTL/cortexm0ds_logic.v(1637)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I0opw6 ;  // ../RTL/cortexm0ds_logic.v(1595)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I0wiu6 ;  // ../RTL/cortexm0ds_logic.v(731)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I13iu6 ;  // ../RTL/cortexm0ds_logic.v(344)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I1lpw6 ;  // ../RTL/cortexm0ds_logic.v(1589)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I1phu6 ;  // ../RTL/cortexm0ds_logic.v(157)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I28ju6 ;  // ../RTL/cortexm0ds_logic.v(893)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I2vhu6 ;  // ../RTL/cortexm0ds_logic.v(237)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I2zax6 ;  // ../RTL/cortexm0ds_logic.v(1678)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I30ju6_lutinv ;  // ../RTL/cortexm0ds_logic.v(786)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I3fiu6 ;  // ../RTL/cortexm0ds_logic.v(505)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I3lhu6 ;  // ../RTL/cortexm0ds_logic.v(138)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I40iu6 ;  // ../RTL/cortexm0ds_logic.v(305)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I45bx6 ;  // ../RTL/cortexm0ds_logic.v(1688)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I46ju6 ;  // ../RTL/cortexm0ds_logic.v(867)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I4eiu6 ;  // ../RTL/cortexm0ds_logic.v(492)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I4epw6 ;  // ../RTL/cortexm0ds_logic.v(1517)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I4rpw6 ;  // ../RTL/cortexm0ds_logic.v(1601)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I55ju6 ;  // ../RTL/cortexm0ds_logic.v(854)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I5nhu6 ;  // ../RTL/cortexm0ds_logic.v(144)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I5xax6 ;  // ../RTL/cortexm0ds_logic.v(1674)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I6row6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1210)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I6yhu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(279)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I74bx6 ;  // ../RTL/cortexm0ds_logic.v(1687)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I74iu6 ;  // ../RTL/cortexm0ds_logic.v(360)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I7cow6 ;  // ../RTL/cortexm0ds_logic.v(1010)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I7xhu6 ;  // ../RTL/cortexm0ds_logic.v(266)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I82ju6 ;  // ../RTL/cortexm0ds_logic.v(815)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I8lax6 ;  // ../RTL/cortexm0ds_logic.v(1653)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I8phu6 ;  // ../RTL/cortexm0ds_logic.v(159)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I98ju6_lutinv ;  // ../RTL/cortexm0ds_logic.v(895)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I9ihu6 ;  // ../RTL/cortexm0ds_logic.v(130)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ia0ju6 ;  // ../RTL/cortexm0ds_logic.v(789)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ia8iu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(414)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iauhu6 ;  // ../RTL/cortexm0ds_logic.v(227)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ib0iu6 ;  // ../RTL/cortexm0ds_logic.v(308)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ibliu6 ;  // ../RTL/cortexm0ds_logic.v(588)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ibqpw6 ;  // ../RTL/cortexm0ds_logic.v(1599)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ibsiu6 ;  // ../RTL/cortexm0ds_logic.v(682)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ickiu6 ;  // ../RTL/cortexm0ds_logic.v(575)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Id4ju6 ;  // ../RTL/cortexm0ds_logic.v(843)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iddax6 ;  // ../RTL/cortexm0ds_logic.v(1638)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idkow6 ;  // ../RTL/cortexm0ds_logic.v(1119)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idqpw6 ;  // ../RTL/cortexm0ds_logic.v(1599)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iecow6 ;  // ../RTL/cortexm0ds_logic.v(1012)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iekax6 ;  // ../RTL/cortexm0ds_logic.v(1651)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iexow6 ;  // ../RTL/cortexm0ds_logic.v(1293)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/If3pw6 ;  // ../RTL/cortexm0ds_logic.v(1374)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ifoiu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(630)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ifphu6 ;  // ../RTL/cortexm0ds_logic.v(162)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ig2bx6 ;  // ../RTL/cortexm0ds_logic.v(1684)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Igohu6 ;  // ../RTL/cortexm0ds_logic.v(149)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ih0bx6 ;  // ../RTL/cortexm0ds_logic.v(1680)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iiliu6 ;  // ../RTL/cortexm0ds_logic.v(591)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iimow6 ;  // ../RTL/cortexm0ds_logic.v(1147)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iithu6 ;  // ../RTL/cortexm0ds_logic.v(217)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iixpw6 ;  // ../RTL/cortexm0ds_logic.v(1612)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ikhbx6 ;  // ../RTL/cortexm0ds_logic.v(1711)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ilwiu6 ;  // ../RTL/cortexm0ds_logic.v(739)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Im2ju6 ;  // ../RTL/cortexm0ds_logic.v(820)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Im9ax6 ;  // ../RTL/cortexm0ds_logic.v(1630)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Imhbx6 ;  // ../RTL/cortexm0ds_logic.v(1711)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Inniu6 ;  // ../RTL/cortexm0ds_logic.v(620)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Inohu6 ;  // ../RTL/cortexm0ds_logic.v(152)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Io9ow6 ;  // ../RTL/cortexm0ds_logic.v(976)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ipliu6 ;  // ../RTL/cortexm0ds_logic.v(594)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ipthu6 ;  // ../RTL/cortexm0ds_logic.v(219)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iqihu6 ;  // ../RTL/cortexm0ds_logic.v(132)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iqriu6 ;  // ../RTL/cortexm0ds_logic.v(674)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iqsow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1231)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iqzhu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(300)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ir6ow6 ;  // ../RTL/cortexm0ds_logic.v(937)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Irmpw6 ;  // ../RTL/cortexm0ds_logic.v(1593)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Irrhu6 ;  // ../RTL/cortexm0ds_logic.v(193)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Irrow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1218)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Isbpw6 ;  // ../RTL/cortexm0ds_logic.v(1485)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Isjpw6 ;  // ../RTL/cortexm0ds_logic.v(1587)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/It3iu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(354)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Itbow6 ;  // ../RTL/cortexm0ds_logic.v(1004)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Itcbx6 ;  // ../RTL/cortexm0ds_logic.v(1702)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iugiu6 ;  // ../RTL/cortexm0ds_logic.v(529)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iuohu6 ;  // ../RTL/cortexm0ds_logic.v(154)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iv1iu6 ;  // ../RTL/cortexm0ds_logic.v(328)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ivfiu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(516)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ivmiu6 ;  // ../RTL/cortexm0ds_logic.v(609)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iwtow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1246)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ixzhu6 ;  // ../RTL/cortexm0ds_logic.v(302)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Izxhu6 ;  // ../RTL/cortexm0ds_logic.v(276)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J0fiu6 ;  // ../RTL/cortexm0ds_logic.v(504)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J0gax6 ;  // ../RTL/cortexm0ds_logic.v(1643)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J0iax6 ;  // ../RTL/cortexm0ds_logic.v(1647)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J10iu6 ;  // ../RTL/cortexm0ds_logic.v(304)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J17iu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(397)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J1epw6 ;  // ../RTL/cortexm0ds_logic.v(1515)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J2sow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1222)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J39bx6 ;  // ../RTL/cortexm0ds_logic.v(1695)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J3row6 ;  // ../RTL/cortexm0ds_logic.v(1209)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J3xiu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(746)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J3yhu6 ;  // ../RTL/cortexm0ds_logic.v(278)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J43ju6_lutinv ;  // ../RTL/cortexm0ds_logic.v(826)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J44iu6 ;  // ../RTL/cortexm0ds_logic.v(358)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J4cbx6 ;  // ../RTL/cortexm0ds_logic.v(1701)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J4xhu6 ;  // ../RTL/cortexm0ds_logic.v(265)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J59ax6 ;  // ../RTL/cortexm0ds_logic.v(1630)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J5eax6 ;  // ../RTL/cortexm0ds_logic.v(1639)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J5jbx6 ;  // ../RTL/cortexm0ds_logic.v(1714)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J5phu6 ;  // ../RTL/cortexm0ds_logic.v(158)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J5pow6 ;  // ../RTL/cortexm0ds_logic.v(1183)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J6ebx6 ;  // ../RTL/cortexm0ds_logic.v(1705)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J6vhu6 ;  // ../RTL/cortexm0ds_logic.v(239)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J6zax6 ;  // ../RTL/cortexm0ds_logic.v(1678)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J71iu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(319)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J77ju6 ;  // ../RTL/cortexm0ds_logic.v(881)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J7xax6 ;  // ../RTL/cortexm0ds_logic.v(1674)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J80iu6 ;  // ../RTL/cortexm0ds_logic.v(306)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J8cax6 ;  // ../RTL/cortexm0ds_logic.v(1636)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J8eiu6 ;  // ../RTL/cortexm0ds_logic.v(494)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J8fow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1050)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J8ziu6 ;  // ../RTL/cortexm0ds_logic.v(774)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J9eow6 ;  // ../RTL/cortexm0ds_logic.v(1037)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J9kiu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(574)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J9zhu6 ;  // ../RTL/cortexm0ds_logic.v(293)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ja5iu6 ;  // ../RTL/cortexm0ds_logic.v(374)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jajiu6 ;  // ../RTL/cortexm0ds_logic.v(561)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jaqiu6 ;  // ../RTL/cortexm0ds_logic.v(655)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jb3ju6_lutinv ;  // ../RTL/cortexm0ds_logic.v(829)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jbjow6 ;  // ../RTL/cortexm0ds_logic.v(1105)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jc3pw6 ;  // ../RTL/cortexm0ds_logic.v(1372)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jckax6 ;  // ../RTL/cortexm0ds_logic.v(1651)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jcphu6 ;  // ../RTL/cortexm0ds_logic.v(161)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jcpow6 ;  // ../RTL/cortexm0ds_logic.v(1185)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jdgbx6 ;  // ../RTL/cortexm0ds_logic.v(1709)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jdohu6 ;  // ../RTL/cortexm0ds_logic.v(148)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jeuhu6 ;  // ../RTL/cortexm0ds_logic.v(228)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jf6ju6 ;  // ../RTL/cortexm0ds_logic.v(871)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jf7iu6 ;  // ../RTL/cortexm0ds_logic.v(403)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jfdbx6 ;  // ../RTL/cortexm0ds_logic.v(1703)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jflpw6 ;  // ../RTL/cortexm0ds_logic.v(1590)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jfmow6 ;  // ../RTL/cortexm0ds_logic.v(1146)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jfthu6 ;  // ../RTL/cortexm0ds_logic.v(215)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jgeow6 ;  // ../RTL/cortexm0ds_logic.v(1040)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jgkiu6 ;  // ../RTL/cortexm0ds_logic.v(577)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jgxpw6 ;  // ../RTL/cortexm0ds_logic.v(1612)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jhebx6 ;  // ../RTL/cortexm0ds_logic.v(1705)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jhyow6 ;  // ../RTL/cortexm0ds_logic.v(1307)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jieax6 ;  // ../RTL/cortexm0ds_logic.v(1640)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jj0bx6 ;  // ../RTL/cortexm0ds_logic.v(1680)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jjoiu6 ;  // ../RTL/cortexm0ds_logic.v(631)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jjwow6 ;  // ../RTL/cortexm0ds_logic.v(1281)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jkhow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1081)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jkniu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(618)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jkohu6 ;  // ../RTL/cortexm0ds_logic.v(150)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jl3qw6 ;  // ../RTL/cortexm0ds_logic.v(1624)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jl8iu6 ;  // ../RTL/cortexm0ds_logic.v(418)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jlmiu6 ;  // ../RTL/cortexm0ds_logic.v(605)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jn7ow6 ;  // ../RTL/cortexm0ds_logic.v(949)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jo4ju6_lutinv ;  // ../RTL/cortexm0ds_logic.v(847)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Johbx6 ;  // ../RTL/cortexm0ds_logic.v(1711)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jp9bx6 ;  // ../RTL/cortexm0ds_logic.v(1697)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jpmpw6 ;  // ../RTL/cortexm0ds_logic.v(1593)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jq3iu6 ;  // ../RTL/cortexm0ds_logic.v(353)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jr1ju6_lutinv ;  // ../RTL/cortexm0ds_logic.v(808)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jraax6 ;  // ../RTL/cortexm0ds_logic.v(1633)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jrhow6 ;  // ../RTL/cortexm0ds_logic.v(1084)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jrohu6 ;  // ../RTL/cortexm0ds_logic.v(153)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jrvow6 ;  // ../RTL/cortexm0ds_logic.v(1271)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jrypw6 ;  // ../RTL/cortexm0ds_logic.v(1615)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jsmiu6 ;  // ../RTL/cortexm0ds_logic.v(608)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jsuhu6 ;  // ../RTL/cortexm0ds_logic.v(234)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jvdow6 ;  // ../RTL/cortexm0ds_logic.v(1032)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jvkpw6 ;  // ../RTL/cortexm0ds_logic.v(1589)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jvvpw6 ;  // ../RTL/cortexm0ds_logic.v(1609)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jwxhu6 ;  // ../RTL/cortexm0ds_logic.v(275)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jwxow6 ;  // ../RTL/cortexm0ds_logic.v(1300)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jx1bx6 ;  // ../RTL/cortexm0ds_logic.v(1683)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jxaiu6 ;  // ../RTL/cortexm0ds_logic.v(449)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jxgax6 ;  // ../RTL/cortexm0ds_logic.v(1645)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jy2pw6 ;  // ../RTL/cortexm0ds_logic.v(1367)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jy9iu6 ;  // ../RTL/cortexm0ds_logic.v(436)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jyohu6 ;  // ../RTL/cortexm0ds_logic.v(156)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jz2bx6 ;  // ../RTL/cortexm0ds_logic.v(1684)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jz8iu6 ;  // ../RTL/cortexm0ds_logic.v(423)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jzfiu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(517)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jzmiu6 ;  // ../RTL/cortexm0ds_logic.v(611)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jzuhu6 ;  // ../RTL/cortexm0ds_logic.v(236)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K0qiu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(651)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K0xiu6 ;  // ../RTL/cortexm0ds_logic.v(745)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K0yhu6 ;  // ../RTL/cortexm0ds_logic.v(277)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K1cow6 ;  // ../RTL/cortexm0ds_logic.v(1007)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K2phu6 ;  // ../RTL/cortexm0ds_logic.v(157)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K39iu6 ;  // ../RTL/cortexm0ds_logic.v(425)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K3niu6 ;  // ../RTL/cortexm0ds_logic.v(612)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K3vhu6 ;  // ../RTL/cortexm0ds_logic.v(238)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K49ow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(968)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K50iu6 ;  // ../RTL/cortexm0ds_logic.v(305)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K5eiu6 ;  // ../RTL/cortexm0ds_logic.v(493)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K5hbx6 ;  // ../RTL/cortexm0ds_logic.v(1710)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K5ihu6 ;  // ../RTL/cortexm0ds_logic.v(130)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K65bx6 ;  // ../RTL/cortexm0ds_logic.v(1688)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K66iu6 ;  // ../RTL/cortexm0ds_logic.v(386)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K6gax6 ;  // ../RTL/cortexm0ds_logic.v(1643)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K75iu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(373)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K7row6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1210)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K84iu6 ;  // ../RTL/cortexm0ds_logic.v(360)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K8iiu6 ;  // ../RTL/cortexm0ds_logic.v(547)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K8qhu6 ;  // ../RTL/cortexm0ds_logic.v(173)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K8xhu6 ;  // ../RTL/cortexm0ds_logic.v(266)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K94bx6 ;  // ../RTL/cortexm0ds_logic.v(1687)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K9phu6 ;  // ../RTL/cortexm0ds_logic.v(160)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ka8ju6 ;  // ../RTL/cortexm0ds_logic.v(896)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kadbx6 ;  // ../RTL/cortexm0ds_logic.v(1703)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kakax6 ;  // ../RTL/cortexm0ds_logic.v(1651)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kalpw6 ;  // ../RTL/cortexm0ds_logic.v(1590)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kavhu6 ;  // ../RTL/cortexm0ds_logic.v(240)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kb9ow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(971)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kbuhu6 ;  // ../RTL/cortexm0ds_logic.v(227)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kc6ju6 ;  // ../RTL/cortexm0ds_logic.v(870)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kcaax6 ;  // ../RTL/cortexm0ds_logic.v(1632)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kctow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1239)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kdkiu6 ;  // ../RTL/cortexm0ds_logic.v(576)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ke1qw6 ;  // ../RTL/cortexm0ds_logic.v(1619)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kfcow6 ;  // ../RTL/cortexm0ds_logic.v(1013)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kgoiu6 ;  // ../RTL/cortexm0ds_logic.v(630)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Khgax6 ;  // ../RTL/cortexm0ds_logic.v(1644)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Khniu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(617)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Khohu6 ;  // ../RTL/cortexm0ds_logic.v(149)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Khvhu6 ;  // ../RTL/cortexm0ds_logic.v(243)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kikhu6 ;  // ../RTL/cortexm0ds_logic.v(137)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kjthu6 ;  // ../RTL/cortexm0ds_logic.v(217)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kjziu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(779)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kkkiu6 ;  // ../RTL/cortexm0ds_logic.v(578)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kkriu6 ;  // ../RTL/cortexm0ds_logic.v(672)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kl0bx6 ;  // ../RTL/cortexm0ds_logic.v(1680)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kl4ju6_lutinv ;  // ../RTL/cortexm0ds_logic.v(846)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kl8ax6 ;  // ../RTL/cortexm0ds_logic.v(1628)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kldow6 ;  // ../RTL/cortexm0ds_logic.v(1028)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kmihu6 ;  // ../RTL/cortexm0ds_logic.v(131)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kmiiu6 ;  // ../RTL/cortexm0ds_logic.v(552)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kmqow6 ;  // ../RTL/cortexm0ds_logic.v(1202)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kn1qw6 ;  // ../RTL/cortexm0ds_logic.v(1620)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kn2qw6 ;  // ../RTL/cortexm0ds_logic.v(1622)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Knbbx6 ;  // ../RTL/cortexm0ds_logic.v(1700)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Koabx6 ;  // ../RTL/cortexm0ds_logic.v(1698)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kojpw6 ;  // ../RTL/cortexm0ds_logic.v(1587)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Koohu6 ;  // ../RTL/cortexm0ds_logic.v(152)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kp1pw6 ;  // ../RTL/cortexm0ds_logic.v(1351)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kpfbx6 ;  // ../RTL/cortexm0ds_logic.v(1708)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kpuhu6 ;  // ../RTL/cortexm0ds_logic.v(233)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kq0pw6 ;  // ../RTL/cortexm0ds_logic.v(1338)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kq7iu6 ;  // ../RTL/cortexm0ds_logic.v(407)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kqdax6 ;  // ../RTL/cortexm0ds_logic.v(1638)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kqhbx6 ;  // ../RTL/cortexm0ds_logic.v(1711)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kqthu6 ;  // ../RTL/cortexm0ds_logic.v(220)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Krbax6 ;  // ../RTL/cortexm0ds_logic.v(1635)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Krkiu6 ;  // ../RTL/cortexm0ds_logic.v(581)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Krlpw6 ;  // ../RTL/cortexm0ds_logic.v(1591)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ksgax6 ;  // ../RTL/cortexm0ds_logic.v(1644)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kswpw6 ;  // ../RTL/cortexm0ds_logic.v(1611)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kt4iu6 ;  // ../RTL/cortexm0ds_logic.v(368)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ktwiu6 ;  // ../RTL/cortexm0ds_logic.v(742)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kubow6 ;  // ../RTL/cortexm0ds_logic.v(1005)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kuphu6 ;  // ../RTL/cortexm0ds_logic.v(168)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kupow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1192)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kv9iu6 ;  // ../RTL/cortexm0ds_logic.v(435)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kw1iu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(329)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kwfiu6 ;  // ../RTL/cortexm0ds_logic.v(516)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kwlpw6 ;  // ../RTL/cortexm0ds_logic.v(1591)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kwuhu6 ;  // ../RTL/cortexm0ds_logic.v(235)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kwuow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1260)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kxeax6 ;  // ../RTL/cortexm0ds_logic.v(1641)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kxhpw6 ;  // ../RTL/cortexm0ds_logic.v(1584)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kxziu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(784)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kyzhu6 ;  // ../RTL/cortexm0ds_logic.v(303)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kzabx6 ;  // ../RTL/cortexm0ds_logic.v(1699)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kzkhu6 ;  // ../RTL/cortexm0ds_logic.v(138)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L03qw6 ;  // ../RTL/cortexm0ds_logic.v(1623)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L0how6 ;  // ../RTL/cortexm0ds_logic.v(1074)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L0niu6 ;  // ../RTL/cortexm0ds_logic.v(611)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L0vhu6 ;  // ../RTL/cortexm0ds_logic.v(237)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L0vow6 ;  // ../RTL/cortexm0ds_logic.v(1261)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L0ypw6 ;  // ../RTL/cortexm0ds_logic.v(1613)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L18iu6 ;  // ../RTL/cortexm0ds_logic.v(411)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L1bbx6 ;  // ../RTL/cortexm0ds_logic.v(1699)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L1fiu6 ;  // ../RTL/cortexm0ds_logic.v(504)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L20iu6 ;  // ../RTL/cortexm0ds_logic.v(304)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L27pw6 ;  // ../RTL/cortexm0ds_logic.v(1422)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L2bax6 ;  // ../RTL/cortexm0ds_logic.v(1633)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L2epw6 ;  // ../RTL/cortexm0ds_logic.v(1516)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L3sow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1222)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L45iu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(372)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L4lax6 ;  // ../RTL/cortexm0ds_logic.v(1652)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L4rhu6 ;  // ../RTL/cortexm0ds_logic.v(185)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L54iu6 ;  // ../RTL/cortexm0ds_logic.v(359)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L5lpw6 ;  // ../RTL/cortexm0ds_logic.v(1590)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6lax6 ;  // ../RTL/cortexm0ds_logic.v(1653)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6phu6 ;  // ../RTL/cortexm0ds_logic.v(159)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L8kax6 ;  // ../RTL/cortexm0ds_logic.v(1651)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L8uow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1251)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L8zax6 ;  // ../RTL/cortexm0ds_logic.v(1678)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L90iu6 ;  // ../RTL/cortexm0ds_logic.v(307)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L9bbx6 ;  // ../RTL/cortexm0ds_logic.v(1699)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L9eiu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(494)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L9mow6 ;  // ../RTL/cortexm0ds_logic.v(1144)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L9xax6 ;  // ../RTL/cortexm0ds_logic.v(1674)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lariu6 ;  // ../RTL/cortexm0ds_logic.v(668)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lashu6 ;  // ../RTL/cortexm0ds_logic.v(200)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lbbax6 ;  // ../RTL/cortexm0ds_logic.v(1634)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lbyhu6 ;  // ../RTL/cortexm0ds_logic.v(281)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lclhu6 ;  // ../RTL/cortexm0ds_logic.v(139)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lcqow6 ;  // ../RTL/cortexm0ds_logic.v(1199)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ldiow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1092)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ldoiu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(629)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ldphu6 ;  // ../RTL/cortexm0ds_logic.v(161)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ldvpw6 ;  // ../RTL/cortexm0ds_logic.v(1608)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Le2qw6 ;  // ../RTL/cortexm0ds_logic.v(1621)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Leohu6 ;  // ../RTL/cortexm0ds_logic.v(148)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lf1iu6 ;  // ../RTL/cortexm0ds_logic.v(322)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lf8iu6 ;  // ../RTL/cortexm0ds_logic.v(416)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lfgbx6 ;  // ../RTL/cortexm0ds_logic.v(1709)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lfgow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1066)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lg1bx6 ;  // ../RTL/cortexm0ds_logic.v(1682)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lg7iu6 ;  // ../RTL/cortexm0ds_logic.v(403)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lg9bx6 ;  // ../RTL/cortexm0ds_logic.v(1696)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lgkax6 ;  // ../RTL/cortexm0ds_logic.v(1651)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lgthu6 ;  // ../RTL/cortexm0ds_logic.v(216)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lhbbx6 ;  // ../RTL/cortexm0ds_logic.v(1700)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lhdiu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(484)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Li2bx6 ;  // ../RTL/cortexm0ds_logic.v(1684)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Li5iu6 ;  // ../RTL/cortexm0ds_logic.v(377)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Li7ax6 ;  // ../RTL/cortexm0ds_logic.v(1626)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Liabx6 ;  // ../RTL/cortexm0ds_logic.v(1698)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lj3ju6_lutinv ;  // ../RTL/cortexm0ds_logic.v(832)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljbpw6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1482)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljcax6 ;  // ../RTL/cortexm0ds_logic.v(1636)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljiiu6 ;  // ../RTL/cortexm0ds_logic.v(551)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljqow6 ;  // ../RTL/cortexm0ds_logic.v(1201)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lk9ax6 ;  // ../RTL/cortexm0ds_logic.v(1630)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ll2pw6 ;  // ../RTL/cortexm0ds_logic.v(1362)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Llaow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(988)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Llohu6 ;  // ../RTL/cortexm0ds_logic.v(151)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lm1iu6 ;  // ../RTL/cortexm0ds_logic.v(325)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lmkbx6 ;  // ../RTL/cortexm0ds_logic.v(1717)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lmuhu6 ;  // ../RTL/cortexm0ds_logic.v(231)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ln0bx6 ;  // ../RTL/cortexm0ds_logic.v(1680)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ln0pw6 ;  // ../RTL/cortexm0ds_logic.v(1336)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lokiu6 ;  // ../RTL/cortexm0ds_logic.v(580)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lolow6 ;  // ../RTL/cortexm0ds_logic.v(1136)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Loshu6 ;  // ../RTL/cortexm0ds_logic.v(205)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lp4ju6 ;  // ../RTL/cortexm0ds_logic.v(848)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lqcow6 ;  // ../RTL/cortexm0ds_logic.v(1017)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lr9bx6 ;  // ../RTL/cortexm0ds_logic.v(1697)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lrhiu6 ;  // ../RTL/cortexm0ds_logic.v(541)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ls1ju6 ;  // ../RTL/cortexm0ds_logic.v(809)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ls9pw6 ;  // ../RTL/cortexm0ds_logic.v(1459)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ltmiu6 ;  // ../RTL/cortexm0ds_logic.v(608)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ltuhu6 ;  // ../RTL/cortexm0ds_logic.v(234)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lu0iu6 ;  // ../RTL/cortexm0ds_logic.v(315)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lv7ow6 ;  // ../RTL/cortexm0ds_logic.v(952)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lvzhu6 ;  // ../RTL/cortexm0ds_logic.v(302)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lx9ax6 ;  // ../RTL/cortexm0ds_logic.v(1631)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lxxhu6 ;  // ../RTL/cortexm0ds_logic.v(276)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ly2ju6 ;  // ../RTL/cortexm0ds_logic.v(824)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lycax6 ;  // ../RTL/cortexm0ds_logic.v(1637)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lywpw6 ;  // ../RTL/cortexm0ds_logic.v(1611)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lzohu6 ;  // ../RTL/cortexm0ds_logic.v(156)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M0eow6 ;  // ../RTL/cortexm0ds_logic.v(1034)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M13bx6 ;  // ../RTL/cortexm0ds_logic.v(1685)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M14ju6 ;  // ../RTL/cortexm0ds_logic.v(839)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M15iu6 ;  // ../RTL/cortexm0ds_logic.v(371)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M1ihu6 ;  // ../RTL/cortexm0ds_logic.v(130)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M1jiu6 ;  // ../RTL/cortexm0ds_logic.v(558)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M1xiu6 ;  // ../RTL/cortexm0ds_logic.v(745)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M1yhu6 ;  // ../RTL/cortexm0ds_logic.v(277)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M24iu6 ;  // ../RTL/cortexm0ds_logic.v(358)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M2cow6 ;  // ../RTL/cortexm0ds_logic.v(1008)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M2ebx6 ;  // ../RTL/cortexm0ds_logic.v(1705)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M2xhu6 ;  // ../RTL/cortexm0ds_logic.v(264)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M3phu6 ;  // ../RTL/cortexm0ds_logic.v(158)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M4ebx6 ;  // ../RTL/cortexm0ds_logic.v(1705)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M4vhu6 ;  // ../RTL/cortexm0ds_logic.v(238)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M60iu6 ;  // ../RTL/cortexm0ds_logic.v(306)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6cax6 ;  // ../RTL/cortexm0ds_logic.v(1635)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6eiu6 ;  // ../RTL/cortexm0ds_logic.v(493)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6kax6 ;  // ../RTL/cortexm0ds_logic.v(1651)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6rpw6 ;  // ../RTL/cortexm0ds_logic.v(1601)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M7kiu6 ;  // ../RTL/cortexm0ds_logic.v(574)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M7zhu6 ;  // ../RTL/cortexm0ds_logic.v(293)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M81qw6 ;  // ../RTL/cortexm0ds_logic.v(1619)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M85bx6 ;  // ../RTL/cortexm0ds_logic.v(1688)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M8fax6 ;  // ../RTL/cortexm0ds_logic.v(1641)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M8ipw6 ;  // ../RTL/cortexm0ds_logic.v(1584)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M8row6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1211)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M93ju6_lutinv ;  // ../RTL/cortexm0ds_logic.v(828)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M94iu6 ;  // ../RTL/cortexm0ds_logic.v(360)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Maphu6 ;  // ../RTL/cortexm0ds_logic.v(160)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mb1ju6 ;  // ../RTL/cortexm0ds_logic.v(802)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mb4bx6 ;  // ../RTL/cortexm0ds_logic.v(1687)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mbdax6 ;  // ../RTL/cortexm0ds_logic.v(1638)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mbhow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1078)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mbohu6 ;  // ../RTL/cortexm0ds_logic.v(147)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mbvhu6 ;  // ../RTL/cortexm0ds_logic.v(241)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mcuhu6 ;  // ../RTL/cortexm0ds_logic.v(228)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Md7iu6 ;  // ../RTL/cortexm0ds_logic.v(402)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mdfow6 ;  // ../RTL/cortexm0ds_logic.v(1052)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mekiu6 ;  // ../RTL/cortexm0ds_logic.v(576)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mfjiu6 ;  // ../RTL/cortexm0ds_logic.v(563)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mfyax6 ;  // ../RTL/cortexm0ds_logic.v(1677)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mg3ju6_lutinv ;  // ../RTL/cortexm0ds_logic.v(831)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mgeax6 ;  // ../RTL/cortexm0ds_logic.v(1640)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mh1qw6 ;  // ../RTL/cortexm0ds_logic.v(1620)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mi8ju6_lutinv ;  // ../RTL/cortexm0ds_logic.v(899)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mihow6 ;  // ../RTL/cortexm0ds_logic.v(1081)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Miihu6 ;  // ../RTL/cortexm0ds_logic.v(131)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Miniu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(618)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Miohu6 ;  // ../RTL/cortexm0ds_logic.v(150)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mivhu6 ;  // ../RTL/cortexm0ds_logic.v(243)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mj8iu6 ;  // ../RTL/cortexm0ds_logic.v(418)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mjgow6 ;  // ../RTL/cortexm0ds_logic.v(1068)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mjmiu6 ;  // ../RTL/cortexm0ds_logic.v(605)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mjnow6 ;  // ../RTL/cortexm0ds_logic.v(1161)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mjtiu6 ;  // ../RTL/cortexm0ds_logic.v(698)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mk3bx6 ;  // ../RTL/cortexm0ds_logic.v(1685)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mk6ju6_lutinv ;  // ../RTL/cortexm0ds_logic.v(873)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ml6pw6 ;  // ../RTL/cortexm0ds_logic.v(1416)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mldpw6 ;  // ../RTL/cortexm0ds_logic.v(1510)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mmjiu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(566)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mmqiu6 ;  // ../RTL/cortexm0ds_logic.v(659)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mmyhu6 ;  // ../RTL/cortexm0ds_logic.v(285)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mnmpw6 ;  // ../RTL/cortexm0ds_logic.v(1593)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mnqow6 ;  // ../RTL/cortexm0ds_logic.v(1203)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mp0bx6 ;  // ../RTL/cortexm0ds_logic.v(1681)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mpgiu6 ;  // ../RTL/cortexm0ds_logic.v(527)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mpniu6 ;  // ../RTL/cortexm0ds_logic.v(620)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mpohu6 ;  // ../RTL/cortexm0ds_logic.v(152)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mq1iu6 ;  // ../RTL/cortexm0ds_logic.v(327)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mrfow6 ;  // ../RTL/cortexm0ds_logic.v(1057)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mrthu6 ;  // ../RTL/cortexm0ds_logic.v(220)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ms5bx6 ;  // ../RTL/cortexm0ds_logic.v(1689)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mt4ju6 ;  // ../RTL/cortexm0ds_logic.v(849)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mt6ow6 ;  // ../RTL/cortexm0ds_logic.v(938)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mtrow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1218)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mu3ju6 ;  // ../RTL/cortexm0ds_logic.v(836)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Muhbx6 ;  // ../RTL/cortexm0ds_logic.v(1712)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mx8iu6 ;  // ../RTL/cortexm0ds_logic.v(423)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mxfiu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(516)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mxuhu6 ;  // ../RTL/cortexm0ds_logic.v(236)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/My0iu6 ;  // ../RTL/cortexm0ds_logic.v(316)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mz1bx6 ;  // ../RTL/cortexm0ds_logic.v(1683)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mz6iu6 ;  // ../RTL/cortexm0ds_logic.v(397)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mzihu6 ;  // ../RTL/cortexm0ds_logic.v(132)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mzkiu6 ;  // ../RTL/cortexm0ds_logic.v(584)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mzzhu6 ;  // ../RTL/cortexm0ds_logic.v(303)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N0cbx6 ;  // ../RTL/cortexm0ds_logic.v(1701)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N0phu6 ;  // ../RTL/cortexm0ds_logic.v(156)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N0xpw6 ;  // ../RTL/cortexm0ds_logic.v(1611)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N18ju6_lutinv ;  // ../RTL/cortexm0ds_logic.v(892)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N19bx6 ;  // ../RTL/cortexm0ds_logic.v(1695)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N1vhu6 ;  // ../RTL/cortexm0ds_logic.v(237)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N2fiu6 ;  // ../RTL/cortexm0ds_logic.v(505)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N30iu6 ;  // ../RTL/cortexm0ds_logic.v(305)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N39ax6 ;  // ../RTL/cortexm0ds_logic.v(1629)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N3eax6 ;  // ../RTL/cortexm0ds_logic.v(1639)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N3epw6 ;  // ../RTL/cortexm0ds_logic.v(1516)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N3hbx6 ;  // ../RTL/cortexm0ds_logic.v(1710)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N3jbx6 ;  // ../RTL/cortexm0ds_logic.v(1714)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N3ziu6 ;  // ../RTL/cortexm0ds_logic.v(773)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N45ju6 ;  // ../RTL/cortexm0ds_logic.v(853)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N4gax6 ;  // ../RTL/cortexm0ds_logic.v(1643)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N4kax6 ;  // ../RTL/cortexm0ds_logic.v(1651)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5bbx6 ;  // ../RTL/cortexm0ds_logic.v(1699)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N61qw6 ;  // ../RTL/cortexm0ds_logic.v(1619)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N64iu6 ;  // ../RTL/cortexm0ds_logic.v(359)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N6xhu6 ;  // ../RTL/cortexm0ds_logic.v(266)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N7phu6 ;  // ../RTL/cortexm0ds_logic.v(159)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N7pow6 ;  // ../RTL/cortexm0ds_logic.v(1183)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N8rpw6 ;  // ../RTL/cortexm0ds_logic.v(1601)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N98iu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(414)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N9now6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1157)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N9uhu6 ;  // ../RTL/cortexm0ds_logic.v(227)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Na0iu6 ;  // ../RTL/cortexm0ds_logic.v(307)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Naaax6 ;  // ../RTL/cortexm0ds_logic.v(1632)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nazax6 ;  // ../RTL/cortexm0ds_logic.v(1678)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nbdiu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(481)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nbkiu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(575)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nbxax6 ;  // ../RTL/cortexm0ds_logic.v(1675)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ncjiu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(562)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nckbx6 ;  // ../RTL/cortexm0ds_logic.v(1716)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nd3ju6 ;  // ../RTL/cortexm0ds_logic.v(830)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nd3qw6 ;  // ../RTL/cortexm0ds_logic.v(1623)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ne3iu6 ;  // ../RTL/cortexm0ds_logic.v(349)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nephu6 ;  // ../RTL/cortexm0ds_logic.v(162)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nfgax6 ;  // ../RTL/cortexm0ds_logic.v(1644)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nfohu6 ;  // ../RTL/cortexm0ds_logic.v(149)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nfqpw6 ;  // ../RTL/cortexm0ds_logic.v(1600)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ng8iu6 ;  // ../RTL/cortexm0ds_logic.v(416)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ngmiu6 ;  // ../RTL/cortexm0ds_logic.v(604)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nhgbx6 ;  // ../RTL/cortexm0ds_logic.v(1709)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nhlhu6 ;  // ../RTL/cortexm0ds_logic.v(139)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nhthu6 ;  // ../RTL/cortexm0ds_logic.v(216)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nj2qw6 ;  // ../RTL/cortexm0ds_logic.v(1622)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Njjiu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(565)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nkaju6_lutinv ;  // ../RTL/cortexm0ds_logic.v(926)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nkxow6 ;  // ../RTL/cortexm0ds_logic.v(1295)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nlbbx6 ;  // ../RTL/cortexm0ds_logic.v(1700)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nlcbx6 ;  // ../RTL/cortexm0ds_logic.v(1702)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nmabx6 ;  // ../RTL/cortexm0ds_logic.v(1698)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nmfax6 ;  // ../RTL/cortexm0ds_logic.v(1642)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nmohu6 ;  // ../RTL/cortexm0ds_logic.v(151)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nn8iu6 ;  // ../RTL/cortexm0ds_logic.v(419)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nnfbx6 ;  // ../RTL/cortexm0ds_logic.v(1708)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nnuhu6 ;  // ../RTL/cortexm0ds_logic.v(232)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/No3qw6 ;  // ../RTL/cortexm0ds_logic.v(1624)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nodax6 ;  // ../RTL/cortexm0ds_logic.v(1638)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Np7ow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(949)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Npaax6 ;  // ../RTL/cortexm0ds_logic.v(1633)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Npghu6 ;  // ../RTL/cortexm0ds_logic.v(127)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nq4ju6_lutinv ;  // ../RTL/cortexm0ds_logic.v(848)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nr0bx6 ;  // ../RTL/cortexm0ds_logic.v(1681)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nr4iu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(367)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nr7ax6 ;  // ../RTL/cortexm0ds_logic.v(1627)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nrkpw6 ;  // ../RTL/cortexm0ds_logic.v(1589)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nrqpw6 ;  // ../RTL/cortexm0ds_logic.v(1600)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nrxhu6 ;  // ../RTL/cortexm0ds_logic.v(273)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ns8ax6 ;  // ../RTL/cortexm0ds_logic.v(1629)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nsaiu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(448)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nt9bx6 ;  // ../RTL/cortexm0ds_logic.v(1697)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ntuiu6 ;  // ../RTL/cortexm0ds_logic.v(715)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nu5bx6 ;  // ../RTL/cortexm0ds_logic.v(1689)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nu9ow6 ;  // ../RTL/cortexm0ds_logic.v(978)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Numiu6 ;  // ../RTL/cortexm0ds_logic.v(609)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nv3qw6 ;  // ../RTL/cortexm0ds_logic.v(1624)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nv9bx6 ;  // ../RTL/cortexm0ds_logic.v(1697)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nw6iu6 ;  // ../RTL/cortexm0ds_logic.v(396)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nwbbx6 ;  // ../RTL/cortexm0ds_logic.v(1701)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nwdbx6 ;  // ../RTL/cortexm0ds_logic.v(1704)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nwdpw6 ;  // ../RTL/cortexm0ds_logic.v(1514)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nweow6 ;  // ../RTL/cortexm0ds_logic.v(1046)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nwzhu6 ;  // ../RTL/cortexm0ds_logic.v(302)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxrow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1220)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nybbx6 ;  // ../RTL/cortexm0ds_logic.v(1701)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nycow6 ;  // ../RTL/cortexm0ds_logic.v(1020)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nyhpw6 ;  // ../RTL/cortexm0ds_logic.v(1584)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nyiiu6 ;  // ../RTL/cortexm0ds_logic.v(557)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nyxhu6 ;  // ../RTL/cortexm0ds_logic.v(276)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nyxow6 ;  // ../RTL/cortexm0ds_logic.v(1300)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nz2ju6 ;  // ../RTL/cortexm0ds_logic.v(825)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O00iu6 ;  // ../RTL/cortexm0ds_logic.v(304)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O16iu6 ;  // ../RTL/cortexm0ds_logic.v(384)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O1mpw6 ;  // ../RTL/cortexm0ds_logic.v(1592)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O25iu6 ;  // ../RTL/cortexm0ds_logic.v(371)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O2kax6 ;  // ../RTL/cortexm0ds_logic.v(1651)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O34iu6 ;  // ../RTL/cortexm0ds_logic.v(358)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O3xhu6 ;  // ../RTL/cortexm0ds_logic.v(265)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O4bow6 ;  // ../RTL/cortexm0ds_logic.v(995)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O4phu6 ;  // ../RTL/cortexm0ds_logic.v(158)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O59iu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(426)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O5vhu6 ;  // ../RTL/cortexm0ds_logic.v(239)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O70iu6 ;  // ../RTL/cortexm0ds_logic.v(306)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O8lhu6 ;  // ../RTL/cortexm0ds_logic.v(139)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oa4iu6 ;  // ../RTL/cortexm0ds_logic.v(361)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oa5bx6 ;  // ../RTL/cortexm0ds_logic.v(1688)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oarpw6 ;  // ../RTL/cortexm0ds_logic.v(1601)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oaxow6 ;  // ../RTL/cortexm0ds_logic.v(1292)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Obbow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(998)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Obphu6 ;  // ../RTL/cortexm0ds_logic.v(161)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ocniu6 ;  // ../RTL/cortexm0ds_logic.v(616)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ocohu6 ;  // ../RTL/cortexm0ds_logic.v(148)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Od4bx6 ;  // ../RTL/cortexm0ds_logic.v(1687)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Odfiu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(509)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Odgow6 ;  // ../RTL/cortexm0ds_logic.v(1065)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oduhu6 ;  // ../RTL/cortexm0ds_logic.v(228)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oe7iu6 ;  // ../RTL/cortexm0ds_logic.v(402)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oeihu6 ;  // ../RTL/cortexm0ds_logic.v(131)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oetow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1240)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oeziu6 ;  // ../RTL/cortexm0ds_logic.v(777)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Of5ju6_lutinv ;  // ../RTL/cortexm0ds_logic.v(857)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ofkiu6 ;  // ../RTL/cortexm0ds_logic.v(577)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ofmpw6 ;  // ../RTL/cortexm0ds_logic.v(1592)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ogdow6 ;  // ../RTL/cortexm0ds_logic.v(1026)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ogqiu6 ;  // ../RTL/cortexm0ds_logic.v(657)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oh3ju6 ;  // ../RTL/cortexm0ds_logic.v(831)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oh4iu6 ;  // ../RTL/cortexm0ds_logic.v(363)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oh8ax6 ;  // ../RTL/cortexm0ds_logic.v(1628)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ohqhu6 ;  // ../RTL/cortexm0ds_logic.v(176)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ohyax6 ;  // ../RTL/cortexm0ds_logic.v(1677)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oi9ax6 ;  // ../RTL/cortexm0ds_logic.v(1630)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oikax6 ;  // ../RTL/cortexm0ds_logic.v(1651)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ojebx6 ;  // ../RTL/cortexm0ds_logic.v(1706)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ojohu6 ;  // ../RTL/cortexm0ds_logic.v(150)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ok2bx6 ;  // ../RTL/cortexm0ds_logic.v(1684)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ok7ju6 ;  // ../RTL/cortexm0ds_logic.v(886)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ok8iu6 ;  // ../RTL/cortexm0ds_logic.v(418)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Okfax6 ;  // ../RTL/cortexm0ds_logic.v(1642)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oltow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1242)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Om3bx6 ;  // ../RTL/cortexm0ds_logic.v(1686)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Opbax6 ;  // ../RTL/cortexm0ds_logic.v(1635)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oqohu6 ;  // ../RTL/cortexm0ds_logic.v(153)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Orkhu6 ;  // ../RTL/cortexm0ds_logic.v(137)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oruhu6 ;  // ../RTL/cortexm0ds_logic.v(233)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Osthu6 ;  // ../RTL/cortexm0ds_logic.v(220)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ot0bx6 ;  // ../RTL/cortexm0ds_logic.v(1681)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ot7ow6 ;  // ../RTL/cortexm0ds_logic.v(951)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oulpw6 ;  // ../RTL/cortexm0ds_logic.v(1591)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ov3ju6_lutinv ;  // ../RTL/cortexm0ds_logic.v(837)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oveax6 ;  // ../RTL/cortexm0ds_logic.v(1641)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ovihu6 ;  // ../RTL/cortexm0ds_logic.v(132)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ovpiu6 ;  // ../RTL/cortexm0ds_logic.v(649)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Owcax6 ;  // ../RTL/cortexm0ds_logic.v(1637)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Owhbx6 ;  // ../RTL/cortexm0ds_logic.v(1712)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Owoiu6 ;  // ../RTL/cortexm0ds_logic.v(636)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ox9bx6 ;  // ../RTL/cortexm0ds_logic.v(1697)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oxhhu6 ;  // ../RTL/cortexm0ds_logic.v(129)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oxhow6 ;  // ../RTL/cortexm0ds_logic.v(1086)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oxkpw6 ;  // ../RTL/cortexm0ds_logic.v(1589)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oxohu6 ;  // ../RTL/cortexm0ds_logic.v(155)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oy8iu6 ;  // ../RTL/cortexm0ds_logic.v(423)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oyhbx6 ;  // ../RTL/cortexm0ds_logic.v(1712)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ozeiu6 ;  // ../RTL/cortexm0ds_logic.v(504)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0bax6 ;  // ../RTL/cortexm0ds_logic.v(1633)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0biu6 ;  // ../RTL/cortexm0ds_logic.v(451)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0cow6 ;  // ../RTL/cortexm0ds_logic.v(1007)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0ibx6 ;  // ../RTL/cortexm0ds_logic.v(1712)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 ;  // ../RTL/cortexm0ds_logic.v(1650)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P12bx6 ;  // ../RTL/cortexm0ds_logic.v(1683)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P13iu6 ;  // ../RTL/cortexm0ds_logic.v(344)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P14qw6 ;  // ../RTL/cortexm0ds_logic.v(1625)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P1phu6 ;  // ../RTL/cortexm0ds_logic.v(157)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P22iu6 ;  // ../RTL/cortexm0ds_logic.v(331)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P23qw6 ;  // ../RTL/cortexm0ds_logic.v(1623)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P2vhu6 ;  // ../RTL/cortexm0ds_logic.v(237)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P33bx6 ;  // ../RTL/cortexm0ds_logic.v(1685)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P3fiu6 ;  // ../RTL/cortexm0ds_logic.v(505)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P3uow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1249)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P40iu6 ;  // ../RTL/cortexm0ds_logic.v(305)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P4cax6 ;  // ../RTL/cortexm0ds_logic.v(1635)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P4epw6 ;  // ../RTL/cortexm0ds_logic.v(1517)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P4liu6 ;  // ../RTL/cortexm0ds_logic.v(586)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 ;  // ../RTL/cortexm0ds_logic.v(1608)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P73ju6 ;  // ../RTL/cortexm0ds_logic.v(828)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P74iu6 ;  // ../RTL/cortexm0ds_logic.v(360)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P7biu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(453)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P7xhu6 ;  // ../RTL/cortexm0ds_logic.v(266)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P8aiu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(440)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P8oiu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(627)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P8phu6 ;  // ../RTL/cortexm0ds_logic.v(159)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P8viu6 ;  // ../RTL/cortexm0ds_logic.v(721)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P91ju6 ;  // ../RTL/cortexm0ds_logic.v(802)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P92iu6 ;  // ../RTL/cortexm0ds_logic.v(334)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P93qw6 ;  // ../RTL/cortexm0ds_logic.v(1623)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P9bax6 ;  // ../RTL/cortexm0ds_logic.v(1634)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P9niu6 ;  // ../RTL/cortexm0ds_logic.v(614)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pa7ju6 ;  // ../RTL/cortexm0ds_logic.v(882)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pagow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1064)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Panow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1158)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pauhu6 ;  // ../RTL/cortexm0ds_logic.v(227)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pb0iu6 ;  // ../RTL/cortexm0ds_logic.v(308)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pbbbx6 ;  // ../RTL/cortexm0ds_logic.v(1699)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pckiu6 ;  // ../RTL/cortexm0ds_logic.v(575)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pczax6 ;  // ../RTL/cortexm0ds_logic.v(1678)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pdbbx6 ;  // ../RTL/cortexm0ds_logic.v(1700)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pdrhu6 ;  // ../RTL/cortexm0ds_logic.v(188)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pdxax6 ;  // ../RTL/cortexm0ds_logic.v(1675)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pdyax6 ;  // ../RTL/cortexm0ds_logic.v(1676)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pdyow6 ;  // ../RTL/cortexm0ds_logic.v(1306)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pe7ax6 ;  // ../RTL/cortexm0ds_logic.v(1626)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pe9bx6 ;  // ../RTL/cortexm0ds_logic.v(1696)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Peeax6 ;  // ../RTL/cortexm0ds_logic.v(1640)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Peqow6 ;  // ../RTL/cortexm0ds_logic.v(1199)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pexpw6 ;  // ../RTL/cortexm0ds_logic.v(1612)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pfphu6 ;  // ../RTL/cortexm0ds_logic.v(162)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pg3qw6 ;  // ../RTL/cortexm0ds_logic.v(1623)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pgohu6 ;  // ../RTL/cortexm0ds_logic.v(149)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ph1iu6 ;  // ../RTL/cortexm0ds_logic.v(323)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ph8iu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(417)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Phcax6 ;  // ../RTL/cortexm0ds_logic.v(1636)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Phuow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1254)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pifax6 ;  // ../RTL/cortexm0ds_logic.v(1642)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pithu6 ;  // ../RTL/cortexm0ds_logic.v(217)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Piziu6 ;  // ../RTL/cortexm0ds_logic.v(778)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pj7ow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(947)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pjgbx6 ;  // ../RTL/cortexm0ds_logic.v(1709)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pjyiu6 ;  // ../RTL/cortexm0ds_logic.v(765)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pk4ju6 ;  // ../RTL/cortexm0ds_logic.v(846)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pkdow6 ;  // ../RTL/cortexm0ds_logic.v(1028)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pkkbx6 ;  // ../RTL/cortexm0ds_logic.v(1717)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pl4iu6 ;  // ../RTL/cortexm0ds_logic.v(365)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Plcow6 ;  // ../RTL/cortexm0ds_logic.v(1015)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pmlpw6 ;  // ../RTL/cortexm0ds_logic.v(1591)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pmoiu6 ;  // ../RTL/cortexm0ds_logic.v(633)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pnohu6 ;  // ../RTL/cortexm0ds_logic.v(152)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pouhu6 ;  // ../RTL/cortexm0ds_logic.v(232)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pp7iu6 ;  // ../RTL/cortexm0ds_logic.v(406)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ppthu6 ;  // ../RTL/cortexm0ds_logic.v(219)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pqsow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1231)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Prdow6 ;  // ../RTL/cortexm0ds_logic.v(1030)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Psxhu6 ;  // ../RTL/cortexm0ds_logic.v(274)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pt7ax6 ;  // ../RTL/cortexm0ds_logic.v(1627)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pthiu6 ;  // ../RTL/cortexm0ds_logic.v(542)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pu1ju6_lutinv ;  // ../RTL/cortexm0ds_logic.v(809)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Puohu6 ;  // ../RTL/cortexm0ds_logic.v(154)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Puwpw6 ;  // ../RTL/cortexm0ds_logic.v(1611)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pv0bx6 ;  // ../RTL/cortexm0ds_logic.v(1681)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pv9ax6 ;  // ../RTL/cortexm0ds_logic.v(1631)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pvuhu6 ;  // ../RTL/cortexm0ds_logic.v(235)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pwfow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1059)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pxlow6 ;  // ../RTL/cortexm0ds_logic.v(1140)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pxriu6 ;  // ../RTL/cortexm0ds_logic.v(677)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pxzhu6 ;  // ../RTL/cortexm0ds_logic.v(302)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pyjiu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(570)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pyyhu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(289)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pz4iu6 ;  // ../RTL/cortexm0ds_logic.v(370)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pz9bx6 ;  // ../RTL/cortexm0ds_logic.v(1697)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pzxhu6 ;  // ../RTL/cortexm0ds_logic.v(276)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q07ju6_lutinv ;  // ../RTL/cortexm0ds_logic.v(879)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q0fiu6 ;  // ../RTL/cortexm0ds_logic.v(504)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q10iu6 ;  // ../RTL/cortexm0ds_logic.v(304)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q1epw6 ;  // ../RTL/cortexm0ds_logic.v(1516)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q1fow6 ;  // ../RTL/cortexm0ds_logic.v(1048)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q1hbx6 ;  // ../RTL/cortexm0ds_logic.v(1710)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q2eow6 ;  // ../RTL/cortexm0ds_logic.v(1035)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q2gax6 ;  // ../RTL/cortexm0ds_logic.v(1643)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q2ibx6 ;  // ../RTL/cortexm0ds_logic.v(1712)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q34ju6_lutinv ;  // ../RTL/cortexm0ds_logic.v(840)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q3qiu6 ;  // ../RTL/cortexm0ds_logic.v(652)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q3yhu6 ;  // ../RTL/cortexm0ds_logic.v(278)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q44iu6 ;  // ../RTL/cortexm0ds_logic.v(359)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q4dbx6 ;  // ../RTL/cortexm0ds_logic.v(1703)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q4lhu6 ;  // ../RTL/cortexm0ds_logic.v(138)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q5hiu6 ;  // ../RTL/cortexm0ds_logic.v(533)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q5phu6 ;  // ../RTL/cortexm0ds_logic.v(158)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q6fax6 ;  // ../RTL/cortexm0ds_logic.v(1641)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q6vhu6 ;  // ../RTL/cortexm0ds_logic.v(239)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q7miu6 ;  // ../RTL/cortexm0ds_logic.v(600)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q7uow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1250)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q80iu6 ;  // ../RTL/cortexm0ds_logic.v(307)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q89bx6 ;  // ../RTL/cortexm0ds_logic.v(1696)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q8aax6 ;  // ../RTL/cortexm0ds_logic.v(1632)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q8eiu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(494)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q8tow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1237)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q9dax6 ;  // ../RTL/cortexm0ds_logic.v(1638)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qa1qw6 ;  // ../RTL/cortexm0ds_logic.v(1619)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qa5iu6 ;  // ../RTL/cortexm0ds_logic.v(374)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qaciu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(468)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qaipw6 ;  // ../RTL/cortexm0ds_logic.v(1584)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qakbx6 ;  // ../RTL/cortexm0ds_logic.v(1716)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qaqiu6 ;  // ../RTL/cortexm0ds_logic.v(655)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qb3ju6_lutinv ;  // ../RTL/cortexm0ds_logic.v(829)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qc3pw6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1373)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qc5bx6 ;  // ../RTL/cortexm0ds_logic.v(1689)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qcaiu6 ;  // ../RTL/cortexm0ds_logic.v(442)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qcphu6 ;  // ../RTL/cortexm0ds_logic.v(161)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qdhow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1079)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qdvhu6 ;  // ../RTL/cortexm0ds_logic.v(242)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qe8iu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(416)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qehbx6 ;  // ../RTL/cortexm0ds_logic.v(1711)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qeuhu6 ;  // ../RTL/cortexm0ds_logic.v(229)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qf4bx6 ;  // ../RTL/cortexm0ds_logic.v(1687)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qf7iu6 ;  // ../RTL/cortexm0ds_logic.v(403)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qfthu6 ;  // ../RTL/cortexm0ds_logic.v(216)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qgkiu6 ;  // ../RTL/cortexm0ds_logic.v(577)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qh5iu6 ;  // ../RTL/cortexm0ds_logic.v(377)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qiqow6 ;  // ../RTL/cortexm0ds_logic.v(1201)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qj1qw6 ;  // ../RTL/cortexm0ds_logic.v(1620)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qj2ju6 ;  // ../RTL/cortexm0ds_logic.v(819)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qjbbx6 ;  // ../RTL/cortexm0ds_logic.v(1700)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qjcbx6 ;  // ../RTL/cortexm0ds_logic.v(1702)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qjyax6 ;  // ../RTL/cortexm0ds_logic.v(1677)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qk8ju6_lutinv ;  // ../RTL/cortexm0ds_logic.v(899)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qk9pw6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1456)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qkabx6 ;  // ../RTL/cortexm0ds_logic.v(1698)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qkniu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(619)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qkohu6 ;  // ../RTL/cortexm0ds_logic.v(151)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ql8iu6 ;  // ../RTL/cortexm0ds_logic.v(418)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qlfbx6 ;  // ../RTL/cortexm0ds_logic.v(1707)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qmdax6 ;  // ../RTL/cortexm0ds_logic.v(1638)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qmthu6 ;  // ../RTL/cortexm0ds_logic.v(218)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qnkhu6 ;  // ../RTL/cortexm0ds_logic.v(137)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qo3bx6 ;  // ../RTL/cortexm0ds_logic.v(1686)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qodow6 ;  // ../RTL/cortexm0ds_logic.v(1029)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qoyow6 ;  // ../RTL/cortexm0ds_logic.v(1310)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qq3iu6 ;  // ../RTL/cortexm0ds_logic.v(353)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qqhiu6 ;  // ../RTL/cortexm0ds_logic.v(541)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qqiow6 ;  // ../RTL/cortexm0ds_logic.v(1097)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qrgiu6 ;  // ../RTL/cortexm0ds_logic.v(528)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qrihu6 ;  // ../RTL/cortexm0ds_logic.v(132)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qrohu6 ;  // ../RTL/cortexm0ds_logic.v(153)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qsfax6 ;  // ../RTL/cortexm0ds_logic.v(1642)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qsmiu6 ;  // ../RTL/cortexm0ds_logic.v(608)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qsuhu6 ;  // ../RTL/cortexm0ds_logic.v(234)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qtfow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1058)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qudbx6 ;  // ../RTL/cortexm0ds_logic.v(1704)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Queow6 ;  // ../RTL/cortexm0ds_logic.v(1045)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qufax6 ;  // ../RTL/cortexm0ds_logic.v(1643)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qwfax6 ;  // ../RTL/cortexm0ds_logic.v(1643)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qwfbx6 ;  // ../RTL/cortexm0ds_logic.v(1708)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qwxhu6 ;  // ../RTL/cortexm0ds_logic.v(275)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qx0bx6 ;  // ../RTL/cortexm0ds_logic.v(1681)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qxbow6 ;  // ../RTL/cortexm0ds_logic.v(1006)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qxoiu6 ;  // ../RTL/cortexm0ds_logic.v(637)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qy2pw6 ;  // ../RTL/cortexm0ds_logic.v(1367)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qyjax6 ;  // ../RTL/cortexm0ds_logic.v(1650)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qyniu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(624)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qyohu6 ;  // ../RTL/cortexm0ds_logic.v(156)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qz0ju6 ;  // ../RTL/cortexm0ds_logic.v(798)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qzuhu6 ;  // ../RTL/cortexm0ds_logic.v(236)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R04ju6 ;  // ../RTL/cortexm0ds_logic.v(838)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R05iu6 ;  // ../RTL/cortexm0ds_logic.v(370)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R0ghu6 ;  // ../RTL/cortexm0ds_logic.v(125)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R0yhu6 ;  // ../RTL/cortexm0ds_logic.v(277)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R19ax6 ;  // ../RTL/cortexm0ds_logic.v(1629)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R1abx6 ;  // ../RTL/cortexm0ds_logic.v(1697)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R1eax6 ;  // ../RTL/cortexm0ds_logic.v(1639)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R2phu6 ;  // ../RTL/cortexm0ds_logic.v(157)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3giu6 ;  // ../RTL/cortexm0ds_logic.v(519)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3how6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1075)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vhu6 ;  // ../RTL/cortexm0ds_logic.v(238)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 ;  // ../RTL/cortexm0ds_logic.v(1608)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R47ju6_lutinv ;  // ../RTL/cortexm0ds_logic.v(880)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R4miu6 ;  // ../RTL/cortexm0ds_logic.v(599)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R50iu6 ;  // ../RTL/cortexm0ds_logic.v(305)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R5eiu6 ;  // ../RTL/cortexm0ds_logic.v(493)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R5liu6 ;  // ../RTL/cortexm0ds_logic.v(586)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R7kpw6 ;  // ../RTL/cortexm0ds_logic.v(1588)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R83ju6_lutinv ;  // ../RTL/cortexm0ds_logic.v(828)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R84iu6 ;  // ../RTL/cortexm0ds_logic.v(360)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R8xhu6 ;  // ../RTL/cortexm0ds_logic.v(266)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R9aiu6 ;  // ../RTL/cortexm0ds_logic.v(441)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R9mpw6 ;  // ../RTL/cortexm0ds_logic.v(1592)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R9phu6 ;  // ../RTL/cortexm0ds_logic.v(160)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R9wow6 ;  // ../RTL/cortexm0ds_logic.v(1278)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R9yax6 ;  // ../RTL/cortexm0ds_logic.v(1676)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ra2qw6 ;  // ../RTL/cortexm0ds_logic.v(1621)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rb7ju6 ;  // ../RTL/cortexm0ds_logic.v(883)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rbuhu6 ;  // ../RTL/cortexm0ds_logic.v(227)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rc7iu6 ;  // ../RTL/cortexm0ds_logic.v(402)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rcliu6 ;  // ../RTL/cortexm0ds_logic.v(589)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rcziu6 ;  // ../RTL/cortexm0ds_logic.v(776)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rdkiu6 ;  // ../RTL/cortexm0ds_logic.v(576)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rerow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1213)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rezax6 ;  // ../RTL/cortexm0ds_logic.v(1678)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rfxax6 ;  // ../RTL/cortexm0ds_logic.v(1675)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rfxhu6 ;  // ../RTL/cortexm0ds_logic.v(269)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rg9ax6 ;  // ../RTL/cortexm0ds_logic.v(1630)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rgoiu6 ;  // ../RTL/cortexm0ds_logic.v(630)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rhgiu6 ;  // ../RTL/cortexm0ds_logic.v(524)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rhkpw6 ;  // ../RTL/cortexm0ds_logic.v(1588)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rhniu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(617)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rhohu6 ;  // ../RTL/cortexm0ds_logic.v(149)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rhoow6 ;  // ../RTL/cortexm0ds_logic.v(1174)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rhvhu6 ;  // ../RTL/cortexm0ds_logic.v(243)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rijbx6 ;  // ../RTL/cortexm0ds_logic.v(1715)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rilpw6 ;  // ../RTL/cortexm0ds_logic.v(1590)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rimiu6 ;  // ../RTL/cortexm0ds_logic.v(604)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rjthu6 ;  // ../RTL/cortexm0ds_logic.v(217)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rjtow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1241)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rjziu6 ;  // ../RTL/cortexm0ds_logic.v(779)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rk1bx6 ;  // ../RTL/cortexm0ds_logic.v(1682)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rk5ju6 ;  // ../RTL/cortexm0ds_logic.v(859)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rkbax6 ;  // ../RTL/cortexm0ds_logic.v(1634)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rkkax6 ;  // ../RTL/cortexm0ds_logic.v(1651)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rkkiu6 ;  // ../RTL/cortexm0ds_logic.v(578)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rksow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1228)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rkzhu6 ;  // ../RTL/cortexm0ds_logic.v(298)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rlgbx6 ;  // ../RTL/cortexm0ds_logic.v(1709)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rm2bx6 ;  // ../RTL/cortexm0ds_logic.v(1684)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rmbpw6 ;  // ../RTL/cortexm0ds_logic.v(1483)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rmcow6 ;  // ../RTL/cortexm0ds_logic.v(1015)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rmiiu6 ;  // ../RTL/cortexm0ds_logic.v(552)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rnaax6 ;  // ../RTL/cortexm0ds_logic.v(1632)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rnbow6 ;  // ../RTL/cortexm0ds_logic.v(1002)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ro1ju6 ;  // ../RTL/cortexm0ds_logic.v(807)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ro2pw6 ;  // ../RTL/cortexm0ds_logic.v(1364)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ro8ax6 ;  // ../RTL/cortexm0ds_logic.v(1629)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Roohu6 ;  // ../RTL/cortexm0ds_logic.v(152)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rpuhu6 ;  // ../RTL/cortexm0ds_logic.v(233)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rq0qw6 ;  // ../RTL/cortexm0ds_logic.v(1618)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rqthu6 ;  // ../RTL/cortexm0ds_logic.v(220)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rr3qw6 ;  // ../RTL/cortexm0ds_logic.v(1624)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rs4ju6_lutinv ;  // ../RTL/cortexm0ds_logic.v(849)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rs5pw6 ;  // ../RTL/cortexm0ds_logic.v(1405)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rskax6 ;  // ../RTL/cortexm0ds_logic.v(1652)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rsyhu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(287)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rt4pw6 ;  // ../RTL/cortexm0ds_logic.v(1392)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rteax6 ;  // ../RTL/cortexm0ds_logic.v(1641)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rtxhu6 ;  // ../RTL/cortexm0ds_logic.v(274)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ru2ju6 ;  // ../RTL/cortexm0ds_logic.v(823)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rucax6 ;  // ../RTL/cortexm0ds_logic.v(1637)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rupow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1192)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rv7ax6 ;  // ../RTL/cortexm0ds_logic.v(1627)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rvniu6 ;  // ../RTL/cortexm0ds_logic.v(623)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rw1iu6 ;  // ../RTL/cortexm0ds_logic.v(329)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rw8iu6 ;  // ../RTL/cortexm0ds_logic.v(422)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rwgow6 ;  // ../RTL/cortexm0ds_logic.v(1072)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rwjax6 ;  // ../RTL/cortexm0ds_logic.v(1650)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rwuhu6 ;  // ../RTL/cortexm0ds_logic.v(235)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ry2qw6 ;  // ../RTL/cortexm0ds_logic.v(1622)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ryfax6 ;  // ../RTL/cortexm0ds_logic.v(1643)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ryzhu6 ;  // ../RTL/cortexm0ds_logic.v(303)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rz0bx6 ;  // ../RTL/cortexm0ds_logic.v(1681)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rz8bx6 ;  // ../RTL/cortexm0ds_logic.v(1695)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rzciu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(477)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S02iu6 ;  // ../RTL/cortexm0ds_logic.v(330)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S0kbx6 ;  // ../RTL/cortexm0ds_logic.v(1716)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S0lhu6 ;  // ../RTL/cortexm0ds_logic.v(138)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S0vhu6 ;  // ../RTL/cortexm0ds_logic.v(237)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S11bx6 ;  // ../RTL/cortexm0ds_logic.v(1681)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S18iu6 ;  // ../RTL/cortexm0ds_logic.v(411)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S1fiu6 ;  // ../RTL/cortexm0ds_logic.v(505)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S1tiu6 ;  // ../RTL/cortexm0ds_logic.v(692)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S20iu6 ;  // ../RTL/cortexm0ds_logic.v(304)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S2cax6 ;  // ../RTL/cortexm0ds_logic.v(1635)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S2cbx6 ;  // ../RTL/cortexm0ds_logic.v(1701)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S2epw6 ;  // ../RTL/cortexm0ds_logic.v(1516)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S2ziu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(772)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S32bx6 ;  // ../RTL/cortexm0ds_logic.v(1683)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S3kiu6 ;  // ../RTL/cortexm0ds_logic.v(572)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S3mpw6 ;  // ../RTL/cortexm0ds_logic.v(1592)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S4kbx6 ;  // ../RTL/cortexm0ds_logic.v(1716)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S53bx6 ;  // ../RTL/cortexm0ds_logic.v(1685)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S54iu6 ;  // ../RTL/cortexm0ds_logic.v(359)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S5biu6 ;  // ../RTL/cortexm0ds_logic.v(453)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S63iu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(346)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S6ihu6 ;  // ../RTL/cortexm0ds_logic.v(130)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S6phu6 ;  // ../RTL/cortexm0ds_logic.v(159)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S7mpw6 ;  // ../RTL/cortexm0ds_logic.v(1592)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S7vhu6 ;  // ../RTL/cortexm0ds_logic.v(239)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S88iu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(414)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S8uhu6 ;  // ../RTL/cortexm0ds_logic.v(226)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S90iu6 ;  // ../RTL/cortexm0ds_logic.v(307)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S98ow6 ;  // ../RTL/cortexm0ds_logic.v(957)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sb8ax6 ;  // ../RTL/cortexm0ds_logic.v(1628)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sbfax6 ;  // ../RTL/cortexm0ds_logic.v(1642)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sbrow6 ;  // ../RTL/cortexm0ds_logic.v(1212)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sbyhu6 ;  // ../RTL/cortexm0ds_logic.v(281)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Scbiu6 ;  // ../RTL/cortexm0ds_logic.v(455)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sd8ax6 ;  // ../RTL/cortexm0ds_logic.v(1628)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sddbx6 ;  // ../RTL/cortexm0ds_logic.v(1703)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sdlhu6 ;  // ../RTL/cortexm0ds_logic.v(139)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sdlpw6 ;  // ../RTL/cortexm0ds_logic.v(1590)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sdoiu6 ;  // ../RTL/cortexm0ds_logic.v(629)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sdphu6 ;  // ../RTL/cortexm0ds_logic.v(161)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sdwow6 ;  // ../RTL/cortexm0ds_logic.v(1279)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sejax6 ;  // ../RTL/cortexm0ds_logic.v(1649)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Seohu6 ;  // ../RTL/cortexm0ds_logic.v(148)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sf1iu6 ;  // ../RTL/cortexm0ds_logic.v(323)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sf8iu6 ;  // ../RTL/cortexm0ds_logic.v(416)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sg7iu6 ;  // ../RTL/cortexm0ds_logic.v(403)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sgjax6 ;  // ../RTL/cortexm0ds_logic.v(1649)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sgthu6 ;  // ../RTL/cortexm0ds_logic.v(216)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sh4bx6 ;  // ../RTL/cortexm0ds_logic.v(1687)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sh7ow6 ;  // ../RTL/cortexm0ds_logic.v(947)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Shopw6 ;  // ../RTL/cortexm0ds_logic.v(1596)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sijax6 ;  // ../RTL/cortexm0ds_logic.v(1650)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sjkhu6 ;  // ../RTL/cortexm0ds_logic.v(137)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sjqow6 ;  // ../RTL/cortexm0ds_logic.v(1201)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Skjax6 ;  // ../RTL/cortexm0ds_logic.v(1650)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Slohu6 ;  // ../RTL/cortexm0ds_logic.v(151)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Slyax6 ;  // ../RTL/cortexm0ds_logic.v(1677)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Smjax6 ;  // ../RTL/cortexm0ds_logic.v(1650)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Smnow6 ;  // ../RTL/cortexm0ds_logic.v(1162)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Smuhu6 ;  // ../RTL/cortexm0ds_logic.v(232)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sn4bx6 ;  // ../RTL/cortexm0ds_logic.v(1687)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sn7iu6 ;  // ../RTL/cortexm0ds_logic.v(406)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Snihu6 ;  // ../RTL/cortexm0ds_logic.v(131)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Snthu6 ;  // ../RTL/cortexm0ds_logic.v(219)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 ;  // ../RTL/cortexm0ds_logic.v(1650)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sokiu6 ;  // ../RTL/cortexm0ds_logic.v(580)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Spyhu6 ;  // ../RTL/cortexm0ds_logic.v(286)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sq3bx6 ;  // ../RTL/cortexm0ds_logic.v(1686)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sq3ju6 ;  // ../RTL/cortexm0ds_logic.v(835)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sq4iu6 ;  // ../RTL/cortexm0ds_logic.v(367)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sqfax6 ;  // ../RTL/cortexm0ds_logic.v(1642)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sqjax6 ;  // ../RTL/cortexm0ds_logic.v(1650)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sqkax6 ;  // ../RTL/cortexm0ds_logic.v(1652)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sqqhu6 ;  // ../RTL/cortexm0ds_logic.v(180)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sqwpw6 ;  // ../RTL/cortexm0ds_logic.v(1611)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Srbow6 ;  // ../RTL/cortexm0ds_logic.v(1004)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ss0qw6 ;  // ../RTL/cortexm0ds_logic.v(1618)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6 ;  // ../RTL/cortexm0ds_logic.v(1650)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssohu6 ;  // ../RTL/cortexm0ds_logic.v(154)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/St1iu6 ;  // ../RTL/cortexm0ds_logic.v(328)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Stkpw6 ;  // ../RTL/cortexm0ds_logic.v(1589)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Stmiu6 ;  // ../RTL/cortexm0ds_logic.v(609)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Stuhu6 ;  // ../RTL/cortexm0ds_logic.v(234)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Stuow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1259)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Su8ax6 ;  // ../RTL/cortexm0ds_logic.v(1629)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sujax6 ;  // ../RTL/cortexm0ds_logic.v(1650)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Svzhu6 ;  // ../RTL/cortexm0ds_logic.v(302)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Swjbx6 ;  // ../RTL/cortexm0ds_logic.v(1715)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Swyhu6 ;  // ../RTL/cortexm0ds_logic.v(289)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sx3qw6 ;  // ../RTL/cortexm0ds_logic.v(1624)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sxxhu6 ;  // ../RTL/cortexm0ds_logic.v(276)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sy2ju6 ;  // ../RTL/cortexm0ds_logic.v(824)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Syjbx6 ;  // ../RTL/cortexm0ds_logic.v(1715)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sz3qw6 ;  // ../RTL/cortexm0ds_logic.v(1625)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Szohu6 ;  // ../RTL/cortexm0ds_logic.v(156)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T05ju6 ;  // ../RTL/cortexm0ds_logic.v(852)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T0ipw6 ;  // ../RTL/cortexm0ds_logic.v(1584)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T0zhu6 ;  // ../RTL/cortexm0ds_logic.v(290)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T0zow6 ;  // ../RTL/cortexm0ds_logic.v(1315)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T14ju6 ;  // ../RTL/cortexm0ds_logic.v(839)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1jiu6 ;  // ../RTL/cortexm0ds_logic.v(558)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 ;  // ../RTL/cortexm0ds_logic.v(1608)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1yhu6 ;  // ../RTL/cortexm0ds_logic.v(277)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T23ju6_lutinv ;  // ../RTL/cortexm0ds_logic.v(826)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T24iu6 ;  // ../RTL/cortexm0ds_logic.v(358)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T2dbx6 ;  // ../RTL/cortexm0ds_logic.v(1703)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T2kbx6 ;  // ../RTL/cortexm0ds_logic.v(1716)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T2xhu6 ;  // ../RTL/cortexm0ds_logic.v(264)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T33iu6 ;  // ../RTL/cortexm0ds_logic.v(345)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T3abx6 ;  // ../RTL/cortexm0ds_logic.v(1697)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T3opw6 ;  // ../RTL/cortexm0ds_logic.v(1595)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T3phu6 ;  // ../RTL/cortexm0ds_logic.v(158)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T41ju6 ;  // ../RTL/cortexm0ds_logic.v(800)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T4vhu6 ;  // ../RTL/cortexm0ds_logic.v(238)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T5mpw6 ;  // ../RTL/cortexm0ds_logic.v(1592)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T5yax6 ;  // ../RTL/cortexm0ds_logic.v(1676)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T6aax6 ;  // ../RTL/cortexm0ds_logic.v(1632)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T6kbx6 ;  // ../RTL/cortexm0ds_logic.v(1716)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T6ziu6 ;  // ../RTL/cortexm0ds_logic.v(774)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T75ju6 ;  // ../RTL/cortexm0ds_logic.v(854)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T7bax6 ;  // ../RTL/cortexm0ds_logic.v(1634)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T82qw6 ;  // ../RTL/cortexm0ds_logic.v(1621)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T8kbx6 ;  // ../RTL/cortexm0ds_logic.v(1716)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T94iu6 ;  // ../RTL/cortexm0ds_logic.v(360)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T9kpw6 ;  // ../RTL/cortexm0ds_logic.v(1588)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T9qow6 ;  // ../RTL/cortexm0ds_logic.v(1198)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tajax6 ;  // ../RTL/cortexm0ds_logic.v(1649)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Taphu6 ;  // ../RTL/cortexm0ds_logic.v(160)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tb3qw6 ;  // ../RTL/cortexm0ds_logic.v(1623)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tbohu6 ;  // ../RTL/cortexm0ds_logic.v(147)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tbvhu6 ;  // ../RTL/cortexm0ds_logic.v(241)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tc8iu6 ;  // ../RTL/cortexm0ds_logic.v(415)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tc9bx6 ;  // ../RTL/cortexm0ds_logic.v(1696)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tceax6 ;  // ../RTL/cortexm0ds_logic.v(1640)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tchbx6 ;  // ../RTL/cortexm0ds_logic.v(1711)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tcipw6 ;  // ../RTL/cortexm0ds_logic.v(1585)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tcjax6 ;  // ../RTL/cortexm0ds_logic.v(1649)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tcjbx6 ;  // ../RTL/cortexm0ds_logic.v(1714)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tcuhu6 ;  // ../RTL/cortexm0ds_logic.v(228)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Td7iu6 ;  // ../RTL/cortexm0ds_logic.v(402)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tdtow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1239)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tekiu6 ;  // ../RTL/cortexm0ds_logic.v(576)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tezhu6 ;  // ../RTL/cortexm0ds_logic.v(295)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tfcax6 ;  // ../RTL/cortexm0ds_logic.v(1636)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgcow6 ;  // ../RTL/cortexm0ds_logic.v(1013)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgkbx6 ;  // ../RTL/cortexm0ds_logic.v(1716)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgzax6 ;  // ../RTL/cortexm0ds_logic.v(1678)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Thcbx6 ;  // ../RTL/cortexm0ds_logic.v(1702)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Thiax6 ;  // ../RTL/cortexm0ds_logic.v(1648)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Thxax6 ;  // ../RTL/cortexm0ds_logic.v(1675)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tikbx6 ;  // ../RTL/cortexm0ds_logic.v(1716)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tivhu6 ;  // ../RTL/cortexm0ds_logic.v(243)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tj1iu6 ;  // ../RTL/cortexm0ds_logic.v(324)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tjfbx6 ;  // ../RTL/cortexm0ds_logic.v(1707)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tjkpw6 ;  // ../RTL/cortexm0ds_logic.v(1589)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tkdax6 ;  // ../RTL/cortexm0ds_logic.v(1638)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tkfow6 ;  // ../RTL/cortexm0ds_logic.v(1055)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tkjbx6 ;  // ../RTL/cortexm0ds_logic.v(1715)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tktow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1242)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tl4bx6 ;  // ../RTL/cortexm0ds_logic.v(1687)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tlebx6 ;  // ../RTL/cortexm0ds_logic.v(1706)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tmjbx6 ;  // ../RTL/cortexm0ds_logic.v(1715)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tmqiu6 ;  // ../RTL/cortexm0ds_logic.v(659)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tmrow6 ;  // ../RTL/cortexm0ds_logic.v(1216)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tngbx6 ;  // ../RTL/cortexm0ds_logic.v(1709)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/To2ju6_lutinv ;  // ../RTL/cortexm0ds_logic.v(821)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tokax6 ;  // ../RTL/cortexm0ds_logic.v(1652)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tpohu6 ;  // ../RTL/cortexm0ds_logic.v(152)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tptpw6 ;  // ../RTL/cortexm0ds_logic.v(1605)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tquhu6 ;  // ../RTL/cortexm0ds_logic.v(233)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tsdbx6 ;  // ../RTL/cortexm0ds_logic.v(1704)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tsriu6 ;  // ../RTL/cortexm0ds_logic.v(675)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tszhu6 ;  // ../RTL/cortexm0ds_logic.v(301)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tt4ju6_lutinv ;  // ../RTL/cortexm0ds_logic.v(849)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tt9ax6 ;  // ../RTL/cortexm0ds_logic.v(1631)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ttmhu6 ;  // ../RTL/cortexm0ds_logic.v(143)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tu3ju6 ;  // ../RTL/cortexm0ds_logic.v(836)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tu4iu6 ;  // ../RTL/cortexm0ds_logic.v(368)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tucow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1018)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tujbx6 ;  // ../RTL/cortexm0ds_logic.v(1715)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tw2iu6 ;  // ../RTL/cortexm0ds_logic.v(342)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Twohu6 ;  // ../RTL/cortexm0ds_logic.v(155)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tx8iu6 ;  // ../RTL/cortexm0ds_logic.v(423)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tyaax6 ;  // ../RTL/cortexm0ds_logic.v(1633)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tyipw6 ;  // ../RTL/cortexm0ds_logic.v(1586)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tzdiu6 ;  // ../RTL/cortexm0ds_logic.v(490)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tzgbx6 ;  // ../RTL/cortexm0ds_logic.v(1710)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tzsow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1234)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tzzhu6 ;  // ../RTL/cortexm0ds_logic.v(303)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U03iu6 ;  // ../RTL/cortexm0ds_logic.v(344)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U0oiu6 ;  // ../RTL/cortexm0ds_logic.v(625)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U0phu6 ;  // ../RTL/cortexm0ds_logic.v(157)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U19iu6 ;  // ../RTL/cortexm0ds_logic.v(424)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U1kpw6 ;  // ../RTL/cortexm0ds_logic.v(1588)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U1uiu6 ;  // ../RTL/cortexm0ds_logic.v(705)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U1vhu6 ;  // ../RTL/cortexm0ds_logic.v(237)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U28iu6 ;  // ../RTL/cortexm0ds_logic.v(411)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U2fiu6 ;  // ../RTL/cortexm0ds_logic.v(505)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U30iu6 ;  // ../RTL/cortexm0ds_logic.v(305)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U31bx6 ;  // ../RTL/cortexm0ds_logic.v(1681)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U3epw6 ;  // ../RTL/cortexm0ds_logic.v(1516)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U4fax6 ;  // ../RTL/cortexm0ds_logic.v(1641)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U5yhu6 ;  // ../RTL/cortexm0ds_logic.v(279)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U64iu6 ;  // ../RTL/cortexm0ds_logic.v(359)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U6wiu6 ;  // ../RTL/cortexm0ds_logic.v(734)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U6xhu6 ;  // ../RTL/cortexm0ds_logic.v(266)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U73iu6 ;  // ../RTL/cortexm0ds_logic.v(346)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U7dax6 ;  // ../RTL/cortexm0ds_logic.v(1637)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U7phu6 ;  // ../RTL/cortexm0ds_logic.v(159)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U8jax6 ;  // ../RTL/cortexm0ds_logic.v(1649)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U8uiu6 ;  // ../RTL/cortexm0ds_logic.v(708)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U8vhu6 ;  // ../RTL/cortexm0ds_logic.v(240)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U98iu6 ;  // ../RTL/cortexm0ds_logic.v(414)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U99ow6 ;  // ../RTL/cortexm0ds_logic.v(970)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9now6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1158)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9uhu6 ;  // ../RTL/cortexm0ds_logic.v(227)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9ypw6 ;  // ../RTL/cortexm0ds_logic.v(1614)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ua0iu6 ;  // ../RTL/cortexm0ds_logic.v(307)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ua9bx6 ;  // ../RTL/cortexm0ds_logic.v(1696)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ubypw6 ;  // ../RTL/cortexm0ds_logic.v(1614)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uc4ju6 ;  // ../RTL/cortexm0ds_logic.v(843)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ud4iu6 ;  // ../RTL/cortexm0ds_logic.v(362)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ue9ax6 ;  // ../RTL/cortexm0ds_logic.v(1630)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ueapw6 ;  // ../RTL/cortexm0ds_logic.v(1467)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uehiu6 ;  // ../RTL/cortexm0ds_logic.v(536)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uephu6 ;  // ../RTL/cortexm0ds_logic.v(162)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uf9iu6 ;  // ../RTL/cortexm0ds_logic.v(430)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufbbx6 ;  // ../RTL/cortexm0ds_logic.v(1700)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufebx6 ;  // ../RTL/cortexm0ds_logic.v(1705)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufkhu6 ;  // ../RTL/cortexm0ds_logic.v(136)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufohu6 ;  // ../RTL/cortexm0ds_logic.v(149)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 ;  // ../RTL/cortexm0ds_logic.v(1596)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufvhu6 ;  // ../RTL/cortexm0ds_logic.v(242)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ug8iu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(417)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ugmiu6 ;  // ../RTL/cortexm0ds_logic.v(604)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uh2qw6 ;  // ../RTL/cortexm0ds_logic.v(1622)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uhthu6 ;  // ../RTL/cortexm0ds_logic.v(216)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uilhu6 ;  // ../RTL/cortexm0ds_logic.v(139)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uizax6 ;  // ../RTL/cortexm0ds_logic.v(1678)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uj4bx6 ;  // ../RTL/cortexm0ds_logic.v(1687)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uj4ju6 ;  // ../RTL/cortexm0ds_logic.v(846)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ujihu6 ;  // ../RTL/cortexm0ds_logic.v(131)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ujjiu6 ;  // ../RTL/cortexm0ds_logic.v(565)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ujspw6 ;  // ../RTL/cortexm0ds_logic.v(1603)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ujxax6 ;  // ../RTL/cortexm0ds_logic.v(1675)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ukbpw6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1483)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ukcow6 ;  // ../RTL/cortexm0ds_logic.v(1015)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Umkax6 ;  // ../RTL/cortexm0ds_logic.v(1652)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Umniu6 ;  // ../RTL/cortexm0ds_logic.v(619)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Umohu6 ;  // ../RTL/cortexm0ds_logic.v(151)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Umuiu6 ;  // ../RTL/cortexm0ds_logic.v(713)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Unyax6 ;  // ../RTL/cortexm0ds_logic.v(1677)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uo2bx6 ;  // ../RTL/cortexm0ds_logic.v(1684)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uofax6 ;  // ../RTL/cortexm0ds_logic.v(1642)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uojbx6 ;  // ../RTL/cortexm0ds_logic.v(1715)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uoliu6 ;  // ../RTL/cortexm0ds_logic.v(593)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uosiu6 ;  // ../RTL/cortexm0ds_logic.v(687)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Up4bx6 ;  // ../RTL/cortexm0ds_logic.v(1687)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Upsow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1230)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uqyow6 ;  // ../RTL/cortexm0ds_logic.v(1311)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ur4iu6 ;  // ../RTL/cortexm0ds_logic.v(367)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ureax6 ;  // ../RTL/cortexm0ds_logic.v(1640)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Urgbx6 ;  // ../RTL/cortexm0ds_logic.v(1710)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Urxhu6 ;  // ../RTL/cortexm0ds_logic.v(274)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Us2ju6 ;  // ../RTL/cortexm0ds_logic.v(822)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Us3bx6 ;  // ../RTL/cortexm0ds_logic.v(1686)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Usaiu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(448)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uscax6 ;  // ../RTL/cortexm0ds_logic.v(1637)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Usipw6 ;  // ../RTL/cortexm0ds_logic.v(1585)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Usjbx6 ;  // ../RTL/cortexm0ds_logic.v(1715)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Usnpw6 ;  // ../RTL/cortexm0ds_logic.v(1595)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Utgiu6 ;  // ../RTL/cortexm0ds_logic.v(528)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Utniu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(622)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Utohu6 ;  // ../RTL/cortexm0ds_logic.v(154)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Utqpw6 ;  // ../RTL/cortexm0ds_logic.v(1600)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uu1iu6 ;  // ../RTL/cortexm0ds_logic.v(328)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uu8iu6 ;  // ../RTL/cortexm0ds_logic.v(422)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uu9ow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(978)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uunpw6 ;  // ../RTL/cortexm0ds_logic.v(1595)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uuuhu6 ;  // ../RTL/cortexm0ds_logic.v(235)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uvliu6 ;  // ../RTL/cortexm0ds_logic.v(596)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uvsiu6 ;  // ../RTL/cortexm0ds_logic.v(690)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uwdpw6 ;  // ../RTL/cortexm0ds_logic.v(1514)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uwkhu6 ;  // ../RTL/cortexm0ds_logic.v(138)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uwzhu6 ;  // ../RTL/cortexm0ds_logic.v(302)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uwzow6 ;  // ../RTL/cortexm0ds_logic.v(1327)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ux5iu6 ;  // ../RTL/cortexm0ds_logic.v(383)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ux8bx6 ;  // ../RTL/cortexm0ds_logic.v(1695)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uy4iu6 ;  // ../RTL/cortexm0ds_logic.v(370)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uybpw6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1488)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uyiiu6 ;  // ../RTL/cortexm0ds_logic.v(557)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uyxhu6 ;  // ../RTL/cortexm0ds_logic.v(276)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uzaiu6 ;  // ../RTL/cortexm0ds_logic.v(450)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V00iu6 ;  // ../RTL/cortexm0ds_logic.v(304)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V0cax6 ;  // ../RTL/cortexm0ds_logic.v(1635)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V0jpw6 ;  // ../RTL/cortexm0ds_logic.v(1586)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V17ow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(941)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V1low6 ;  // ../RTL/cortexm0ds_logic.v(1128)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V1sow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1221)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V2kow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1115)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V2row6 ;  // ../RTL/cortexm0ds_logic.v(1208)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V34iu6 ;  // ../RTL/cortexm0ds_logic.v(358)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V3cow6 ;  // ../RTL/cortexm0ds_logic.v(1008)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V3qhu6 ;  // ../RTL/cortexm0ds_logic.v(171)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V3xhu6 ;  // ../RTL/cortexm0ds_logic.v(265)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V4phu6 ;  // ../RTL/cortexm0ds_logic.v(158)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V52bx6 ;  // ../RTL/cortexm0ds_logic.v(1683)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V52iu6 ;  // ../RTL/cortexm0ds_logic.v(332)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V53qw6 ;  // ../RTL/cortexm0ds_logic.v(1623)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V59iu6 ;  // ../RTL/cortexm0ds_logic.v(426)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V5abx6 ;  // ../RTL/cortexm0ds_logic.v(1697)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V5oow6 ;  // ../RTL/cortexm0ds_logic.v(1169)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V5vhu6 ;  // ../RTL/cortexm0ds_logic.v(239)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V6jax6 ;  // ../RTL/cortexm0ds_logic.v(1649)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V6now6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1156)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V70iu6 ;  // ../RTL/cortexm0ds_logic.v(306)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V73bx6 ;  // ../RTL/cortexm0ds_logic.v(1685)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V77pw6 ;  // ../RTL/cortexm0ds_logic.v(1424)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Va7ax6 ;  // ../RTL/cortexm0ds_logic.v(1626)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vacow6 ;  // ../RTL/cortexm0ds_logic.v(1011)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vbiow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1091)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vbphu6 ;  // ../RTL/cortexm0ds_logic.v(161)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vbspw6 ;  // ../RTL/cortexm0ds_logic.v(1603)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vcohu6 ;  // ../RTL/cortexm0ds_logic.v(148)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vdmiu6 ;  // ../RTL/cortexm0ds_logic.v(603)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vduhu6 ;  // ../RTL/cortexm0ds_logic.v(228)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ve7iu6 ;  // ../RTL/cortexm0ds_logic.v(402)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vefax6 ;  // ../RTL/cortexm0ds_logic.v(1642)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Veziu6 ;  // ../RTL/cortexm0ds_logic.v(777)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vfkiu6 ;  // ../RTL/cortexm0ds_logic.v(577)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vgjpw6 ;  // ../RTL/cortexm0ds_logic.v(1587)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vhcow6 ;  // ../RTL/cortexm0ds_logic.v(1013)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vhspw6 ;  // ../RTL/cortexm0ds_logic.v(1603)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vibax6 ;  // ../RTL/cortexm0ds_logic.v(1634)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vihiu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(538)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vioiu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(631)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vj3qw6 ;  // ../RTL/cortexm0ds_logic.v(1624)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vjniu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(618)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vjohu6 ;  // ../RTL/cortexm0ds_logic.v(150)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vk1iu6 ;  // ../RTL/cortexm0ds_logic.v(324)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vkzax6 ;  // ../RTL/cortexm0ds_logic.v(1679)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vlaax6 ;  // ../RTL/cortexm0ds_logic.v(1632)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vlxax6 ;  // ../RTL/cortexm0ds_logic.v(1675)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vmipw6 ;  // ../RTL/cortexm0ds_logic.v(1585)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vn9bx6 ;  // ../RTL/cortexm0ds_logic.v(1696)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vo3ju6_lutinv ;  // ../RTL/cortexm0ds_logic.v(834)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vobiu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(460)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Voqow6 ;  // ../RTL/cortexm0ds_logic.v(1203)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vowiu6 ;  // ../RTL/cortexm0ds_logic.v(740)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Voxow6 ;  // ../RTL/cortexm0ds_logic.v(1297)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vpgbx6 ;  // ../RTL/cortexm0ds_logic.v(1709)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vpkpw6 ;  // ../RTL/cortexm0ds_logic.v(1589)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vplpw6 ;  // ../RTL/cortexm0ds_logic.v(1591)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vpoiu6 ;  // ../RTL/cortexm0ds_logic.v(634)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vpphu6 ;  // ../RTL/cortexm0ds_logic.v(166)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vqgax6 ;  // ../RTL/cortexm0ds_logic.v(1644)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vqjbx6 ;  // ../RTL/cortexm0ds_logic.v(1715)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vqohu6 ;  // ../RTL/cortexm0ds_logic.v(153)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vr1iu6 ;  // ../RTL/cortexm0ds_logic.v(327)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vrmiu6 ;  // ../RTL/cortexm0ds_logic.v(608)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vrtpw6 ;  // ../RTL/cortexm0ds_logic.v(1606)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vruhu6 ;  // ../RTL/cortexm0ds_logic.v(233)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vs0iu6 ;  // ../RTL/cortexm0ds_logic.v(314)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vs7pw6 ;  // ../RTL/cortexm0ds_logic.v(1432)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vsthu6 ;  // ../RTL/cortexm0ds_logic.v(220)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vtzhu6 ;  // ../RTL/cortexm0ds_logic.v(301)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vu5iu6 ;  // ../RTL/cortexm0ds_logic.v(382)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vuciu6 ;  // ../RTL/cortexm0ds_logic.v(475)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vviiu6 ;  // ../RTL/cortexm0ds_logic.v(556)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vvpiu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(649)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vvxhu6 ;  // ../RTL/cortexm0ds_logic.v(275)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vwapw6 ;  // ../RTL/cortexm0ds_logic.v(1474)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vx9iu6 ;  // ../RTL/cortexm0ds_logic.v(436)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vxniu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(623)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vyfbx6 ;  // ../RTL/cortexm0ds_logic.v(1708)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vygax6 ;  // ../RTL/cortexm0ds_logic.v(1645)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vynow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1167)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vyuhu6 ;  // ../RTL/cortexm0ds_logic.v(236)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vz8ax6 ;  // ../RTL/cortexm0ds_logic.v(1629)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzdax6 ;  // ../RTL/cortexm0ds_logic.v(1639)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzeiu6 ;  // ../RTL/cortexm0ds_logic.v(504)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzjpw6 ;  // ../RTL/cortexm0ds_logic.v(1588)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ;  // ../RTL/cortexm0ds_logic.v(1608)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W0dbx6 ;  // ../RTL/cortexm0ds_logic.v(1703)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W0jax6 ;  // ../RTL/cortexm0ds_logic.v(1649)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W0piu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(638)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W13iu6 ;  // ../RTL/cortexm0ds_logic.v(344)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W1phu6 ;  // ../RTL/cortexm0ds_logic.v(157)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W1wow6 ;  // ../RTL/cortexm0ds_logic.v(1275)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W2jax6 ;  // ../RTL/cortexm0ds_logic.v(1649)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W2vhu6 ;  // ../RTL/cortexm0ds_logic.v(238)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W38pw6 ;  // ../RTL/cortexm0ds_logic.v(1436)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W40iu6 ;  // ../RTL/cortexm0ds_logic.v(305)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W48ow6 ;  // ../RTL/cortexm0ds_logic.v(955)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4aax6 ;  // ../RTL/cortexm0ds_logic.v(1631)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4epw6 ;  // ../RTL/cortexm0ds_logic.v(1517)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4fow6 ;  // ../RTL/cortexm0ds_logic.v(1049)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4jax6 ;  // ../RTL/cortexm0ds_logic.v(1649)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4siu6 ;  // ../RTL/cortexm0ds_logic.v(680)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W51bx6 ;  // ../RTL/cortexm0ds_logic.v(1681)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W5shu6 ;  // ../RTL/cortexm0ds_logic.v(199)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W5ypw6 ;  // ../RTL/cortexm0ds_logic.v(1614)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W6ipw6 ;  // ../RTL/cortexm0ds_logic.v(1584)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W74iu6 ;  // ../RTL/cortexm0ds_logic.v(360)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W7biu6 ;  // ../RTL/cortexm0ds_logic.v(453)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W7cow6 ;  // ../RTL/cortexm0ds_logic.v(1010)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W7iiu6 ;  // ../RTL/cortexm0ds_logic.v(547)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W7xhu6 ;  // ../RTL/cortexm0ds_logic.v(266)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W8hbx6 ;  // ../RTL/cortexm0ds_logic.v(1710)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W8phu6 ;  // ../RTL/cortexm0ds_logic.v(160)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W9lhu6 ;  // ../RTL/cortexm0ds_logic.v(139)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wa0ju6 ;  // ../RTL/cortexm0ds_logic.v(789)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wahbx6 ;  // ../RTL/cortexm0ds_logic.v(1711)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wamiu6 ;  // ../RTL/cortexm0ds_logic.v(602)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wanow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1158)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wauhu6 ;  // ../RTL/cortexm0ds_logic.v(227)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wb0iu6 ;  // ../RTL/cortexm0ds_logic.v(308)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wbkhu6 ;  // ../RTL/cortexm0ds_logic.v(136)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wc2qw6 ;  // ../RTL/cortexm0ds_logic.v(1621)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wc5ju6_lutinv ;  // ../RTL/cortexm0ds_logic.v(856)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wckiu6 ;  // ../RTL/cortexm0ds_logic.v(576)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Webiu6 ;  // ../RTL/cortexm0ds_logic.v(456)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wfcbx6 ;  // ../RTL/cortexm0ds_logic.v(1702)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wfihu6 ;  // ../RTL/cortexm0ds_logic.v(131)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wfphu6 ;  // ../RTL/cortexm0ds_logic.v(162)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wfspw6 ;  // ../RTL/cortexm0ds_logic.v(1603)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wfviu6 ;  // ../RTL/cortexm0ds_logic.v(724)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wgipw6 ;  // ../RTL/cortexm0ds_logic.v(1585)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wgohu6 ;  // ../RTL/cortexm0ds_logic.v(149)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wgvhu6 ;  // ../RTL/cortexm0ds_logic.v(243)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wh0ju6 ;  // ../RTL/cortexm0ds_logic.v(791)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wh9ow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(973)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Whgow6 ;  // ../RTL/cortexm0ds_logic.v(1067)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Widax6 ;  // ../RTL/cortexm0ds_logic.v(1638)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Withu6 ;  // ../RTL/cortexm0ds_logic.v(217)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wjshu6 ;  // ../RTL/cortexm0ds_logic.v(204)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wjyiu6 ;  // ../RTL/cortexm0ds_logic.v(765)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wk5pw6 ;  // ../RTL/cortexm0ds_logic.v(1402)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wkciu6 ;  // ../RTL/cortexm0ds_logic.v(472)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wkipw6 ;  // ../RTL/cortexm0ds_logic.v(1585)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wkjiu6 ;  // ../RTL/cortexm0ds_logic.v(565)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wlcow6 ;  // ../RTL/cortexm0ds_logic.v(1015)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wlspw6 ;  // ../RTL/cortexm0ds_logic.v(1603)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wlxow6 ;  // ../RTL/cortexm0ds_logic.v(1296)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wmviu6 ;  // ../RTL/cortexm0ds_logic.v(726)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wmzax6 ;  // ../RTL/cortexm0ds_logic.v(1679)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wnohu6 ;  // ../RTL/cortexm0ds_logic.v(152)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wnxax6 ;  // ../RTL/cortexm0ds_logic.v(1675)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Womiu6 ;  // ../RTL/cortexm0ds_logic.v(607)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wouhu6 ;  // ../RTL/cortexm0ds_logic.v(232)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wpthu6 ;  // ../RTL/cortexm0ds_logic.v(219)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wpyax6 ;  // ../RTL/cortexm0ds_logic.v(1677)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wq8ax6 ;  // ../RTL/cortexm0ds_logic.v(1629)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wqdbx6 ;  // ../RTL/cortexm0ds_logic.v(1704)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wqzhu6 ;  // ../RTL/cortexm0ds_logic.v(300)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wr4bx6 ;  // ../RTL/cortexm0ds_logic.v(1688)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wr4ju6_lutinv ;  // ../RTL/cortexm0ds_logic.v(849)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wr6ow6 ;  // ../RTL/cortexm0ds_logic.v(937)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wrcpw6 ;  // ../RTL/cortexm0ds_logic.v(1499)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ws4iu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(368)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wskhu6 ;  // ../RTL/cortexm0ds_logic.v(137)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wsxhu6 ;  // ../RTL/cortexm0ds_logic.v(274)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wt3qw6 ;  // ../RTL/cortexm0ds_logic.v(1624)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wtbow6 ;  // ../RTL/cortexm0ds_logic.v(1005)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wtviu6 ;  // ../RTL/cortexm0ds_logic.v(729)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wtxax6 ;  // ../RTL/cortexm0ds_logic.v(1675)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wu3bx6 ;  // ../RTL/cortexm0ds_logic.v(1686)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wv8pw6 ;  // ../RTL/cortexm0ds_logic.v(1447)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wv9ow6 ;  // ../RTL/cortexm0ds_logic.v(979)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wvgax6 ;  // ../RTL/cortexm0ds_logic.v(1645)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wvuhu6 ;  // ../RTL/cortexm0ds_logic.v(235)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ww6ju6 ;  // ../RTL/cortexm0ds_logic.v(877)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wwiax6 ;  // ../RTL/cortexm0ds_logic.v(1648)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wwihu6 ;  // ../RTL/cortexm0ds_logic.v(132)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wxgbx6 ;  // ../RTL/cortexm0ds_logic.v(1710)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wxjpw6 ;  // ../RTL/cortexm0ds_logic.v(1587)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wxlow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1140)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wxyiu6 ;  // ../RTL/cortexm0ds_logic.v(771)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wxzhu6 ;  // ../RTL/cortexm0ds_logic.v(303)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wy4ju6 ;  // ../RTL/cortexm0ds_logic.v(851)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wydow6 ;  // ../RTL/cortexm0ds_logic.v(1033)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wyhhu6 ;  // ../RTL/cortexm0ds_logic.v(130)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wyiax6 ;  // ../RTL/cortexm0ds_logic.v(1649)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wyqiu6 ;  // ../RTL/cortexm0ds_logic.v(664)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wz4iu6 ;  // ../RTL/cortexm0ds_logic.v(370)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wzpiu6 ;  // ../RTL/cortexm0ds_logic.v(651)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wzqhu6 ;  // ../RTL/cortexm0ds_logic.v(183)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wzxhu6 ;  // ../RTL/cortexm0ds_logic.v(277)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X0fiu6 ;  // ../RTL/cortexm0ds_logic.v(504)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X10iu6 ;  // ../RTL/cortexm0ds_logic.v(304)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X1epw6 ;  // ../RTL/cortexm0ds_logic.v(1516)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X1liu6 ;  // ../RTL/cortexm0ds_logic.v(585)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X2zhu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(291)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X42qw6 ;  // ../RTL/cortexm0ds_logic.v(1621)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X44iu6 ;  // ../RTL/cortexm0ds_logic.v(359)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X4xhu6 ;  // ../RTL/cortexm0ds_logic.v(265)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X53pw6 ;  // ../RTL/cortexm0ds_logic.v(1370)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X5bax6 ;  // ../RTL/cortexm0ds_logic.v(1633)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X5opw6 ;  // ../RTL/cortexm0ds_logic.v(1595)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X5phu6 ;  // ../RTL/cortexm0ds_logic.v(158)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X5upw6 ;  // ../RTL/cortexm0ds_logic.v(1606)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X62pw6 ;  // ../RTL/cortexm0ds_logic.v(1357)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X6jpw6 ;  // ../RTL/cortexm0ds_logic.v(1586)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X6niu6 ;  // ../RTL/cortexm0ds_logic.v(613)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X6vhu6 ;  // ../RTL/cortexm0ds_logic.v(239)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X71pw6 ;  // ../RTL/cortexm0ds_logic.v(1344)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X7abx6 ;  // ../RTL/cortexm0ds_logic.v(1697)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X7miu6 ;  // ../RTL/cortexm0ds_logic.v(600)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X7now6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1157)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X7ypw6 ;  // ../RTL/cortexm0ds_logic.v(1614)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X80iu6 ;  // ../RTL/cortexm0ds_logic.v(307)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X80pw6 ;  // ../RTL/cortexm0ds_logic.v(1331)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X87iu6 ;  // ../RTL/cortexm0ds_logic.v(400)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X87pw6 ;  // ../RTL/cortexm0ds_logic.v(1425)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xa4ju6_lutinv ;  // ../RTL/cortexm0ds_logic.v(842)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xaeax6 ;  // ../RTL/cortexm0ds_logic.v(1640)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xajbx6 ;  // ../RTL/cortexm0ds_logic.v(1714)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xbcow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1011)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xbiiu6 ;  // ../RTL/cortexm0ds_logic.v(548)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xc2ju6_lutinv ;  // ../RTL/cortexm0ds_logic.v(816)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xc9ax6 ;  // ../RTL/cortexm0ds_logic.v(1630)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xcphu6 ;  // ../RTL/cortexm0ds_logic.v(161)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xdcax6 ;  // ../RTL/cortexm0ds_logic.v(1636)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xdebx6 ;  // ../RTL/cortexm0ds_logic.v(1705)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xdspw6 ;  // ../RTL/cortexm0ds_logic.v(1603)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xeuhu6 ;  // ../RTL/cortexm0ds_logic.v(229)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xf7iu6 ;  // ../RTL/cortexm0ds_logic.v(403)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xf8ax6 ;  // ../RTL/cortexm0ds_logic.v(1628)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xfliu6 ;  // ../RTL/cortexm0ds_logic.v(590)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xg6iu6 ;  // ../RTL/cortexm0ds_logic.v(390)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xi4iu6 ;  // ../RTL/cortexm0ds_logic.v(364)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xiaju6 ;  // ../RTL/cortexm0ds_logic.v(925)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xibiu6 ;  // ../RTL/cortexm0ds_logic.v(457)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xiipw6 ;  // ../RTL/cortexm0ds_logic.v(1585)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xipiu6 ;  // ../RTL/cortexm0ds_logic.v(645)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xkohu6 ;  // ../RTL/cortexm0ds_logic.v(151)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xl1iu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(325)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xmthu6 ;  // ../RTL/cortexm0ds_logic.v(218)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xn7ax6 ;  // ../RTL/cortexm0ds_logic.v(1627)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xnbax6 ;  // ../RTL/cortexm0ds_logic.v(1634)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xneow6 ;  // ../RTL/cortexm0ds_logic.v(1042)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xo1bx6 ;  // ../RTL/cortexm0ds_logic.v(1682)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xozax6 ;  // ../RTL/cortexm0ds_logic.v(1679)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xpeax6 ;  // ../RTL/cortexm0ds_logic.v(1640)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xpqow6 ;  // ../RTL/cortexm0ds_logic.v(1204)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xpxax6 ;  // ../RTL/cortexm0ds_logic.v(1675)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xq2bx6 ;  // ../RTL/cortexm0ds_logic.v(1684)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xq3pw6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1378)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xqcax6 ;  // ../RTL/cortexm0ds_logic.v(1637)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xqoiu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(634)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xqpow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1191)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xr9ax6 ;  // ../RTL/cortexm0ds_logic.v(1631)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xrgiu6 ;  // ../RTL/cortexm0ds_logic.v(528)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xrohu6 ;  // ../RTL/cortexm0ds_logic.v(153)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xrxax6 ;  // ../RTL/cortexm0ds_logic.v(1675)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xs1iu6 ;  // ../RTL/cortexm0ds_logic.v(327)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xsmiu6 ;  // ../RTL/cortexm0ds_logic.v(608)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xsuhu6 ;  // ../RTL/cortexm0ds_logic.v(234)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xttow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1245)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xu2qw6 ;  // ../RTL/cortexm0ds_logic.v(1622)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuiax6 ;  // ../RTL/cortexm0ds_logic.v(1648)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuyiu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(769)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 ;  // ../RTL/cortexm0ds_logic.v(301)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xv6ow6 ;  // ../RTL/cortexm0ds_logic.v(938)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xv8bx6 ;  // ../RTL/cortexm0ds_logic.v(1695)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xvqpw6 ;  // ../RTL/cortexm0ds_logic.v(1600)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xwaax6 ;  // ../RTL/cortexm0ds_logic.v(1633)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xwxhu6 ;  // ../RTL/cortexm0ds_logic.v(275)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xx6bx6 ;  // ../RTL/cortexm0ds_logic.v(1691)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxaiu6 ;  // ../RTL/cortexm0ds_logic.v(450)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxqpw6 ;  // ../RTL/cortexm0ds_logic.v(1600)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 ;  // ../RTL/cortexm0ds_logic.v(1608)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xyohu6 ;  // ../RTL/cortexm0ds_logic.v(156)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xz9ow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(980)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xznow6 ;  // ../RTL/cortexm0ds_logic.v(1167)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xzuhu6 ;  // ../RTL/cortexm0ds_logic.v(236)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y0gbx6 ;  // ../RTL/cortexm0ds_logic.v(1708)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y0jiu6 ;  // ../RTL/cortexm0ds_logic.v(558)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y0yhu6 ;  // ../RTL/cortexm0ds_logic.v(277)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y1qow6 ;  // ../RTL/cortexm0ds_logic.v(1195)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y1xhu6 ;  // ../RTL/cortexm0ds_logic.v(264)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y1xow6 ;  // ../RTL/cortexm0ds_logic.v(1288)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y2fax6 ;  // ../RTL/cortexm0ds_logic.v(1641)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y2hiu6 ;  // ../RTL/cortexm0ds_logic.v(532)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y2phu6 ;  // ../RTL/cortexm0ds_logic.v(157)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y32pw6 ;  // ../RTL/cortexm0ds_logic.v(1356)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y3niu6 ;  // ../RTL/cortexm0ds_logic.v(612)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y3vhu6 ;  // ../RTL/cortexm0ds_logic.v(238)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y40ju6 ;  // ../RTL/cortexm0ds_logic.v(787)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y41pw6 ;  // ../RTL/cortexm0ds_logic.v(1343)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y48iu6 ;  // ../RTL/cortexm0ds_logic.v(412)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y4miu6 ;  // ../RTL/cortexm0ds_logic.v(599)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y50iu6 ;  // ../RTL/cortexm0ds_logic.v(306)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y50pw6 ;  // ../RTL/cortexm0ds_logic.v(1330)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y5dax6 ;  // ../RTL/cortexm0ds_logic.v(1637)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y5lhu6 ;  // ../RTL/cortexm0ds_logic.v(138)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y5liu6 ;  // ../RTL/cortexm0ds_logic.v(586)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y72bx6 ;  // ../RTL/cortexm0ds_logic.v(1683)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y7cpw6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1491)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y7jiu6 ;  // ../RTL/cortexm0ds_logic.v(560)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y7opw6 ;  // ../RTL/cortexm0ds_logic.v(1596)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y7yow6 ;  // ../RTL/cortexm0ds_logic.v(1304)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y84iu6 ;  // ../RTL/cortexm0ds_logic.v(360)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y8lpw6 ;  // ../RTL/cortexm0ds_logic.v(1590)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y8xhu6 ;  // ../RTL/cortexm0ds_logic.v(267)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y93bx6 ;  // ../RTL/cortexm0ds_logic.v(1685)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y93iu6 ;  // ../RTL/cortexm0ds_logic.v(347)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y9phu6 ;  // ../RTL/cortexm0ds_logic.v(160)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ya1ju6_lutinv ;  // ../RTL/cortexm0ds_logic.v(802)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yaohu6 ;  // ../RTL/cortexm0ds_logic.v(147)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yavhu6 ;  // ../RTL/cortexm0ds_logic.v(241)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yavow6 ;  // ../RTL/cortexm0ds_logic.v(1265)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yb8iu6 ;  // ../RTL/cortexm0ds_logic.v(415)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ybuhu6 ;  // ../RTL/cortexm0ds_logic.v(228)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yc0pw6 ;  // ../RTL/cortexm0ds_logic.v(1333)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yc7iu6 ;  // ../RTL/cortexm0ds_logic.v(402)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ycliu6 ;  // ../RTL/cortexm0ds_logic.v(589)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yctow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1239)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yd7ow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(945)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydgax6 ;  // ../RTL/cortexm0ds_logic.v(1644)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydkiu6 ;  // ../RTL/cortexm0ds_logic.v(576)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 ;  // ../RTL/cortexm0ds_logic.v(1596)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yecpw6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1494)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yf1qw6 ;  // ../RTL/cortexm0ds_logic.v(1620)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yfcow6 ;  // ../RTL/cortexm0ds_logic.v(1013)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yfiiu6 ;  // ../RTL/cortexm0ds_logic.v(550)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yfqow6 ;  // ../RTL/cortexm0ds_logic.v(1200)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yfxhu6 ;  // ../RTL/cortexm0ds_logic.v(269)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yg3iu6 ;  // ../RTL/cortexm0ds_logic.v(350)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yh8ju6_lutinv ;  // ../RTL/cortexm0ds_logic.v(898)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yhvhu6 ;  // ../RTL/cortexm0ds_logic.v(243)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yi1iu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(324)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yi7ju6_lutinv ;  // ../RTL/cortexm0ds_logic.v(885)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yi8iu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(417)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yj8ow6 ;  // ../RTL/cortexm0ds_logic.v(961)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yjaax6 ;  // ../RTL/cortexm0ds_logic.v(1632)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yjliu6 ;  // ../RTL/cortexm0ds_logic.v(592)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yjtow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1242)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yjupw6 ;  // ../RTL/cortexm0ds_logic.v(1607)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ykkiu6 ;  // ../RTL/cortexm0ds_logic.v(579)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yklpw6 ;  // ../RTL/cortexm0ds_logic.v(1591)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yksow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1229)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yljiu6 ;  // ../RTL/cortexm0ds_logic.v(566)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ym3qw6 ;  // ../RTL/cortexm0ds_logic.v(1624)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ym4iu6 ;  // ../RTL/cortexm0ds_logic.v(365)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ymwiu6 ;  // ../RTL/cortexm0ds_logic.v(740)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ymwpw6 ;  // ../RTL/cortexm0ds_logic.v(1611)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yn3iu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(352)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ynwow6 ;  // ../RTL/cortexm0ds_logic.v(1283)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yo1ju6 ;  // ../RTL/cortexm0ds_logic.v(807)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yogax6 ;  // ../RTL/cortexm0ds_logic.v(1644)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yogiu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(527)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yokhu6 ;  // ../RTL/cortexm0ds_logic.v(137)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yoniu6 ;  // ../RTL/cortexm0ds_logic.v(620)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ypuhu6 ;  // ../RTL/cortexm0ds_logic.v(233)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yqzax6 ;  // ../RTL/cortexm0ds_logic.v(1679)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yqziu6 ;  // ../RTL/cortexm0ds_logic.v(781)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yryax6 ;  // ../RTL/cortexm0ds_logic.v(1677)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ys4ju6 ;  // ../RTL/cortexm0ds_logic.v(849)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ysiax6 ;  // ../RTL/cortexm0ds_logic.v(1648)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ysihu6 ;  // ../RTL/cortexm0ds_logic.v(132)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yt3ju6 ;  // ../RTL/cortexm0ds_logic.v(836)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yt4bx6 ;  // ../RTL/cortexm0ds_logic.v(1688)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yubbx6 ;  // ../RTL/cortexm0ds_logic.v(1700)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yuiow6 ;  // ../RTL/cortexm0ds_logic.v(1099)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yv1ju6 ;  // ../RTL/cortexm0ds_logic.v(810)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yv9pw6 ;  // ../RTL/cortexm0ds_logic.v(1460)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvabx6 ;  // ../RTL/cortexm0ds_logic.v(1699)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvgiu6 ;  // ../RTL/cortexm0ds_logic.v(529)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 ;  // ../RTL/cortexm0ds_logic.v(1587)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yw1iu6 ;  // ../RTL/cortexm0ds_logic.v(329)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yw3bx6 ;  // ../RTL/cortexm0ds_logic.v(1686)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ywuhu6 ;  // ../RTL/cortexm0ds_logic.v(235)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yxdax6 ;  // ../RTL/cortexm0ds_logic.v(1639)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yxrpw6 ;  // ../RTL/cortexm0ds_logic.v(1602)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yy7ow6 ;  // ../RTL/cortexm0ds_logic.v(953)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yybax6 ;  // ../RTL/cortexm0ds_logic.v(1635)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yyzhu6 ;  // ../RTL/cortexm0ds_logic.v(303)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yzlpw6 ;  // ../RTL/cortexm0ds_logic.v(1591)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yzqiu6 ;  // ../RTL/cortexm0ds_logic.v(664)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yzqpw6 ;  // ../RTL/cortexm0ds_logic.v(1601)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yzspw6 ;  // ../RTL/cortexm0ds_logic.v(1604)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z08ju6_lutinv ;  // ../RTL/cortexm0ds_logic.v(892)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z0niu6 ;  // ../RTL/cortexm0ds_logic.v(611)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z0vhu6 ;  // ../RTL/cortexm0ds_logic.v(237)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z18iu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(411)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z18pw6 ;  // ../RTL/cortexm0ds_logic.v(1435)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z1fiu6 ;  // ../RTL/cortexm0ds_logic.v(505)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z1miu6 ;  // ../RTL/cortexm0ds_logic.v(598)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z20iu6 ;  // ../RTL/cortexm0ds_logic.v(304)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z2aax6 ;  // ../RTL/cortexm0ds_logic.v(1631)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z2epw6 ;  // ../RTL/cortexm0ds_logic.v(1516)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z2fow6 ;  // ../RTL/cortexm0ds_logic.v(1048)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z37ow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(941)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z3sow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1222)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z47ax6 ;  // ../RTL/cortexm0ds_logic.v(1626)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z4kow6 ;  // ../RTL/cortexm0ds_logic.v(1116)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z54iu6 ;  // ../RTL/cortexm0ds_logic.v(359)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z67ax6 ;  // ../RTL/cortexm0ds_logic.v(1626)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z6iow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1090)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z6phu6 ;  // ../RTL/cortexm0ds_logic.v(159)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z71bx6 ;  // ../RTL/cortexm0ds_logic.v(1681)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z71ju6 ;  // ../RTL/cortexm0ds_logic.v(801)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z73qw6 ;  // ../RTL/cortexm0ds_logic.v(1623)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z7vhu6 ;  // ../RTL/cortexm0ds_logic.v(239)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z8jpw6 ;  // ../RTL/cortexm0ds_logic.v(1586)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z8uhu6 ;  // ../RTL/cortexm0ds_logic.v(226)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z90iu6 ;  // ../RTL/cortexm0ds_logic.v(307)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z9abx6 ;  // ../RTL/cortexm0ds_logic.v(1698)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z9opw6 ;  // ../RTL/cortexm0ds_logic.v(1596)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Za6pw6 ;  // ../RTL/cortexm0ds_logic.v(1412)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zbjiu6 ;  // ../RTL/cortexm0ds_logic.v(562)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zccow6 ;  // ../RTL/cortexm0ds_logic.v(1012)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zcqhu6 ;  // ../RTL/cortexm0ds_logic.v(174)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zdcbx6 ;  // ../RTL/cortexm0ds_logic.v(1701)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zdiax6 ;  // ../RTL/cortexm0ds_logic.v(1647)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zdphu6 ;  // ../RTL/cortexm0ds_logic.v(161)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zdtpw6 ;  // ../RTL/cortexm0ds_logic.v(1605)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zelhu6 ;  // ../RTL/cortexm0ds_logic.v(139)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zeohu6 ;  // ../RTL/cortexm0ds_logic.v(148)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zf7ju6 ;  // ../RTL/cortexm0ds_logic.v(884)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zf8iu6 ;  // ../RTL/cortexm0ds_logic.v(416)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zfgow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1066)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zfmiu6 ;  // ../RTL/cortexm0ds_logic.v(603)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zg7iu6 ;  // ../RTL/cortexm0ds_logic.v(403)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgbax6 ;  // ../RTL/cortexm0ds_logic.v(1634)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgfax6 ;  // ../RTL/cortexm0ds_logic.v(1642)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgthu6 ;  // ../RTL/cortexm0ds_logic.v(216)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgziu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(778)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zi5iu6 ;  // ../RTL/cortexm0ds_logic.v(377)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zkphu6 ;  // ../RTL/cortexm0ds_logic.v(164)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zl9bx6 ;  // ../RTL/cortexm0ds_logic.v(1696)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zlohu6 ;  // ../RTL/cortexm0ds_logic.v(151)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zm8ax6 ;  // ../RTL/cortexm0ds_logic.v(1629)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zmuhu6 ;  // ../RTL/cortexm0ds_logic.v(232)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zodbx6 ;  // ../RTL/cortexm0ds_logic.v(1704)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zokiu6 ;  // ../RTL/cortexm0ds_logic.v(580)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zp6ow6 ;  // ../RTL/cortexm0ds_logic.v(936)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zpkow6 ;  // ../RTL/cortexm0ds_logic.v(1123)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zqiax6 ;  // ../RTL/cortexm0ds_logic.v(1648)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zqxhu6 ;  // ../RTL/cortexm0ds_logic.v(273)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zrhiu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(541)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zslpw6 ;  // ../RTL/cortexm0ds_logic.v(1591)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsohu6 ;  // ../RTL/cortexm0ds_logic.v(154)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zszax6 ;  // ../RTL/cortexm0ds_logic.v(1679)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zt1iu6 ;  // ../RTL/cortexm0ds_logic.v(328)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztgbx6 ;  // ../RTL/cortexm0ds_logic.v(1710)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztmiu6 ;  // ../RTL/cortexm0ds_logic.v(609)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztuhu6 ;  // ../RTL/cortexm0ds_logic.v(234)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztupw6 ;  // ../RTL/cortexm0ds_logic.v(1607)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zuliu6 ;  // ../RTL/cortexm0ds_logic.v(596)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zvgbx6 ;  // ../RTL/cortexm0ds_logic.v(1710)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zvkiu6 ;  // ../RTL/cortexm0ds_logic.v(583)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zvzhu6 ;  // ../RTL/cortexm0ds_logic.v(302)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zwcpw6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1500)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zwnpw6 ;  // ../RTL/cortexm0ds_logic.v(1595)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zx8ax6 ;  // ../RTL/cortexm0ds_logic.v(1629)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zxxhu6 ;  // ../RTL/cortexm0ds_logic.v(276)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zycbx6 ;  // ../RTL/cortexm0ds_logic.v(1703)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zyoiu6 ;  // ../RTL/cortexm0ds_logic.v(637)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zzniu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(624)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zzohu6 ;  // ../RTL/cortexm0ds_logic.v(156)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add0/c0 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add0/c1 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add0/c2 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add0/c3 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add0/c4 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add0/c5 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add0/c6 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add0/c7 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add0/c8 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add0/c9 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c0 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c1 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c10 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c11 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c12 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c13 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c14 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c15 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c16 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c17 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c18 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c19 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c2 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c20 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c21 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c22 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c23 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c24 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c25 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c26 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c27 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c28 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c29 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c3 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c30 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c4 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c5 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c6 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c7 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c8 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c9 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c0 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c1 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c10 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c11 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c12 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c13 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c14 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c15 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c16 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c17 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c18 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c19 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c2 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c20 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c21 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c22 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c23 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c24 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c25 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c26 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c27 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c28 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c29 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c3 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c4 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c5 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c6 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c7 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c8 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c9 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c0 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c1 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c10 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c11 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c12 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c13 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c14 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c15 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c16 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c17 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c18 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c19 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c2 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c20 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c21 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c22 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c23 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c24 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c25 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c26 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c27 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c28 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c29 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c3 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c30 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c31 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c32 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c4 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c5 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c6 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c7 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c8 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c9 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/eq0/xor_i0[12]_i1[12]_o_lutinv ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/eq0/xor_i0[16]_i1[16]_o_lutinv ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/eq0/xor_i0[1]_i1[1]_o_lutinv ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/eq0/xor_i0[21]_i1[21]_o_lutinv ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/eq0/xor_i0[27]_i1[27]_o_lutinv ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/eq0/xor_i0[3]_i1[3]_o_lutinv ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/eq0/xor_i0[5]_i1[5]_o_lutinv ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/eq1/xor_i0[12]_i1[12]_o_lutinv ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/eq1/xor_i0[15]_i1[15]_o_lutinv ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/eq1/xor_i0[1]_i1[1]_o_lutinv ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/eq1/xor_i0[5]_i1[5]_o_lutinv ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_0 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_1 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_10 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_11 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_12 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_13 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_14 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_15 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_16 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_17 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_18 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_19 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_2 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_20 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_21 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_22 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_23 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_24 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_25 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_26 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_27 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_28 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_29 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_3 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_30 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_31 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_4 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_5 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_6 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_7 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_8 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_9 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_1_0 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_1_1 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_1_10 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_1_11 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_1_12 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_1_13 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_1_2 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_1_3 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_1_4 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_1_5 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_1_6 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_1_7 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_1_8 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_1_9 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_1_0_0 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_1_0_1 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_1_0_10 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_1_0_11 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_1_0_12 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_1_0_13 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_1_0_2 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_1_0_3 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_1_0_4 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_1_0_5 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_1_0_6 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_1_0_7 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_1_0_8 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_1_0_9 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n1465 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n1552 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n265 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n267 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n3436 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n3685 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n382 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n590 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n5992_lutinv ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n5995_lutinv ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n5997_lutinv ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n6006_lutinv ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n6018_lutinv ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n6021_lutinv ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n6023_lutinv ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n689 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n853 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/c0 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/c1 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/c10 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/c11 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/c12 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/c13 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/c14 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/c15 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/c16 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/c17 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/c18 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/c19 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/c2 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/c20 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/c21 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/c22 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/c23 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/c3 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/c4 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/c5 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/c6 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/c7 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/c8 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/c9 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub1/c0 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub1/c1 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub1/c2 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub1/c3 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub1/c4 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub1/c5 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub1/c6 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub1/c7 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub1/c8 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_apsr_o[0] ;  // ../RTL/cortexm0ds_logic.v(70)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_apsr_o[1] ;  // ../RTL/cortexm0ds_logic.v(70)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_apsr_o[2] ;  // ../RTL/cortexm0ds_logic.v(70)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_apsr_o[3] ;  // ../RTL/cortexm0ds_logic.v(70)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_control_o ;  // ../RTL/cortexm0ds_logic.v(117)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[0] ;  // ../RTL/cortexm0ds_logic.v(71)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[1] ;  // ../RTL/cortexm0ds_logic.v(71)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[2] ;  // ../RTL/cortexm0ds_logic.v(71)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[3] ;  // ../RTL/cortexm0ds_logic.v(71)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[4] ;  // ../RTL/cortexm0ds_logic.v(71)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[5] ;  // ../RTL/cortexm0ds_logic.v(71)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[0] ;  // ../RTL/cortexm0ds_logic.v(67)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[10] ;  // ../RTL/cortexm0ds_logic.v(67)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[11] ;  // ../RTL/cortexm0ds_logic.v(67)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[12] ;  // ../RTL/cortexm0ds_logic.v(67)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[13] ;  // ../RTL/cortexm0ds_logic.v(67)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[14] ;  // ../RTL/cortexm0ds_logic.v(67)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[15] ;  // ../RTL/cortexm0ds_logic.v(67)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[16] ;  // ../RTL/cortexm0ds_logic.v(67)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[17] ;  // ../RTL/cortexm0ds_logic.v(67)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[18] ;  // ../RTL/cortexm0ds_logic.v(67)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[19] ;  // ../RTL/cortexm0ds_logic.v(67)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[1] ;  // ../RTL/cortexm0ds_logic.v(67)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[20] ;  // ../RTL/cortexm0ds_logic.v(67)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[21] ;  // ../RTL/cortexm0ds_logic.v(67)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[22] ;  // ../RTL/cortexm0ds_logic.v(67)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[23] ;  // ../RTL/cortexm0ds_logic.v(67)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[24] ;  // ../RTL/cortexm0ds_logic.v(67)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[25] ;  // ../RTL/cortexm0ds_logic.v(67)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[26] ;  // ../RTL/cortexm0ds_logic.v(67)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[27] ;  // ../RTL/cortexm0ds_logic.v(67)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[28] ;  // ../RTL/cortexm0ds_logic.v(67)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[29] ;  // ../RTL/cortexm0ds_logic.v(67)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[2] ;  // ../RTL/cortexm0ds_logic.v(67)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[3] ;  // ../RTL/cortexm0ds_logic.v(67)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[4] ;  // ../RTL/cortexm0ds_logic.v(67)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[5] ;  // ../RTL/cortexm0ds_logic.v(67)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[6] ;  // ../RTL/cortexm0ds_logic.v(67)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[7] ;  // ../RTL/cortexm0ds_logic.v(67)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[8] ;  // ../RTL/cortexm0ds_logic.v(67)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[9] ;  // ../RTL/cortexm0ds_logic.v(67)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[0] ;  // ../RTL/cortexm0ds_logic.v(69)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[10] ;  // ../RTL/cortexm0ds_logic.v(69)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[11] ;  // ../RTL/cortexm0ds_logic.v(69)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[12] ;  // ../RTL/cortexm0ds_logic.v(69)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[13] ;  // ../RTL/cortexm0ds_logic.v(69)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[14] ;  // ../RTL/cortexm0ds_logic.v(69)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[15] ;  // ../RTL/cortexm0ds_logic.v(69)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[16] ;  // ../RTL/cortexm0ds_logic.v(69)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[17] ;  // ../RTL/cortexm0ds_logic.v(69)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[18] ;  // ../RTL/cortexm0ds_logic.v(69)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[19] ;  // ../RTL/cortexm0ds_logic.v(69)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[1] ;  // ../RTL/cortexm0ds_logic.v(69)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[20] ;  // ../RTL/cortexm0ds_logic.v(69)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[21] ;  // ../RTL/cortexm0ds_logic.v(69)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[22] ;  // ../RTL/cortexm0ds_logic.v(69)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[23] ;  // ../RTL/cortexm0ds_logic.v(69)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[24] ;  // ../RTL/cortexm0ds_logic.v(69)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[25] ;  // ../RTL/cortexm0ds_logic.v(69)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[26] ;  // ../RTL/cortexm0ds_logic.v(69)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[27] ;  // ../RTL/cortexm0ds_logic.v(69)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[28] ;  // ../RTL/cortexm0ds_logic.v(69)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[29] ;  // ../RTL/cortexm0ds_logic.v(69)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[2] ;  // ../RTL/cortexm0ds_logic.v(69)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[30] ;  // ../RTL/cortexm0ds_logic.v(69)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[3] ;  // ../RTL/cortexm0ds_logic.v(69)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[4] ;  // ../RTL/cortexm0ds_logic.v(69)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[5] ;  // ../RTL/cortexm0ds_logic.v(69)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[6] ;  // ../RTL/cortexm0ds_logic.v(69)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[7] ;  // ../RTL/cortexm0ds_logic.v(69)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[8] ;  // ../RTL/cortexm0ds_logic.v(69)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[9] ;  // ../RTL/cortexm0ds_logic.v(69)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_primask_o ;  // ../RTL/cortexm0ds_logic.v(118)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[0] ;  // ../RTL/cortexm0ds_logic.v(68)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[10] ;  // ../RTL/cortexm0ds_logic.v(68)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[11] ;  // ../RTL/cortexm0ds_logic.v(68)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[12] ;  // ../RTL/cortexm0ds_logic.v(68)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[13] ;  // ../RTL/cortexm0ds_logic.v(68)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[14] ;  // ../RTL/cortexm0ds_logic.v(68)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[15] ;  // ../RTL/cortexm0ds_logic.v(68)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[16] ;  // ../RTL/cortexm0ds_logic.v(68)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[17] ;  // ../RTL/cortexm0ds_logic.v(68)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[18] ;  // ../RTL/cortexm0ds_logic.v(68)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[19] ;  // ../RTL/cortexm0ds_logic.v(68)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[1] ;  // ../RTL/cortexm0ds_logic.v(68)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[20] ;  // ../RTL/cortexm0ds_logic.v(68)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[21] ;  // ../RTL/cortexm0ds_logic.v(68)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[22] ;  // ../RTL/cortexm0ds_logic.v(68)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[23] ;  // ../RTL/cortexm0ds_logic.v(68)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[24] ;  // ../RTL/cortexm0ds_logic.v(68)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[25] ;  // ../RTL/cortexm0ds_logic.v(68)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[26] ;  // ../RTL/cortexm0ds_logic.v(68)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[27] ;  // ../RTL/cortexm0ds_logic.v(68)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[28] ;  // ../RTL/cortexm0ds_logic.v(68)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[29] ;  // ../RTL/cortexm0ds_logic.v(68)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[2] ;  // ../RTL/cortexm0ds_logic.v(68)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[3] ;  // ../RTL/cortexm0ds_logic.v(68)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[4] ;  // ../RTL/cortexm0ds_logic.v(68)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[5] ;  // ../RTL/cortexm0ds_logic.v(68)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[6] ;  // ../RTL/cortexm0ds_logic.v(68)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[7] ;  // ../RTL/cortexm0ds_logic.v(68)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[8] ;  // ../RTL/cortexm0ds_logic.v(68)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[9] ;  // ../RTL/cortexm0ds_logic.v(68)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[0] ;  // ../RTL/cortexm0ds_logic.v(53)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[10] ;  // ../RTL/cortexm0ds_logic.v(53)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[11] ;  // ../RTL/cortexm0ds_logic.v(53)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[12] ;  // ../RTL/cortexm0ds_logic.v(53)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[13] ;  // ../RTL/cortexm0ds_logic.v(53)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[14] ;  // ../RTL/cortexm0ds_logic.v(53)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[15] ;  // ../RTL/cortexm0ds_logic.v(53)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[16] ;  // ../RTL/cortexm0ds_logic.v(53)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[17] ;  // ../RTL/cortexm0ds_logic.v(53)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[18] ;  // ../RTL/cortexm0ds_logic.v(53)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[19] ;  // ../RTL/cortexm0ds_logic.v(53)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[1] ;  // ../RTL/cortexm0ds_logic.v(53)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[20] ;  // ../RTL/cortexm0ds_logic.v(53)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[21] ;  // ../RTL/cortexm0ds_logic.v(53)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[22] ;  // ../RTL/cortexm0ds_logic.v(53)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[23] ;  // ../RTL/cortexm0ds_logic.v(53)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[24] ;  // ../RTL/cortexm0ds_logic.v(53)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[25] ;  // ../RTL/cortexm0ds_logic.v(53)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[26] ;  // ../RTL/cortexm0ds_logic.v(53)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[27] ;  // ../RTL/cortexm0ds_logic.v(53)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[28] ;  // ../RTL/cortexm0ds_logic.v(53)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[29] ;  // ../RTL/cortexm0ds_logic.v(53)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[2] ;  // ../RTL/cortexm0ds_logic.v(53)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[30] ;  // ../RTL/cortexm0ds_logic.v(53)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[31] ;  // ../RTL/cortexm0ds_logic.v(53)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[3] ;  // ../RTL/cortexm0ds_logic.v(53)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[4] ;  // ../RTL/cortexm0ds_logic.v(53)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[5] ;  // ../RTL/cortexm0ds_logic.v(53)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[6] ;  // ../RTL/cortexm0ds_logic.v(53)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[7] ;  // ../RTL/cortexm0ds_logic.v(53)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[8] ;  // ../RTL/cortexm0ds_logic.v(53)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[9] ;  // ../RTL/cortexm0ds_logic.v(53)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[0] ;  // ../RTL/cortexm0ds_logic.v(63)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[10] ;  // ../RTL/cortexm0ds_logic.v(63)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[11] ;  // ../RTL/cortexm0ds_logic.v(63)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[12] ;  // ../RTL/cortexm0ds_logic.v(63)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[13] ;  // ../RTL/cortexm0ds_logic.v(63)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[14] ;  // ../RTL/cortexm0ds_logic.v(63)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[15] ;  // ../RTL/cortexm0ds_logic.v(63)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[16] ;  // ../RTL/cortexm0ds_logic.v(63)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[17] ;  // ../RTL/cortexm0ds_logic.v(63)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[18] ;  // ../RTL/cortexm0ds_logic.v(63)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[19] ;  // ../RTL/cortexm0ds_logic.v(63)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[1] ;  // ../RTL/cortexm0ds_logic.v(63)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[20] ;  // ../RTL/cortexm0ds_logic.v(63)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[21] ;  // ../RTL/cortexm0ds_logic.v(63)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[22] ;  // ../RTL/cortexm0ds_logic.v(63)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[23] ;  // ../RTL/cortexm0ds_logic.v(63)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[24] ;  // ../RTL/cortexm0ds_logic.v(63)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[25] ;  // ../RTL/cortexm0ds_logic.v(63)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[26] ;  // ../RTL/cortexm0ds_logic.v(63)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[27] ;  // ../RTL/cortexm0ds_logic.v(63)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[28] ;  // ../RTL/cortexm0ds_logic.v(63)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[29] ;  // ../RTL/cortexm0ds_logic.v(63)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[2] ;  // ../RTL/cortexm0ds_logic.v(63)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[30] ;  // ../RTL/cortexm0ds_logic.v(63)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[31] ;  // ../RTL/cortexm0ds_logic.v(63)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[3] ;  // ../RTL/cortexm0ds_logic.v(63)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[4] ;  // ../RTL/cortexm0ds_logic.v(63)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[5] ;  // ../RTL/cortexm0ds_logic.v(63)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[6] ;  // ../RTL/cortexm0ds_logic.v(63)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[7] ;  // ../RTL/cortexm0ds_logic.v(63)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[8] ;  // ../RTL/cortexm0ds_logic.v(63)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[9] ;  // ../RTL/cortexm0ds_logic.v(63)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[0] ;  // ../RTL/cortexm0ds_logic.v(64)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[10] ;  // ../RTL/cortexm0ds_logic.v(64)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[11] ;  // ../RTL/cortexm0ds_logic.v(64)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[12] ;  // ../RTL/cortexm0ds_logic.v(64)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[13] ;  // ../RTL/cortexm0ds_logic.v(64)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[14] ;  // ../RTL/cortexm0ds_logic.v(64)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[15] ;  // ../RTL/cortexm0ds_logic.v(64)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[16] ;  // ../RTL/cortexm0ds_logic.v(64)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[17] ;  // ../RTL/cortexm0ds_logic.v(64)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[18] ;  // ../RTL/cortexm0ds_logic.v(64)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[19] ;  // ../RTL/cortexm0ds_logic.v(64)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[1] ;  // ../RTL/cortexm0ds_logic.v(64)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[20] ;  // ../RTL/cortexm0ds_logic.v(64)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[21] ;  // ../RTL/cortexm0ds_logic.v(64)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[22] ;  // ../RTL/cortexm0ds_logic.v(64)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[23] ;  // ../RTL/cortexm0ds_logic.v(64)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[24] ;  // ../RTL/cortexm0ds_logic.v(64)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[25] ;  // ../RTL/cortexm0ds_logic.v(64)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[26] ;  // ../RTL/cortexm0ds_logic.v(64)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[27] ;  // ../RTL/cortexm0ds_logic.v(64)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[28] ;  // ../RTL/cortexm0ds_logic.v(64)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[29] ;  // ../RTL/cortexm0ds_logic.v(64)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[2] ;  // ../RTL/cortexm0ds_logic.v(64)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[30] ;  // ../RTL/cortexm0ds_logic.v(64)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[31] ;  // ../RTL/cortexm0ds_logic.v(64)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[3] ;  // ../RTL/cortexm0ds_logic.v(64)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[4] ;  // ../RTL/cortexm0ds_logic.v(64)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[5] ;  // ../RTL/cortexm0ds_logic.v(64)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[6] ;  // ../RTL/cortexm0ds_logic.v(64)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[7] ;  // ../RTL/cortexm0ds_logic.v(64)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[8] ;  // ../RTL/cortexm0ds_logic.v(64)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[9] ;  // ../RTL/cortexm0ds_logic.v(64)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[0] ;  // ../RTL/cortexm0ds_logic.v(65)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[10] ;  // ../RTL/cortexm0ds_logic.v(65)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[11] ;  // ../RTL/cortexm0ds_logic.v(65)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[12] ;  // ../RTL/cortexm0ds_logic.v(65)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[13] ;  // ../RTL/cortexm0ds_logic.v(65)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[14] ;  // ../RTL/cortexm0ds_logic.v(65)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[15] ;  // ../RTL/cortexm0ds_logic.v(65)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[16] ;  // ../RTL/cortexm0ds_logic.v(65)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[17] ;  // ../RTL/cortexm0ds_logic.v(65)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[18] ;  // ../RTL/cortexm0ds_logic.v(65)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[19] ;  // ../RTL/cortexm0ds_logic.v(65)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[1] ;  // ../RTL/cortexm0ds_logic.v(65)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[20] ;  // ../RTL/cortexm0ds_logic.v(65)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[21] ;  // ../RTL/cortexm0ds_logic.v(65)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[22] ;  // ../RTL/cortexm0ds_logic.v(65)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[23] ;  // ../RTL/cortexm0ds_logic.v(65)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[24] ;  // ../RTL/cortexm0ds_logic.v(65)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[25] ;  // ../RTL/cortexm0ds_logic.v(65)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[26] ;  // ../RTL/cortexm0ds_logic.v(65)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[27] ;  // ../RTL/cortexm0ds_logic.v(65)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[28] ;  // ../RTL/cortexm0ds_logic.v(65)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[29] ;  // ../RTL/cortexm0ds_logic.v(65)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[2] ;  // ../RTL/cortexm0ds_logic.v(65)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[30] ;  // ../RTL/cortexm0ds_logic.v(65)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[31] ;  // ../RTL/cortexm0ds_logic.v(65)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[3] ;  // ../RTL/cortexm0ds_logic.v(65)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[4] ;  // ../RTL/cortexm0ds_logic.v(65)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[5] ;  // ../RTL/cortexm0ds_logic.v(65)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[6] ;  // ../RTL/cortexm0ds_logic.v(65)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[7] ;  // ../RTL/cortexm0ds_logic.v(65)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[8] ;  // ../RTL/cortexm0ds_logic.v(65)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[9] ;  // ../RTL/cortexm0ds_logic.v(65)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[0] ;  // ../RTL/cortexm0ds_logic.v(66)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[10] ;  // ../RTL/cortexm0ds_logic.v(66)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[11] ;  // ../RTL/cortexm0ds_logic.v(66)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[12] ;  // ../RTL/cortexm0ds_logic.v(66)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[13] ;  // ../RTL/cortexm0ds_logic.v(66)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[14] ;  // ../RTL/cortexm0ds_logic.v(66)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[15] ;  // ../RTL/cortexm0ds_logic.v(66)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[16] ;  // ../RTL/cortexm0ds_logic.v(66)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[17] ;  // ../RTL/cortexm0ds_logic.v(66)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[18] ;  // ../RTL/cortexm0ds_logic.v(66)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[19] ;  // ../RTL/cortexm0ds_logic.v(66)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[1] ;  // ../RTL/cortexm0ds_logic.v(66)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[20] ;  // ../RTL/cortexm0ds_logic.v(66)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[21] ;  // ../RTL/cortexm0ds_logic.v(66)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[22] ;  // ../RTL/cortexm0ds_logic.v(66)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[23] ;  // ../RTL/cortexm0ds_logic.v(66)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[24] ;  // ../RTL/cortexm0ds_logic.v(66)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[25] ;  // ../RTL/cortexm0ds_logic.v(66)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[26] ;  // ../RTL/cortexm0ds_logic.v(66)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[27] ;  // ../RTL/cortexm0ds_logic.v(66)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[28] ;  // ../RTL/cortexm0ds_logic.v(66)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[29] ;  // ../RTL/cortexm0ds_logic.v(66)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[2] ;  // ../RTL/cortexm0ds_logic.v(66)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[30] ;  // ../RTL/cortexm0ds_logic.v(66)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[31] ;  // ../RTL/cortexm0ds_logic.v(66)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[3] ;  // ../RTL/cortexm0ds_logic.v(66)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[4] ;  // ../RTL/cortexm0ds_logic.v(66)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[5] ;  // ../RTL/cortexm0ds_logic.v(66)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[6] ;  // ../RTL/cortexm0ds_logic.v(66)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[7] ;  // ../RTL/cortexm0ds_logic.v(66)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[8] ;  // ../RTL/cortexm0ds_logic.v(66)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[9] ;  // ../RTL/cortexm0ds_logic.v(66)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[0] ;  // ../RTL/cortexm0ds_logic.v(54)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[10] ;  // ../RTL/cortexm0ds_logic.v(54)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[11] ;  // ../RTL/cortexm0ds_logic.v(54)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[12] ;  // ../RTL/cortexm0ds_logic.v(54)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[13] ;  // ../RTL/cortexm0ds_logic.v(54)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[14] ;  // ../RTL/cortexm0ds_logic.v(54)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[15] ;  // ../RTL/cortexm0ds_logic.v(54)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[16] ;  // ../RTL/cortexm0ds_logic.v(54)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[17] ;  // ../RTL/cortexm0ds_logic.v(54)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[18] ;  // ../RTL/cortexm0ds_logic.v(54)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[19] ;  // ../RTL/cortexm0ds_logic.v(54)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[1] ;  // ../RTL/cortexm0ds_logic.v(54)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[20] ;  // ../RTL/cortexm0ds_logic.v(54)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[21] ;  // ../RTL/cortexm0ds_logic.v(54)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[22] ;  // ../RTL/cortexm0ds_logic.v(54)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[23] ;  // ../RTL/cortexm0ds_logic.v(54)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[24] ;  // ../RTL/cortexm0ds_logic.v(54)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[25] ;  // ../RTL/cortexm0ds_logic.v(54)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[26] ;  // ../RTL/cortexm0ds_logic.v(54)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[27] ;  // ../RTL/cortexm0ds_logic.v(54)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[28] ;  // ../RTL/cortexm0ds_logic.v(54)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[29] ;  // ../RTL/cortexm0ds_logic.v(54)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[2] ;  // ../RTL/cortexm0ds_logic.v(54)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[30] ;  // ../RTL/cortexm0ds_logic.v(54)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[31] ;  // ../RTL/cortexm0ds_logic.v(54)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[3] ;  // ../RTL/cortexm0ds_logic.v(54)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[4] ;  // ../RTL/cortexm0ds_logic.v(54)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[5] ;  // ../RTL/cortexm0ds_logic.v(54)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[6] ;  // ../RTL/cortexm0ds_logic.v(54)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[7] ;  // ../RTL/cortexm0ds_logic.v(54)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[8] ;  // ../RTL/cortexm0ds_logic.v(54)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[9] ;  // ../RTL/cortexm0ds_logic.v(54)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[0] ;  // ../RTL/cortexm0ds_logic.v(55)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[10] ;  // ../RTL/cortexm0ds_logic.v(55)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[11] ;  // ../RTL/cortexm0ds_logic.v(55)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[12] ;  // ../RTL/cortexm0ds_logic.v(55)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[13] ;  // ../RTL/cortexm0ds_logic.v(55)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[14] ;  // ../RTL/cortexm0ds_logic.v(55)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[15] ;  // ../RTL/cortexm0ds_logic.v(55)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[16] ;  // ../RTL/cortexm0ds_logic.v(55)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[17] ;  // ../RTL/cortexm0ds_logic.v(55)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[18] ;  // ../RTL/cortexm0ds_logic.v(55)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[19] ;  // ../RTL/cortexm0ds_logic.v(55)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[1] ;  // ../RTL/cortexm0ds_logic.v(55)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[20] ;  // ../RTL/cortexm0ds_logic.v(55)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[21] ;  // ../RTL/cortexm0ds_logic.v(55)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[22] ;  // ../RTL/cortexm0ds_logic.v(55)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[23] ;  // ../RTL/cortexm0ds_logic.v(55)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[24] ;  // ../RTL/cortexm0ds_logic.v(55)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[25] ;  // ../RTL/cortexm0ds_logic.v(55)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[26] ;  // ../RTL/cortexm0ds_logic.v(55)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[27] ;  // ../RTL/cortexm0ds_logic.v(55)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[28] ;  // ../RTL/cortexm0ds_logic.v(55)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[29] ;  // ../RTL/cortexm0ds_logic.v(55)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[2] ;  // ../RTL/cortexm0ds_logic.v(55)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[30] ;  // ../RTL/cortexm0ds_logic.v(55)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[31] ;  // ../RTL/cortexm0ds_logic.v(55)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[3] ;  // ../RTL/cortexm0ds_logic.v(55)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[4] ;  // ../RTL/cortexm0ds_logic.v(55)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[5] ;  // ../RTL/cortexm0ds_logic.v(55)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[6] ;  // ../RTL/cortexm0ds_logic.v(55)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[7] ;  // ../RTL/cortexm0ds_logic.v(55)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[8] ;  // ../RTL/cortexm0ds_logic.v(55)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[9] ;  // ../RTL/cortexm0ds_logic.v(55)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[0] ;  // ../RTL/cortexm0ds_logic.v(56)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[10] ;  // ../RTL/cortexm0ds_logic.v(56)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[11] ;  // ../RTL/cortexm0ds_logic.v(56)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[12] ;  // ../RTL/cortexm0ds_logic.v(56)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[13] ;  // ../RTL/cortexm0ds_logic.v(56)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[14] ;  // ../RTL/cortexm0ds_logic.v(56)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[15] ;  // ../RTL/cortexm0ds_logic.v(56)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[16] ;  // ../RTL/cortexm0ds_logic.v(56)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[17] ;  // ../RTL/cortexm0ds_logic.v(56)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[18] ;  // ../RTL/cortexm0ds_logic.v(56)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[19] ;  // ../RTL/cortexm0ds_logic.v(56)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[1] ;  // ../RTL/cortexm0ds_logic.v(56)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[20] ;  // ../RTL/cortexm0ds_logic.v(56)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[21] ;  // ../RTL/cortexm0ds_logic.v(56)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[22] ;  // ../RTL/cortexm0ds_logic.v(56)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[23] ;  // ../RTL/cortexm0ds_logic.v(56)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[24] ;  // ../RTL/cortexm0ds_logic.v(56)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[25] ;  // ../RTL/cortexm0ds_logic.v(56)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[26] ;  // ../RTL/cortexm0ds_logic.v(56)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[27] ;  // ../RTL/cortexm0ds_logic.v(56)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[28] ;  // ../RTL/cortexm0ds_logic.v(56)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[29] ;  // ../RTL/cortexm0ds_logic.v(56)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[2] ;  // ../RTL/cortexm0ds_logic.v(56)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[30] ;  // ../RTL/cortexm0ds_logic.v(56)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[31] ;  // ../RTL/cortexm0ds_logic.v(56)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[3] ;  // ../RTL/cortexm0ds_logic.v(56)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[4] ;  // ../RTL/cortexm0ds_logic.v(56)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[5] ;  // ../RTL/cortexm0ds_logic.v(56)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[6] ;  // ../RTL/cortexm0ds_logic.v(56)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[7] ;  // ../RTL/cortexm0ds_logic.v(56)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[8] ;  // ../RTL/cortexm0ds_logic.v(56)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[9] ;  // ../RTL/cortexm0ds_logic.v(56)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[0] ;  // ../RTL/cortexm0ds_logic.v(57)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[10] ;  // ../RTL/cortexm0ds_logic.v(57)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[11] ;  // ../RTL/cortexm0ds_logic.v(57)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[12] ;  // ../RTL/cortexm0ds_logic.v(57)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[13] ;  // ../RTL/cortexm0ds_logic.v(57)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[14] ;  // ../RTL/cortexm0ds_logic.v(57)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[15] ;  // ../RTL/cortexm0ds_logic.v(57)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[16] ;  // ../RTL/cortexm0ds_logic.v(57)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[17] ;  // ../RTL/cortexm0ds_logic.v(57)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[18] ;  // ../RTL/cortexm0ds_logic.v(57)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[19] ;  // ../RTL/cortexm0ds_logic.v(57)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[1] ;  // ../RTL/cortexm0ds_logic.v(57)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[20] ;  // ../RTL/cortexm0ds_logic.v(57)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[21] ;  // ../RTL/cortexm0ds_logic.v(57)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[22] ;  // ../RTL/cortexm0ds_logic.v(57)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[23] ;  // ../RTL/cortexm0ds_logic.v(57)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[24] ;  // ../RTL/cortexm0ds_logic.v(57)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[25] ;  // ../RTL/cortexm0ds_logic.v(57)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[26] ;  // ../RTL/cortexm0ds_logic.v(57)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[27] ;  // ../RTL/cortexm0ds_logic.v(57)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[28] ;  // ../RTL/cortexm0ds_logic.v(57)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[29] ;  // ../RTL/cortexm0ds_logic.v(57)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[2] ;  // ../RTL/cortexm0ds_logic.v(57)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[30] ;  // ../RTL/cortexm0ds_logic.v(57)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[31] ;  // ../RTL/cortexm0ds_logic.v(57)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[3] ;  // ../RTL/cortexm0ds_logic.v(57)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[4] ;  // ../RTL/cortexm0ds_logic.v(57)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[5] ;  // ../RTL/cortexm0ds_logic.v(57)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[6] ;  // ../RTL/cortexm0ds_logic.v(57)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[7] ;  // ../RTL/cortexm0ds_logic.v(57)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[8] ;  // ../RTL/cortexm0ds_logic.v(57)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[9] ;  // ../RTL/cortexm0ds_logic.v(57)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[0] ;  // ../RTL/cortexm0ds_logic.v(58)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[10] ;  // ../RTL/cortexm0ds_logic.v(58)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[11] ;  // ../RTL/cortexm0ds_logic.v(58)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[12] ;  // ../RTL/cortexm0ds_logic.v(58)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[13] ;  // ../RTL/cortexm0ds_logic.v(58)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[14] ;  // ../RTL/cortexm0ds_logic.v(58)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[15] ;  // ../RTL/cortexm0ds_logic.v(58)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[16] ;  // ../RTL/cortexm0ds_logic.v(58)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[17] ;  // ../RTL/cortexm0ds_logic.v(58)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[18] ;  // ../RTL/cortexm0ds_logic.v(58)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[19] ;  // ../RTL/cortexm0ds_logic.v(58)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[1] ;  // ../RTL/cortexm0ds_logic.v(58)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[20] ;  // ../RTL/cortexm0ds_logic.v(58)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[21] ;  // ../RTL/cortexm0ds_logic.v(58)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[22] ;  // ../RTL/cortexm0ds_logic.v(58)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[23] ;  // ../RTL/cortexm0ds_logic.v(58)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[24] ;  // ../RTL/cortexm0ds_logic.v(58)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[25] ;  // ../RTL/cortexm0ds_logic.v(58)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[26] ;  // ../RTL/cortexm0ds_logic.v(58)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[27] ;  // ../RTL/cortexm0ds_logic.v(58)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[28] ;  // ../RTL/cortexm0ds_logic.v(58)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[29] ;  // ../RTL/cortexm0ds_logic.v(58)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[2] ;  // ../RTL/cortexm0ds_logic.v(58)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[30] ;  // ../RTL/cortexm0ds_logic.v(58)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[31] ;  // ../RTL/cortexm0ds_logic.v(58)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[3] ;  // ../RTL/cortexm0ds_logic.v(58)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[4] ;  // ../RTL/cortexm0ds_logic.v(58)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[5] ;  // ../RTL/cortexm0ds_logic.v(58)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[6] ;  // ../RTL/cortexm0ds_logic.v(58)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[7] ;  // ../RTL/cortexm0ds_logic.v(58)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[8] ;  // ../RTL/cortexm0ds_logic.v(58)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[9] ;  // ../RTL/cortexm0ds_logic.v(58)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[0] ;  // ../RTL/cortexm0ds_logic.v(59)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[10] ;  // ../RTL/cortexm0ds_logic.v(59)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[11] ;  // ../RTL/cortexm0ds_logic.v(59)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[12] ;  // ../RTL/cortexm0ds_logic.v(59)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[13] ;  // ../RTL/cortexm0ds_logic.v(59)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[14] ;  // ../RTL/cortexm0ds_logic.v(59)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[15] ;  // ../RTL/cortexm0ds_logic.v(59)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[16] ;  // ../RTL/cortexm0ds_logic.v(59)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[17] ;  // ../RTL/cortexm0ds_logic.v(59)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[18] ;  // ../RTL/cortexm0ds_logic.v(59)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[19] ;  // ../RTL/cortexm0ds_logic.v(59)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[1] ;  // ../RTL/cortexm0ds_logic.v(59)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[20] ;  // ../RTL/cortexm0ds_logic.v(59)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[21] ;  // ../RTL/cortexm0ds_logic.v(59)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[22] ;  // ../RTL/cortexm0ds_logic.v(59)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[23] ;  // ../RTL/cortexm0ds_logic.v(59)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[24] ;  // ../RTL/cortexm0ds_logic.v(59)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[25] ;  // ../RTL/cortexm0ds_logic.v(59)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[26] ;  // ../RTL/cortexm0ds_logic.v(59)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[27] ;  // ../RTL/cortexm0ds_logic.v(59)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[28] ;  // ../RTL/cortexm0ds_logic.v(59)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[29] ;  // ../RTL/cortexm0ds_logic.v(59)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[2] ;  // ../RTL/cortexm0ds_logic.v(59)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[30] ;  // ../RTL/cortexm0ds_logic.v(59)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[31] ;  // ../RTL/cortexm0ds_logic.v(59)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[3] ;  // ../RTL/cortexm0ds_logic.v(59)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[4] ;  // ../RTL/cortexm0ds_logic.v(59)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[5] ;  // ../RTL/cortexm0ds_logic.v(59)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[6] ;  // ../RTL/cortexm0ds_logic.v(59)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[7] ;  // ../RTL/cortexm0ds_logic.v(59)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[8] ;  // ../RTL/cortexm0ds_logic.v(59)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[9] ;  // ../RTL/cortexm0ds_logic.v(59)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[0] ;  // ../RTL/cortexm0ds_logic.v(60)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[10] ;  // ../RTL/cortexm0ds_logic.v(60)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[11] ;  // ../RTL/cortexm0ds_logic.v(60)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[12] ;  // ../RTL/cortexm0ds_logic.v(60)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[13] ;  // ../RTL/cortexm0ds_logic.v(60)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[14] ;  // ../RTL/cortexm0ds_logic.v(60)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[15] ;  // ../RTL/cortexm0ds_logic.v(60)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[16] ;  // ../RTL/cortexm0ds_logic.v(60)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[17] ;  // ../RTL/cortexm0ds_logic.v(60)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[18] ;  // ../RTL/cortexm0ds_logic.v(60)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[19] ;  // ../RTL/cortexm0ds_logic.v(60)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[1] ;  // ../RTL/cortexm0ds_logic.v(60)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[20] ;  // ../RTL/cortexm0ds_logic.v(60)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[21] ;  // ../RTL/cortexm0ds_logic.v(60)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[22] ;  // ../RTL/cortexm0ds_logic.v(60)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[23] ;  // ../RTL/cortexm0ds_logic.v(60)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[24] ;  // ../RTL/cortexm0ds_logic.v(60)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[25] ;  // ../RTL/cortexm0ds_logic.v(60)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[26] ;  // ../RTL/cortexm0ds_logic.v(60)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[27] ;  // ../RTL/cortexm0ds_logic.v(60)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[28] ;  // ../RTL/cortexm0ds_logic.v(60)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[29] ;  // ../RTL/cortexm0ds_logic.v(60)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[2] ;  // ../RTL/cortexm0ds_logic.v(60)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[30] ;  // ../RTL/cortexm0ds_logic.v(60)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[31] ;  // ../RTL/cortexm0ds_logic.v(60)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[3] ;  // ../RTL/cortexm0ds_logic.v(60)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[4] ;  // ../RTL/cortexm0ds_logic.v(60)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[5] ;  // ../RTL/cortexm0ds_logic.v(60)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[6] ;  // ../RTL/cortexm0ds_logic.v(60)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[7] ;  // ../RTL/cortexm0ds_logic.v(60)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[8] ;  // ../RTL/cortexm0ds_logic.v(60)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[9] ;  // ../RTL/cortexm0ds_logic.v(60)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[0] ;  // ../RTL/cortexm0ds_logic.v(61)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[10] ;  // ../RTL/cortexm0ds_logic.v(61)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[11] ;  // ../RTL/cortexm0ds_logic.v(61)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[12] ;  // ../RTL/cortexm0ds_logic.v(61)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[13] ;  // ../RTL/cortexm0ds_logic.v(61)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[14] ;  // ../RTL/cortexm0ds_logic.v(61)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[15] ;  // ../RTL/cortexm0ds_logic.v(61)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[16] ;  // ../RTL/cortexm0ds_logic.v(61)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[17] ;  // ../RTL/cortexm0ds_logic.v(61)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[18] ;  // ../RTL/cortexm0ds_logic.v(61)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[19] ;  // ../RTL/cortexm0ds_logic.v(61)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[1] ;  // ../RTL/cortexm0ds_logic.v(61)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[20] ;  // ../RTL/cortexm0ds_logic.v(61)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[21] ;  // ../RTL/cortexm0ds_logic.v(61)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[22] ;  // ../RTL/cortexm0ds_logic.v(61)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[23] ;  // ../RTL/cortexm0ds_logic.v(61)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[24] ;  // ../RTL/cortexm0ds_logic.v(61)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[25] ;  // ../RTL/cortexm0ds_logic.v(61)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[26] ;  // ../RTL/cortexm0ds_logic.v(61)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[27] ;  // ../RTL/cortexm0ds_logic.v(61)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[28] ;  // ../RTL/cortexm0ds_logic.v(61)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[29] ;  // ../RTL/cortexm0ds_logic.v(61)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[2] ;  // ../RTL/cortexm0ds_logic.v(61)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[30] ;  // ../RTL/cortexm0ds_logic.v(61)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[31] ;  // ../RTL/cortexm0ds_logic.v(61)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[3] ;  // ../RTL/cortexm0ds_logic.v(61)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[4] ;  // ../RTL/cortexm0ds_logic.v(61)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[5] ;  // ../RTL/cortexm0ds_logic.v(61)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[6] ;  // ../RTL/cortexm0ds_logic.v(61)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[7] ;  // ../RTL/cortexm0ds_logic.v(61)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[8] ;  // ../RTL/cortexm0ds_logic.v(61)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[9] ;  // ../RTL/cortexm0ds_logic.v(61)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[0] ;  // ../RTL/cortexm0ds_logic.v(62)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[10] ;  // ../RTL/cortexm0ds_logic.v(62)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[11] ;  // ../RTL/cortexm0ds_logic.v(62)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[12] ;  // ../RTL/cortexm0ds_logic.v(62)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[13] ;  // ../RTL/cortexm0ds_logic.v(62)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[14] ;  // ../RTL/cortexm0ds_logic.v(62)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[15] ;  // ../RTL/cortexm0ds_logic.v(62)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[16] ;  // ../RTL/cortexm0ds_logic.v(62)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[17] ;  // ../RTL/cortexm0ds_logic.v(62)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[18] ;  // ../RTL/cortexm0ds_logic.v(62)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[19] ;  // ../RTL/cortexm0ds_logic.v(62)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[1] ;  // ../RTL/cortexm0ds_logic.v(62)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[20] ;  // ../RTL/cortexm0ds_logic.v(62)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[21] ;  // ../RTL/cortexm0ds_logic.v(62)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[22] ;  // ../RTL/cortexm0ds_logic.v(62)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[23] ;  // ../RTL/cortexm0ds_logic.v(62)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[24] ;  // ../RTL/cortexm0ds_logic.v(62)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[25] ;  // ../RTL/cortexm0ds_logic.v(62)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[26] ;  // ../RTL/cortexm0ds_logic.v(62)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[27] ;  // ../RTL/cortexm0ds_logic.v(62)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[28] ;  // ../RTL/cortexm0ds_logic.v(62)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[29] ;  // ../RTL/cortexm0ds_logic.v(62)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[2] ;  // ../RTL/cortexm0ds_logic.v(62)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[30] ;  // ../RTL/cortexm0ds_logic.v(62)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[31] ;  // ../RTL/cortexm0ds_logic.v(62)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[3] ;  // ../RTL/cortexm0ds_logic.v(62)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[4] ;  // ../RTL/cortexm0ds_logic.v(62)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[5] ;  // ../RTL/cortexm0ds_logic.v(62)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[6] ;  // ../RTL/cortexm0ds_logic.v(62)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[7] ;  // ../RTL/cortexm0ds_logic.v(62)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[8] ;  // ../RTL/cortexm0ds_logic.v(62)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[9] ;  // ../RTL/cortexm0ds_logic.v(62)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_tbit_o ;  // ../RTL/cortexm0ds_logic.v(116)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/trans_valid ;  // ../RTL/cmsdk_ahb_cs_rom_table.v(157)
  wire uart0_txd_pad;  // ../RTL/M0demo.v(20)
  wire uart0_txen_pad;  // ../RTL/M0demo.v(21)

  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("INV"))
    _al_u100 (
    .do({open_n1,open_n2,open_n3,\u_cmsdk_mcu/p0_out [10]}),
    .ts(\u_cmsdk_mcu/p0_outen [10]),
    .opad(P0[10]));  // ../RTL/cmsdk_mcu_pin_mux.v(136)
  AL_MAP_LUT4 #(
    .EQN("(~D*~(~A*~(C*B)))"),
    .INIT(16'h00ea))
    _al_u1000 (
    .a(_al_u996_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_raw_intstatus [2]),
    .c(_al_u999_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[5] ),
    .o(_al_u1000_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~A*~(C*B))"),
    .INIT(16'h1500))
    _al_u1001 (
    .a(_al_u1000_o),
    .b(_al_u945_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/int_gpio_ls_sync [2]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[6] ),
    .o(_al_u1001_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h3ff5))
    _al_u1002 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inten [2]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_int_polarity [2]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] ),
    .o(_al_u1002_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf35f))
    _al_u1003 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_intmask [2]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inttype_level [2]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] ),
    .o(_al_u1003_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u1004 (
    .a(_al_u566_o),
    .b(_al_u1002_o),
    .c(_al_u1003_o),
    .o(_al_u1004_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'h00ac))
    _al_u1005 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_ddr [2]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_dr [2]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/sel0_b2/B1_0 ));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(~C*~B*A))"),
    .INIT(16'h00fd))
    _al_u1006 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/sel0_b2/B1_0 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[4] ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[5] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[6] ),
    .o(_al_u1006_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u1007 (
    .a(_al_u1001_o),
    .b(_al_u1004_o),
    .c(_al_u1006_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n81 [2]));
  AL_MAP_LUT4 #(
    .EQN("(A*(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C))"),
    .INIT(16'ha808))
    _al_u1008 (
    .a(_al_u470_o),
    .b(b_pad_gpio_porta_pad[1]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_ddr [1]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_dr [1]),
    .o(_al_u1008_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*(A*~(D)*~(C)+A*D*~(C)+~(A)*D*C+A*D*C))"),
    .INIT(16'h3202))
    _al_u1009 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/gpio_ext_porta_int [1]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_ddr [1]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_ls_sync ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/int_pre_in [1]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/ls_int_in [1]));
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("INV"))
    _al_u101 (
    .do({open_n17,open_n18,open_n19,\u_cmsdk_mcu/p0_out [9]}),
    .ts(\u_cmsdk_mcu/p0_outen [9]),
    .opad(P0[9]));  // ../RTL/cmsdk_mcu_pin_mux.v(135)
  AL_MAP_LUT4 #(
    .EQN("(~(~C*B)*~(~D*A))"),
    .INIT(16'hf351))
    _al_u1010 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_intmask [1]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inttype_level [1]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/gpio_intr_ed_pm [1]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] ),
    .o(_al_u1010_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    _al_u1011 (
    .a(_al_u1010_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inten [1]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[4] ),
    .o(_al_u1011_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(C*~(~D*~B)))"),
    .INIT(16'h0515))
    _al_u1012 (
    .a(_al_u1008_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/ls_int_in [1]),
    .c(_al_u1011_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inttype_level [1]),
    .o(_al_u1012_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B*A))"),
    .INIT(8'h70))
    _al_u1013 (
    .a(_al_u945_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/int_gpio_ls_sync [1]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[6] ),
    .o(_al_u1013_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'h00ac))
    _al_u1014 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_ddr [1]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_dr [1]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/sel0_b1/B1_0 ));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(~C*~B*A))"),
    .INIT(16'h00fd))
    _al_u1015 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/sel0_b1/B1_0 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[4] ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[5] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[6] ),
    .o(_al_u1015_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h3ff5))
    _al_u1016 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inten [1]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_int_polarity [1]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] ),
    .o(_al_u1016_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf35f))
    _al_u1017 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_intmask [1]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inttype_level [1]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] ),
    .o(_al_u1017_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*~(D*C)))"),
    .INIT(16'ha222))
    _al_u1018 (
    .a(_al_u1015_o),
    .b(_al_u566_o),
    .c(_al_u1016_o),
    .d(_al_u1017_o),
    .o(_al_u1018_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(B*~(~D*~A)))"),
    .INIT(16'h0307))
    _al_u1019 (
    .a(_al_u1012_o),
    .b(_al_u1013_o),
    .c(_al_u1018_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[5] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n81 [1]));
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("INV"))
    _al_u102 (
    .do({open_n33,open_n34,open_n35,\u_cmsdk_mcu/p0_out [8]}),
    .ts(\u_cmsdk_mcu/p0_outen [8]),
    .opad(P0[8]));  // ../RTL/cmsdk_mcu_pin_mux.v(134)
  AL_MAP_LUT4 #(
    .EQN("(A*(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C))"),
    .INIT(16'ha808))
    _al_u1020 (
    .a(_al_u470_o),
    .b(b_pad_gpio_porta_pad[0]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_ddr [0]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_dr [0]),
    .o(_al_u1020_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*(A*~(D)*~(C)+A*D*~(C)+~(A)*D*C+A*D*C))"),
    .INIT(16'h3202))
    _al_u1021 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/gpio_ext_porta_int [0]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_ddr [0]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_ls_sync ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/int_pre_in [0]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/ls_int_in [0]));
  AL_MAP_LUT4 #(
    .EQN("(B*(A*~(D)*~(C)+A*D*~(C)+~(A)*D*C+A*D*C))"),
    .INIT(16'hc808))
    _al_u1022 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/ls_int_in [0]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inten [0]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inttype_level [0]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/gpio_intr_ed_pm [0]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_raw_intstatus [0]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~(~B*A))"),
    .INIT(16'h000d))
    _al_u1023 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_intmask [0]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[4] ),
    .o(_al_u1023_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(~A*~(C*B)))"),
    .INIT(16'h00ea))
    _al_u1024 (
    .a(_al_u1020_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_raw_intstatus [0]),
    .c(_al_u1023_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[5] ),
    .o(_al_u1024_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~A*~(C*B))"),
    .INIT(16'h1500))
    _al_u1025 (
    .a(_al_u1024_o),
    .b(_al_u945_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_ls_sync ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[6] ),
    .o(_al_u1025_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h3ff5))
    _al_u1026 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inten [0]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_int_polarity [0]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] ),
    .o(_al_u1026_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf35f))
    _al_u1027 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_intmask [0]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inttype_level [0]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] ),
    .o(_al_u1027_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u1028 (
    .a(_al_u566_o),
    .b(_al_u1026_o),
    .c(_al_u1027_o),
    .o(_al_u1028_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'h00ac))
    _al_u1029 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_ddr [0]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_dr [0]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/sel0_b0/B1_0 ));
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("INV"))
    _al_u103 (
    .do({open_n49,open_n50,open_n51,\u_cmsdk_mcu/p0_out [7]}),
    .ts(\u_cmsdk_mcu/p0_outen [7]),
    .opad(P0[7]));  // ../RTL/cmsdk_mcu_pin_mux.v(133)
  AL_MAP_LUT4 #(
    .EQN("(~D*~(~C*~B*A))"),
    .INIT(16'h00fd))
    _al_u1030 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/sel0_b0/B1_0 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[4] ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[5] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[6] ),
    .o(_al_u1030_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u1031 (
    .a(_al_u1025_o),
    .b(_al_u1028_o),
    .c(_al_u1030_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n81 [0]));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*B*~A)"),
    .INIT(16'h0400))
    _al_u1032 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_state_inc ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/lt2/o_1_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_state [2]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_state [3]),
    .o(_al_u1032_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    _al_u1033 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/lt2/o_1_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_state [2]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_state [3]),
    .o(_al_u1033_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u1034 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_state [0]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_state [1]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_state [2]),
    .o(_al_u1034_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*~B))"),
    .INIT(8'h54))
    _al_u1035 (
    .a(_al_u1033_o),
    .b(_al_u1034_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_state [3]),
    .o(_al_u1035_o));
  AL_MAP_LUT3 #(
    .EQN("~(~A*~(C*~B))"),
    .INIT(8'hba))
    _al_u1036 (
    .a(_al_u1032_o),
    .b(_al_u1035_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n67 [3]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_tx_state [3]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u1037 (
    .a(_al_u1035_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n67 [2]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_tx_state [2]));
  AL_MAP_LUT4 #(
    .EQN("~(~C*~A*~(D*~B))"),
    .INIT(16'hfbfa))
    _al_u1038 (
    .a(_al_u1032_o),
    .b(_al_u1035_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n63 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n67 [1]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_tx_state [1]));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(A*~(D*B)))"),
    .INIT(16'h0d05))
    _al_u1039 (
    .a(_al_u1034_o),
    .b(uart0_txen_pad),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_state [3]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_buf_full ),
    .o(_al_u1039_o));
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("INV"))
    _al_u104 (
    .do({open_n65,open_n66,open_n67,\u_cmsdk_mcu/p0_out [6]}),
    .ts(\u_cmsdk_mcu/p0_outen [6]),
    .opad(P0[6]));  // ../RTL/cmsdk_mcu_pin_mux.v(132)
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*~(B)*C*D)"),
    .INIT(16'h113f))
    _al_u1040 (
    .a(_al_u1033_o),
    .b(_al_u1039_o),
    .c(_al_u1034_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n67 [0]),
    .o(_al_u1040_o));
  AL_MAP_LUT2 #(
    .EQN("~(B*~A)"),
    .INIT(4'hb))
    _al_u1041 (
    .a(_al_u1032_o),
    .b(_al_u1040_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_tx_state [0]));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*A)"),
    .INIT(16'h0080))
    _al_u1042 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n6 ),
    .b(_al_u472_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n43 ));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u1043 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n6 ),
    .b(_al_u692_o),
    .c(_al_u571_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n55 ));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*A)"),
    .INIT(16'h0080))
    _al_u1044 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n6 ),
    .b(_al_u692_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n52 ));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*~A))"),
    .INIT(8'hdc))
    _al_u1045 (
    .a(_al_u650_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rxbuf_sample ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_buf_full ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_rx_buf_full ));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*~A)"),
    .INIT(8'h04))
    _al_u1046 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V3xhu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_tbit_o ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sz3qw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vobiu6_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("~(~B*A)"),
    .INIT(4'hd))
    _al_u1047 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vobiu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pexpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wz4iu6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u1048 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] ),
    .o(_al_u1048_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u1049 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n6 ),
    .b(_al_u692_o),
    .c(_al_u1048_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n58 ));
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("INV"))
    _al_u105 (
    .do({open_n81,open_n82,open_n83,\u_cmsdk_mcu/p0_out [5]}),
    .ts(\u_cmsdk_mcu/p0_outen [5]),
    .opad(P0[5]));  // ../RTL/cmsdk_mcu_pin_mux.v(131)
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*~A)"),
    .INIT(16'h0040))
    _al_u1050 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Htmpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iixpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vhspw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vmipw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xpqow6 ));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*A)"),
    .INIT(16'h0080))
    _al_u1051 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Htmpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iixpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vhspw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vmipw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eqqow6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1052 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xpqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eqqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[0] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[0] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X53pw6 ));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u1053 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Htmpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iixpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vhspw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vmipw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cpqow6 ));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*A)"),
    .INIT(16'h0002))
    _al_u1054 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Htmpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iixpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vhspw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vmipw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mnqow6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1055 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cpqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mnqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[0] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[0] ),
    .o(_al_u1055_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*~B*A)"),
    .INIT(16'h0020))
    _al_u1056 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Htmpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iixpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vhspw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vmipw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fnqow6 ));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*~B*~A)"),
    .INIT(16'h0010))
    _al_u1057 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Htmpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iixpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vhspw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vmipw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Voqow6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1058 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fnqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Voqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[0] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[0] ),
    .o(_al_u1058_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    _al_u1059 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Htmpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iixpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vhspw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vmipw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kmqow6 ));
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("INV"))
    _al_u106 (
    .do({open_n97,open_n98,open_n99,\u_cmsdk_mcu/p0_out [4]}),
    .ts(\u_cmsdk_mcu/p0_outen [4]),
    .opad(P0[4]));  // ../RTL/cmsdk_mcu_pin_mux.v(130)
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*~A)"),
    .INIT(16'h0004))
    _al_u1060 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Htmpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iixpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vhspw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vmipw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dmqow6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1061 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kmqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dmqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[0] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[0] ),
    .o(_al_u1061_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u1062 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X53pw6 ),
    .b(_al_u1055_o),
    .c(_al_u1058_o),
    .d(_al_u1061_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N30iu6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u1063 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N30iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgfpw6 [0]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1064 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cpqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Voqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[2] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[2] ),
    .o(_al_u1064_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1065 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eqqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kmqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[2] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[2] ),
    .o(_al_u1065_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1066 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xpqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dmqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[2] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[2] ),
    .o(_al_u1066_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1067 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mnqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fnqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[2] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[2] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bu2pw6 ));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u1068 (
    .a(_al_u1064_o),
    .b(_al_u1065_o),
    .c(_al_u1066_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bu2pw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pxzhu6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u1069 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pxzhu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgfpw6 [2]));
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("INV"))
    _al_u107 (
    .do({open_n113,open_n114,open_n115,\u_cmsdk_mcu/p0_out [3]}),
    .ts(\u_cmsdk_mcu/p0_outen [3]),
    .opad(P0[3]));  // ../RTL/cmsdk_mcu_pin_mux.v(129)
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1070 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Voqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kmqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[10] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[10] ),
    .o(_al_u1070_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1071 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fnqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dmqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[10] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[10] ),
    .o(_al_u1071_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1072 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xpqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eqqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[10] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[10] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ll2pw6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1073 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cpqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mnqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[10] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[10] ),
    .o(_al_u1073_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u1074 (
    .a(_al_u1070_o),
    .b(_al_u1071_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ll2pw6 ),
    .d(_al_u1073_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G30iu6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u1075 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G30iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgfpw6 [10]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1076 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xpqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dmqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[3] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[3] ),
    .o(_al_u1076_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1077 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eqqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mnqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[3] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[3] ),
    .o(_al_u1077_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1078 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fnqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kmqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[3] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[3] ),
    .o(_al_u1078_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1079 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cpqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Voqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[3] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[3] ),
    .o(_al_u1079_o));
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("INV"))
    _al_u108 (
    .do({open_n129,open_n130,open_n131,\u_cmsdk_mcu/p0_out [2]}),
    .ts(\u_cmsdk_mcu/p0_outen [2]),
    .opad(P0[2]));  // ../RTL/cmsdk_mcu_pin_mux.v(128)
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u1080 (
    .a(_al_u1076_o),
    .b(_al_u1077_o),
    .c(_al_u1078_o),
    .d(_al_u1079_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uwzhu6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u1081 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uwzhu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgfpw6 [3]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1082 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Voqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kmqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[11] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[11] ),
    .o(_al_u1082_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1083 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fnqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dmqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[11] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[11] ),
    .o(_al_u1083_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1084 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xpqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eqqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[11] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[11] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y32pw6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1085 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cpqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mnqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[11] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[11] ),
    .o(_al_u1085_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u1086 (
    .a(_al_u1082_o),
    .b(_al_u1083_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y32pw6 ),
    .d(_al_u1085_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z20iu6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u1087 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z20iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgfpw6 [11]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1088 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xpqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dmqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[4] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[4] ),
    .o(_al_u1088_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1089 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eqqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mnqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[4] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[4] ),
    .o(_al_u1089_o));
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("INV"))
    _al_u109 (
    .do({open_n145,open_n146,open_n147,\u_cmsdk_mcu/p0_out [1]}),
    .ts(\u_cmsdk_mcu/p0_outen [1]),
    .opad(P0[1]));  // ../RTL/cmsdk_mcu_pin_mux.v(127)
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1090 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fnqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kmqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[4] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[4] ),
    .o(_al_u1090_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1091 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cpqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Voqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[4] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[4] ),
    .o(_al_u1091_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u1092 (
    .a(_al_u1088_o),
    .b(_al_u1089_o),
    .c(_al_u1090_o),
    .d(_al_u1091_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nwzhu6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u1093 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nwzhu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgfpw6 [4]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1094 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xpqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dmqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[12] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[12] ),
    .o(_al_u1094_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1095 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eqqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mnqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[12] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[12] ),
    .o(_al_u1095_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1096 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fnqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kmqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[12] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[12] ),
    .o(_al_u1096_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1097 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cpqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Voqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[12] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[12] ),
    .o(_al_u1097_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u1098 (
    .a(_al_u1094_o),
    .b(_al_u1095_o),
    .c(_al_u1096_o),
    .d(_al_u1097_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S20iu6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u1099 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S20iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgfpw6 [12]));
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("INV"))
    _al_u110 (
    .do({open_n161,open_n162,open_n163,\u_cmsdk_mcu/p0_out [0]}),
    .ts(\u_cmsdk_mcu/p0_outen [0]),
    .opad(P0[0]));  // ../RTL/cmsdk_mcu_pin_mux.v(126)
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1100 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cpqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Voqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[5] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[5] ),
    .o(_al_u1100_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1101 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mnqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kmqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[5] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[5] ),
    .o(_al_u1101_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1102 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xpqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dmqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[5] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[5] ),
    .o(_al_u1102_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1103 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eqqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fnqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[5] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[5] ),
    .o(_al_u1103_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u1104 (
    .a(_al_u1100_o),
    .b(_al_u1101_o),
    .c(_al_u1102_o),
    .d(_al_u1103_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gwzhu6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u1105 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gwzhu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgfpw6 [5]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1106 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Voqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dmqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[13] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[13] ),
    .o(_al_u1106_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1107 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fnqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kmqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[13] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[13] ),
    .o(_al_u1107_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1108 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xpqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eqqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[13] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[13] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y41pw6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1109 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cpqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mnqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[13] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[13] ),
    .o(_al_u1109_o));
  EG_PHY_PAD #(
    //.LOCATION("A8"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u111 (
    .ipad(SWCLKTCK),
    .di(SWCLKTCK_pad));  // ../RTL/M0demo.v(15)
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u1110 (
    .a(_al_u1106_o),
    .b(_al_u1107_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y41pw6 ),
    .d(_al_u1109_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L20iu6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u1111 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L20iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgfpw6 [13]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1112 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xpqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dmqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[6] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[6] ),
    .o(_al_u1112_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1113 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eqqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mnqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[6] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[6] ),
    .o(_al_u1113_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1114 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fnqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kmqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[6] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[6] ),
    .o(_al_u1114_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1115 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cpqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Voqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[6] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[6] ),
    .o(_al_u1115_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u1116 (
    .a(_al_u1112_o),
    .b(_al_u1113_o),
    .c(_al_u1114_o),
    .d(_al_u1115_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zvzhu6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u1117 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zvzhu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgfpw6 [6]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1118 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fnqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Voqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[14] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[14] ),
    .o(_al_u1118_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1119 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mnqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kmqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[14] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[14] ),
    .o(_al_u1119_o));
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u112 (
    .ipad(TDI));  // ../RTL/M0demo.v(12)
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1120 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xpqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eqqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[14] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[14] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ln0pw6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1121 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cpqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dmqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[14] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[14] ),
    .o(_al_u1121_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u1122 (
    .a(_al_u1118_o),
    .b(_al_u1119_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ln0pw6 ),
    .d(_al_u1121_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E20iu6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u1123 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E20iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgfpw6 [14]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1124 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cpqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kmqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[7] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[7] ),
    .o(_al_u1124_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1125 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eqqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Voqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[7] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[7] ),
    .o(_al_u1125_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1126 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xpqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dmqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[7] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[7] ),
    .o(_al_u1126_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1127 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mnqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fnqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[7] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[7] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yc0pw6 ));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u1128 (
    .a(_al_u1124_o),
    .b(_al_u1125_o),
    .c(_al_u1126_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yc0pw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Svzhu6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u1129 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Svzhu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgfpw6 [7]));
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("INV"))
    _al_u113 (
    .do({open_n212,open_n213,open_n214,1'b0}),
    .ts(1'b1),
    .opad(TDO));  // ../RTL/cmsdk_mcu_pin_mux.v(211)
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1130 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xpqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eqqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[15] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[15] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y50pw6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1131 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mnqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dmqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[15] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[15] ),
    .o(_al_u1131_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1132 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cpqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fnqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[15] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[15] ),
    .o(_al_u1132_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1133 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Voqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kmqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[15] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[15] ),
    .o(_al_u1133_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u1134 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y50pw6 ),
    .b(_al_u1131_o),
    .c(_al_u1132_o),
    .d(_al_u1133_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X10iu6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u1135 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X10iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgfpw6 [15]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1136 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xpqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eqqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[17] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[17] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uwzow6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1137 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mnqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kmqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[17] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[17] ),
    .o(_al_u1137_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1138 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cpqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fnqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[17] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[17] ),
    .o(_al_u1138_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1139 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Voqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dmqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[17] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[17] ),
    .o(_al_u1139_o));
  EG_PHY_PAD #(
    //.LOCATION("K14"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u114 (
    .ipad(XTAL1),
    .di(XTAL1_pad));  // ../RTL/M0demo.v(5)
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u1140 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uwzow6 ),
    .b(_al_u1137_o),
    .c(_al_u1138_o),
    .d(_al_u1139_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J10iu6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u1141 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J10iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgfpw6 [17]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1142 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cpqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Voqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[1] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[1] ),
    .o(_al_u1142_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1143 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fnqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kmqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[1] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[1] ),
    .o(_al_u1143_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1144 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xpqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dmqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[1] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[1] ),
    .o(_al_u1144_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1145 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eqqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mnqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[1] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[1] ),
    .o(_al_u1145_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u1146 (
    .a(_al_u1142_o),
    .b(_al_u1143_o),
    .c(_al_u1144_o),
    .d(_al_u1145_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O00iu6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u1147 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O00iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgfpw6 [1]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1148 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xpqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fnqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[18] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[18] ),
    .o(_al_u1148_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1149 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eqqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dmqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[18] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[18] ),
    .o(_al_u1149_o));
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u115 (
    .do({open_n245,open_n246,open_n247,XTAL2_pad}),
    .opad(XTAL2));  // ../RTL/M0demo.v(6)
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1150 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cpqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kmqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[18] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[18] ),
    .o(_al_u1150_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1151 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mnqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Voqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[18] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[18] ),
    .o(_al_u1151_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u1152 (
    .a(_al_u1148_o),
    .b(_al_u1149_o),
    .c(_al_u1150_o),
    .d(_al_u1151_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C10iu6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u1153 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C10iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgfpw6 [18]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1154 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cpqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mnqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[19] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[19] ),
    .o(_al_u1154_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1155 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Voqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kmqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[19] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[19] ),
    .o(_al_u1155_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1156 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xpqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fnqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[19] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[19] ),
    .o(_al_u1156_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1157 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eqqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dmqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[19] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[19] ),
    .o(_al_u1157_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u1158 (
    .a(_al_u1154_o),
    .b(_al_u1155_o),
    .c(_al_u1156_o),
    .d(_al_u1157_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V00iu6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u1159 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V00iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgfpw6 [19]));
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("BI"),
    .TSMUX("INV"))
    _al_u116 (
    .do({open_n262,open_n263,open_n264,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_dr [7]}),
    .ts(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_ddr [7]),
    .di(b_pad_gpio_porta_pad[7]),
    .bpad(b_pad_gpio_porta[7]));  // ../RTL/gpio.v(182)
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1160 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xpqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fnqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[20] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[20] ),
    .o(_al_u1160_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1161 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eqqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dmqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[20] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[20] ),
    .o(_al_u1161_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1162 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Voqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kmqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[20] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[20] ),
    .o(_al_u1162_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1163 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cpqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mnqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[20] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[20] ),
    .o(_al_u1163_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u1164 (
    .a(_al_u1160_o),
    .b(_al_u1161_o),
    .c(_al_u1162_o),
    .d(_al_u1163_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H00iu6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u1165 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H00iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgfpw6 [20]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1166 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mnqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Voqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[21] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[21] ),
    .o(_al_u1166_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1167 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cpqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dmqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[21] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[21] ),
    .o(_al_u1167_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1168 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xpqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fnqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[21] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[21] ),
    .o(_al_u1168_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1169 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eqqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kmqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[21] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[21] ),
    .o(_al_u1169_o));
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("BI"),
    .TSMUX("INV"))
    _al_u117 (
    .do({open_n277,open_n278,open_n279,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_dr [6]}),
    .ts(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_ddr [6]),
    .di(b_pad_gpio_porta_pad[6]),
    .bpad(b_pad_gpio_porta[6]));  // ../RTL/gpio.v(178)
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u1170 (
    .a(_al_u1166_o),
    .b(_al_u1167_o),
    .c(_al_u1168_o),
    .d(_al_u1169_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A00iu6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u1171 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A00iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgfpw6 [21]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1172 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xpqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eqqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[22] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[22] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pdyow6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1173 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mnqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dmqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[22] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[22] ),
    .o(_al_u1173_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1174 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cpqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kmqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[22] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[22] ),
    .o(_al_u1174_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1175 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fnqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Voqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[22] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[22] ),
    .o(_al_u1175_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u1176 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pdyow6 ),
    .b(_al_u1173_o),
    .c(_al_u1174_o),
    .d(_al_u1175_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tzzhu6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u1177 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tzzhu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgfpw6 [22]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1178 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Voqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kmqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[23] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[23] ),
    .o(_al_u1178_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1179 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fnqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dmqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[23] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[23] ),
    .o(_al_u1179_o));
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("BI"),
    .TSMUX("INV"))
    _al_u118 (
    .do({open_n292,open_n293,open_n294,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_dr [5]}),
    .ts(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_ddr [5]),
    .di(b_pad_gpio_porta_pad[5]),
    .bpad(b_pad_gpio_porta[5]));  // ../RTL/gpio.v(174)
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1180 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xpqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eqqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[23] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[23] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E4yow6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1181 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cpqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mnqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[23] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[23] ),
    .o(_al_u1181_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u1182 (
    .a(_al_u1178_o),
    .b(_al_u1179_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E4yow6 ),
    .d(_al_u1181_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mzzhu6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u1183 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mzzhu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgfpw6 [23]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1184 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xpqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fnqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[24] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[24] ),
    .o(_al_u1184_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1185 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eqqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dmqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[24] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[24] ),
    .o(_al_u1185_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1186 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Voqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kmqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[24] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[24] ),
    .o(_al_u1186_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1187 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cpqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mnqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[24] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[24] ),
    .o(_al_u1187_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u1188 (
    .a(_al_u1184_o),
    .b(_al_u1185_o),
    .c(_al_u1186_o),
    .d(_al_u1187_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fzzhu6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u1189 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fzzhu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgfpw6 [24]));
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("BI"),
    .TSMUX("INV"))
    _al_u119 (
    .do({open_n307,open_n308,open_n309,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_dr [4]}),
    .ts(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_ddr [4]),
    .di(b_pad_gpio_porta_pad[4]),
    .bpad(b_pad_gpio_porta[4]));  // ../RTL/gpio.v(170)
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1190 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fnqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Voqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[8] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[8] ),
    .o(_al_u1190_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1191 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kmqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dmqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[8] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[8] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nkxow6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1192 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xpqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eqqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[8] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[8] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wlxow6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1193 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cpqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mnqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[8] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[8] ),
    .o(_al_u1193_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u1194 (
    .a(_al_u1190_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nkxow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wlxow6 ),
    .d(_al_u1193_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lvzhu6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u1195 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lvzhu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgfpw6 [8]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1196 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mnqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Voqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[25] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[25] ),
    .o(_al_u1196_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1197 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eqqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cpqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[25] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[25] ),
    .o(_al_u1197_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1198 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xpqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fnqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[25] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[25] ),
    .o(_al_u1198_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1199 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kmqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dmqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[25] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[25] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oaxow6 ));
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("BI"),
    .TSMUX("INV"))
    _al_u120 (
    .do({open_n322,open_n323,open_n324,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_dr [3]}),
    .ts(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_ddr [3]),
    .di(b_pad_gpio_porta_pad[3]),
    .bpad(b_pad_gpio_porta[3]));  // ../RTL/gpio.v(166)
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u1200 (
    .a(_al_u1196_o),
    .b(_al_u1197_o),
    .c(_al_u1198_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oaxow6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yyzhu6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u1201 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yyzhu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgfpw6 [25]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1202 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cpqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kmqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[9] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[9] ),
    .o(_al_u1202_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1203 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eqqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Voqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[9] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[9] ),
    .o(_al_u1203_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1204 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xpqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dmqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[9] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[9] ),
    .o(_al_u1204_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1205 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mnqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fnqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[9] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[9] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y1xow6 ));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u1206 (
    .a(_al_u1202_o),
    .b(_al_u1203_o),
    .c(_al_u1204_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y1xow6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Evzhu6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u1207 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Evzhu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgfpw6 [9]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1208 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xpqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fnqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[26] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[26] ),
    .o(_al_u1208_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1209 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eqqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kmqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[26] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[26] ),
    .o(_al_u1209_o));
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("BI"),
    .TSMUX("INV"))
    _al_u121 (
    .do({open_n337,open_n338,open_n339,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_dr [2]}),
    .ts(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_ddr [2]),
    .di(b_pad_gpio_porta_pad[2]),
    .bpad(b_pad_gpio_porta[2]));  // ../RTL/gpio.v(162)
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1210 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Voqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dmqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[26] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[26] ),
    .o(_al_u1210_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1211 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cpqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mnqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[26] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[26] ),
    .o(_al_u1211_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u1212 (
    .a(_al_u1208_o),
    .b(_al_u1209_o),
    .c(_al_u1210_o),
    .d(_al_u1211_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ryzhu6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u1213 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ryzhu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgfpw6 [26]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1214 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xpqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eqqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[27] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[27] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jjwow6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1215 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mnqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kmqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[27] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[27] ),
    .o(_al_u1215_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1216 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cpqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fnqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[27] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[27] ),
    .o(_al_u1216_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1217 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Voqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dmqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[27] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[27] ),
    .o(_al_u1217_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u1218 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jjwow6 ),
    .b(_al_u1215_o),
    .c(_al_u1216_o),
    .d(_al_u1217_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kyzhu6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u1219 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kyzhu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgfpw6 [27]));
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("BI"),
    .TSMUX("INV"))
    _al_u122 (
    .do({open_n352,open_n353,open_n354,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_dr [1]}),
    .ts(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_ddr [1]),
    .di(b_pad_gpio_porta_pad[1]),
    .bpad(b_pad_gpio_porta[1]));  // ../RTL/gpio.v(158)
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1220 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kmqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dmqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[28] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[28] ),
    .o(_al_u1220_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1221 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cpqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fnqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[28] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[28] ),
    .o(_al_u1221_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1222 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xpqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eqqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[28] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[28] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R9wow6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1223 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mnqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Voqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[28] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[28] ),
    .o(_al_u1223_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u1224 (
    .a(_al_u1220_o),
    .b(_al_u1221_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R9wow6 ),
    .d(_al_u1223_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dyzhu6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u1225 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dyzhu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgfpw6 [28]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1226 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cpqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Voqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[30] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[30] ),
    .o(_al_u1226_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1227 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fnqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kmqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[30] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[30] ),
    .o(_al_u1227_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1228 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xpqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dmqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[30] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[30] ),
    .o(_al_u1228_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1229 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eqqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mnqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[30] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[30] ),
    .o(_al_u1229_o));
  EG_PHY_PAD #(
    //.LOCATION("N3"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("BI"),
    .TSMUX("INV"))
    _al_u123 (
    .do({open_n367,open_n368,open_n369,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_dr [0]}),
    .ts(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_ddr [0]),
    .di(b_pad_gpio_porta_pad[0]),
    .bpad(b_pad_gpio_porta[0]));  // ../RTL/gpio.v(154)
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u1230 (
    .a(_al_u1226_o),
    .b(_al_u1227_o),
    .c(_al_u1228_o),
    .d(_al_u1229_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ixzhu6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u1231 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ixzhu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgfpw6 [30]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1232 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cpqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mnqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[31] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[31] ),
    .o(_al_u1232_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1233 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Voqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kmqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[31] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[31] ),
    .o(_al_u1233_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1234 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xpqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fnqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[31] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[31] ),
    .o(_al_u1234_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1235 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eqqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dmqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[31] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[31] ),
    .o(_al_u1235_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u1236 (
    .a(_al_u1232_o),
    .b(_al_u1233_o),
    .c(_al_u1234_o),
    .d(_al_u1235_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bxzhu6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u1237 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bxzhu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgfpw6 [31]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1238 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xpqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fnqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[29] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[29] ),
    .o(_al_u1238_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1239 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eqqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dmqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[29] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[29] ),
    .o(_al_u1239_o));
  EG_PHY_PAD #(
    //.LOCATION("R5"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u124 (
    .ipad(nTRST));  // ../RTL/M0demo.v(11)
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1240 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cpqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kmqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[29] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[29] ),
    .o(_al_u1240_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1241 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mnqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Voqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[29] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[29] ),
    .o(_al_u1241_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u1242 (
    .a(_al_u1238_o),
    .b(_al_u1239_o),
    .c(_al_u1240_o),
    .d(_al_u1241_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wxzhu6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u1243 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wxzhu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgfpw6 [29]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1244 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xpqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fnqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[16] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[16] ),
    .o(_al_u1244_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1245 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eqqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dmqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[16] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[16] ),
    .o(_al_u1245_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1246 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cpqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kmqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[16] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[16] ),
    .o(_al_u1246_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1247 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mnqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Voqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[16] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[16] ),
    .o(_al_u1247_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u1248 (
    .a(_al_u1244_o),
    .b(_al_u1245_o),
    .c(_al_u1246_o),
    .d(_al_u1247_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q10iu6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u1249 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q10iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgfpw6 [16]));
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u125 (
    .do({open_n400,open_n401,open_n402,uart0_txd_pad}),
    .opad(uart0_txd));  // ../RTL/M0demo.v(20)
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u1250 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kalpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yklpw6 ),
    .o(_al_u1250_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u1251 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bclpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sdlpw6 ),
    .o(_al_u1251_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u1252 (
    .a(_al_u1250_o),
    .b(_al_u1251_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jflpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Agyhu6 ));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u1253 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Agyhu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U5yhu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rilpw6 ),
    .o(_al_u1253_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u1254 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Golpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vplpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pyyhu6_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u1255 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pyyhu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zslpw6 ),
    .o(_al_u1255_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u1256 (
    .a(_al_u1253_o),
    .b(_al_u1255_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Krlpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U73iu6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u1257 (
    .a(_al_u903_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ),
    .o(_al_u1257_o));
  AL_MAP_LUT4 #(
    .EQN("~(~C*~(D*~(B*A)))"),
    .INIT(16'hf7f0))
    _al_u1258 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Scbiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O34iu6 ),
    .c(_al_u1257_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xnbax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X6vhu6 ));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    _al_u1259 (
    .a(_al_u650_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rxbuf_sample ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_buf_full ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_overrun ));
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u126 (
    .do({open_n417,open_n418,open_n419,uart0_txen_pad}),
    .opad(uart0_txen));  // ../RTL/M0demo.v(21)
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u1260 (
    .a(_al_u473_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/write_enable ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n9_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    _al_u1261 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_overrun ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n9_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n17 ));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u1262 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n6 ),
    .b(_al_u945_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[6] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n61 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u1263 (
    .a(_al_u681_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qe8iu6_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u1264 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 ),
    .o(_al_u1264_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*B*A))"),
    .INIT(16'h070f))
    _al_u1265 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qe8iu6_lutinv ),
    .b(_al_u606_o),
    .c(_al_u1264_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lv7ow6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u1266 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 ),
    .o(_al_u1266_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u1267 (
    .a(_al_u1266_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Us2ju6 ));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u1268 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Us2ju6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 ),
    .o(_al_u1268_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u1269 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vygax6 ),
    .o(_al_u1269_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(~C*~(D*B)))"),
    .INIT(16'ha8a0))
    _al_u1270 (
    .a(_al_u1268_o),
    .b(_al_u1269_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 ),
    .o(_al_u1270_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u1271 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 ),
    .o(_al_u1271_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u1272 (
    .a(_al_u1269_o),
    .b(_al_u1271_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kwuow6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(C*B*~(~D*~A))"),
    .INIT(16'hc080))
    _al_u1273 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kwuow6_lutinv ),
    .b(_al_u604_o),
    .c(_al_u609_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 ),
    .o(_al_u1273_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u1274 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Llaow6_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u1275 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Llaow6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vygax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Apaiu6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*A)"),
    .INIT(16'h0002))
    _al_u1276 (
    .a(_al_u681_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 ),
    .o(_al_u1276_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(~D*C*A))"),
    .INIT(16'h3313))
    _al_u1277 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Apaiu6_lutinv ),
    .b(_al_u1276_o),
    .c(_al_u682_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yavow6 ));
  AL_MAP_LUT4 #(
    .EQN("~(D*~C*~B*A)"),
    .INIT(16'hfdff))
    _al_u1278 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lv7ow6 ),
    .b(_al_u1270_o),
    .c(_al_u1273_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yavow6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fnpiu6 ));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u1279 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/write_enable00 ),
    .b(_al_u637_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_buf_full ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_overrun ));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    _al_u1280 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_overrun ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n9_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n20 ));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u1281 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/haddr_reg [7]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/haddr_reg [8]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/haddr_reg [9]),
    .o(_al_u1281_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*A)"),
    .INIT(16'h0002))
    _al_u1282 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [8]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/haddr_reg [4]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/haddr_reg [5]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/haddr_reg [6]),
    .o(_al_u1282_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    _al_u1283 (
    .a(_al_u1281_o),
    .b(_al_u1282_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/haddr_reg [2]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/haddr_reg [3]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n37 [1]));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u1284 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n37 [1]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/haddr_reg [0]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/haddr_reg [1]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n37 [14]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1285 (
    .a(\u_cmsdk_mcu/sram_hrdata [30]),
    .b(\u_cmsdk_mcu/flash_hrdata [30]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [0]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [1]),
    .o(_al_u1285_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u1286 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n37 [14]),
    .b(_al_u1285_o),
    .o(_al_u1286_o));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(B*~A))"),
    .INIT(8'hf4))
    _al_u1287 (
    .a(_al_u1286_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vobiu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pexpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rw8iu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u1288 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ujxax6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uojbx6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V0jpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vrtpw6 ),
    .o(_al_u1288_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*A)"),
    .INIT(16'h0002))
    _al_u1289 (
    .a(_al_u1288_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wlspw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y7opw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z8jpw6 ),
    .o(_al_u1289_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u1290 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rv7ax6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ss0qw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T9kpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tjkpw6 ),
    .o(_al_u1290_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u1291 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oarpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0ibx6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pt7ax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rfxax6 ),
    .o(_al_u1291_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u1292 (
    .a(_al_u1289_o),
    .b(_al_u1290_o),
    .c(_al_u1291_o),
    .o(_al_u1292_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u1293 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kzabx6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N0xpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nbxax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nr7ax6 ),
    .o(_al_u1293_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u1294 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Amupw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Coupw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F9gbx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Johbx6 ),
    .o(_al_u1294_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u1295 (
    .a(_al_u1292_o),
    .b(_al_u1293_o),
    .c(_al_u1294_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Azeiu6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u1296 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 ),
    .o(_al_u1296_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u1297 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D6kiu6_lutinv ),
    .b(_al_u1296_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 ),
    .o(_al_u1297_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u1298 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mfjiu6 ));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u1299 (
    .a(_al_u1297_o),
    .b(_al_u604_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mfjiu6 ),
    .o(_al_u1299_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u1300 (
    .a(_al_u1299_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zszax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ozeiu6 ));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u1301 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Azeiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ozeiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N8rpw6 ),
    .o(_al_u1301_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u1302 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vowiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cvciu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ur4iu6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u1303 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jcpow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vynow6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvgiu6 ));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B*A))"),
    .INIT(8'h70))
    _al_u1304 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvgiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C1wpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T2kbx6 ),
    .o(_al_u1304_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~D*C*A))"),
    .INIT(16'hcc4c))
    _al_u1305 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ur4iu6 ),
    .b(_al_u1304_o),
    .c(_al_u405_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C1wpw6 ),
    .o(_al_u1305_o));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    _al_u1306 (
    .a(_al_u1301_o),
    .b(_al_u1305_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kjthu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~B*(~A*~(C)*~(D)+~A*C*~(D)+~(~A)*C*D+~A*C*D))"),
    .INIT(16'h3011))
    _al_u1307 (
    .a(_al_u530_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahlpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Krlpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pmlpw6 ),
    .o(_al_u1307_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u1308 (
    .a(_al_u1250_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jflpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sdlpw6 ),
    .o(_al_u1308_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*~A))"),
    .INIT(8'h32))
    _al_u1309 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bclpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jflpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Krlpw6 ),
    .o(_al_u1309_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u1310 (
    .a(_al_u1250_o),
    .b(_al_u1309_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sdlpw6 ),
    .o(_al_u1310_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~A*~(~D*C))"),
    .INIT(16'h1101))
    _al_u1311 (
    .a(_al_u1308_o),
    .b(_al_u1310_o),
    .c(_al_u1251_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jflpw6 ),
    .o(_al_u1311_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u1312 (
    .a(_al_u529_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kalpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yklpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rsyhu6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(A*~(~D*~(~C*B)))"),
    .INIT(16'haa08))
    _al_u1313 (
    .a(_al_u1307_o),
    .b(_al_u1311_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rsyhu6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pmlpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tw2iu6 ));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u1314 (
    .a(_al_u702_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dzvpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6kax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ds4ju6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*B*A)"),
    .INIT(16'h0800))
    _al_u1315 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dzvpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6kax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Shopw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wxjpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jo4ju6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1316 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ds4ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jo4ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[0] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[0] ),
    .o(_al_u1316_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    _al_u1317 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dzvpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6kax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Shopw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wxjpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gq4ju6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*~A)"),
    .INIT(16'h0004))
    _al_u1318 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dzvpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6kax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Shopw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wxjpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rs4ju6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1319 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gq4ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rs4ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[0] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[0] ),
    .o(_al_u1319_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*~A)"),
    .INIT(16'h4000))
    _al_u1320 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dzvpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6kax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Shopw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wxjpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nq4ju6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*B*~A)"),
    .INIT(16'h0400))
    _al_u1321 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dzvpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6kax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Shopw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wxjpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wr4ju6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1322 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nq4ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wr4ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[0] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[0] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ls9pw6 ));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u1323 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dc0iu6 ),
    .b(_al_u1316_o),
    .c(_al_u1319_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ls9pw6 ),
    .o(_al_u1323_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u1324 (
    .a(_al_u1266_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xc2ju6_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u1325 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Frziu6_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u1326 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Frziu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yqziu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1327 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xc2ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yqziu6 ),
    .c(_al_u914_o),
    .d(_al_u1271_o),
    .o(_al_u1327_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u1328 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dzvpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6kax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Shopw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wxjpw6 ),
    .o(_al_u1328_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u1329 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 ),
    .o(_al_u1329_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u1330 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Btoiu6_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u1331 (
    .a(_al_u1328_o),
    .b(_al_u1329_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Btoiu6_lutinv ),
    .o(_al_u1331_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*A)"),
    .INIT(16'h0002))
    _al_u1332 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Frziu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ),
    .o(_al_u1332_o));
  AL_MAP_LUT4 #(
    .EQN("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'ha088))
    _al_u1333 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ),
    .o(_al_u1333_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    _al_u1334 (
    .a(_al_u1327_o),
    .b(_al_u1331_o),
    .c(_al_u1332_o),
    .d(_al_u1333_o),
    .o(_al_u1334_o));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    _al_u1335 (
    .a(_al_u1323_o),
    .b(_al_u1334_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I1lpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Go0iu6_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u1336 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 ),
    .o(_al_u1336_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    _al_u1337 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xc2ju6_lutinv ),
    .b(_al_u1336_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vgjpw6 ),
    .o(_al_u1337_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u1338 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T23ju6_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*B))"),
    .INIT(8'ha2))
    _al_u1339 (
    .a(_al_u1337_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T23ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 ),
    .o(_al_u1339_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u1340 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ldoiu6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u1341 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ldoiu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ),
    .o(_al_u1341_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u1342 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 ),
    .o(_al_u1342_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(~D*~(~C*~B)))"),
    .INIT(16'h5501))
    _al_u1343 (
    .a(_al_u1341_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Np7ow6_lutinv ),
    .c(_al_u1342_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 ),
    .o(_al_u1343_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u1344 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 ),
    .o(_al_u1344_o));
  AL_MAP_LUT4 #(
    .EQN("~(A*~((C*B))*~(D)+A*(C*B)*~(D)+~(A)*(C*B)*D+A*(C*B)*D)"),
    .INIT(16'h3f55))
    _al_u1345 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Us2ju6 ),
    .b(_al_u696_o),
    .c(_al_u1344_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 ),
    .o(_al_u1345_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u1346 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 ),
    .o(_al_u1346_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(~A*~(~D*C)))"),
    .INIT(16'h2232))
    _al_u1347 (
    .a(_al_u1346_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ),
    .o(_al_u1347_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*A)"),
    .INIT(16'h0080))
    _al_u1348 (
    .a(_al_u1339_o),
    .b(_al_u1343_o),
    .c(_al_u1345_o),
    .d(_al_u1347_o),
    .o(_al_u1348_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u1349 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Go0iu6_lutinv ),
    .b(_al_u1348_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [0]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1350 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ds4ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nq4ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[1] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[1] ),
    .o(_al_u1350_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1351 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rs4ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wr4ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[1] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[1] ),
    .o(_al_u1351_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1352 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jo4ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gq4ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[1] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[1] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X87pw6 ));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u1353 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E90iu6 ),
    .b(_al_u1350_o),
    .c(_al_u1351_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X87pw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V77pw6 ));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    _al_u1354 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V77pw6 ),
    .b(_al_u1334_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nu5bx6 ),
    .o(_al_u1354_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u1355 (
    .a(_al_u1354_o),
    .b(_al_u1348_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [1]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u1356 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ia8iu6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u1357 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P14qw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Skjax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9ypw6 ),
    .o(_al_u1357_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u1358 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ia8iu6_lutinv ),
    .b(_al_u1357_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Srbow6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u1359 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 ),
    .o(_al_u1359_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u1360 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Srbow6 ),
    .b(_al_u1359_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wkipw6 ),
    .o(_al_u1360_o));
  AL_MAP_LUT4 #(
    .EQN("(A*(~(B)*C*~(D)+B*~(C)*D+B*C*D))"),
    .INIT(16'h8820))
    _al_u1361 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Llaow6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P14qw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9ypw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fb1ju6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u1362 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Skjax6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9ypw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ya1ju6_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u1363 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ya1ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P14qw6 ),
    .o(_al_u1363_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u1364 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Llaow6_lutinv ),
    .b(_al_u1363_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 ),
    .o(_al_u1364_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u1365 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fb1ju6 ),
    .b(_al_u1364_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rwjax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B91ju6 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*~A))"),
    .INIT(8'h8c))
    _al_u1366 (
    .a(_al_u1360_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B91ju6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S7mpw6 ),
    .o(_al_u1366_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u1367 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Skjax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9ypw6 ),
    .o(_al_u1367_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*~A)"),
    .INIT(8'h04))
    _al_u1368 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv ),
    .b(_al_u1367_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hs8ow6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u1369 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rwjax6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qxoiu6 ));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(B*A))"),
    .INIT(8'h07))
    _al_u1370 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qxoiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 ),
    .o(_al_u1370_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u1371 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S7mpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wfspw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R9aiu6 ));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u1372 (
    .a(_al_u1359_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R9aiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wkipw6 ),
    .o(_al_u1372_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~B*~(~C*A))"),
    .INIT(16'h0031))
    _al_u1373 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Srbow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hs8ow6 ),
    .c(_al_u1370_o),
    .d(_al_u1372_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mb1ju6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u1374 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Skjax6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9ypw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujiu6 ));
  AL_MAP_LUT4 #(
    .EQN("(C*~(~B*~(D*A)))"),
    .INIT(16'he0c0))
    _al_u1375 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P14qw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rwjax6 ),
    .o(_al_u1375_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(A*~(D)*~(C)+A*D*~(C)+~(A)*D*C+A*D*C))"),
    .INIT(16'h0131))
    _al_u1376 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P14qw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Skjax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9ypw6 ),
    .o(_al_u1376_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*~B))"),
    .INIT(8'ha8))
    _al_u1377 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Llaow6_lutinv ),
    .b(_al_u1375_o),
    .c(_al_u1376_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P91ju6 ));
  AL_MAP_LUT4 #(
    .EQN("~(B*A*~(D*C))"),
    .INIT(16'hf777))
    _al_u1378 (
    .a(_al_u1366_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mb1ju6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P91ju6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jgxpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z71ju6 ));
  AL_MAP_LUT4 #(
    .EQN("(~B*A*~(D*C))"),
    .INIT(16'h0222))
    _al_u1379 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F85iu6 ),
    .b(_al_u908_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K75iu6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jgxpw6 ),
    .o(_al_u1379_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1380 (
    .a(_al_u912_o),
    .b(_al_u696_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lgkax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N4kax6 ),
    .o(_al_u1380_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u1381 (
    .a(_al_u1379_o),
    .b(_al_u1380_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A95iu6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S7mpw6 ),
    .o(_al_u1381_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u1382 (
    .a(_al_u916_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iekax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lgkax6 ),
    .o(_al_u1382_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u1383 (
    .a(_al_u916_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fkrpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ubypw6 ),
    .o(_al_u1383_o));
  AL_MAP_LUT4 #(
    .EQN("~(A*~(B*~(~D*~C)))"),
    .INIT(16'hddd5))
    _al_u1384 (
    .a(_al_u1381_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L45iu6_lutinv ),
    .c(_al_u1382_o),
    .d(_al_u1383_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H25iu6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u1385 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gr2qw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Isjpw6 ),
    .o(_al_u1385_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u1386 (
    .a(_al_u1299_o),
    .b(_al_u1385_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/HALTED ));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u1387 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vuciu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cvciu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dg2qw6 ),
    .o(_al_u1387_o));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*C)*~(B*A))"),
    .INIT(16'hf888))
    _al_u1388 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/HALTED ),
    .b(_al_u1387_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M8fax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Czuhu6 ));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*B*A)"),
    .INIT(16'h0800))
    _al_u1389 (
    .a(_al_u702_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dzvpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jrypw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6kax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lp4ju6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1390 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nq4ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wr4ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[12] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[12] ),
    .o(_al_u1390_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u1391 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lp4ju6 ),
    .b(_al_u1390_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[10] ),
    .o(_al_u1391_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u1392 (
    .a(_al_u702_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dzvpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jrypw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6kax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ep4ju6 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u1393 (
    .a(_al_u1391_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ep4ju6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[10] ),
    .o(_al_u1393_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1394 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ds4ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jo4ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[12] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[12] ),
    .o(_al_u1394_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1395 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gq4ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rs4ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[12] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[12] ),
    .o(_al_u1395_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u1396 (
    .a(_al_u1393_o),
    .b(_al_u1394_o),
    .c(_al_u1395_o),
    .o(_al_u1396_o));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~((B*A))*~(C)+~D*(B*A)*~(C)+~(~D)*(B*A)*C+~D*(B*A)*C)"),
    .INIT(16'h7f70))
    _al_u1397 (
    .a(_al_u1396_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ib0iu6 ),
    .c(_al_u1334_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dm6bx6 ),
    .o(_al_u1397_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u1398 (
    .a(_al_u1397_o),
    .b(_al_u1348_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [12]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1399 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rs4ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wr4ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[13] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[13] ),
    .o(_al_u1399_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u1400 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lp4ju6 ),
    .b(_al_u1399_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[11] ),
    .o(_al_u1400_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u1401 (
    .a(_al_u1400_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ep4ju6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[11] ),
    .o(_al_u1401_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1402 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ds4ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nq4ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[13] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[13] ),
    .o(_al_u1402_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1403 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jo4ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gq4ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[13] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[13] ),
    .o(_al_u1403_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u1404 (
    .a(_al_u1401_o),
    .b(_al_u1402_o),
    .c(_al_u1403_o),
    .o(_al_u1404_o));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~((B*A))*~(C)+~D*(B*A)*~(C)+~(~D)*(B*A)*C+~D*(B*A)*C)"),
    .INIT(16'h7f70))
    _al_u1405 (
    .a(_al_u1404_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bb0iu6 ),
    .c(_al_u1334_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xpxax6 ),
    .o(_al_u1405_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u1406 (
    .a(_al_u1405_o),
    .b(_al_u1348_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [13]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1407 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jo4ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wr4ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[14] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[14] ),
    .o(_al_u1407_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u1408 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lp4ju6 ),
    .b(_al_u1407_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[12] ),
    .o(_al_u1408_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u1409 (
    .a(_al_u1408_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ep4ju6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[12] ),
    .o(_al_u1409_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1410 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ds4ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gq4ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[14] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[14] ),
    .o(_al_u1410_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1411 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rs4ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nq4ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[14] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[14] ),
    .o(_al_u1411_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u1412 (
    .a(_al_u1409_o),
    .b(_al_u1410_o),
    .c(_al_u1411_o),
    .o(_al_u1412_o));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~((B*A))*~(C)+~D*(B*A)*~(C)+~(~D)*(B*A)*C+~D*(B*A)*C)"),
    .INIT(16'h7f70))
    _al_u1413 (
    .a(_al_u1412_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ua0iu6 ),
    .c(_al_u1334_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sb8ax6 ),
    .o(_al_u1413_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u1414 (
    .a(_al_u1413_o),
    .b(_al_u1348_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [14]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1415 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rs4ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wr4ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[15] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[15] ),
    .o(_al_u1415_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u1416 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ep4ju6 ),
    .b(_al_u1415_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[13] ),
    .o(_al_u1416_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u1417 (
    .a(_al_u1416_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lp4ju6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[13] ),
    .o(_al_u1417_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1418 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ds4ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nq4ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[15] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[15] ),
    .o(_al_u1418_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1419 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jo4ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gq4ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[15] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[15] ),
    .o(_al_u1419_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u1420 (
    .a(_al_u1417_o),
    .b(_al_u1418_o),
    .c(_al_u1419_o),
    .o(_al_u1420_o));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~((B*A))*~(C)+~D*(B*A)*~(C)+~(~D)*(B*A)*C+~D*(B*A)*C)"),
    .INIT(16'h7f70))
    _al_u1421 (
    .a(_al_u1420_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Na0iu6 ),
    .c(_al_u1334_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z47ax6 ),
    .o(_al_u1421_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u1422 (
    .a(_al_u1421_o),
    .b(_al_u1348_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [15]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1423 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jo4ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rs4ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[16] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[16] ),
    .o(_al_u1423_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u1424 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lp4ju6 ),
    .b(_al_u1423_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[14] ),
    .o(_al_u1424_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u1425 (
    .a(_al_u1424_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ep4ju6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[14] ),
    .o(_al_u1425_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1426 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ds4ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nq4ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[16] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[16] ),
    .o(_al_u1426_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1427 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gq4ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wr4ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[16] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[16] ),
    .o(_al_u1427_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u1428 (
    .a(_al_u1425_o),
    .b(_al_u1426_o),
    .c(_al_u1427_o),
    .o(_al_u1428_o));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~((B*A))*~(C)+~D*(B*A)*~(C)+~(~D)*(B*A)*C+~D*(B*A)*C)"),
    .INIT(16'h7f70))
    _al_u1429 (
    .a(_al_u1428_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ga0iu6 ),
    .c(_al_u1334_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Chwpw6 ),
    .o(_al_u1429_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u1430 (
    .a(_al_u1429_o),
    .b(_al_u1348_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [16]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1431 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rs4ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nq4ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[17] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[17] ),
    .o(_al_u1431_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u1432 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ep4ju6 ),
    .b(_al_u1431_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[15] ),
    .o(_al_u1432_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u1433 (
    .a(_al_u1432_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lp4ju6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[15] ),
    .o(_al_u1433_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1434 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ds4ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wr4ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[17] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[17] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z18pw6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1435 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jo4ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gq4ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[17] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[17] ),
    .o(_al_u1435_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u1436 (
    .a(_al_u1433_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z18pw6 ),
    .c(_al_u1435_o),
    .o(_al_u1436_o));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~((B*A))*~(C)+~D*(B*A)*~(C)+~(~D)*(B*A)*C+~D*(B*A)*C)"),
    .INIT(16'h7f70))
    _al_u1437 (
    .a(_al_u1436_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z90iu6 ),
    .c(_al_u1334_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pbbbx6 ),
    .o(_al_u1437_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u1438 (
    .a(_al_u1437_o),
    .b(_al_u1348_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [17]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1439 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rs4ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nq4ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[18] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[18] ),
    .o(_al_u1439_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u1440 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lp4ju6 ),
    .b(_al_u1439_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[16] ),
    .o(_al_u1440_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u1441 (
    .a(_al_u1440_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ep4ju6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[16] ),
    .o(_al_u1441_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1442 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ds4ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wr4ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[18] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[18] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vs7pw6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1443 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jo4ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gq4ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[18] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[18] ),
    .o(_al_u1443_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u1444 (
    .a(_al_u1441_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vs7pw6 ),
    .c(_al_u1443_o),
    .o(_al_u1444_o));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~((B*A))*~(C)+~D*(B*A)*~(C)+~(~D)*(B*A)*C+~D*(B*A)*C)"),
    .INIT(16'h7f70))
    _al_u1445 (
    .a(_al_u1444_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S90iu6 ),
    .c(_al_u1334_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Syjbx6 ),
    .o(_al_u1445_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u1446 (
    .a(_al_u1445_o),
    .b(_al_u1348_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [18]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1447 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rs4ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wr4ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[19] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[19] ),
    .o(_al_u1447_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u1448 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ep4ju6 ),
    .b(_al_u1447_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[17] ),
    .o(_al_u1448_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u1449 (
    .a(_al_u1448_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lp4ju6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[17] ),
    .o(_al_u1449_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1450 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ds4ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gq4ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[19] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[19] ),
    .o(_al_u1450_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1451 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jo4ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nq4ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[19] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[19] ),
    .o(_al_u1451_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u1452 (
    .a(_al_u1449_o),
    .b(_al_u1450_o),
    .c(_al_u1451_o),
    .o(_al_u1452_o));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~((B*A))*~(C)+~D*(B*A)*~(C)+~(~D)*(B*A)*C+~D*(B*A)*C)"),
    .INIT(16'h7f70))
    _al_u1453 (
    .a(_al_u1452_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L90iu6 ),
    .c(_al_u1334_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T6kbx6 ),
    .o(_al_u1453_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u1454 (
    .a(_al_u1453_o),
    .b(_al_u1348_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [19]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1455 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gq4ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wr4ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[20] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[20] ),
    .o(_al_u1455_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u1456 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ep4ju6 ),
    .b(_al_u1455_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[18] ),
    .o(_al_u1456_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u1457 (
    .a(_al_u1456_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lp4ju6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[18] ),
    .o(_al_u1457_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1458 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ds4ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rs4ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[20] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[20] ),
    .o(_al_u1458_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1459 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jo4ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nq4ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[20] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[20] ),
    .o(_al_u1459_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u1460 (
    .a(_al_u1457_o),
    .b(_al_u1458_o),
    .c(_al_u1459_o),
    .o(_al_u1460_o));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~((B*A))*~(C)+~D*(B*A)*~(C)+~(~D)*(B*A)*C+~D*(B*A)*C)"),
    .INIT(16'h7f70))
    _al_u1461 (
    .a(_al_u1460_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X80iu6 ),
    .c(_al_u1334_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fjdbx6 ),
    .o(_al_u1461_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u1462 (
    .a(_al_u1461_o),
    .b(_al_u1348_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [20]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1463 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jo4ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rs4ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[21] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[21] ),
    .o(_al_u1463_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u1464 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lp4ju6 ),
    .b(_al_u1463_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[19] ),
    .o(_al_u1464_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u1465 (
    .a(_al_u1464_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ep4ju6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[19] ),
    .o(_al_u1465_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1466 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ds4ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nq4ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[21] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[21] ),
    .o(_al_u1466_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1467 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gq4ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wr4ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[21] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[21] ),
    .o(_al_u1467_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u1468 (
    .a(_al_u1465_o),
    .b(_al_u1466_o),
    .c(_al_u1467_o),
    .o(_al_u1468_o));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~((B*A))*~(C)+~D*(B*A)*~(C)+~(~D)*(B*A)*C+~D*(B*A)*C)"),
    .INIT(16'h7f70))
    _al_u1469 (
    .a(_al_u1468_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q80iu6 ),
    .c(_al_u1334_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M2ebx6 ),
    .o(_al_u1469_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u1470 (
    .a(_al_u1469_o),
    .b(_al_u1348_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [21]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1471 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nq4ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wr4ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[22] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[22] ),
    .o(_al_u1471_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u1472 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lp4ju6 ),
    .b(_al_u1471_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[20] ),
    .o(_al_u1472_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u1473 (
    .a(_al_u1472_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ep4ju6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[20] ),
    .o(_al_u1473_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1474 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ds4ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rs4ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[22] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[22] ),
    .o(_al_u1474_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1475 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jo4ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gq4ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[22] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[22] ),
    .o(_al_u1475_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u1476 (
    .a(_al_u1473_o),
    .b(_al_u1474_o),
    .c(_al_u1475_o),
    .o(_al_u1476_o));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~((B*A))*~(C)+~D*(B*A)*~(C)+~(~D)*(B*A)*C+~D*(B*A)*C)"),
    .INIT(16'h7f70))
    _al_u1477 (
    .a(_al_u1476_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J80iu6 ),
    .c(_al_u1334_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tlebx6 ),
    .o(_al_u1477_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u1478 (
    .a(_al_u1477_o),
    .b(_al_u1348_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [22]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1479 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jo4ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nq4ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[23] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[23] ),
    .o(_al_u1479_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u1480 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lp4ju6 ),
    .b(_al_u1479_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[21] ),
    .o(_al_u1480_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u1481 (
    .a(_al_u1480_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ep4ju6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[21] ),
    .o(_al_u1481_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1482 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ds4ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wr4ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[23] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[23] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C96pw6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1483 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gq4ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rs4ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[23] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[23] ),
    .o(_al_u1483_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u1484 (
    .a(_al_u1481_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C96pw6 ),
    .c(_al_u1483_o),
    .o(_al_u1484_o));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~((B*A))*~(C)+~D*(B*A)*~(C)+~(~D)*(B*A)*C+~D*(B*A)*C)"),
    .INIT(16'h7f70))
    _al_u1485 (
    .a(_al_u1484_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C80iu6 ),
    .c(_al_u1334_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztgbx6 ),
    .o(_al_u1485_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u1486 (
    .a(_al_u1485_o),
    .b(_al_u1348_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [23]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1487 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jo4ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wr4ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[24] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[24] ),
    .o(_al_u1487_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u1488 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lp4ju6 ),
    .b(_al_u1487_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[22] ),
    .o(_al_u1488_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u1489 (
    .a(_al_u1488_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ep4ju6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[22] ),
    .o(_al_u1489_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1490 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ds4ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gq4ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[24] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[24] ),
    .o(_al_u1490_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1491 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rs4ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nq4ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[24] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[24] ),
    .o(_al_u1491_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u1492 (
    .a(_al_u1489_o),
    .b(_al_u1490_o),
    .c(_al_u1491_o),
    .o(_al_u1492_o));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~((B*A))*~(C)+~D*(B*A)*~(C)+~(~D)*(B*A)*C+~D*(B*A)*C)"),
    .INIT(16'h7f70))
    _al_u1493 (
    .a(_al_u1492_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V70iu6 ),
    .c(_al_u1334_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgkbx6 ),
    .o(_al_u1493_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u1494 (
    .a(_al_u1493_o),
    .b(_al_u1348_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [24]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1495 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jo4ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rs4ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[25] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[25] ),
    .o(_al_u1495_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u1496 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lp4ju6 ),
    .b(_al_u1495_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[23] ),
    .o(_al_u1496_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u1497 (
    .a(_al_u1496_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ep4ju6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[23] ),
    .o(_al_u1497_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1498 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ds4ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nq4ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[25] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[25] ),
    .o(_al_u1498_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1499 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gq4ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wr4ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[25] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[25] ),
    .o(_al_u1499_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u1500 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O70iu6 ),
    .b(_al_u1497_o),
    .c(_al_u1498_o),
    .d(_al_u1499_o),
    .o(_al_u1500_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h8b))
    _al_u1501 (
    .a(_al_u1500_o),
    .b(_al_u1334_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nwbbx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mi8ju6_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u1502 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mi8ju6_lutinv ),
    .b(_al_u1348_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [25]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1503 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jo4ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wr4ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[26] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[26] ),
    .o(_al_u1503_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u1504 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lp4ju6 ),
    .b(_al_u1503_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[24] ),
    .o(_al_u1504_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u1505 (
    .a(_al_u1504_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ep4ju6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[24] ),
    .o(_al_u1505_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1506 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ds4ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nq4ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[26] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[26] ),
    .o(_al_u1506_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1507 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gq4ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rs4ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[26] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[26] ),
    .o(_al_u1507_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u1508 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H70iu6 ),
    .b(_al_u1505_o),
    .c(_al_u1506_o),
    .d(_al_u1507_o),
    .o(_al_u1508_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h8b))
    _al_u1509 (
    .a(_al_u1508_o),
    .b(_al_u1334_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F8cbx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E17ju6_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u1510 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E17ju6_lutinv ),
    .b(_al_u1348_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [26]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1511 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gq4ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rs4ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[27] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[27] ),
    .o(_al_u1511_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u1512 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ep4ju6 ),
    .b(_al_u1511_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[25] ),
    .o(_al_u1512_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u1513 (
    .a(_al_u1512_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lp4ju6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[25] ),
    .o(_al_u1513_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1514 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ds4ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jo4ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[27] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[27] ),
    .o(_al_u1514_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1515 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nq4ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wr4ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[27] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[27] ),
    .o(_al_u1515_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u1516 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A70iu6 ),
    .b(_al_u1513_o),
    .c(_al_u1514_o),
    .d(_al_u1515_o),
    .o(_al_u1516_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h8b))
    _al_u1517 (
    .a(_al_u1516_o),
    .b(_al_u1334_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nybbx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F57ju6_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u1518 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F57ju6_lutinv ),
    .b(_al_u1348_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [27]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1519 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rs4ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wr4ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[28] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[28] ),
    .o(_al_u1519_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u1520 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ep4ju6 ),
    .b(_al_u1519_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[26] ),
    .o(_al_u1520_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u1521 (
    .a(_al_u1520_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lp4ju6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[26] ),
    .o(_al_u1521_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1522 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ds4ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nq4ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[28] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[28] ),
    .o(_al_u1522_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1523 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jo4ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gq4ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[28] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[28] ),
    .o(_al_u1523_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u1524 (
    .a(_al_u1521_o),
    .b(_al_u1522_o),
    .c(_al_u1523_o),
    .o(_al_u1524_o));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~((B*A))*~(C)+~D*(B*A)*~(C)+~(~D)*(B*A)*C+~D*(B*A)*C)"),
    .INIT(16'h7f70))
    _al_u1525 (
    .a(_al_u1524_o),
    .b(_al_u823_o),
    .c(_al_u1334_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ibqpw6 ),
    .o(_al_u1525_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u1526 (
    .a(_al_u1525_o),
    .b(_al_u1348_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [28]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1527 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rs4ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nq4ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[29] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[29] ),
    .o(_al_u1527_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u1528 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ep4ju6 ),
    .b(_al_u1527_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[27] ),
    .o(_al_u1528_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u1529 (
    .a(_al_u1528_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lp4ju6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[27] ),
    .o(_al_u1529_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1530 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ds4ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wr4ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[29] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[29] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eq4pw6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1531 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jo4ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gq4ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[29] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[29] ),
    .o(_al_u1531_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u1532 (
    .a(_al_u1529_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eq4pw6 ),
    .c(_al_u1531_o),
    .o(_al_u1532_o));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~((B*A))*~(C)+~D*(B*A)*~(C)+~(~D)*(B*A)*C+~D*(B*A)*C)"),
    .INIT(16'h7f70))
    _al_u1533 (
    .a(_al_u1532_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M60iu6 ),
    .c(_al_u1334_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sx3qw6 ),
    .o(_al_u1533_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u1534 (
    .a(_al_u1533_o),
    .b(_al_u1348_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [29]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1535 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gq4ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wr4ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[30] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[30] ),
    .o(_al_u1535_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u1536 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lp4ju6 ),
    .b(_al_u1535_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[28] ),
    .o(_al_u1536_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u1537 (
    .a(_al_u1536_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ep4ju6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[28] ),
    .o(_al_u1537_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1538 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ds4ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rs4ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[30] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[30] ),
    .o(_al_u1538_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1539 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jo4ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nq4ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[30] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[30] ),
    .o(_al_u1539_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u1540 (
    .a(_al_u1537_o),
    .b(_al_u1538_o),
    .c(_al_u1539_o),
    .o(_al_u1540_o));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~((B*A))*~(C)+~D*(B*A)*~(C)+~(~D)*(B*A)*C+~D*(B*A)*C)"),
    .INIT(16'h7f70))
    _al_u1541 (
    .a(_al_u1540_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y50iu6 ),
    .c(_al_u1334_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F6dbx6 ),
    .o(_al_u1541_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u1542 (
    .a(_al_u1541_o),
    .b(_al_u1348_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [30]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1543 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gq4ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wr4ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[6] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[6] ),
    .o(_al_u1543_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u1544 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lp4ju6 ),
    .b(_al_u1543_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[4] ),
    .o(_al_u1544_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u1545 (
    .a(_al_u1544_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ep4ju6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[4] ),
    .o(_al_u1545_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1546 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ds4ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jo4ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[6] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[6] ),
    .o(_al_u1546_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1547 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rs4ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nq4ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[6] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[6] ),
    .o(_al_u1547_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u1548 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P40iu6 ),
    .b(_al_u1545_o),
    .c(_al_u1546_o),
    .d(_al_u1547_o),
    .o(_al_u1548_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h8b))
    _al_u1549 (
    .a(_al_u1548_o),
    .b(_al_u1334_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ua9bx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mk6ju6_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u1550 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mk6ju6_lutinv ),
    .b(_al_u1348_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [6]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1551 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jo4ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nq4ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[9] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[9] ),
    .o(_al_u1551_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u1552 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lp4ju6 ),
    .b(_al_u1551_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[7] ),
    .o(_al_u1552_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u1553 (
    .a(_al_u1552_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ep4ju6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[7] ),
    .o(_al_u1553_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1554 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ds4ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rs4ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[9] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[9] ),
    .o(_al_u1554_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1555 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gq4ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wr4ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[9] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[9] ),
    .o(_al_u1555_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u1556 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U30iu6 ),
    .b(_al_u1553_o),
    .c(_al_u1554_o),
    .d(_al_u1555_o),
    .o(_al_u1556_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h8b))
    _al_u1557 (
    .a(_al_u1556_o),
    .b(_al_u1334_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kn1qw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N18ju6_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u1558 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N18ju6_lutinv ),
    .b(_al_u1348_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [9]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1559 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rs4ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wr4ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[31] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[31] ),
    .o(_al_u1559_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u1560 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lp4ju6 ),
    .b(_al_u1559_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[29] ),
    .o(_al_u1560_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u1561 (
    .a(_al_u1560_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ep4ju6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[29] ),
    .o(_al_u1561_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1562 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ds4ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gq4ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[31] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[31] ),
    .o(_al_u1562_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1563 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jo4ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nq4ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[31] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[31] ),
    .o(_al_u1563_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u1564 (
    .a(_al_u1561_o),
    .b(_al_u1562_o),
    .c(_al_u1563_o),
    .o(_al_u1564_o));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~((B*A))*~(C)+~D*(B*A)*~(C)+~(~D)*(B*A)*C+~D*(B*A)*C)"),
    .INIT(16'h7f70))
    _al_u1565 (
    .a(_al_u1564_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R50iu6 ),
    .c(_al_u1334_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Usnpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/To2ju6_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u1566 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/To2ju6_lutinv ),
    .b(_al_u1348_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [31]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1567 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jo4ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wr4ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[4] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[4] ),
    .o(_al_u1567_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u1568 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lp4ju6 ),
    .b(_al_u1567_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[2] ),
    .o(_al_u1568_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u1569 (
    .a(_al_u1568_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ep4ju6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[2] ),
    .o(_al_u1569_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1570 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ds4ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nq4ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[4] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[4] ),
    .o(_al_u1570_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1571 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gq4ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rs4ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[4] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[4] ),
    .o(_al_u1571_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u1572 (
    .a(_al_u1569_o),
    .b(_al_u1570_o),
    .c(_al_u1571_o),
    .o(_al_u1572_o));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~((B*A))*~(C)+~D*(B*A)*~(C)+~(~D)*(B*A)*C+~D*(B*A)*C)"),
    .INIT(16'h7f70))
    _al_u1573 (
    .a(_al_u1572_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D50iu6 ),
    .c(_al_u1334_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wtxax6 ),
    .o(_al_u1573_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u1574 (
    .a(_al_u1573_o),
    .b(_al_u1348_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [4]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1575 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jo4ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wr4ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[2] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[2] ),
    .o(_al_u1575_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u1576 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lp4ju6 ),
    .b(_al_u1575_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[0] ),
    .o(_al_u1576_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u1577 (
    .a(_al_u1576_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ep4ju6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[0] ),
    .o(_al_u1577_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1578 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ds4ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gq4ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[2] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[2] ),
    .o(_al_u1578_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1579 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rs4ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nq4ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[2] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[2] ),
    .o(_al_u1579_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u1580 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F60iu6 ),
    .b(_al_u1577_o),
    .c(_al_u1578_o),
    .d(_al_u1579_o),
    .o(_al_u1580_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h8b))
    _al_u1581 (
    .a(_al_u1580_o),
    .b(_al_u1334_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xrxax6 ),
    .o(_al_u1581_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u1582 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 ),
    .o(_al_u1582_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u1583 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ),
    .o(_al_u1583_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u1584 (
    .a(_al_u1582_o),
    .b(_al_u1583_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vgjpw6 ),
    .o(_al_u1584_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u1585 (
    .a(_al_u1581_o),
    .b(_al_u1348_o),
    .c(_al_u1584_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [2]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1586 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jo4ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wr4ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[3] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[3] ),
    .o(_al_u1586_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u1587 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lp4ju6 ),
    .b(_al_u1586_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[1] ),
    .o(_al_u1587_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u1588 (
    .a(_al_u1587_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ep4ju6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[1] ),
    .o(_al_u1588_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1589 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ds4ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nq4ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[3] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[3] ),
    .o(_al_u1589_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1590 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gq4ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rs4ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[3] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[3] ),
    .o(_al_u1590_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u1591 (
    .a(_al_u1588_o),
    .b(_al_u1589_o),
    .c(_al_u1590_o),
    .o(_al_u1591_o));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~((B*A))*~(C)+~D*(B*A)*~(C)+~(~D)*(B*A)*C+~D*(B*A)*C)"),
    .INIT(16'h7f70))
    _al_u1592 (
    .a(_al_u1591_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K50iu6 ),
    .c(_al_u1334_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T5yax6 ),
    .o(_al_u1592_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u1593 (
    .a(_al_u1592_o),
    .b(_al_u1348_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [3]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1594 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nq4ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wr4ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[5] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[5] ),
    .o(_al_u1594_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u1595 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lp4ju6 ),
    .b(_al_u1594_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[3] ),
    .o(_al_u1595_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u1596 (
    .a(_al_u1595_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ep4ju6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[3] ),
    .o(_al_u1596_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1597 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ds4ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rs4ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[5] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[5] ),
    .o(_al_u1597_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1598 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jo4ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gq4ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[5] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[5] ),
    .o(_al_u1598_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u1599 (
    .a(_al_u1596_o),
    .b(_al_u1597_o),
    .c(_al_u1598_o),
    .o(_al_u1599_o));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~((B*A))*~(C)+~D*(B*A)*~(C)+~(~D)*(B*A)*C+~D*(B*A)*C)"),
    .INIT(16'h7f70))
    _al_u1600 (
    .a(_al_u1599_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W40iu6 ),
    .c(_al_u1334_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qc5bx6 ),
    .o(_al_u1600_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u1601 (
    .a(_al_u1600_o),
    .b(_al_u1348_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [5]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1602 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jo4ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nq4ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[8] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[8] ),
    .o(_al_u1602_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u1603 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lp4ju6 ),
    .b(_al_u1602_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[6] ),
    .o(_al_u1603_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u1604 (
    .a(_al_u1603_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ep4ju6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[6] ),
    .o(_al_u1604_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1605 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ds4ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rs4ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[8] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[8] ),
    .o(_al_u1605_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1606 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gq4ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wr4ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[8] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[8] ),
    .o(_al_u1606_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u1607 (
    .a(_al_u1604_o),
    .b(_al_u1605_o),
    .c(_al_u1606_o),
    .o(_al_u1607_o));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~((B*A))*~(C)+~D*(B*A)*~(C)+~(~D)*(B*A)*C+~D*(B*A)*C)"),
    .INIT(16'h7f70))
    _al_u1608 (
    .a(_al_u1607_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B40iu6 ),
    .c(_al_u1334_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N61qw6 ),
    .o(_al_u1608_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u1609 (
    .a(_al_u1608_o),
    .b(_al_u1348_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [8]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1610 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jo4ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wr4ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[7] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[7] ),
    .o(_al_u1610_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u1611 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lp4ju6 ),
    .b(_al_u1610_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[5] ),
    .o(_al_u1611_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u1612 (
    .a(_al_u1611_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ep4ju6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[5] ),
    .o(_al_u1612_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1613 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ds4ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gq4ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[7] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[7] ),
    .o(_al_u1613_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1614 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rs4ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nq4ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[7] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[7] ),
    .o(_al_u1614_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u1615 (
    .a(_al_u1612_o),
    .b(_al_u1613_o),
    .c(_al_u1614_o),
    .o(_al_u1615_o));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~((B*A))*~(C)+~D*(B*A)*~(C)+~(~D)*(B*A)*C+~D*(B*A)*C)"),
    .INIT(16'h7f70))
    _al_u1616 (
    .a(_al_u1615_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I40iu6 ),
    .c(_al_u1334_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Asupw6 ),
    .o(_al_u1616_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u1617 (
    .a(_al_u1616_o),
    .b(_al_u1348_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [7]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1618 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nq4ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wr4ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[10] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[10] ),
    .o(_al_u1618_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u1619 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lp4ju6 ),
    .b(_al_u1618_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[8] ),
    .o(_al_u1619_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u1620 (
    .a(_al_u1619_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ep4ju6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[8] ),
    .o(_al_u1620_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1621 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ds4ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jo4ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[10] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[10] ),
    .o(_al_u1621_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1622 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gq4ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rs4ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[10] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[10] ),
    .o(_al_u1622_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u1623 (
    .a(_al_u1620_o),
    .b(_al_u1621_o),
    .c(_al_u1622_o),
    .o(_al_u1623_o));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~((B*A))*~(C)+~D*(B*A)*~(C)+~(~D)*(B*A)*C+~D*(B*A)*C)"),
    .INIT(16'h7f70))
    _al_u1624 (
    .a(_al_u1623_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wb0iu6 ),
    .c(_al_u1334_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gwxpw6 ),
    .o(_al_u1624_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u1625 (
    .a(_al_u1624_o),
    .b(_al_u1348_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [10]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1626 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jo4ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wr4ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[11] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[11] ),
    .o(_al_u1626_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u1627 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lp4ju6 ),
    .b(_al_u1626_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[9] ),
    .o(_al_u1627_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u1628 (
    .a(_al_u1627_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ep4ju6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[9] ),
    .o(_al_u1628_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1629 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ds4ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gq4ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[11] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[11] ),
    .o(_al_u1629_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1630 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rs4ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nq4ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[11] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[11] ),
    .o(_al_u1630_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u1631 (
    .a(_al_u1628_o),
    .b(_al_u1629_o),
    .c(_al_u1630_o),
    .o(_al_u1631_o));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~((B*A))*~(C)+~D*(B*A)*~(C)+~(~D)*(B*A)*C+~D*(B*A)*C)"),
    .INIT(16'h7f70))
    _al_u1632 (
    .a(_al_u1631_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pb0iu6 ),
    .c(_al_u1334_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C07bx6 ),
    .o(_al_u1632_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u1633 (
    .a(_al_u1632_o),
    .b(_al_u1348_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [11]));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(B*~(~D*C)))"),
    .INIT(16'h1151))
    _al_u1634 (
    .a(_al_u1363_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wkipw6 ),
    .o(_al_u1634_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u1635 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 ),
    .o(_al_u1635_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u1636 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P14qw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rwjax6 ),
    .o(_al_u1636_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    _al_u1637 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mb1ju6 ),
    .b(_al_u1634_o),
    .c(_al_u1635_o),
    .d(_al_u1636_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ir6ow6 ));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u1638 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Srbow6 ),
    .b(_al_u1359_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6 ),
    .o(_al_u1638_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*~B))"),
    .INIT(8'h75))
    _al_u1639 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ir6ow6 ),
    .b(_al_u1638_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N4kax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jrhow6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u1640 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[0] ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[1] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ukbpw6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    _al_u1641 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M8row6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ukbpw6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[4] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[5] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hlliu6 ));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u1642 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[27] ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[28] ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zdiax6 ),
    .o(_al_u1642_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*~A)"),
    .INIT(16'h4000))
    _al_u1643 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hlliu6 ),
    .b(_al_u1642_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[29] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[30] ),
    .o(_al_u1643_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u1644 (
    .a(_al_u1643_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_control_o ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[1] ),
    .o(_al_u1644_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u1645 (
    .a(_al_u903_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wkipw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xqoiu6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*A)"),
    .INIT(16'h0080))
    _al_u1646 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xqoiu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S7mpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wfspw6 ),
    .o(_al_u1646_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(D*~C*B))"),
    .INIT(16'h5155))
    _al_u1647 (
    .a(_al_u1646_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Llaow6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wfspw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G7aiu6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .INIT(16'h5140))
    _al_u1648 (
    .a(_al_u1635_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wkipw6 ),
    .o(_al_u1648_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+A*~(B)*C*D+A*B*C*D)"),
    .INIT(16'haf30))
    _al_u1649 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R9aiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P8aiu6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("~(B*~(~A*~(~D*C)))"),
    .INIT(16'h7737))
    _al_u1650 (
    .a(_al_u1644_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G7aiu6_lutinv ),
    .c(_al_u1648_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P8aiu6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cy9iu6 ));
  AL_MAP_LUT2 #(
    .EQN("~(~B*A)"),
    .INIT(4'hd))
    _al_u1651 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/DBGRESTARTED ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vyuhu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*~A))"),
    .INIT(16'h23af))
    _al_u1652 (
    .a(_al_u1360_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fb1ju6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Irmpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6 ),
    .o(_al_u1652_o));
  AL_MAP_LUT4 #(
    .EQN("~(B*A*~(D*C))"),
    .INIT(16'hf777))
    _al_u1653 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ir6ow6 ),
    .b(_al_u1652_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P91ju6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jckax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rnbow6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*~A))"),
    .INIT(16'h2a3f))
    _al_u1654 (
    .a(_al_u1360_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fb1ju6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wfspw6 ),
    .o(_al_u1654_o));
  AL_MAP_LUT4 #(
    .EQN("~(B*A*~(D*C))"),
    .INIT(16'hf777))
    _al_u1655 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ir6ow6 ),
    .b(_al_u1654_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P91ju6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wkipw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zp6ow6 ));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u1656 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ldoiu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 ),
    .o(_al_u1656_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    _al_u1657 (
    .a(_al_u1656_o),
    .b(_al_u604_o),
    .c(_al_u1346_o),
    .o(_al_u1657_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u1658 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 ),
    .o(_al_u1658_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u1659 (
    .a(_al_u1658_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 ),
    .o(_al_u1659_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*~A)"),
    .INIT(8'h04))
    _al_u1660 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 ),
    .o(_al_u1660_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~A*~(C*B))"),
    .INIT(16'h0015))
    _al_u1661 (
    .a(_al_u1659_o),
    .b(_al_u679_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D6kiu6_lutinv ),
    .d(_al_u1660_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lu0iu6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u1662 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 ),
    .o(_al_u1662_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u1663 (
    .a(_al_u1662_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 ),
    .o(_al_u1663_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(~D*C))"),
    .INIT(16'h4404))
    _al_u1664 (
    .a(_al_u1657_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lu0iu6 ),
    .c(_al_u1663_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 ),
    .o(_al_u1664_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u1665 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S2ziu6_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u1666 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S2ziu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vs0iu6 ));
  AL_MAP_LUT4 #(
    .EQN("~(B*~((~D*A))*~(C)+B*(~D*A)*~(C)+~(B)*(~D*A)*C+B*(~D*A)*C)"),
    .INIT(16'hf353))
    _al_u1667 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T23ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 ),
    .o(_al_u1667_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(~A*~(C*~B)))"),
    .INIT(16'hba00))
    _al_u1668 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vs0iu6 ),
    .b(_al_u1667_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_apsr_o[1] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 ),
    .o(_al_u1668_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(~B*A))"),
    .INIT(8'hd0))
    _al_u1669 (
    .a(_al_u1664_o),
    .b(_al_u1668_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vgjpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dqfhu6 ));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    _al_u1670 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B7lpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P13iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ryfax6 ),
    .o(_al_u1670_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D@C))"),
    .INIT(16'h8008))
    _al_u1671 (
    .a(_al_u1253_o),
    .b(_al_u1670_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qwfax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Utqpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gf1ju6 ));
  AL_MAP_LUT4 #(
    .EQN("(A*~(~D*~(C*B)))"),
    .INIT(16'haa80))
    _al_u1672 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gf1ju6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pyyhu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Krlpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zslpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vk1iu6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u1673 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Golpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zslpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yn3iu6_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u1674 (
    .a(_al_u1253_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yn3iu6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y93iu6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u1675 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y93iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vplpw6 ),
    .o(_al_u1675_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u1676 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahlpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pmlpw6 ),
    .o(_al_u1676_o));
  AL_MAP_LUT4 #(
    .EQN("~((D*~A)*~(C)*~(B)+(D*~A)*C*~(B)+~((D*~A))*C*B+(D*~A)*C*B)"),
    .INIT(16'h2e3f))
    _al_u1677 (
    .a(_al_u1253_o),
    .b(_al_u1676_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bx2qw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Li7ax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yg3iu6 ));
  AL_MAP_LUT4 #(
    .EQN("~(C*~B*~(D*A))"),
    .INIT(16'hefcf))
    _al_u1678 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vk1iu6 ),
    .b(_al_u1675_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yg3iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hg7ax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Urxhu6 ));
  AL_MAP_LUT4 #(
    .EQN("~((C*~A)*~(D)*~(B)+(C*~A)*D*~(B)+~((C*~A))*D*B+(C*~A)*D*B)"),
    .INIT(16'h23ef))
    _al_u1679 (
    .a(_al_u1253_o),
    .b(_al_u1676_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bx2qw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z73qw6 ),
    .o(_al_u1679_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C*A))"),
    .INIT(8'hb3))
    _al_u1680 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vk1iu6 ),
    .b(_al_u1679_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xu2qw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bsxhu6 ));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u1681 (
    .a(_al_u1675_o),
    .b(_al_u1676_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D2opw6 ),
    .o(_al_u1681_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u1682 (
    .a(_al_u1253_o),
    .b(_al_u1676_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xl1iu6_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u1683 (
    .a(_al_u1681_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xl1iu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z73qw6 ),
    .o(_al_u1683_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*B))"),
    .INIT(8'hd5))
    _al_u1684 (
    .a(_al_u1683_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vk1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V53qw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Psxhu6 ));
  AL_MAP_LUT4 #(
    .EQN("~((C*~A)*~(D)*~(B)+(C*~A)*D*~(B)+~((C*~A))*D*B+(C*~A)*D*B)"),
    .INIT(16'h23ef))
    _al_u1685 (
    .a(_al_u1253_o),
    .b(_al_u1676_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qa1qw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qj1qw6 ),
    .o(_al_u1685_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C*A))"),
    .INIT(8'hb3))
    _al_u1686 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vk1iu6 ),
    .b(_al_u1685_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M81qw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vvxhu6 ));
  AL_MAP_LUT4 #(
    .EQN("~((D*~A)*~(C)*~(B)+(D*~A)*C*~(B)+~((D*~A))*C*B+(D*~A)*C*B)"),
    .INIT(16'h2e3f))
    _al_u1687 (
    .a(_al_u1253_o),
    .b(_al_u1676_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L0ypw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qj1qw6 ),
    .o(_al_u1687_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C*A))"),
    .INIT(8'hb3))
    _al_u1688 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vk1iu6 ),
    .b(_al_u1687_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mh1qw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cwxhu6 ));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u1689 (
    .a(_al_u1675_o),
    .b(_al_u1676_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gw6bx6 ),
    .o(_al_u1689_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u1690 (
    .a(_al_u1689_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xl1iu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L0ypw6 ),
    .o(_al_u1690_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*B))"),
    .INIT(8'hd5))
    _al_u1691 (
    .a(_al_u1690_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vk1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gyxpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jwxhu6 ));
  AL_MAP_LUT4 #(
    .EQN("~((C*~A)*~(D)*~(B)+(C*~A)*D*~(B)+~((C*~A))*D*B+(C*~A)*D*B)"),
    .INIT(16'h23ef))
    _al_u1692 (
    .a(_al_u1253_o),
    .b(_al_u1676_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gw6bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wq8ax6 ),
    .o(_al_u1692_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C*A))"),
    .INIT(8'hb3))
    _al_u1693 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vk1iu6 ),
    .b(_al_u1692_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bu6bx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qwxhu6 ));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u1694 (
    .a(_al_u1675_o),
    .b(_al_u1676_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oh8ax6 ),
    .o(_al_u1694_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u1695 (
    .a(_al_u1694_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xl1iu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wq8ax6 ),
    .o(_al_u1695_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*B))"),
    .INIT(8'hd5))
    _al_u1696 (
    .a(_al_u1695_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vk1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ro8ax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xwxhu6 ));
  AL_MAP_LUT4 #(
    .EQN("~((C*~A)*~(D)*~(B)+(C*~A)*D*~(B)+~((C*~A))*D*B+(C*~A)*D*B)"),
    .INIT(16'h23ef))
    _al_u1697 (
    .a(_al_u1253_o),
    .b(_al_u1676_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oh8ax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xf8ax6 ),
    .o(_al_u1697_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C*A))"),
    .INIT(8'hb3))
    _al_u1698 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vk1iu6 ),
    .b(_al_u1697_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ggabx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Exxhu6 ));
  AL_MAP_LUT4 #(
    .EQN("~((D*~A)*~(C)*~(B)+(D*~A)*C*~(B)+~((D*~A))*C*B+(D*~A)*C*B)"),
    .INIT(16'h2e3f))
    _al_u1699 (
    .a(_al_u1253_o),
    .b(_al_u1676_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E97ax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xf8ax6 ),
    .o(_al_u1699_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C*A))"),
    .INIT(8'hb3))
    _al_u1700 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vk1iu6 ),
    .b(_al_u1699_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sd8ax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lxxhu6 ));
  AL_MAP_LUT4 #(
    .EQN("~((C*~A)*~(D)*~(B)+(C*~A)*D*~(B)+~((C*~A))*D*B+(C*~A)*D*B)"),
    .INIT(16'h23ef))
    _al_u1701 (
    .a(_al_u1253_o),
    .b(_al_u1676_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E97ax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hlwpw6 ),
    .o(_al_u1701_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C*A))"),
    .INIT(8'hb3))
    _al_u1702 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vk1iu6 ),
    .b(_al_u1701_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z67ax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sxxhu6 ));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u1703 (
    .a(_al_u1675_o),
    .b(_al_u1676_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufbbx6 ),
    .o(_al_u1703_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u1704 (
    .a(_al_u1703_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xl1iu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hlwpw6 ),
    .o(_al_u1704_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*B))"),
    .INIT(8'hd5))
    _al_u1705 (
    .a(_al_u1704_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vk1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cjwpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zxxhu6 ));
  AL_MAP_LUT4 #(
    .EQN("~((D*~A)*~(C)*~(B)+(D*~A)*C*~(B)+~((D*~A))*C*B+(D*~A)*C*B)"),
    .INIT(16'h2e3f))
    _al_u1706 (
    .a(_al_u1253_o),
    .b(_al_u1676_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Puwpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufbbx6 ),
    .o(_al_u1706_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C*A))"),
    .INIT(8'hb3))
    _al_u1707 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vk1iu6 ),
    .b(_al_u1706_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pdbbx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gyxhu6 ));
  AL_MAP_LUT4 #(
    .EQN("~((D*~A)*~(C)*~(B)+(D*~A)*C*~(B)+~((D*~A))*C*B+(D*~A)*C*B)"),
    .INIT(16'h2e3f))
    _al_u1708 (
    .a(_al_u1253_o),
    .b(_al_u1676_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ldvpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Puwpw6 ),
    .o(_al_u1708_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C*A))"),
    .INIT(8'hb3))
    _al_u1709 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vk1iu6 ),
    .b(_al_u1708_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kswpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nyxhu6 ));
  AL_MAP_LUT4 #(
    .EQN("~((D*~A)*~(C)*~(B)+(D*~A)*C*~(B)+~((D*~A))*C*B+(D*~A)*C*B)"),
    .INIT(16'h2e3f))
    _al_u1710 (
    .a(_al_u1253_o),
    .b(_al_u1676_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jfdbx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ldvpw6 ),
    .o(_al_u1710_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C*A))"),
    .INIT(8'hb3))
    _al_u1711 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vk1iu6 ),
    .b(_al_u1710_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gbvpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uyxhu6 ));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u1712 (
    .a(_al_u1675_o),
    .b(_al_u1676_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sddbx6 ),
    .o(_al_u1712_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u1713 (
    .a(_al_u1712_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xl1iu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jfdbx6 ),
    .o(_al_u1713_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*B))"),
    .INIT(8'hd5))
    _al_u1714 (
    .a(_al_u1713_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vk1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cydbx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bzxhu6 ));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u1715 (
    .a(_al_u1675_o),
    .b(_al_u1676_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bcdbx6 ),
    .o(_al_u1715_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u1716 (
    .a(_al_u1715_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xl1iu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sddbx6 ),
    .o(_al_u1716_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*B))"),
    .INIT(8'hd5))
    _al_u1717 (
    .a(_al_u1716_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vk1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jhebx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Izxhu6 ));
  AL_MAP_LUT4 #(
    .EQN("~((C*~A)*~(D)*~(B)+(C*~A)*D*~(B)+~((C*~A))*D*B+(C*~A)*D*B)"),
    .INIT(16'h23ef))
    _al_u1718 (
    .a(_al_u1253_o),
    .b(_al_u1676_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bcdbx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kadbx6 ),
    .o(_al_u1718_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C*A))"),
    .INIT(8'hb3))
    _al_u1719 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vk1iu6 ),
    .b(_al_u1718_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qwfbx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pzxhu6 ));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u1720 (
    .a(_al_u1675_o),
    .b(_al_u1676_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Stkpw6 ),
    .o(_al_u1720_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u1721 (
    .a(_al_u1720_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xl1iu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kadbx6 ),
    .o(_al_u1721_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*B))"),
    .INIT(8'hd5))
    _al_u1722 (
    .a(_al_u1721_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vk1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F8dbx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wzxhu6 ));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u1723 (
    .a(_al_u1675_o),
    .b(_al_u1676_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kn2qw6 ),
    .o(_al_u1723_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u1724 (
    .a(_al_u1723_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xl1iu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Stkpw6 ),
    .o(_al_u1724_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*B))"),
    .INIT(8'hd5))
    _al_u1725 (
    .a(_al_u1724_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vk1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nrkpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D0yhu6 ));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u1726 (
    .a(_al_u1675_o),
    .b(_al_u1676_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J4cbx6 ),
    .o(_al_u1726_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u1727 (
    .a(_al_u1726_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xl1iu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kn2qw6 ),
    .o(_al_u1727_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*B))"),
    .INIT(8'hd5))
    _al_u1728 (
    .a(_al_u1727_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vk1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fl2qw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K0yhu6 ));
  AL_MAP_LUT4 #(
    .EQN("~((C*~A)*~(D)*~(B)+(C*~A)*D*~(B)+~((C*~A))*D*B+(C*~A)*D*B)"),
    .INIT(16'h23ef))
    _al_u1729 (
    .a(_al_u1253_o),
    .b(_al_u1676_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J4cbx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S2cbx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P92iu6 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u1730 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vk1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P92iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cncbx6 ),
    .o(_al_u1730_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u1731 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y93iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oulpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vplpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cl1iu6 ));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*B))"),
    .INIT(8'hd5))
    _al_u1732 (
    .a(_al_u1730_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cl1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hpcbx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R0yhu6 ));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u1733 (
    .a(_al_u1675_o),
    .b(_al_u1676_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nfqpw6 ),
    .o(_al_u1733_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u1734 (
    .a(_al_u1733_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xl1iu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S2cbx6 ),
    .o(_al_u1734_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*B))"),
    .INIT(8'hd5))
    _al_u1735 (
    .a(_al_u1734_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vk1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N0cbx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y0yhu6 ));
  AL_MAP_LUT4 #(
    .EQN("~((C*~A)*~(D)*~(B)+(C*~A)*D*~(B)+~((C*~A))*D*B+(C*~A)*D*B)"),
    .INIT(16'h23ef))
    _al_u1736 (
    .a(_al_u1253_o),
    .b(_al_u1676_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nfqpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wt3qw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V52iu6 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u1737 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vk1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V52iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idqpw6 ),
    .o(_al_u1737_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*B))"),
    .INIT(8'hd5))
    _al_u1738 (
    .a(_al_u1737_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cl1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ehqpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F1yhu6 ));
  AL_MAP_LUT4 #(
    .EQN("~((D*~A)*~(C)*~(B)+(D*~A)*C*~(B)+~((D*~A))*C*B+(D*~A)*C*B)"),
    .INIT(16'h2e3f))
    _al_u1739 (
    .a(_al_u1253_o),
    .b(_al_u1676_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C72qw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wt3qw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P22iu6 ));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B*~(D*A)))"),
    .INIT(16'hb030))
    _al_u1740 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cjqpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ehqpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T0ipw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/cpu0cdbgpwrupreq ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F42iu6 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u1741 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cl1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P22iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F42iu6 ),
    .o(_al_u1741_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*B))"),
    .INIT(8'hd5))
    _al_u1742 (
    .a(_al_u1741_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vk1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rr3qw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M1yhu6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u1743 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cl1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T82qw6 ),
    .o(_al_u1743_o));
  AL_MAP_LUT4 #(
    .EQN("~((C*~A)*~(D)*~(B)+(C*~A)*D*~(B)+~((C*~A))*D*B+(C*~A)*D*B)"),
    .INIT(16'h23ef))
    _al_u1744 (
    .a(_al_u1253_o),
    .b(_al_u1676_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C72qw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zwnpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S02iu6 ));
  AL_MAP_LUT4 #(
    .EQN("~(C*~A*~(D*B))"),
    .INIT(16'hefaf))
    _al_u1745 (
    .a(_al_u1743_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vk1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S02iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X42qw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1yhu6 ));
  AL_MAP_LUT4 #(
    .EQN("~((D*~A)*~(C)*~(B)+(D*~A)*C*~(B)+~((D*~A))*C*B+(D*~A)*C*B)"),
    .INIT(16'h2e3f))
    _al_u1746 (
    .a(_al_u1253_o),
    .b(_al_u1676_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rilpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zwnpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ay1iu6 ));
  AL_MAP_LUT4 #(
    .EQN("~(C*~A*~(D*B))"),
    .INIT(16'hefaf))
    _al_u1747 (
    .a(_al_u1743_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vk1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ay1iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uunpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A2yhu6 ));
  AL_MAP_LUT4 #(
    .EQN("~((D*~A)*~(C)*~(B)+(D*~A)*C*~(B)+~((D*~A))*C*B+(D*~A)*C*B)"),
    .INIT(16'h2e3f))
    _al_u1748 (
    .a(_al_u1253_o),
    .b(_al_u1676_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qa1qw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yzlpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tj1iu6 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u1749 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cl1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tj1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ry2qw6 ),
    .o(_al_u1749_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*B))"),
    .INIT(8'hd5))
    _al_u1750 (
    .a(_al_u1749_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vk1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nckbx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C3yhu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1751 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vk1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cl1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gylpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vefax6 ),
    .o(_al_u1751_o));
  AL_MAP_LUT4 #(
    .EQN("~((D*~A)*~(C)*~(B)+(D*~A)*C*~(B)+~((D*~A))*C*B+(D*~A)*C*B)"),
    .INIT(16'h2e3f))
    _al_u1752 (
    .a(_al_u1253_o),
    .b(_al_u1676_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yzlpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgfax6 ),
    .o(_al_u1752_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(A*~(D*~C)))"),
    .INIT(16'h4c44))
    _al_u1753 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y93iu6 ),
    .b(_al_u1752_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oulpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vplpw6 ),
    .o(_al_u1753_o));
  AL_MAP_LUT2 #(
    .EQN("~(B*A)"),
    .INIT(4'h7))
    _al_u1754 (
    .a(_al_u1751_o),
    .b(_al_u1753_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dtxhu6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u1755 (
    .a(_al_u529_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kalpw6 ),
    .o(_al_u1755_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u1756 (
    .a(_al_u1755_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jflpw6 ),
    .o(_al_u1756_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u1757 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jflpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kalpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sdlpw6 ),
    .o(_al_u1757_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(D*C*B))"),
    .INIT(16'h1555))
    _al_u1758 (
    .a(_al_u1756_o),
    .b(_al_u1757_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bclpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Krlpw6 ),
    .o(_al_u1758_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*~A)"),
    .INIT(8'h04))
    _al_u1759 (
    .a(_al_u1758_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U5yhu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yklpw6 ),
    .o(_al_u1759_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u1760 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pmlpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sdlpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yklpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cayhu6 ));
  AL_MAP_LUT4 #(
    .EQN("~(C*~((D*~A))*~(B)+C*(D*~A)*~(B)+~(C)*(D*~A)*B+C*(D*~A)*B)"),
    .INIT(16'h8bcf))
    _al_u1761 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cayhu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahlpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pmlpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rilpw6 ),
    .o(_al_u1761_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*(C@(D*A)))"),
    .INIT(16'h1230))
    _al_u1762 (
    .a(_al_u1756_o),
    .b(_al_u1761_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pmlpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yklpw6 ),
    .o(_al_u1762_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u1763 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cayhu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahlpw6 ),
    .o(_al_u1763_o));
  AL_MAP_LUT4 #(
    .EQN("~(~B*~A*~(D*C))"),
    .INIT(16'hfeee))
    _al_u1764 (
    .a(_al_u1759_o),
    .b(_al_u1762_o),
    .c(_al_u1763_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rilpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zehpw6 [5]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u1765 (
    .a(_al_u1383_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Umkax6 ),
    .o(_al_u1765_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u1766 (
    .a(_al_u1765_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V6jax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eoyiu6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(D*C*B))"),
    .INIT(16'h1555))
    _al_u1767 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eoyiu6_lutinv ),
    .b(_al_u916_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ubypw6 ),
    .o(_al_u1767_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1768 (
    .a(_al_u696_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A95iu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rkkax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wkipw6 ),
    .o(_al_u1768_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u1769 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4jax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 ),
    .o(_al_u1769_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*~(D*~C)))"),
    .INIT(16'h2a22))
    _al_u1770 (
    .a(_al_u1768_o),
    .b(_al_u1769_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P14qw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Skjax6 ),
    .o(_al_u1770_o));
  AL_MAP_LUT4 #(
    .EQN("~(C*B*~(D*~A))"),
    .INIT(16'h7f3f))
    _al_u1771 (
    .a(_al_u1767_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gpyiu6 ),
    .c(_al_u1770_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L45iu6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Flyiu6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u1772 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[0] ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[1] ),
    .o(_al_u1772_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u1773 (
    .a(_al_u1772_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[4] ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[5] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F8row6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u1774 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F8row6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M8row6_lutinv ),
    .o(_al_u1774_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u1775 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D6kiu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ),
    .o(_al_u1775_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u1776 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yecpw6_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u1777 (
    .a(_al_u1775_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yecpw6_lutinv ),
    .o(_al_u1777_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u1778 (
    .a(_al_u1774_o),
    .b(_al_u1777_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hdfax6 ),
    .o(_al_u1778_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(~A*~(C*B)))"),
    .INIT(16'hea00))
    _al_u1779 (
    .a(_al_u1778_o),
    .b(_al_u933_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eafax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gr2qw6 ),
    .o(_al_u1779_o));
  AL_MAP_LUT4 #(
    .EQN("~(~A*~(D*~(C*B)))"),
    .INIT(16'hbfaa))
    _al_u1780 (
    .a(_al_u1779_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Scbiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Df4iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Thiax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Frthu6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u1781 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 ),
    .o(_al_u1781_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u1782 (
    .a(_al_u1781_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 ),
    .o(_al_u1782_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u1783 (
    .a(_al_u1782_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Daiax6 ),
    .o(_al_u1783_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u1784 (
    .a(_al_u1783_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 ),
    .o(_al_u1784_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    _al_u1785 (
    .a(_al_u606_o),
    .b(_al_u607_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ),
    .o(_al_u1785_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u1786 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pu1ju6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(~B*~A*~(D*C))"),
    .INIT(16'h0111))
    _al_u1787 (
    .a(_al_u906_o),
    .b(_al_u1785_o),
    .c(_al_u932_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pu1ju6_lutinv ),
    .o(_al_u1787_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D*C*B))"),
    .INIT(16'h2aaa))
    _al_u1788 (
    .a(_al_u1787_o),
    .b(_al_u1775_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yecpw6_lutinv ),
    .o(_al_u1788_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u1789 (
    .a(_al_u1784_o),
    .b(_al_u1788_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uzaiu6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u1790 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[0] ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[1] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A9row6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    _al_u1791 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M8row6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A9row6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[4] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[5] ),
    .o(_al_u1791_o));
  AL_MAP_LUT4 #(
    .EQN("~((B*A)*~(C)*~(D)+(B*A)*C*~(D)+~((B*A))*C*D+(B*A)*C*D)"),
    .INIT(16'h0f77))
    _al_u1792 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uzaiu6 ),
    .b(_al_u1791_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F9vpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I8lax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bofiu6_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    _al_u1793 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bofiu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n3685 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vygax6 ),
    .o(_al_u1793_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u1794 (
    .a(_al_u1299_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 ),
    .o(_al_u1794_o));
  AL_MAP_LUT3 #(
    .EQN("~(~A*~(C*~B))"),
    .INIT(8'hba))
    _al_u1795 (
    .a(_al_u1793_o),
    .b(_al_u1794_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qakbx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rqthu6 ));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~((C*B))*~(A)+~D*(C*B)*~(A)+~(~D)*(C*B)*A+~D*(C*B)*A)"),
    .INIT(16'h7f2a))
    _al_u1796 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uzaiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B0biu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[0] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[1] ),
    .o(_al_u1796_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    _al_u1797 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n3685 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I8lax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vygax6 ),
    .o(_al_u1797_o));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*~B)*~(C*~A))"),
    .INIT(16'h7350))
    _al_u1798 (
    .a(_al_u1796_o),
    .b(_al_u1794_o),
    .c(_al_u1797_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Halax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z7vhu6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u1799 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ya1ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 ),
    .o(_al_u1799_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u1800 (
    .a(_al_u1799_o),
    .b(_al_u909_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nu9ow6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u1801 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nu9ow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 ),
    .o(_al_u1801_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u1802 (
    .a(_al_u1643_o),
    .b(_al_u1635_o),
    .o(_al_u1802_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u1803 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 ),
    .o(_al_u1803_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*~B*A)"),
    .INIT(16'h0020))
    _al_u1804 (
    .a(_al_u1803_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 ),
    .o(_al_u1804_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u1805 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yljiu6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u1806 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yljiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ),
    .o(_al_u1806_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u1807 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vo3ju6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(D*C*B))"),
    .INIT(16'h1555))
    _al_u1808 (
    .a(_al_u1804_o),
    .b(_al_u1806_o),
    .c(_al_u607_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vo3ju6_lutinv ),
    .o(_al_u1808_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u1809 (
    .a(_al_u1296_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pu1ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 ),
    .o(_al_u1809_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u1810 (
    .a(_al_u1808_o),
    .b(_al_u1809_o),
    .o(_al_u1810_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~B*~(D*A))"),
    .INIT(16'h1030))
    _al_u1811 (
    .a(_al_u1801_o),
    .b(_al_u1802_o),
    .c(_al_u1810_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wkipw6 ),
    .o(_al_u1811_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u1812 (
    .a(_al_u1385_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/SLEEPHOLDACKn ),
    .o(_al_u1812_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u1813 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 ),
    .o(_al_u1813_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u1814 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D6kiu6_lutinv ),
    .b(_al_u1813_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M8fax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uu9ow6_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u1815 (
    .a(_al_u1812_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uu9ow6_lutinv ),
    .o(_al_u1815_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u1816 (
    .a(_al_u903_o),
    .b(_al_u1582_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 ),
    .o(_al_u1816_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u1817 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 ),
    .o(_al_u1817_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u1818 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pu1ju6_lutinv ),
    .b(_al_u1817_o),
    .o(_al_u1818_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~A*~(D*C))"),
    .INIT(16'h0111))
    _al_u1819 (
    .a(_al_u1816_o),
    .b(_al_u1818_o),
    .c(_al_u604_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mfjiu6 ),
    .o(_al_u1819_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*A)"),
    .INIT(16'h0080))
    _al_u1820 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ldoiu6_lutinv ),
    .b(_al_u1658_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vo3ju6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 ),
    .o(_al_u1820_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(~D*C))"),
    .INIT(16'h4404))
    _al_u1821 (
    .a(_al_u1815_o),
    .b(_al_u1819_o),
    .c(_al_u1820_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ),
    .o(_al_u1821_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(B*A))"),
    .INIT(8'h07))
    _al_u1822 (
    .a(_al_u1811_o),
    .b(_al_u1821_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jy9iu6 ));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u1823 (
    .a(_al_u1675_o),
    .b(_al_u1676_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W6ipw6 ),
    .o(_al_u1823_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1824 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vk1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cl1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H3lpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kwlpw6 ),
    .o(_al_u1824_o));
  AL_MAP_LUT4 #(
    .EQN("~(B*A*~(D*C))"),
    .INIT(16'hf777))
    _al_u1825 (
    .a(_al_u1823_o),
    .b(_al_u1824_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xl1iu6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L5lpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zqxhu6 ));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u1826 (
    .a(_al_u1675_o),
    .b(_al_u1676_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Li7ax6 ),
    .o(_al_u1826_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1827 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vk1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cl1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A5ipw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L9bbx6 ),
    .o(_al_u1827_o));
  AL_MAP_LUT4 #(
    .EQN("~(B*A*~(D*C))"),
    .INIT(16'hf777))
    _al_u1828 (
    .a(_al_u1826_o),
    .b(_al_u1827_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xl1iu6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W6ipw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Grxhu6 ));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u1829 (
    .a(_al_u1675_o),
    .b(_al_u1676_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgfax6 ),
    .o(_al_u1829_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1830 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vk1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cl1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ceabx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I0opw6 ),
    .o(_al_u1830_o));
  AL_MAP_LUT4 #(
    .EQN("~(B*A*~(D*C))"),
    .INIT(16'hf777))
    _al_u1831 (
    .a(_al_u1829_o),
    .b(_al_u1830_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xl1iu6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D2opw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wsxhu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1832 (
    .a(\u_cmsdk_mcu/sram_hrdata [17]),
    .b(\u_cmsdk_mcu/flash_hrdata [17]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [0]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [1]),
    .o(_al_u1832_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(D*C))"),
    .INIT(16'h0444))
    _al_u1833 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n37 [14]),
    .b(_al_u1832_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [4]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/rwdata_reg [17]),
    .o(_al_u1833_o));
  AL_MAP_LUT4 #(
    .EQN("((~B*~A)*~(D)*~(C)+(~B*~A)*D*~(C)+~((~B*~A))*D*C+(~B*~A)*D*C)"),
    .INIT(16'hf101))
    _al_u1834 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wz4iu6 ),
    .b(_al_u1833_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qqhiu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tujbx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mbohu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1835 (
    .a(\u_cmsdk_mcu/sram_hrdata [18]),
    .b(\u_cmsdk_mcu/flash_hrdata [18]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [0]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [1]),
    .o(_al_u1835_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(D*C))"),
    .INIT(16'h0444))
    _al_u1836 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n37 [14]),
    .b(_al_u1835_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [4]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/rwdata_reg [18]),
    .o(_al_u1836_o));
  AL_MAP_LUT4 #(
    .EQN("((~B*~A)*~(D)*~(C)+(~B*~A)*D*~(C)+~((~B*~A))*D*C+(~B*~A)*D*C)"),
    .INIT(16'hf101))
    _al_u1837 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wz4iu6 ),
    .b(_al_u1836_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qqhiu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Usjbx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tbohu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1838 (
    .a(\u_cmsdk_mcu/sram_hrdata [19]),
    .b(\u_cmsdk_mcu/flash_hrdata [19]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [0]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [1]),
    .o(_al_u1838_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(D*C))"),
    .INIT(16'h0444))
    _al_u1839 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n37 [14]),
    .b(_al_u1838_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [4]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/rwdata_reg [19]),
    .o(_al_u1839_o));
  AL_MAP_LUT4 #(
    .EQN("((~B*~A)*~(D)*~(C)+(~B*~A)*D*~(C)+~((~B*~A))*D*C+(~B*~A)*D*C)"),
    .INIT(16'hf101))
    _al_u1840 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wz4iu6 ),
    .b(_al_u1839_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qqhiu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vqjbx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Acohu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1841 (
    .a(\u_cmsdk_mcu/sram_hrdata [20]),
    .b(\u_cmsdk_mcu/flash_hrdata [20]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [0]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [1]),
    .o(_al_u1841_o));
  AL_MAP_LUT4 #(
    .EQN("((~C*~A)*~(D)*~(B)+(~C*~A)*D*~(B)+~((~C*~A))*D*B+(~C*~A)*D*B)"),
    .INIT(16'hcd01))
    _al_u1842 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wz4iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qqhiu6 ),
    .c(_al_u1841_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tokax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eeohu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1843 (
    .a(\u_cmsdk_mcu/sram_hrdata [21]),
    .b(\u_cmsdk_mcu/flash_hrdata [21]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [0]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [1]),
    .o(_al_u1843_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~D*C*A))"),
    .INIT(16'hcc4c))
    _al_u1844 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n37 [1]),
    .b(_al_u1843_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/haddr_reg [0]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/haddr_reg [1]),
    .o(_al_u1844_o));
  AL_MAP_LUT4 #(
    .EQN("((~B*~A)*~(D)*~(C)+(~B*~A)*D*~(C)+~((~B*~A))*D*C+(~B*~A)*D*C)"),
    .INIT(16'hf101))
    _al_u1845 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wz4iu6 ),
    .b(_al_u1844_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qqhiu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kakax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Seohu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1846 (
    .a(\u_cmsdk_mcu/sram_hrdata [22]),
    .b(\u_cmsdk_mcu/flash_hrdata [22]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [0]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [1]),
    .o(_al_u1846_o));
  AL_MAP_LUT4 #(
    .EQN("((~C*~A)*~(D)*~(B)+(~C*~A)*D*~(B)+~((~C*~A))*D*B+(~C*~A)*D*B)"),
    .INIT(16'hcd01))
    _al_u1847 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wz4iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qqhiu6 ),
    .c(_al_u1846_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L8kax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zeohu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1848 (
    .a(\u_cmsdk_mcu/sram_hrdata [23]),
    .b(\u_cmsdk_mcu/flash_hrdata [23]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [0]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [1]),
    .o(_al_u1848_o));
  AL_MAP_LUT4 #(
    .EQN("((~C*~A)*~(D)*~(B)+(~C*~A)*D*~(B)+~((~C*~A))*D*B+(~C*~A)*D*B)"),
    .INIT(16'hcd01))
    _al_u1849 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wz4iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qqhiu6 ),
    .c(_al_u1848_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O2kax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nfohu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1850 (
    .a(\u_cmsdk_mcu/sram_hrdata [24]),
    .b(\u_cmsdk_mcu/flash_hrdata [24]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [0]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [1]),
    .o(_al_u1850_o));
  AL_MAP_LUT4 #(
    .EQN("((~C*~A)*~(D)*~(B)+(~C*~A)*D*~(B)+~((~C*~A))*D*B+(~C*~A)*D*B)"),
    .INIT(16'hcd01))
    _al_u1851 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wz4iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qqhiu6 ),
    .c(_al_u1850_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qyjax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufohu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1852 (
    .a(\u_cmsdk_mcu/sram_hrdata [25]),
    .b(\u_cmsdk_mcu/flash_hrdata [25]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [0]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [1]),
    .o(_al_u1852_o));
  AL_MAP_LUT4 #(
    .EQN("((~C*~A)*~(D)*~(B)+(~C*~A)*D*~(B)+~((~C*~A))*D*B+(~C*~A)*D*B)"),
    .INIT(16'hcd01))
    _al_u1853 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wz4iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qqhiu6 ),
    .c(_al_u1852_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sujax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bgohu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1854 (
    .a(\u_cmsdk_mcu/sram_hrdata [26]),
    .b(\u_cmsdk_mcu/flash_hrdata [26]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [0]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [1]),
    .o(_al_u1854_o));
  AL_MAP_LUT4 #(
    .EQN("((~C*~A)*~(D)*~(B)+(~C*~A)*D*~(B)+~((~C*~A))*D*B+(~C*~A)*D*B)"),
    .INIT(16'hcd01))
    _al_u1855 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wz4iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qqhiu6 ),
    .c(_al_u1854_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sqjax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Igohu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1856 (
    .a(\u_cmsdk_mcu/sram_hrdata [27]),
    .b(\u_cmsdk_mcu/flash_hrdata [27]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [0]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [1]),
    .o(_al_u1856_o));
  AL_MAP_LUT4 #(
    .EQN("((~C*~A)*~(D)*~(B)+(~C*~A)*D*~(B)+~((~C*~A))*D*B+(~C*~A)*D*B)"),
    .INIT(16'hcd01))
    _al_u1857 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wz4iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qqhiu6 ),
    .c(_al_u1856_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Smjax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pgohu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1858 (
    .a(\u_cmsdk_mcu/sram_hrdata [28]),
    .b(\u_cmsdk_mcu/flash_hrdata [28]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [0]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [1]),
    .o(_al_u1858_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(A*~(~D*C)))"),
    .INIT(16'h44c4))
    _al_u1859 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n37 [1]),
    .b(_al_u1858_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/haddr_reg [0]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/haddr_reg [1]),
    .o(_al_u1859_o));
  AL_MAP_LUT4 #(
    .EQN("((~B*~A)*~(D)*~(C)+(~B*~A)*D*~(C)+~((~B*~A))*D*C+(~B*~A)*D*C)"),
    .INIT(16'hf101))
    _al_u1860 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wz4iu6 ),
    .b(_al_u1859_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qqhiu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sijax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wgohu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1861 (
    .a(\u_cmsdk_mcu/sram_hrdata [29]),
    .b(\u_cmsdk_mcu/flash_hrdata [29]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [0]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [1]),
    .o(_al_u1861_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u1862 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n37 [14]),
    .b(_al_u1861_o),
    .o(_al_u1862_o));
  AL_MAP_LUT4 #(
    .EQN("((~B*~A)*~(D)*~(C)+(~B*~A)*D*~(C)+~((~B*~A))*D*C+(~B*~A)*D*C)"),
    .INIT(16'hf101))
    _al_u1863 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wz4iu6 ),
    .b(_al_u1862_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qqhiu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sgjax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dhohu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1864 (
    .a(\u_cmsdk_mcu/sram_hrdata [31]),
    .b(\u_cmsdk_mcu/flash_hrdata [31]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [0]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [1]),
    .o(_al_u1864_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u1865 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n37 [14]),
    .b(_al_u1864_o),
    .o(_al_u1865_o));
  AL_MAP_LUT4 #(
    .EQN("((~B*~A)*~(D)*~(C)+(~B*~A)*D*~(C)+~((~B*~A))*D*C+(~B*~A)*D*C)"),
    .INIT(16'hf101))
    _al_u1866 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wz4iu6 ),
    .b(_al_u1865_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qqhiu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sejax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Khohu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1867 (
    .a(\u_cmsdk_mcu/sram_hrdata [16]),
    .b(\u_cmsdk_mcu/flash_hrdata [16]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [0]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [1]),
    .o(_al_u1867_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(D*C))"),
    .INIT(16'h0444))
    _al_u1868 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n37 [14]),
    .b(_al_u1867_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [4]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/rwdata_reg [16]),
    .o(_al_u1868_o));
  AL_MAP_LUT4 #(
    .EQN("((~B*~A)*~(D)*~(C)+(~B*~A)*D*~(C)+~((~B*~A))*D*C+(~B*~A)*D*C)"),
    .INIT(16'hf101))
    _al_u1869 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wz4iu6 ),
    .b(_al_u1868_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qqhiu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tcjax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rhohu6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u1870 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Htmpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vmipw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aq2pw6_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u1871 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aq2pw6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iixpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vhspw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hhqow6 ));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*~A)"),
    .INIT(16'h4000))
    _al_u1872 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Htmpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iixpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vhspw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vmipw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljqow6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1873 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hhqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[0] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[0] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jy2pw6 ));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*~A)"),
    .INIT(16'h1000))
    _al_u1874 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Htmpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iixpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vhspw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vmipw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qiqow6 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u1875 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jy2pw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qiqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[0] ),
    .o(_al_u1875_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u1876 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aq2pw6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iixpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vhspw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dfqow6 ));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u1877 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aq2pw6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iixpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vhspw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahqow6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1878 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dfqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I1lpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[0] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qy2pw6 ));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*~A)"),
    .INIT(16'h0100))
    _al_u1879 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Htmpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iixpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vhspw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vmipw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gkqow6 ));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*B*~A)"),
    .INIT(16'h0400))
    _al_u1880 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Htmpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iixpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vhspw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vmipw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sjqow6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1881 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gkqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sjqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[0] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[0] ),
    .o(_al_u1881_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u1882 (
    .a(_al_u1875_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N30iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qy2pw6 ),
    .d(_al_u1881_o),
    .o(_al_u1882_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*~A)"),
    .INIT(8'h04))
    _al_u1883 (
    .a(_al_u1882_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I8lax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wvgax6 ),
    .o(_al_u1883_o));
  AL_MAP_LUT3 #(
    .EQN("~(~A*~(C*B))"),
    .INIT(8'hea))
    _al_u1884 (
    .a(_al_u1883_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T24iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wvgax6 ),
    .o(\u_cmsdk_mcu/HWDATA [0]));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*~B))"),
    .INIT(8'h54))
    _al_u1885 (
    .a(_al_u914_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 ),
    .o(_al_u1885_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u1886 (
    .a(_al_u1885_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sq3ju6 ),
    .c(_al_u1296_o),
    .o(_al_u1886_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u1887 (
    .a(_al_u1658_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 ),
    .o(_al_u1887_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u1888 (
    .a(_al_u1886_o),
    .b(_al_u1887_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ),
    .o(_al_u1888_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u1889 (
    .a(_al_u604_o),
    .b(_al_u678_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Frziu6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qk9pw6_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u1890 (
    .a(_al_u1888_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qk9pw6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J71iu6_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u1891 (
    .a(_al_u1883_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J71iu6_lutinv ),
    .o(_al_u1891_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(B*A))"),
    .INIT(8'h07))
    _al_u1892 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J71iu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I8lax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wvgax6 ),
    .o(_al_u1892_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1893 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qiqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sjqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[8] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[8] ),
    .o(_al_u1893_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u1894 (
    .a(_al_u1893_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gkqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[8] ),
    .o(_al_u1894_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1895 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hhqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dfqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[8] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N61qw6 ),
    .o(_al_u1895_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1896 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[8] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[8] ),
    .o(_al_u1896_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*A)"),
    .INIT(16'h0200))
    _al_u1897 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aq2pw6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iixpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jrypw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vhspw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fgqow6 ));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u1898 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aq2pw6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iixpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jrypw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vhspw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yfqow6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1899 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fgqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yfqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[6] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[6] ),
    .o(_al_u1899_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u1900 (
    .a(_al_u1894_o),
    .b(_al_u1895_o),
    .c(_al_u1896_o),
    .d(_al_u1899_o),
    .o(_al_u1900_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u1901 (
    .a(_al_u1900_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lvzhu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cz7ju6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u1902 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pl4iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wvgax6 ),
    .o(_al_u1902_o));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~A*~(~C*B))"),
    .INIT(16'hffae))
    _al_u1903 (
    .a(_al_u1891_o),
    .b(_al_u1892_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cz7ju6 ),
    .d(_al_u1902_o),
    .o(\u_cmsdk_mcu/HWDATA [8]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u1904 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Llaow6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Obbow6_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u1905 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mfjiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ),
    .o(_al_u1905_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(~D*C*A))"),
    .INIT(16'h3313))
    _al_u1906 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Obbow6_lutinv ),
    .b(_al_u1905_o),
    .c(_al_u607_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 ),
    .o(_al_u1906_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u1907 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 ),
    .o(_al_u1907_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u1908 (
    .a(_al_u681_o),
    .b(_al_u1907_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Stuow6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*C)*~(~B*~A))"),
    .INIT(16'hf111))
    _al_u1909 (
    .a(_al_u1882_o),
    .b(_al_u1906_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Stuow6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iixpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oy8iu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1910 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qiqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[2] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[2] ),
    .o(_al_u1910_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u1911 (
    .a(_al_u1910_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sjqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[2] ),
    .o(_al_u1911_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1912 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dfqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gkqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[2] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xrxax6 ),
    .o(_al_u1912_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1913 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hhqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[2] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[2] ),
    .o(_al_u1913_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1914 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fgqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yfqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[0] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[0] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ro2pw6 ));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u1915 (
    .a(_al_u1911_o),
    .b(_al_u1912_o),
    .c(_al_u1913_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ro2pw6 ),
    .o(_al_u1915_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u1916 (
    .a(_al_u1915_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pxzhu6 ),
    .o(_al_u1916_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*~A)"),
    .INIT(8'h04))
    _al_u1917 (
    .a(_al_u1916_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I8lax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wvgax6 ),
    .o(_al_u1917_o));
  AL_MAP_LUT3 #(
    .EQN("~(~A*~(C*B))"),
    .INIT(8'hea))
    _al_u1918 (
    .a(_al_u1917_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ud4iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wvgax6 ),
    .o(\u_cmsdk_mcu/HWDATA [2]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1919 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hhqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dfqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[3] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T5yax6 ),
    .o(_al_u1919_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u1920 (
    .a(_al_u1919_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qiqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[3] ),
    .o(_al_u1920_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1921 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[3] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[3] ),
    .o(_al_u1921_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1922 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fgqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yfqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[1] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[1] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X62pw6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1923 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gkqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sjqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[3] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[3] ),
    .o(_al_u1923_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u1924 (
    .a(_al_u1920_o),
    .b(_al_u1921_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X62pw6 ),
    .d(_al_u1923_o),
    .o(_al_u1924_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u1925 (
    .a(_al_u1924_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uwzhu6 ),
    .o(_al_u1925_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*~A)"),
    .INIT(8'h04))
    _al_u1926 (
    .a(_al_u1925_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I8lax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wvgax6 ),
    .o(_al_u1926_o));
  AL_MAP_LUT3 #(
    .EQN("~(~A*~(C*B))"),
    .INIT(8'hea))
    _al_u1927 (
    .a(_al_u1926_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Df4iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wvgax6 ),
    .o(\u_cmsdk_mcu/HWDATA [3]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1928 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hhqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dfqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[4] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wtxax6 ),
    .o(_al_u1928_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u1929 (
    .a(_al_u1928_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qiqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[4] ),
    .o(_al_u1929_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1930 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sjqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[4] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[4] ),
    .o(_al_u1930_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1931 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fgqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yfqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[2] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[2] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kp1pw6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1932 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gkqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[4] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[4] ),
    .o(_al_u1932_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u1933 (
    .a(_al_u1929_o),
    .b(_al_u1930_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kp1pw6 ),
    .d(_al_u1932_o),
    .o(_al_u1933_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u1934 (
    .a(_al_u1933_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nwzhu6 ),
    .o(_al_u1934_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*~A)"),
    .INIT(8'h04))
    _al_u1935 (
    .a(_al_u1934_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I8lax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wvgax6 ),
    .o(_al_u1935_o));
  AL_MAP_LUT3 #(
    .EQN("~(~A*~(C*B))"),
    .INIT(8'hea))
    _al_u1936 (
    .a(_al_u1935_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H34iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wvgax6 ),
    .o(\u_cmsdk_mcu/HWDATA [4]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1937 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hhqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qiqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[5] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[5] ),
    .o(_al_u1937_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u1938 (
    .a(_al_u1937_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dfqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qc5bx6 ),
    .o(_al_u1938_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1939 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sjqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[5] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[5] ),
    .o(_al_u1939_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1940 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fgqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yfqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[3] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[3] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X71pw6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1941 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gkqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[5] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[5] ),
    .o(_al_u1941_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u1942 (
    .a(_al_u1938_o),
    .b(_al_u1939_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X71pw6 ),
    .d(_al_u1941_o),
    .o(_al_u1942_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u1943 (
    .a(_al_u1942_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gwzhu6 ),
    .o(_al_u1943_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*~A)"),
    .INIT(8'h04))
    _al_u1944 (
    .a(_al_u1943_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I8lax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wvgax6 ),
    .o(_al_u1944_o));
  AL_MAP_LUT3 #(
    .EQN("~(~A*~(C*B))"),
    .INIT(8'hea))
    _al_u1945 (
    .a(_al_u1944_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oh4iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wvgax6 ),
    .o(\u_cmsdk_mcu/HWDATA [5]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1946 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hhqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qiqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[6] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[6] ),
    .o(_al_u1946_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u1947 (
    .a(_al_u1946_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sjqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[6] ),
    .o(_al_u1947_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1948 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dfqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[6] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ua9bx6 ),
    .o(_al_u1948_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1949 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fgqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yfqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[4] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[4] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kq0pw6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1950 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gkqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[6] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[6] ),
    .o(_al_u1950_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u1951 (
    .a(_al_u1947_o),
    .b(_al_u1948_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kq0pw6 ),
    .d(_al_u1950_o),
    .o(_al_u1951_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u1952 (
    .a(_al_u1951_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zvzhu6 ),
    .o(_al_u1952_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*~A)"),
    .INIT(8'h04))
    _al_u1953 (
    .a(_al_u1952_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I8lax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wvgax6 ),
    .o(_al_u1953_o));
  AL_MAP_LUT3 #(
    .EQN("~(~A*~(C*B))"),
    .INIT(8'hea))
    _al_u1954 (
    .a(_al_u1953_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xi4iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wvgax6 ),
    .o(\u_cmsdk_mcu/HWDATA [6]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1955 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hhqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qiqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[7] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[7] ),
    .o(_al_u1955_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u1956 (
    .a(_al_u1955_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dfqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Asupw6 ),
    .o(_al_u1956_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1957 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[7] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[7] ),
    .o(_al_u1957_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1958 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fgqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yfqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[5] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[5] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X80pw6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1959 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gkqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sjqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[7] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[7] ),
    .o(_al_u1959_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u1960 (
    .a(_al_u1956_o),
    .b(_al_u1957_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X80pw6 ),
    .d(_al_u1959_o),
    .o(_al_u1960_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u1961 (
    .a(_al_u1960_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Svzhu6 ),
    .o(_al_u1961_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*~A)"),
    .INIT(8'h04))
    _al_u1962 (
    .a(_al_u1961_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I8lax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wvgax6 ),
    .o(_al_u1962_o));
  AL_MAP_LUT3 #(
    .EQN("~(~A*~(C*B))"),
    .INIT(8'hea))
    _al_u1963 (
    .a(_al_u1962_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gk4iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wvgax6 ),
    .o(\u_cmsdk_mcu/HWDATA [7]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1964 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dfqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gkqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nu5bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[1] ),
    .o(_al_u1964_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u1965 (
    .a(_al_u1964_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qiqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[1] ),
    .o(_al_u1965_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1966 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hhqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sjqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[1] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[1] ),
    .o(_al_u1966_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1967 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[1] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[1] ),
    .o(_al_u1967_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u1968 (
    .a(_al_u1965_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O00iu6 ),
    .c(_al_u1966_o),
    .d(_al_u1967_o),
    .o(_al_u1968_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*~A)"),
    .INIT(8'h04))
    _al_u1969 (
    .a(_al_u1968_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I8lax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wvgax6 ),
    .o(_al_u1969_o));
  AL_MAP_LUT3 #(
    .EQN("~(~A*~(C*B))"),
    .INIT(8'hea))
    _al_u1970 (
    .a(_al_u1969_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O34iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wvgax6 ),
    .o(\u_cmsdk_mcu/HWDATA [1]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u1971 (
    .a(_al_u1969_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J71iu6_lutinv ),
    .o(_al_u1971_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1972 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dfqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qiqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[9] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kn1qw6 ),
    .o(_al_u1972_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u1973 (
    .a(_al_u1972_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gkqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[9] ),
    .o(_al_u1973_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1974 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hhqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[9] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[9] ),
    .o(_al_u1974_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u1975 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fgqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yfqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[7] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[7] ),
    .o(_al_u1975_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1976 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sjqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[9] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[9] ),
    .o(_al_u1976_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u1977 (
    .a(_al_u1973_o),
    .b(_al_u1974_o),
    .c(_al_u1975_o),
    .d(_al_u1976_o),
    .o(_al_u1977_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u1978 (
    .a(_al_u1977_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Evzhu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I28ju6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u1979 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ym4iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wvgax6 ),
    .o(_al_u1979_o));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~A*~(~C*B))"),
    .INIT(16'hffae))
    _al_u1980 (
    .a(_al_u1971_o),
    .b(_al_u1892_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I28ju6 ),
    .d(_al_u1979_o),
    .o(\u_cmsdk_mcu/HWDATA [9]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u1981 (
    .a(_al_u581_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [6]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/mux4_b10_sel_is_4_o ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u1982 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [5]),
    .o(_al_u1982_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u1983 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/mux4_b10_sel_is_4_o ),
    .b(_al_u1982_o),
    .o(_al_u1983_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    _al_u1984 (
    .a(_al_u1983_o),
    .b(_al_u588_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n223 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u1985 (
    .a(\u_cmsdk_mcu/HWDATA [0]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n223 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpolset [0]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u1986 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [5]),
    .o(_al_u1986_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u1987 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/mux4_b10_sel_is_4_o ),
    .b(_al_u1986_o),
    .o(_al_u1987_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u1988 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .o(_al_u1988_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u1989 (
    .a(_al_u1987_o),
    .b(_al_u588_o),
    .c(_al_u1988_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n178 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u1990 (
    .a(\u_cmsdk_mcu/HWDATA [0]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n178 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttypeset [0]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    _al_u1991 (
    .a(_al_u1987_o),
    .b(_al_u588_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n133 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u1992 (
    .a(\u_cmsdk_mcu/HWDATA [0]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n133 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intenset [0]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    _al_u1993 (
    .a(_al_u581_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [5]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [6]),
    .o(_al_u1993_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u1994 (
    .a(_al_u1993_o),
    .b(_al_u588_o),
    .c(_al_u1988_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n88 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u1995 (
    .a(\u_cmsdk_mcu/HWDATA [0]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n88 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_altfuncset [0]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    _al_u1996 (
    .a(_al_u1993_o),
    .b(_al_u588_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n43 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u1997 (
    .a(\u_cmsdk_mcu/HWDATA [0]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n43 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_doutenset [0]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    _al_u1998 (
    .a(_al_u1983_o),
    .b(_al_u593_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n223 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u1999 (
    .a(\u_cmsdk_mcu/HWDATA [0]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n223 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpolset [0]));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u2000 (
    .a(_al_u1987_o),
    .b(_al_u593_o),
    .c(_al_u1988_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n178 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2001 (
    .a(\u_cmsdk_mcu/HWDATA [0]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n178 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttypeset [0]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    _al_u2002 (
    .a(_al_u1987_o),
    .b(_al_u593_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n133 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2003 (
    .a(\u_cmsdk_mcu/HWDATA [0]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n133 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intenset [0]));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u2004 (
    .a(_al_u1993_o),
    .b(_al_u593_o),
    .c(_al_u1988_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n88 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2005 (
    .a(\u_cmsdk_mcu/HWDATA [0]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n88 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_altfuncset [0]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    _al_u2006 (
    .a(_al_u1993_o),
    .b(_al_u593_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n43 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2007 (
    .a(\u_cmsdk_mcu/HWDATA [0]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n43 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_doutenset [0]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u2008 (
    .a(\u_cmsdk_mcu/HWDATA [0]),
    .b(\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [0]),
    .c(\u_cmsdk_mcu/flash_hrdata [0]),
    .o(\u_cmsdk_mcu/u_ahb_rom/n13 [0]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2009 (
    .a(\u_cmsdk_mcu/HWDATA [0]),
    .b(\u_cmsdk_mcu/sram_hrdata [0]),
    .c(\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [0]),
    .o(\u_cmsdk_mcu/u_ahb_ram/n13 [0]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    _al_u2010 (
    .a(_al_u1983_o),
    .b(_al_u585_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n226 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2011 (
    .a(\u_cmsdk_mcu/HWDATA [8]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n226 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpolset [8]));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u2012 (
    .a(_al_u1987_o),
    .b(_al_u585_o),
    .c(_al_u1988_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n181 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2013 (
    .a(\u_cmsdk_mcu/HWDATA [8]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n181 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttypeset [8]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    _al_u2014 (
    .a(_al_u1987_o),
    .b(_al_u585_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n136 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2015 (
    .a(\u_cmsdk_mcu/HWDATA [8]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n136 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intenset [8]));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u2016 (
    .a(_al_u1993_o),
    .b(_al_u585_o),
    .c(_al_u1988_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n91 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2017 (
    .a(\u_cmsdk_mcu/HWDATA [8]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n91 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_altfuncset [8]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    _al_u2018 (
    .a(_al_u1993_o),
    .b(_al_u585_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n46 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2019 (
    .a(\u_cmsdk_mcu/HWDATA [8]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n46 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_doutenset [8]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    _al_u2020 (
    .a(_al_u1983_o),
    .b(_al_u591_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n226 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2021 (
    .a(\u_cmsdk_mcu/HWDATA [8]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n226 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpolset [8]));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u2022 (
    .a(_al_u1987_o),
    .b(_al_u591_o),
    .c(_al_u1988_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n181 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2023 (
    .a(\u_cmsdk_mcu/HWDATA [8]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n181 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttypeset [8]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    _al_u2024 (
    .a(_al_u1987_o),
    .b(_al_u591_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n136 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2025 (
    .a(\u_cmsdk_mcu/HWDATA [8]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n136 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intenset [8]));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u2026 (
    .a(_al_u1993_o),
    .b(_al_u591_o),
    .c(_al_u1988_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n91 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2027 (
    .a(\u_cmsdk_mcu/HWDATA [8]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n91 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_altfuncset [8]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    _al_u2028 (
    .a(_al_u1993_o),
    .b(_al_u591_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n46 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2029 (
    .a(\u_cmsdk_mcu/HWDATA [8]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n46 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_doutenset [8]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u2030 (
    .a(\u_cmsdk_mcu/HWDATA [8]),
    .b(\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [10]),
    .c(\u_cmsdk_mcu/flash_hrdata [8]),
    .o(\u_cmsdk_mcu/u_ahb_rom/n13 [8]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2031 (
    .a(\u_cmsdk_mcu/HWDATA [8]),
    .b(\u_cmsdk_mcu/sram_hrdata [8]),
    .c(\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [10]),
    .o(\u_cmsdk_mcu/u_ahb_ram/n13 [8]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2032 (
    .a(_al_u1917_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J71iu6_lutinv ),
    .o(_al_u2032_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u2033 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sjqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[10] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[10] ),
    .o(_al_u2033_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u2034 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dfqow6 ),
    .b(_al_u2033_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gwxpw6 ),
    .o(_al_u2034_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u2035 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hhqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qiqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[10] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[10] ),
    .o(_al_u2035_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u2036 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gkqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[10] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[10] ),
    .o(_al_u2036_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u2037 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fgqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yfqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[8] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[8] ),
    .o(_al_u2037_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u2038 (
    .a(_al_u2034_o),
    .b(_al_u2035_o),
    .c(_al_u2036_o),
    .d(_al_u2037_o),
    .o(_al_u2038_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2039 (
    .a(_al_u2038_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G30iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ka8ju6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2040 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J44iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wvgax6 ),
    .o(_al_u2040_o));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~A*~(~C*B))"),
    .INIT(16'hffae))
    _al_u2041 (
    .a(_al_u2032_o),
    .b(_al_u1892_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ka8ju6 ),
    .d(_al_u2040_o),
    .o(\u_cmsdk_mcu/HWDATA [10]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2042 (
    .a(\u_cmsdk_mcu/HWDATA [2]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C1wpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G3eiu6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2043 (
    .a(\u_cmsdk_mcu/HWDATA [2]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n223 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpolset [2]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2044 (
    .a(\u_cmsdk_mcu/HWDATA [2]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n178 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttypeset [2]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2045 (
    .a(\u_cmsdk_mcu/HWDATA [2]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n133 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intenset [2]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2046 (
    .a(\u_cmsdk_mcu/HWDATA [2]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n88 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_altfuncset [2]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2047 (
    .a(\u_cmsdk_mcu/HWDATA [2]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n43 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_doutenset [2]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2048 (
    .a(\u_cmsdk_mcu/HWDATA [2]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n223 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpolset [2]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2049 (
    .a(\u_cmsdk_mcu/HWDATA [2]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n178 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttypeset [2]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2050 (
    .a(\u_cmsdk_mcu/HWDATA [2]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n133 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intenset [2]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2051 (
    .a(\u_cmsdk_mcu/HWDATA [2]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n88 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_altfuncset [2]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2052 (
    .a(\u_cmsdk_mcu/HWDATA [2]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n43 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_doutenset [2]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u2053 (
    .a(\u_cmsdk_mcu/HWDATA [2]),
    .b(\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [0]),
    .c(\u_cmsdk_mcu/flash_hrdata [2]),
    .o(\u_cmsdk_mcu/u_ahb_rom/n13 [2]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2054 (
    .a(\u_cmsdk_mcu/HWDATA [2]),
    .b(\u_cmsdk_mcu/sram_hrdata [2]),
    .c(\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [0]),
    .o(\u_cmsdk_mcu/u_ahb_ram/n13 [2]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2055 (
    .a(_al_u1926_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J71iu6_lutinv ),
    .o(_al_u2055_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u2056 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sjqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[11] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[11] ),
    .o(_al_u2056_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u2057 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hhqow6 ),
    .b(_al_u2056_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[11] ),
    .o(_al_u2057_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u2058 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dfqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qiqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C07bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[11] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hy1pw6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u2059 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gkqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[11] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[11] ),
    .o(_al_u2059_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u2060 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fgqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yfqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[9] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[9] ),
    .o(_al_u2060_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u2061 (
    .a(_al_u2057_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hy1pw6 ),
    .c(_al_u2059_o),
    .d(_al_u2060_o),
    .o(_al_u2061_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2062 (
    .a(_al_u2061_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z20iu6 ),
    .o(_al_u2062_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2063 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q44iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wvgax6 ),
    .o(_al_u2063_o));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~A*~(~C*B))"),
    .INIT(16'hffae))
    _al_u2064 (
    .a(_al_u2055_o),
    .b(_al_u1892_o),
    .c(_al_u2062_o),
    .d(_al_u2063_o),
    .o(\u_cmsdk_mcu/HWDATA [11]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2065 (
    .a(\u_cmsdk_mcu/HWDATA [3]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n223 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpolset [3]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2066 (
    .a(\u_cmsdk_mcu/HWDATA [3]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n178 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttypeset [3]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2067 (
    .a(\u_cmsdk_mcu/HWDATA [3]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n133 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intenset [3]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2068 (
    .a(\u_cmsdk_mcu/HWDATA [3]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n88 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_altfuncset [3]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2069 (
    .a(\u_cmsdk_mcu/HWDATA [3]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n43 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_doutenset [3]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2070 (
    .a(\u_cmsdk_mcu/HWDATA [3]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n223 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpolset [3]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2071 (
    .a(\u_cmsdk_mcu/HWDATA [3]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n178 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttypeset [3]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2072 (
    .a(\u_cmsdk_mcu/HWDATA [3]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n133 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intenset [3]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2073 (
    .a(\u_cmsdk_mcu/HWDATA [3]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n88 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_altfuncset [3]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2074 (
    .a(\u_cmsdk_mcu/HWDATA [3]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n43 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_doutenset [3]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u2075 (
    .a(\u_cmsdk_mcu/HWDATA [3]),
    .b(\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [0]),
    .c(\u_cmsdk_mcu/flash_hrdata [3]),
    .o(\u_cmsdk_mcu/u_ahb_rom/n13 [3]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2076 (
    .a(\u_cmsdk_mcu/HWDATA [3]),
    .b(\u_cmsdk_mcu/sram_hrdata [3]),
    .c(\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [0]),
    .o(\u_cmsdk_mcu/u_ahb_ram/n13 [3]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2077 (
    .a(_al_u1935_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J71iu6_lutinv ),
    .o(_al_u2077_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u2078 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dfqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qiqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dm6bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[12] ),
    .o(_al_u2078_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u2079 (
    .a(_al_u2078_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gkqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[12] ),
    .o(_al_u2079_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u2080 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hhqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[12] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[12] ),
    .o(_al_u2080_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u2081 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fgqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yfqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[10] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[10] ),
    .o(_al_u2081_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u2082 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sjqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[12] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[12] ),
    .o(_al_u2082_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u2083 (
    .a(_al_u2079_o),
    .b(_al_u2080_o),
    .c(_al_u2081_o),
    .d(_al_u2082_o),
    .o(_al_u2083_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2084 (
    .a(_al_u2083_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S20iu6 ),
    .o(_al_u2084_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2085 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X44iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wvgax6 ),
    .o(_al_u2085_o));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~A*~(~C*B))"),
    .INIT(16'hffae))
    _al_u2086 (
    .a(_al_u2077_o),
    .b(_al_u1892_o),
    .c(_al_u2084_o),
    .d(_al_u2085_o),
    .o(\u_cmsdk_mcu/HWDATA [12]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2087 (
    .a(\u_cmsdk_mcu/HWDATA [4]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n223 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpolset [4]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2088 (
    .a(\u_cmsdk_mcu/HWDATA [4]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n178 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttypeset [4]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2089 (
    .a(\u_cmsdk_mcu/HWDATA [4]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n133 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intenset [4]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2090 (
    .a(\u_cmsdk_mcu/HWDATA [4]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n88 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_altfuncset [4]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2091 (
    .a(\u_cmsdk_mcu/HWDATA [4]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n43 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_doutenset [4]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2092 (
    .a(\u_cmsdk_mcu/HWDATA [4]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n223 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpolset [4]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2093 (
    .a(\u_cmsdk_mcu/HWDATA [4]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n178 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttypeset [4]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2094 (
    .a(\u_cmsdk_mcu/HWDATA [4]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n133 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intenset [4]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2095 (
    .a(\u_cmsdk_mcu/HWDATA [4]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n88 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_altfuncset [4]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2096 (
    .a(\u_cmsdk_mcu/HWDATA [4]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n43 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_doutenset [4]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u2097 (
    .a(\u_cmsdk_mcu/HWDATA [4]),
    .b(\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [0]),
    .c(\u_cmsdk_mcu/flash_hrdata [4]),
    .o(\u_cmsdk_mcu/u_ahb_rom/n13 [4]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2098 (
    .a(\u_cmsdk_mcu/HWDATA [4]),
    .b(\u_cmsdk_mcu/sram_hrdata [4]),
    .c(\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [0]),
    .o(\u_cmsdk_mcu/u_ahb_ram/n13 [4]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2099 (
    .a(_al_u1944_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J71iu6_lutinv ),
    .o(_al_u2099_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u2100 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hhqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qiqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[13] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[13] ),
    .o(_al_u2100_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u2101 (
    .a(_al_u2100_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[13] ),
    .o(_al_u2101_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u2102 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dfqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[13] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xpxax6 ),
    .o(_al_u2102_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u2103 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fgqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yfqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[11] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[11] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hz0pw6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u2104 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gkqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sjqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[13] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[13] ),
    .o(_al_u2104_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u2105 (
    .a(_al_u2101_o),
    .b(_al_u2102_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hz0pw6 ),
    .d(_al_u2104_o),
    .o(_al_u2105_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2106 (
    .a(_al_u2105_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L20iu6 ),
    .o(_al_u2106_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2107 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E54iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wvgax6 ),
    .o(_al_u2107_o));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~A*~(~C*B))"),
    .INIT(16'hffae))
    _al_u2108 (
    .a(_al_u2099_o),
    .b(_al_u1892_o),
    .c(_al_u2106_o),
    .d(_al_u2107_o),
    .o(\u_cmsdk_mcu/HWDATA [13]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2109 (
    .a(\u_cmsdk_mcu/HWDATA [5]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n223 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpolset [5]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2110 (
    .a(\u_cmsdk_mcu/HWDATA [5]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n178 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttypeset [5]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2111 (
    .a(\u_cmsdk_mcu/HWDATA [5]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n133 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intenset [5]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2112 (
    .a(\u_cmsdk_mcu/HWDATA [5]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n88 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_altfuncset [5]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2113 (
    .a(\u_cmsdk_mcu/HWDATA [5]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n43 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_doutenset [5]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2114 (
    .a(\u_cmsdk_mcu/HWDATA [5]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n223 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpolset [5]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2115 (
    .a(\u_cmsdk_mcu/HWDATA [5]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n178 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttypeset [5]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2116 (
    .a(\u_cmsdk_mcu/HWDATA [5]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n133 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intenset [5]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2117 (
    .a(\u_cmsdk_mcu/HWDATA [5]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n88 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_altfuncset [5]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2118 (
    .a(\u_cmsdk_mcu/HWDATA [5]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n43 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_doutenset [5]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u2119 (
    .a(\u_cmsdk_mcu/HWDATA [5]),
    .b(\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [0]),
    .c(\u_cmsdk_mcu/flash_hrdata [5]),
    .o(\u_cmsdk_mcu/u_ahb_rom/n13 [5]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2120 (
    .a(\u_cmsdk_mcu/HWDATA [5]),
    .b(\u_cmsdk_mcu/sram_hrdata [5]),
    .c(\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [0]),
    .o(\u_cmsdk_mcu/u_ahb_ram/n13 [5]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2121 (
    .a(_al_u1953_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J71iu6_lutinv ),
    .o(_al_u2121_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u2122 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qiqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sjqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[14] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[14] ),
    .o(_al_u2122_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u2123 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hhqow6 ),
    .b(_al_u2122_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[14] ),
    .o(_al_u2123_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u2124 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dfqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gkqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[14] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sb8ax6 ),
    .o(_al_u2124_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u2125 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[14] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[14] ),
    .o(_al_u2125_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u2126 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fgqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yfqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[12] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[12] ),
    .o(_al_u2126_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u2127 (
    .a(_al_u2123_o),
    .b(_al_u2124_o),
    .c(_al_u2125_o),
    .d(_al_u2126_o),
    .o(_al_u2127_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2128 (
    .a(_al_u2127_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E20iu6 ),
    .o(_al_u2128_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2129 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L54iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wvgax6 ),
    .o(_al_u2129_o));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~A*~(~C*B))"),
    .INIT(16'hffae))
    _al_u2130 (
    .a(_al_u2121_o),
    .b(_al_u1892_o),
    .c(_al_u2128_o),
    .d(_al_u2129_o),
    .o(\u_cmsdk_mcu/HWDATA [14]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2131 (
    .a(\u_cmsdk_mcu/HWDATA [6]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n223 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpolset [6]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2132 (
    .a(\u_cmsdk_mcu/HWDATA [6]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n178 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttypeset [6]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2133 (
    .a(\u_cmsdk_mcu/HWDATA [6]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n133 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intenset [6]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2134 (
    .a(\u_cmsdk_mcu/HWDATA [6]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n88 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_altfuncset [6]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2135 (
    .a(\u_cmsdk_mcu/HWDATA [6]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n43 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_doutenset [6]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2136 (
    .a(\u_cmsdk_mcu/HWDATA [6]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n223 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpolset [6]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2137 (
    .a(\u_cmsdk_mcu/HWDATA [6]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n178 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttypeset [6]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2138 (
    .a(\u_cmsdk_mcu/HWDATA [6]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n133 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intenset [6]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2139 (
    .a(\u_cmsdk_mcu/HWDATA [6]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n88 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_altfuncset [6]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2140 (
    .a(\u_cmsdk_mcu/HWDATA [6]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n43 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_doutenset [6]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u2141 (
    .a(\u_cmsdk_mcu/HWDATA [6]),
    .b(\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [0]),
    .c(\u_cmsdk_mcu/flash_hrdata [6]),
    .o(\u_cmsdk_mcu/u_ahb_rom/n13 [6]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2142 (
    .a(\u_cmsdk_mcu/HWDATA [6]),
    .b(\u_cmsdk_mcu/sram_hrdata [6]),
    .c(\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [0]),
    .o(\u_cmsdk_mcu/u_ahb_ram/n13 [6]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2143 (
    .a(_al_u1962_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J71iu6_lutinv ),
    .o(_al_u2143_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u2144 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hhqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dfqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z47ax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[15] ),
    .o(_al_u2144_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u2145 (
    .a(_al_u2144_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qiqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[15] ),
    .o(_al_u2145_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u2146 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sjqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[15] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[15] ),
    .o(_al_u2146_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u2147 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fgqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yfqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[13] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[13] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H00pw6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u2148 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gkqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[15] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[15] ),
    .o(_al_u2148_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u2149 (
    .a(_al_u2145_o),
    .b(_al_u2146_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H00pw6 ),
    .d(_al_u2148_o),
    .o(_al_u2149_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2150 (
    .a(_al_u2149_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X10iu6 ),
    .o(_al_u2150_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2151 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S54iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wvgax6 ),
    .o(_al_u2151_o));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~A*~(~C*B))"),
    .INIT(16'hffae))
    _al_u2152 (
    .a(_al_u2143_o),
    .b(_al_u1892_o),
    .c(_al_u2150_o),
    .d(_al_u2151_o),
    .o(\u_cmsdk_mcu/HWDATA [15]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2153 (
    .a(\u_cmsdk_mcu/HWDATA [7]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n223 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpolset [7]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2154 (
    .a(\u_cmsdk_mcu/HWDATA [7]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n178 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttypeset [7]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2155 (
    .a(\u_cmsdk_mcu/HWDATA [7]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n133 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intenset [7]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2156 (
    .a(\u_cmsdk_mcu/HWDATA [7]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n88 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_altfuncset [7]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2157 (
    .a(\u_cmsdk_mcu/HWDATA [7]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n43 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_doutenset [7]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2158 (
    .a(\u_cmsdk_mcu/HWDATA [7]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n223 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpolset [7]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2159 (
    .a(\u_cmsdk_mcu/HWDATA [7]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n178 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttypeset [7]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2160 (
    .a(\u_cmsdk_mcu/HWDATA [7]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n133 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intenset [7]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2161 (
    .a(\u_cmsdk_mcu/HWDATA [7]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n88 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_altfuncset [7]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2162 (
    .a(\u_cmsdk_mcu/HWDATA [7]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n43 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_doutenset [7]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u2163 (
    .a(\u_cmsdk_mcu/HWDATA [7]),
    .b(\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [0]),
    .c(\u_cmsdk_mcu/flash_hrdata [7]),
    .o(\u_cmsdk_mcu/u_ahb_rom/n13 [7]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2164 (
    .a(\u_cmsdk_mcu/HWDATA [7]),
    .b(\u_cmsdk_mcu/sram_hrdata [7]),
    .c(\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [0]),
    .o(\u_cmsdk_mcu/u_ahb_ram/n13 [7]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u2165 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qiqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[17] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[17] ),
    .o(_al_u2165_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u2166 (
    .a(_al_u2165_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sjqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[17] ),
    .o(_al_u2166_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u2167 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dfqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gkqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[17] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pbbbx6 ),
    .o(_al_u2167_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u2168 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hhqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[17] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[17] ),
    .o(_al_u2168_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u2169 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fgqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yfqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[15] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[15] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Drzow6 ));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u2170 (
    .a(_al_u2166_o),
    .b(_al_u2167_o),
    .c(_al_u2168_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Drzow6 ),
    .o(_al_u2170_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2171 (
    .a(_al_u2170_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J10iu6 ),
    .o(_al_u2171_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(B*~A))"),
    .INIT(8'h0b))
    _al_u2172 (
    .a(_al_u1888_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I8lax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wvgax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lcqow6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*C)*~(B*~A))"),
    .INIT(16'h0bbb))
    _al_u2173 (
    .a(_al_u1968_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lcqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G64iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wvgax6 ),
    .o(_al_u2173_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*~A)"),
    .INIT(8'h04))
    _al_u2174 (
    .a(_al_u1888_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I8lax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wvgax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gdqow6 ));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C*~A))"),
    .INIT(8'h73))
    _al_u2175 (
    .a(_al_u2171_o),
    .b(_al_u2173_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gdqow6 ),
    .o(\u_cmsdk_mcu/HWDATA [17]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2176 (
    .a(\u_cmsdk_mcu/HWDATA [1]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C1wpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I4eiu6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2177 (
    .a(\u_cmsdk_mcu/HWDATA [1]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n223 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpolset [1]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2178 (
    .a(\u_cmsdk_mcu/HWDATA [1]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n178 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttypeset [1]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2179 (
    .a(\u_cmsdk_mcu/HWDATA [1]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n133 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intenset [1]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2180 (
    .a(\u_cmsdk_mcu/HWDATA [1]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n88 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_altfuncset [1]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2181 (
    .a(\u_cmsdk_mcu/HWDATA [1]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n43 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_doutenset [1]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2182 (
    .a(\u_cmsdk_mcu/HWDATA [1]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n223 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpolset [1]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2183 (
    .a(\u_cmsdk_mcu/HWDATA [1]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n178 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttypeset [1]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2184 (
    .a(\u_cmsdk_mcu/HWDATA [1]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n133 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intenset [1]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2185 (
    .a(\u_cmsdk_mcu/HWDATA [1]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n88 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_altfuncset [1]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2186 (
    .a(\u_cmsdk_mcu/HWDATA [1]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n43 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_doutenset [1]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u2187 (
    .a(\u_cmsdk_mcu/HWDATA [1]),
    .b(\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [0]),
    .c(\u_cmsdk_mcu/flash_hrdata [1]),
    .o(\u_cmsdk_mcu/u_ahb_rom/n13 [1]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2188 (
    .a(\u_cmsdk_mcu/HWDATA [1]),
    .b(\u_cmsdk_mcu/sram_hrdata [1]),
    .c(\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [0]),
    .o(\u_cmsdk_mcu/u_ahb_ram/n13 [1]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2189 (
    .a(\u_cmsdk_mcu/HWDATA [9]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n226 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpolset [9]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2190 (
    .a(\u_cmsdk_mcu/HWDATA [9]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n181 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttypeset [9]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2191 (
    .a(\u_cmsdk_mcu/HWDATA [9]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n136 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intenset [9]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2192 (
    .a(\u_cmsdk_mcu/HWDATA [9]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n91 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_altfuncset [9]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2193 (
    .a(\u_cmsdk_mcu/HWDATA [9]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n46 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_doutenset [9]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2194 (
    .a(\u_cmsdk_mcu/HWDATA [9]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n226 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpolset [9]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2195 (
    .a(\u_cmsdk_mcu/HWDATA [9]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n181 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttypeset [9]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2196 (
    .a(\u_cmsdk_mcu/HWDATA [9]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n136 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intenset [9]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2197 (
    .a(\u_cmsdk_mcu/HWDATA [9]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n91 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_altfuncset [9]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2198 (
    .a(\u_cmsdk_mcu/HWDATA [9]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n46 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_doutenset [9]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u2199 (
    .a(\u_cmsdk_mcu/HWDATA [9]),
    .b(\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [10]),
    .c(\u_cmsdk_mcu/flash_hrdata [9]),
    .o(\u_cmsdk_mcu/u_ahb_rom/n13 [9]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2200 (
    .a(\u_cmsdk_mcu/HWDATA [9]),
    .b(\u_cmsdk_mcu/sram_hrdata [9]),
    .c(\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [10]),
    .o(\u_cmsdk_mcu/u_ahb_ram/n13 [9]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*C)*~(B*~A))"),
    .INIT(16'h0bbb))
    _al_u2201 (
    .a(_al_u1916_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lcqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N64iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wvgax6 ),
    .o(_al_u2201_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u2202 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qiqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[18] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[18] ),
    .o(_al_u2202_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u2203 (
    .a(_al_u2202_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[18] ),
    .o(_al_u2203_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u2204 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dfqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gkqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[18] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Syjbx6 ),
    .o(_al_u2204_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u2205 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hhqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sjqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[18] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[18] ),
    .o(_al_u2205_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u2206 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fgqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yfqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[16] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[16] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eazow6 ));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u2207 (
    .a(_al_u2203_o),
    .b(_al_u2204_o),
    .c(_al_u2205_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eazow6 ),
    .o(_al_u2207_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2208 (
    .a(_al_u2207_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C10iu6 ),
    .o(_al_u2208_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*~B))"),
    .INIT(8'h75))
    _al_u2209 (
    .a(_al_u2201_o),
    .b(_al_u2208_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gdqow6 ),
    .o(\u_cmsdk_mcu/HWDATA [18]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*C)*~(B*~A))"),
    .INIT(16'h0bbb))
    _al_u2210 (
    .a(_al_u1925_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lcqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U64iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wvgax6 ),
    .o(_al_u2210_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u2211 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qiqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[19] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[19] ),
    .o(_al_u2211_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u2212 (
    .a(_al_u2211_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sjqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[19] ),
    .o(_al_u2212_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u2213 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hhqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dfqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[19] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T6kbx6 ),
    .o(_al_u2213_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u2214 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fgqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yfqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[17] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[17] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T0zow6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u2215 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gkqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[19] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[19] ),
    .o(_al_u2215_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u2216 (
    .a(_al_u2212_o),
    .b(_al_u2213_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T0zow6 ),
    .d(_al_u2215_o),
    .o(_al_u2216_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2217 (
    .a(_al_u2216_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V00iu6 ),
    .o(_al_u2217_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*~B))"),
    .INIT(8'h75))
    _al_u2218 (
    .a(_al_u2210_o),
    .b(_al_u2217_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gdqow6 ),
    .o(\u_cmsdk_mcu/HWDATA [19]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u2219 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qiqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[20] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[20] ),
    .o(_al_u2219_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u2220 (
    .a(_al_u2219_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sjqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[20] ),
    .o(_al_u2220_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u2221 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hhqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dfqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[20] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fjdbx6 ),
    .o(_al_u2221_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u2222 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fgqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yfqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[18] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[18] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uqyow6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u2223 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gkqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[20] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[20] ),
    .o(_al_u2223_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u2224 (
    .a(_al_u2220_o),
    .b(_al_u2221_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uqyow6 ),
    .d(_al_u2223_o),
    .o(_al_u2224_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2225 (
    .a(_al_u2224_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H00iu6 ),
    .o(_al_u2225_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*C)*~(B*~A))"),
    .INIT(16'h0bbb))
    _al_u2226 (
    .a(_al_u2225_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gdqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B74iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wvgax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qoyow6 ));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*~B))"),
    .INIT(8'h75))
    _al_u2227 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qoyow6 ),
    .b(_al_u1934_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lcqow6 ),
    .o(\u_cmsdk_mcu/HWDATA [20]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*C)*~(B*~A))"),
    .INIT(16'h0bbb))
    _al_u2228 (
    .a(_al_u1943_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lcqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I74iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wvgax6 ),
    .o(_al_u2228_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u2229 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qiqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[21] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[21] ),
    .o(_al_u2229_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u2230 (
    .a(_al_u2229_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sjqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[21] ),
    .o(_al_u2230_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u2231 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hhqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dfqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[21] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M2ebx6 ),
    .o(_al_u2231_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u2232 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fgqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yfqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[19] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[19] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jhyow6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u2233 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gkqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[21] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[21] ),
    .o(_al_u2233_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u2234 (
    .a(_al_u2230_o),
    .b(_al_u2231_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jhyow6 ),
    .d(_al_u2233_o),
    .o(_al_u2234_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2235 (
    .a(_al_u2234_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A00iu6 ),
    .o(_al_u2235_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*~B))"),
    .INIT(8'h75))
    _al_u2236 (
    .a(_al_u2228_o),
    .b(_al_u2235_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gdqow6 ),
    .o(\u_cmsdk_mcu/HWDATA [21]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*C)*~(B*~A))"),
    .INIT(16'h0bbb))
    _al_u2237 (
    .a(_al_u1952_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lcqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P74iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wvgax6 ),
    .o(_al_u2237_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u2238 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hhqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qiqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[22] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[22] ),
    .o(_al_u2238_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u2239 (
    .a(_al_u2238_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dfqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tlebx6 ),
    .o(_al_u2239_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u2240 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[22] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[22] ),
    .o(_al_u2240_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u2241 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fgqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yfqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[20] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[20] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y7yow6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u2242 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gkqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sjqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[22] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[22] ),
    .o(_al_u2242_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u2243 (
    .a(_al_u2239_o),
    .b(_al_u2240_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y7yow6 ),
    .d(_al_u2242_o),
    .o(_al_u2243_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2244 (
    .a(_al_u2243_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tzzhu6 ),
    .o(_al_u2244_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*~B))"),
    .INIT(8'h75))
    _al_u2245 (
    .a(_al_u2237_o),
    .b(_al_u2244_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gdqow6 ),
    .o(\u_cmsdk_mcu/HWDATA [22]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u2246 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hhqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qiqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[23] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[23] ),
    .o(_al_u2246_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u2247 (
    .a(_al_u2246_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sjqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[23] ),
    .o(_al_u2247_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u2248 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dfqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[23] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztgbx6 ),
    .o(_al_u2248_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u2249 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fgqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yfqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[21] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[21] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nyxow6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u2250 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gkqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[23] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[23] ),
    .o(_al_u2250_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u2251 (
    .a(_al_u2247_o),
    .b(_al_u2248_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nyxow6 ),
    .d(_al_u2250_o),
    .o(_al_u2251_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2252 (
    .a(_al_u2251_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mzzhu6 ),
    .o(_al_u2252_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*C)*~(B*~A))"),
    .INIT(16'h0bbb))
    _al_u2253 (
    .a(_al_u2252_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gdqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W74iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wvgax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jwxow6 ));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*~B))"),
    .INIT(8'h75))
    _al_u2254 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jwxow6 ),
    .b(_al_u1961_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lcqow6 ),
    .o(\u_cmsdk_mcu/HWDATA [23]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u2255 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qiqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[25] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[25] ),
    .o(_al_u2255_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u2256 (
    .a(_al_u2255_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[25] ),
    .o(_al_u2256_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u2257 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hhqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dfqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[25] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nwbbx6 ),
    .o(_al_u2257_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u2258 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fgqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yfqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[23] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[23] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G6xow6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u2259 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gkqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sjqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[25] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[25] ),
    .o(_al_u2259_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u2260 (
    .a(_al_u2256_o),
    .b(_al_u2257_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G6xow6 ),
    .d(_al_u2259_o),
    .o(_al_u2260_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2261 (
    .a(_al_u2260_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yyzhu6 ),
    .o(_al_u2261_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'h0305))
    _al_u2262 (
    .a(_al_u2261_o),
    .b(_al_u1968_o),
    .c(_al_u1906_o),
    .d(_al_u1299_o),
    .o(_al_u2262_o));
  AL_MAP_LUT3 #(
    .EQN("~(~A*~(C*B))"),
    .INIT(8'hea))
    _al_u2263 (
    .a(_al_u2262_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[1] ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zdiax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yjliu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u2264 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hhqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[30] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[30] ),
    .o(_al_u2264_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u2265 (
    .a(_al_u2264_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qiqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[30] ),
    .o(_al_u2265_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u2266 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dfqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F6dbx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[30] ),
    .o(_al_u2266_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u2267 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fgqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yfqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[28] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[28] ),
    .o(_al_u2267_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u2268 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gkqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sjqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[30] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[30] ),
    .o(_al_u2268_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u2269 (
    .a(_al_u2265_o),
    .b(_al_u2266_o),
    .c(_al_u2267_o),
    .d(_al_u2268_o),
    .o(_al_u2269_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2270 (
    .a(_al_u2269_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ixzhu6 ),
    .o(_al_u2270_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*C)*~(B*~A))"),
    .INIT(16'h0bbb))
    _al_u2271 (
    .a(_al_u2270_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gdqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T94iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wvgax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jrvow6 ));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*A)"),
    .INIT(16'h0080))
    _al_u2272 (
    .a(_al_u1888_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qk9pw6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I8lax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wvgax6 ),
    .o(_al_u2272_o));
  AL_MAP_LUT4 #(
    .EQN("~(B*~A*~(D*~C))"),
    .INIT(16'hbfbb))
    _al_u2273 (
    .a(_al_u2121_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jrvow6 ),
    .c(_al_u2128_o),
    .d(_al_u2272_o),
    .o(\u_cmsdk_mcu/HWDATA [30]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*C)*~(B*~A))"),
    .INIT(16'h0bbb))
    _al_u2274 (
    .a(_al_u2150_o),
    .b(_al_u2272_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lm1iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wvgax6 ),
    .o(_al_u2274_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u2275 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sjqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[31] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[31] ),
    .o(_al_u2275_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u2276 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dfqow6 ),
    .b(_al_u2275_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Usnpw6 ),
    .o(_al_u2276_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u2277 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qiqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[31] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[31] ),
    .o(_al_u2277_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u2278 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hhqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gkqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[31] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[31] ),
    .o(_al_u2278_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u2279 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fgqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yfqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[29] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[29] ),
    .o(_al_u2279_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u2280 (
    .a(_al_u2276_o),
    .b(_al_u2277_o),
    .c(_al_u2278_o),
    .d(_al_u2279_o),
    .o(_al_u2280_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2281 (
    .a(_al_u2280_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bxzhu6 ),
    .o(_al_u2281_o));
  AL_MAP_LUT4 #(
    .EQN("~(B*~A*~(~D*C))"),
    .INIT(16'hbbfb))
    _al_u2282 (
    .a(_al_u2143_o),
    .b(_al_u2274_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gdqow6 ),
    .d(_al_u2281_o),
    .o(\u_cmsdk_mcu/HWDATA [31]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u2283 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qiqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[16] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[16] ),
    .o(_al_u2283_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u2284 (
    .a(_al_u2283_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gkqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[16] ),
    .o(_al_u2284_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u2285 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hhqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dfqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Chwpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[16] ),
    .o(_al_u2285_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u2286 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fgqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yfqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[14] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[14] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Peqow6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u2287 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sjqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[16] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[16] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ciqow6 ));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u2288 (
    .a(_al_u2284_o),
    .b(_al_u2285_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Peqow6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ciqow6 ),
    .o(_al_u2288_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2289 (
    .a(_al_u2288_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q10iu6 ),
    .o(_al_u2289_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*C)*~(B*~A))"),
    .INIT(16'h0bbb))
    _al_u2290 (
    .a(_al_u1882_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lcqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z54iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wvgax6 ),
    .o(_al_u2290_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C*~A))"),
    .INIT(8'h73))
    _al_u2291 (
    .a(_al_u2289_o),
    .b(_al_u2290_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gdqow6 ),
    .o(\u_cmsdk_mcu/HWDATA [16]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    _al_u2292 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Golpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Krlpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vplpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zslpw6 ),
    .o(_al_u2292_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C@B))"),
    .INIT(8'h41))
    _al_u2293 (
    .a(_al_u2292_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rilpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y8lpw6 ),
    .o(_al_u2293_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*~B*A)"),
    .INIT(16'h0020))
    _al_u2294 (
    .a(_al_u1250_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bclpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jflpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sdlpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M7zhu6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2295 (
    .a(_al_u2293_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M7zhu6 ),
    .o(_al_u2295_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u2296 (
    .a(_al_u1251_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kalpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yklpw6 ),
    .o(_al_u2296_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*(~(B)*~(C)*~(D)+B*~(C)*~(D)+~(B)*C*~(D)+B*~(C)*D+~(B)*C*D))"),
    .INIT(16'h1415))
    _al_u2297 (
    .a(_al_u2295_o),
    .b(_al_u2296_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jflpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rsyhu6_lutinv ),
    .o(_al_u2297_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u2298 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bclpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sdlpw6 ),
    .o(_al_u2298_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u2299 (
    .a(_al_u1250_o),
    .b(_al_u2298_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jflpw6 ),
    .o(_al_u2299_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2300 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jflpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yklpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Epyhu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(D*C*B))"),
    .INIT(16'h1555))
    _al_u2301 (
    .a(_al_u2299_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Epyhu6 ),
    .c(_al_u1251_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kalpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ffyhu6 ));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u2302 (
    .a(_al_u529_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jflpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kalpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T0zhu6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u2303 (
    .a(_al_u1757_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bclpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A1zhu6_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u2304 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T0zhu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A1zhu6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I6yhu6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    _al_u2305 (
    .a(_al_u1757_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bclpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Krlpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yklpw6 ),
    .o(_al_u2305_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*B*~(~D*~A))"),
    .INIT(16'h0c08))
    _al_u2306 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ffyhu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I6yhu6_lutinv ),
    .c(_al_u2305_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rilpw6 ),
    .o(_al_u2306_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(~C*(D@B)))"),
    .INIT(16'h5451))
    _al_u2307 (
    .a(_al_u1253_o),
    .b(_al_u1755_o),
    .c(_al_u1761_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jflpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Spyhu6 ));
  AL_MAP_LUT4 #(
    .EQN("~(C*~(D*~(B*A)))"),
    .INIT(16'h7f0f))
    _al_u2308 (
    .a(_al_u2297_o),
    .b(_al_u2306_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Spyhu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U5yhu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zehpw6 [3]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u2309 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Azeiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N8rpw6 ),
    .o(_al_u2309_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u2310 (
    .a(_al_u2309_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ozeiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvgiu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C1wpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q8eiu6_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u2311 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ozeiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvgiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C1wpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L9eiu6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u2312 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q8eiu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L9eiu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Coupw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J7xax6 ),
    .o(_al_u2312_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(D*C))"),
    .INIT(16'h0444))
    _al_u2313 (
    .a(_al_u2309_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ozeiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvgiu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C1wpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J8eiu6 ));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*B))"),
    .INIT(8'hd5))
    _al_u2314 (
    .a(_al_u2312_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J8eiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6gpw6 [23]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S8uhu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u2315 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q8eiu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L9eiu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D7gbx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F9gbx6 ),
    .o(_al_u2315_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*B))"),
    .INIT(8'hd5))
    _al_u2316 (
    .a(_al_u2315_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J8eiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6gpw6 [22]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z8uhu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u2317 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J8eiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L9eiu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tjkpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6gpw6 [21]),
    .o(_al_u2317_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*B))"),
    .INIT(8'hd5))
    _al_u2318 (
    .a(_al_u2317_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q8eiu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rhkpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G9uhu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u2319 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J8eiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L9eiu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z8jpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6gpw6 [20]),
    .o(_al_u2319_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*B))"),
    .INIT(8'hd5))
    _al_u2320 (
    .a(_al_u2319_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q8eiu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X6jpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N9uhu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u2321 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q8eiu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L9eiu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hhvpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nr7ax6 ),
    .o(_al_u2321_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*B))"),
    .INIT(8'hd5))
    _al_u2322 (
    .a(_al_u2321_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J8eiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6gpw6 [19]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9uhu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u2323 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J8eiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L9eiu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N0xpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6gpw6 [18]),
    .o(_al_u2323_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*B))"),
    .INIT(8'hd5))
    _al_u2324 (
    .a(_al_u2323_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q8eiu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lywpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bauhu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u2325 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J8eiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L9eiu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Amupw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6gpw6 [17]),
    .o(_al_u2325_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*B))"),
    .INIT(8'hd5))
    _al_u2326 (
    .a(_al_u2325_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q8eiu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yjupw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iauhu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u2327 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J8eiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L9eiu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wlspw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6gpw6 [16]),
    .o(_al_u2327_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*B))"),
    .INIT(8'hd5))
    _al_u2328 (
    .a(_al_u2327_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q8eiu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ujspw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pauhu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u2329 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J8eiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L9eiu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nbxax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6gpw6 [15]),
    .o(_al_u2329_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*B))"),
    .INIT(8'hd5))
    _al_u2330 (
    .a(_al_u2329_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q8eiu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L9xax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wauhu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u2331 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q8eiu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L9eiu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pdxax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rfxax6 ),
    .o(_al_u2331_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*B))"),
    .INIT(8'hd5))
    _al_u2332 (
    .a(_al_u2331_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J8eiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6gpw6 [14]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dbuhu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u2333 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J8eiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L9eiu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T9kpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6gpw6 [13]),
    .o(_al_u2333_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*B))"),
    .INIT(8'hd5))
    _al_u2334 (
    .a(_al_u2333_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q8eiu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R7kpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kbuhu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u2335 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J8eiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L9eiu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V0jpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6gpw6 [12]),
    .o(_al_u2335_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*B))"),
    .INIT(8'hd5))
    _al_u2336 (
    .a(_al_u2335_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q8eiu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tyipw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rbuhu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u2337 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J8eiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L9eiu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pt7ax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6gpw6 [11]),
    .o(_al_u2337_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*B))"),
    .INIT(8'hd5))
    _al_u2338 (
    .a(_al_u2337_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q8eiu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ofmpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ybuhu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u2339 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q8eiu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L9eiu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tptpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vrtpw6 ),
    .o(_al_u2339_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*B))"),
    .INIT(8'hd5))
    _al_u2340 (
    .a(_al_u2339_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J8eiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6gpw6 [10]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fcuhu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u2341 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J8eiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L9eiu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uojbx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6gpw6 [9]),
    .o(_al_u2341_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*B))"),
    .INIT(8'hd5))
    _al_u2342 (
    .a(_al_u2341_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q8eiu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tmjbx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mcuhu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u2343 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q8eiu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L9eiu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rq0qw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ss0qw6 ),
    .o(_al_u2343_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*B))"),
    .INIT(8'hd5))
    _al_u2344 (
    .a(_al_u2343_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J8eiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6gpw6 [8]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tcuhu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u2345 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q8eiu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L9eiu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Thxax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ujxax6 ),
    .o(_al_u2345_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*B))"),
    .INIT(8'hd5))
    _al_u2346 (
    .a(_al_u2345_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J8eiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6gpw6 [7]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aduhu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u2347 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J8eiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L9eiu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rv7ax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6gpw6 [6]),
    .o(_al_u2347_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*B))"),
    .INIT(8'hd5))
    _al_u2348 (
    .a(_al_u2347_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q8eiu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ox9bx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hduhu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u2349 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q8eiu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L9eiu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X5opw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y7opw6 ),
    .o(_al_u2349_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*B))"),
    .INIT(8'hd5))
    _al_u2350 (
    .a(_al_u2349_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J8eiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6gpw6 [5]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oduhu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u2351 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J8eiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L9eiu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Johbx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6gpw6 [4]),
    .o(_al_u2351_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*B))"),
    .INIT(8'hd5))
    _al_u2352 (
    .a(_al_u2351_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q8eiu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Imhbx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vduhu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u2353 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q8eiu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L9eiu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oyhbx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0ibx6 ),
    .o(_al_u2353_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*B))"),
    .INIT(8'hd5))
    _al_u2354 (
    .a(_al_u2353_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J8eiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6gpw6 [3]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ceuhu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u2355 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J8eiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L9eiu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kzabx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6gpw6 [2]),
    .o(_al_u2355_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*B))"),
    .INIT(8'hd5))
    _al_u2356 (
    .a(_al_u2355_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q8eiu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vlxax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jeuhu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u2357 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q8eiu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L9eiu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oarpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wnxax6 ),
    .o(_al_u2357_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*B))"),
    .INIT(8'hd5))
    _al_u2358 (
    .a(_al_u2357_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J8eiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6gpw6 [1]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qeuhu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u2359 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q8eiu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L9eiu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6rpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N8rpw6 ),
    .o(_al_u2359_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*B))"),
    .INIT(8'hd5))
    _al_u2360 (
    .a(_al_u2359_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J8eiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6gpw6 [0]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xeuhu6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u2361 (
    .a(_al_u1812_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hgrpw6 ),
    .o(_al_u2361_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u2362 (
    .a(_al_u2361_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nbkiu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wkjiu6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2363 (
    .a(_al_u1812_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9ypw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W0piu6_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2364 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Skjax6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 ),
    .o(_al_u2364_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u2365 (
    .a(_al_u2364_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P14qw6 ),
    .o(_al_u2365_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~A*~(D*C))"),
    .INIT(16'h0111))
    _al_u2366 (
    .a(_al_u1802_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wkjiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W0piu6_lutinv ),
    .d(_al_u2365_o),
    .o(_al_u2366_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2367 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 ),
    .o(_al_u2367_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2368 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W0piu6_lutinv ),
    .b(_al_u2367_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hviiu6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u2369 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rwjax6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6 ),
    .o(_al_u2369_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*A*~(~D*B))"),
    .INIT(16'h0a02))
    _al_u2370 (
    .a(_al_u2369_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N4kax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4jax6 ),
    .o(_al_u2370_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2371 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rwjax6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6 ),
    .o(_al_u2371_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*~(~D*~C)))"),
    .INIT(16'h222a))
    _al_u2372 (
    .a(_al_u2366_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hviiu6 ),
    .c(_al_u2370_o),
    .d(_al_u2371_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M1jiu6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2373 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Skjax6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 ),
    .o(_al_u2373_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u2374 (
    .a(_al_u2373_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oxhow6 ));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(~D*~C*B))"),
    .INIT(16'h5551))
    _al_u2375 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oxhow6 ),
    .b(_al_u2364_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 ),
    .o(_al_u2375_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u2376 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nbkiu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qxoiu6 ),
    .o(_al_u2376_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*A*~(~D*C))"),
    .INIT(16'h2202))
    _al_u2377 (
    .a(_al_u2375_o),
    .b(_al_u2376_o),
    .c(_al_u2364_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 ),
    .o(_al_u2377_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u2378 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N4kax6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P14qw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 ),
    .o(_al_u2378_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D*~C*~B))"),
    .INIT(16'ha8aa))
    _al_u2379 (
    .a(_al_u2377_o),
    .b(_al_u2378_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9ypw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 ),
    .o(_al_u2379_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u2380 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Irmpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N4kax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S7mpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wfspw6 ),
    .o(_al_u2380_o));
  AL_MAP_LUT4 #(
    .EQN("(C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'ha0c0))
    _al_u2381 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R9aiu6 ),
    .b(_al_u2380_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9ypw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wkipw6 ),
    .o(_al_u2381_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(C*~A))"),
    .INIT(16'haf23))
    _al_u2382 (
    .a(_al_u2379_o),
    .b(_al_u1815_o),
    .c(_al_u2361_o),
    .d(_al_u2381_o),
    .o(_al_u2382_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u2383 (
    .a(_al_u1812_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uyiiu6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2384 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9ypw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J9kiu6_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2385 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uyiiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J9kiu6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vviiu6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u2386 (
    .a(_al_u2364_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 ),
    .o(_al_u2386_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u2387 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 ),
    .o(_al_u2387_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(~B*~(~D*A)))"),
    .INIT(16'hc0e0))
    _al_u2388 (
    .a(_al_u932_o),
    .b(_al_u2387_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 ),
    .o(_al_u2388_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(B*A))"),
    .INIT(8'h07))
    _al_u2389 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W0piu6_lutinv ),
    .b(_al_u2386_o),
    .c(_al_u2388_o),
    .o(_al_u2389_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~D*~C*A))"),
    .INIT(16'hccc4))
    _al_u2390 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vviiu6 ),
    .b(_al_u2389_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6 ),
    .o(_al_u2390_o));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~(C*B*A))"),
    .INIT(16'hff80))
    _al_u2391 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M1jiu6 ),
    .b(_al_u2382_o),
    .c(_al_u2390_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G81ju6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u2392 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 ),
    .o(_al_u2392_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u2393 (
    .a(_al_u1663_o),
    .b(_al_u1583_o),
    .c(_al_u2392_o),
    .o(_al_u2393_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u2394 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nkaju6_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(A*(C@B))"),
    .INIT(8'h28))
    _al_u2395 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nkaju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 ),
    .o(_al_u2395_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u2396 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S2ziu6_lutinv ),
    .b(_al_u1662_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 ),
    .o(_al_u2396_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    _al_u2397 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lu0iu6 ),
    .b(_al_u2393_o),
    .c(_al_u2395_o),
    .d(_al_u2396_o),
    .o(_al_u2397_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2398 (
    .a(_al_u2397_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vgjpw6 ),
    .o(_al_u2398_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u2399 (
    .a(_al_u678_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vgjpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 ),
    .o(_al_u2399_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u2400 (
    .a(_al_u909_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vgjpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zf7ju6 ));
  AL_MAP_LUT3 #(
    .EQN("(C*~(~B*~A))"),
    .INIT(8'he0))
    _al_u2401 (
    .a(_al_u2399_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zf7ju6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rkkax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qk8ju6_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u2402 (
    .a(_al_u2398_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qk8ju6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T75ju6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2403 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 ),
    .o(_al_u2403_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*~B))"),
    .INIT(8'h54))
    _al_u2404 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Np7ow6_lutinv ),
    .b(_al_u2403_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 ),
    .o(_al_u2404_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(~A*~(C*B)))"),
    .INIT(16'hea00))
    _al_u2405 (
    .a(_al_u2404_o),
    .b(_al_u604_o),
    .c(_al_u1344_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ),
    .o(_al_u2405_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u2406 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 ),
    .o(_al_u2406_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u2407 (
    .a(_al_u695_o),
    .b(_al_u2406_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 ),
    .o(_al_u2407_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2408 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N98iu6_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u2409 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N98iu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ),
    .o(_al_u2409_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2410 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Owoiu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(~D*~(~C*~B)))"),
    .INIT(16'h5501))
    _al_u2411 (
    .a(_al_u2409_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Owoiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 ),
    .o(_al_u2411_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C*~B*~A))"),
    .INIT(16'hef00))
    _al_u2412 (
    .a(_al_u2405_o),
    .b(_al_u2407_o),
    .c(_al_u2411_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vgjpw6 ),
    .o(_al_u2412_o));
  AL_MAP_LUT3 #(
    .EQN("(~(A)*~(B)*~(C)+~(A)*B*~(C)+A*B*~(C)+A*~(B)*C+A*B*C)"),
    .INIT(8'had))
    _al_u2413 (
    .a(_al_u2398_o),
    .b(_al_u2412_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qk8ju6_lutinv ),
    .o(_al_u2413_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u2414 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hhqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[28] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[28] ),
    .o(_al_u2414_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u2415 (
    .a(_al_u2414_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[28] ),
    .o(_al_u2415_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u2416 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dfqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qiqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ibqpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[28] ),
    .o(_al_u2416_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u2417 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fgqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yfqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[26] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[26] ),
    .o(_al_u2417_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u2418 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gkqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sjqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[28] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[28] ),
    .o(_al_u2418_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u2419 (
    .a(_al_u2415_o),
    .b(_al_u2416_o),
    .c(_al_u2417_o),
    .d(_al_u2418_o),
    .o(_al_u2419_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2420 (
    .a(_al_u2419_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dyzhu6 ),
    .o(_al_u2420_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2421 (
    .a(_al_u2397_o),
    .b(_al_u2412_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A85ju6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("~(B*~(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    .INIT(16'hbfb3))
    _al_u2422 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T75ju6 ),
    .b(_al_u2413_o),
    .c(_al_u2420_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A85ju6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [28]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u2423 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qiqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sjqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[29] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[29] ),
    .o(_al_u2423_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u2424 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hhqow6 ),
    .b(_al_u2423_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[29] ),
    .o(_al_u2424_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u2425 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dfqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gkqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[29] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sx3qw6 ),
    .o(_al_u2425_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u2426 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[29] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[29] ),
    .o(_al_u2426_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u2427 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fgqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yfqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[27] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[27] ),
    .o(_al_u2427_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u2428 (
    .a(_al_u2424_o),
    .b(_al_u2425_o),
    .c(_al_u2426_o),
    .d(_al_u2427_o),
    .o(_al_u2428_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2429 (
    .a(_al_u2428_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wxzhu6 ),
    .o(_al_u2429_o));
  AL_MAP_LUT4 #(
    .EQN("~(B*~(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D))"),
    .INIT(16'hbbf3))
    _al_u2430 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T75ju6 ),
    .b(_al_u2413_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A85ju6_lutinv ),
    .d(_al_u2429_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [29]));
  AL_MAP_LUT4 #(
    .EQN("~(C*~(D*~(B)*~(A)+D*B*~(A)+~(D)*B*A+D*B*A))"),
    .INIT(16'hdf8f))
    _al_u2431 (
    .a(_al_u2270_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T75ju6 ),
    .c(_al_u2413_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A85ju6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [30]));
  AL_MAP_LUT4 #(
    .EQN("~(C*~(D*~(B)*~(A)+D*B*~(A)+~(D)*B*A+D*B*A))"),
    .INIT(16'hdf8f))
    _al_u2432 (
    .a(_al_u2261_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T75ju6 ),
    .c(_al_u2413_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A85ju6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [25]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u2433 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hhqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dfqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[24] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgkbx6 ),
    .o(_al_u2433_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u2434 (
    .a(_al_u2433_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qiqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[24] ),
    .o(_al_u2434_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u2435 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sjqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[24] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[24] ),
    .o(_al_u2435_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u2436 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fgqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yfqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[22] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[22] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Voxow6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u2437 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gkqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[24] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[24] ),
    .o(_al_u2437_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u2438 (
    .a(_al_u2434_o),
    .b(_al_u2435_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Voxow6 ),
    .d(_al_u2437_o),
    .o(_al_u2438_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2439 (
    .a(_al_u2438_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fzzhu6 ),
    .o(_al_u2439_o));
  AL_MAP_LUT4 #(
    .EQN("~(B*~(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    .INIT(16'hbfb3))
    _al_u2440 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T75ju6 ),
    .b(_al_u2413_o),
    .c(_al_u2439_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A85ju6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [24]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u2441 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hhqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dfqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[27] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nybbx6 ),
    .o(_al_u2441_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u2442 (
    .a(_al_u2441_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[27] ),
    .o(_al_u2442_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u2443 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sjqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[27] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[27] ),
    .o(_al_u2443_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u2444 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fgqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yfqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[25] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[25] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sdwow6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u2445 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qiqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gkqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[27] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[27] ),
    .o(_al_u2445_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u2446 (
    .a(_al_u2442_o),
    .b(_al_u2443_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sdwow6 ),
    .d(_al_u2445_o),
    .o(_al_u2446_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2447 (
    .a(_al_u2446_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kyzhu6 ),
    .o(_al_u2447_o));
  AL_MAP_LUT4 #(
    .EQN("~(B*~(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    .INIT(16'hbfb3))
    _al_u2448 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T75ju6 ),
    .b(_al_u2413_o),
    .c(_al_u2447_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A85ju6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [27]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u2449 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qiqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[26] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[26] ),
    .o(_al_u2449_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u2450 (
    .a(_al_u2449_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[26] ),
    .o(_al_u2450_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u2451 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hhqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dfqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[26] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F8cbx6 ),
    .o(_al_u2451_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u2452 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fgqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yfqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[24] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[24] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ynwow6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u2453 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gkqow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sjqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[26] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[26] ),
    .o(_al_u2453_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u2454 (
    .a(_al_u2450_o),
    .b(_al_u2451_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ynwow6 ),
    .d(_al_u2453_o),
    .o(_al_u2454_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2455 (
    .a(_al_u2454_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ryzhu6 ),
    .o(_al_u2455_o));
  AL_MAP_LUT4 #(
    .EQN("~(B*~(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    .INIT(16'hbfb3))
    _al_u2456 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T75ju6 ),
    .b(_al_u2413_o),
    .c(_al_u2455_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A85ju6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [26]));
  AL_MAP_LUT4 #(
    .EQN("~(B*~(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    .INIT(16'hbfb3))
    _al_u2457 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T75ju6 ),
    .b(_al_u2413_o),
    .c(_al_u2281_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A85ju6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D5epw6 ));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*~A)"),
    .INIT(8'h04))
    _al_u2458 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Np7ow6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D6kiu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ),
    .o(_al_u2458_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D*C*A))"),
    .INIT(16'h1333))
    _al_u2459 (
    .a(_al_u695_o),
    .b(_al_u2458_o),
    .c(_al_u1296_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 ),
    .o(_al_u2459_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(~D*C*B))"),
    .INIT(16'haa2a))
    _al_u2460 (
    .a(_al_u2459_o),
    .b(_al_u1342_o),
    .c(_al_u2403_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 ),
    .o(_al_u2460_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*A*~(D*C))"),
    .INIT(16'h0222))
    _al_u2461 (
    .a(_al_u2460_o),
    .b(_al_u1820_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D6kiu6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 ),
    .o(_al_u2461_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2462 (
    .a(_al_u2461_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vgjpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kc6ju6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u2463 (
    .a(_al_u2399_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zf7ju6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lgkax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 ),
    .o(_al_u2463_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u2464 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kc6ju6 ),
    .b(_al_u2463_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V6jax6 ),
    .o(_al_u2464_o));
  AL_MAP_LUT4 #(
    .EQN("~(C@(A*~(D*~B)))"),
    .INIT(16'h87a5))
    _al_u2465 (
    .a(_al_u2464_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I28ju6 ),
    .c(_al_u2398_o),
    .d(_al_u2412_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q5phu6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2466 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gf1ju6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A3ipw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ph1iu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u2467 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ph1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A5ipw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I0opw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ry2qw6 ),
    .o(_al_u2467_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D*~(~C*B)))"),
    .INIT(16'h08aa))
    _al_u2468 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yn3iu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Krlpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oulpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vplpw6 ),
    .o(_al_u2468_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*B*~(C*A))"),
    .INIT(16'h004c))
    _al_u2469 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pyyhu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B7lpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Krlpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zslpw6 ),
    .o(_al_u2469_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u2470 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qwfax6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P13iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ryfax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Utqpw6 ),
    .o(_al_u2470_o));
  AL_MAP_LUT4 #(
    .EQN("~(~B*~(A*~(D*~C)))"),
    .INIT(16'hecee))
    _al_u2471 (
    .a(_al_u2467_o),
    .b(_al_u2468_o),
    .c(_al_u2469_o),
    .d(_al_u2470_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mmyhu6 ));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u2472 (
    .a(_al_u473_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/write_enable ),
    .c(_al_u1048_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/write_enable0c ));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    _al_u2473 (
    .a(\u_cmsdk_mcu/HWDATA [0]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/intr_stat_set [0]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/write_enable0c ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n114 ));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u2474 (
    .a(_al_u1983_o),
    .b(_al_u588_o),
    .c(_al_u1988_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intclr_normal_write0 ));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(B*A))"),
    .INIT(8'hf8))
    _al_u2475 (
    .a(\u_cmsdk_mcu/HWDATA [0]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intclr_normal_write0 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_masked_int [0]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n271 ));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u2476 (
    .a(_al_u1983_o),
    .b(_al_u588_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .o(_al_u2476_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2477 (
    .a(\u_cmsdk_mcu/HWDATA [0]),
    .b(_al_u2476_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n234 ));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u2478 (
    .a(_al_u1987_o),
    .b(_al_u588_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .o(_al_u2478_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2479 (
    .a(\u_cmsdk_mcu/HWDATA [0]),
    .b(_al_u2478_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n189 ));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u2480 (
    .a(_al_u1987_o),
    .b(_al_u588_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .o(_al_u2480_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2481 (
    .a(\u_cmsdk_mcu/HWDATA [0]),
    .b(_al_u2480_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n144 ));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u2482 (
    .a(_al_u1993_o),
    .b(_al_u588_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .o(_al_u2482_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2483 (
    .a(\u_cmsdk_mcu/HWDATA [0]),
    .b(_al_u2482_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n99 ));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u2484 (
    .a(_al_u1993_o),
    .b(_al_u588_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .o(_al_u2484_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2485 (
    .a(\u_cmsdk_mcu/HWDATA [0]),
    .b(_al_u2484_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n54 ));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u2486 (
    .a(_al_u1983_o),
    .b(_al_u593_o),
    .c(_al_u1988_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intclr_normal_write0 ));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(B*A))"),
    .INIT(8'hf8))
    _al_u2487 (
    .a(\u_cmsdk_mcu/HWDATA [0]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intclr_normal_write0 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/new_masked_int [0]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n271 ));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u2488 (
    .a(_al_u1983_o),
    .b(_al_u593_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .o(_al_u2488_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2489 (
    .a(\u_cmsdk_mcu/HWDATA [0]),
    .b(_al_u2488_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n234 ));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u2490 (
    .a(_al_u1987_o),
    .b(_al_u593_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .o(_al_u2490_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2491 (
    .a(\u_cmsdk_mcu/HWDATA [0]),
    .b(_al_u2490_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n189 ));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u2492 (
    .a(_al_u1987_o),
    .b(_al_u593_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .o(_al_u2492_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2493 (
    .a(\u_cmsdk_mcu/HWDATA [0]),
    .b(_al_u2492_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n144 ));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u2494 (
    .a(_al_u1993_o),
    .b(_al_u593_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .o(_al_u2494_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2495 (
    .a(\u_cmsdk_mcu/HWDATA [0]),
    .b(_al_u2494_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n99 ));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u2496 (
    .a(_al_u1993_o),
    .b(_al_u593_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .o(_al_u2496_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2497 (
    .a(\u_cmsdk_mcu/HWDATA [0]),
    .b(_al_u2496_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n54 ));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u2498 (
    .a(_al_u1983_o),
    .b(_al_u585_o),
    .c(_al_u1988_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intclr_normal_write1 ));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(B*A))"),
    .INIT(8'hf8))
    _al_u2499 (
    .a(\u_cmsdk_mcu/HWDATA [8]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intclr_normal_write1 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_masked_int [8]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n287 ));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u2500 (
    .a(_al_u1983_o),
    .b(_al_u585_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .o(_al_u2500_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2501 (
    .a(\u_cmsdk_mcu/HWDATA [8]),
    .b(_al_u2500_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n250 ));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u2502 (
    .a(_al_u1987_o),
    .b(_al_u585_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .o(_al_u2502_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2503 (
    .a(\u_cmsdk_mcu/HWDATA [8]),
    .b(_al_u2502_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n205 ));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u2504 (
    .a(_al_u1987_o),
    .b(_al_u585_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .o(_al_u2504_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2505 (
    .a(\u_cmsdk_mcu/HWDATA [8]),
    .b(_al_u2504_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n160 ));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u2506 (
    .a(_al_u1993_o),
    .b(_al_u585_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .o(_al_u2506_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2507 (
    .a(\u_cmsdk_mcu/HWDATA [8]),
    .b(_al_u2506_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n115 ));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u2508 (
    .a(_al_u1993_o),
    .b(_al_u585_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .o(_al_u2508_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2509 (
    .a(\u_cmsdk_mcu/HWDATA [8]),
    .b(_al_u2508_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n70 ));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u2510 (
    .a(_al_u1983_o),
    .b(_al_u591_o),
    .c(_al_u1988_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intclr_normal_write1 ));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(B*A))"),
    .INIT(8'hf8))
    _al_u2511 (
    .a(\u_cmsdk_mcu/HWDATA [8]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intclr_normal_write1 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/new_masked_int [8]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n287 ));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u2512 (
    .a(_al_u1983_o),
    .b(_al_u591_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .o(_al_u2512_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2513 (
    .a(\u_cmsdk_mcu/HWDATA [8]),
    .b(_al_u2512_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n250 ));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u2514 (
    .a(_al_u1987_o),
    .b(_al_u591_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .o(_al_u2514_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2515 (
    .a(\u_cmsdk_mcu/HWDATA [8]),
    .b(_al_u2514_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n205 ));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u2516 (
    .a(_al_u1987_o),
    .b(_al_u591_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .o(_al_u2516_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2517 (
    .a(\u_cmsdk_mcu/HWDATA [8]),
    .b(_al_u2516_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n160 ));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u2518 (
    .a(_al_u1993_o),
    .b(_al_u591_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .o(_al_u2518_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2519 (
    .a(\u_cmsdk_mcu/HWDATA [8]),
    .b(_al_u2518_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n115 ));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u2520 (
    .a(_al_u1993_o),
    .b(_al_u591_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .o(_al_u2520_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2521 (
    .a(\u_cmsdk_mcu/HWDATA [8]),
    .b(_al_u2520_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n70 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2522 (
    .a(\u_cmsdk_mcu/HWDATA [10]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n226 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpolset [10]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2523 (
    .a(\u_cmsdk_mcu/HWDATA [10]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n181 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttypeset [10]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2524 (
    .a(\u_cmsdk_mcu/HWDATA [10]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n136 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intenset [10]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2525 (
    .a(\u_cmsdk_mcu/HWDATA [10]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n91 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_altfuncset [10]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2526 (
    .a(\u_cmsdk_mcu/HWDATA [10]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n46 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_doutenset [10]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2527 (
    .a(\u_cmsdk_mcu/HWDATA [10]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n226 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpolset [10]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2528 (
    .a(\u_cmsdk_mcu/HWDATA [10]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n181 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttypeset [10]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2529 (
    .a(\u_cmsdk_mcu/HWDATA [10]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n136 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intenset [10]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2530 (
    .a(\u_cmsdk_mcu/HWDATA [10]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n91 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_altfuncset [10]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2531 (
    .a(\u_cmsdk_mcu/HWDATA [10]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n46 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_doutenset [10]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u2532 (
    .a(\u_cmsdk_mcu/HWDATA [10]),
    .b(\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [10]),
    .c(\u_cmsdk_mcu/flash_hrdata [10]),
    .o(\u_cmsdk_mcu/u_ahb_rom/n13 [10]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2533 (
    .a(\u_cmsdk_mcu/HWDATA [10]),
    .b(\u_cmsdk_mcu/sram_hrdata [10]),
    .c(\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [10]),
    .o(\u_cmsdk_mcu/u_ahb_ram/n13 [10]));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(B*A))"),
    .INIT(8'hf8))
    _al_u2534 (
    .a(\u_cmsdk_mcu/HWDATA [2]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intclr_normal_write0 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_masked_int [2]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n275 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2535 (
    .a(\u_cmsdk_mcu/HWDATA [2]),
    .b(_al_u2476_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n238 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2536 (
    .a(\u_cmsdk_mcu/HWDATA [2]),
    .b(_al_u2478_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n193 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2537 (
    .a(\u_cmsdk_mcu/HWDATA [2]),
    .b(_al_u2480_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n148 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2538 (
    .a(\u_cmsdk_mcu/HWDATA [2]),
    .b(_al_u2482_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n103 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2539 (
    .a(\u_cmsdk_mcu/HWDATA [2]),
    .b(_al_u2484_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n58 ));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(B*A))"),
    .INIT(8'hf8))
    _al_u2540 (
    .a(\u_cmsdk_mcu/HWDATA [2]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intclr_normal_write0 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/new_masked_int [2]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n275 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2541 (
    .a(\u_cmsdk_mcu/HWDATA [2]),
    .b(_al_u2488_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n238 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2542 (
    .a(\u_cmsdk_mcu/HWDATA [2]),
    .b(_al_u2490_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n193 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2543 (
    .a(\u_cmsdk_mcu/HWDATA [2]),
    .b(_al_u2492_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n148 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2544 (
    .a(\u_cmsdk_mcu/HWDATA [2]),
    .b(_al_u2494_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n103 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2545 (
    .a(\u_cmsdk_mcu/HWDATA [2]),
    .b(_al_u2496_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n58 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2546 (
    .a(\u_cmsdk_mcu/HWDATA [11]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n226 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpolset [11]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2547 (
    .a(\u_cmsdk_mcu/HWDATA [11]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n181 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttypeset [11]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2548 (
    .a(\u_cmsdk_mcu/HWDATA [11]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n136 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intenset [11]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2549 (
    .a(\u_cmsdk_mcu/HWDATA [11]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n91 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_altfuncset [11]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2550 (
    .a(\u_cmsdk_mcu/HWDATA [11]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n46 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_doutenset [11]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2551 (
    .a(\u_cmsdk_mcu/HWDATA [11]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n226 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpolset [11]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2552 (
    .a(\u_cmsdk_mcu/HWDATA [11]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n181 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttypeset [11]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2553 (
    .a(\u_cmsdk_mcu/HWDATA [11]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n136 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intenset [11]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2554 (
    .a(\u_cmsdk_mcu/HWDATA [11]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n91 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_altfuncset [11]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2555 (
    .a(\u_cmsdk_mcu/HWDATA [11]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n46 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_doutenset [11]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u2556 (
    .a(\u_cmsdk_mcu/HWDATA [11]),
    .b(\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [10]),
    .c(\u_cmsdk_mcu/flash_hrdata [11]),
    .o(\u_cmsdk_mcu/u_ahb_rom/n13 [11]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2557 (
    .a(\u_cmsdk_mcu/HWDATA [11]),
    .b(\u_cmsdk_mcu/sram_hrdata [11]),
    .c(\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [10]),
    .o(\u_cmsdk_mcu/u_ahb_ram/n13 [11]));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(B*A))"),
    .INIT(8'hf8))
    _al_u2558 (
    .a(\u_cmsdk_mcu/HWDATA [3]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intclr_normal_write0 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_masked_int [3]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n277 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2559 (
    .a(\u_cmsdk_mcu/HWDATA [3]),
    .b(_al_u2476_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n240 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2560 (
    .a(\u_cmsdk_mcu/HWDATA [3]),
    .b(_al_u2478_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n195 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2561 (
    .a(\u_cmsdk_mcu/HWDATA [3]),
    .b(_al_u2480_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n150 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2562 (
    .a(\u_cmsdk_mcu/HWDATA [3]),
    .b(_al_u2482_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n105 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2563 (
    .a(\u_cmsdk_mcu/HWDATA [3]),
    .b(_al_u2484_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n60 ));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(B*A))"),
    .INIT(8'hf8))
    _al_u2564 (
    .a(\u_cmsdk_mcu/HWDATA [3]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intclr_normal_write0 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/new_masked_int [3]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n277 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2565 (
    .a(\u_cmsdk_mcu/HWDATA [3]),
    .b(_al_u2488_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n240 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2566 (
    .a(\u_cmsdk_mcu/HWDATA [3]),
    .b(_al_u2490_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n195 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2567 (
    .a(\u_cmsdk_mcu/HWDATA [3]),
    .b(_al_u2492_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n150 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2568 (
    .a(\u_cmsdk_mcu/HWDATA [3]),
    .b(_al_u2494_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n105 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2569 (
    .a(\u_cmsdk_mcu/HWDATA [3]),
    .b(_al_u2496_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n60 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2570 (
    .a(\u_cmsdk_mcu/HWDATA [12]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n226 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpolset [12]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2571 (
    .a(\u_cmsdk_mcu/HWDATA [12]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n181 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttypeset [12]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2572 (
    .a(\u_cmsdk_mcu/HWDATA [12]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n136 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intenset [12]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2573 (
    .a(\u_cmsdk_mcu/HWDATA [12]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n91 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_altfuncset [12]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2574 (
    .a(\u_cmsdk_mcu/HWDATA [12]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n46 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_doutenset [12]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2575 (
    .a(\u_cmsdk_mcu/HWDATA [12]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n226 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpolset [12]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2576 (
    .a(\u_cmsdk_mcu/HWDATA [12]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n181 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttypeset [12]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2577 (
    .a(\u_cmsdk_mcu/HWDATA [12]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n136 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intenset [12]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2578 (
    .a(\u_cmsdk_mcu/HWDATA [12]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n91 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_altfuncset [12]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2579 (
    .a(\u_cmsdk_mcu/HWDATA [12]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n46 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_doutenset [12]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u2580 (
    .a(\u_cmsdk_mcu/HWDATA [12]),
    .b(\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [10]),
    .c(\u_cmsdk_mcu/flash_hrdata [12]),
    .o(\u_cmsdk_mcu/u_ahb_rom/n13 [12]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2581 (
    .a(\u_cmsdk_mcu/HWDATA [12]),
    .b(\u_cmsdk_mcu/sram_hrdata [12]),
    .c(\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [10]),
    .o(\u_cmsdk_mcu/u_ahb_ram/n13 [12]));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(B*A))"),
    .INIT(8'hf8))
    _al_u2582 (
    .a(\u_cmsdk_mcu/HWDATA [4]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intclr_normal_write0 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_masked_int [4]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n279 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2583 (
    .a(\u_cmsdk_mcu/HWDATA [4]),
    .b(_al_u2476_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n242 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2584 (
    .a(\u_cmsdk_mcu/HWDATA [4]),
    .b(_al_u2478_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n197 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2585 (
    .a(\u_cmsdk_mcu/HWDATA [4]),
    .b(_al_u2480_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n152 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2586 (
    .a(\u_cmsdk_mcu/HWDATA [4]),
    .b(_al_u2482_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n107 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2587 (
    .a(\u_cmsdk_mcu/HWDATA [4]),
    .b(_al_u2484_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n62 ));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(B*A))"),
    .INIT(8'hf8))
    _al_u2588 (
    .a(\u_cmsdk_mcu/HWDATA [4]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intclr_normal_write0 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/new_masked_int [4]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n279 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2589 (
    .a(\u_cmsdk_mcu/HWDATA [4]),
    .b(_al_u2488_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n242 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2590 (
    .a(\u_cmsdk_mcu/HWDATA [4]),
    .b(_al_u2490_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n197 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2591 (
    .a(\u_cmsdk_mcu/HWDATA [4]),
    .b(_al_u2492_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n152 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2592 (
    .a(\u_cmsdk_mcu/HWDATA [4]),
    .b(_al_u2494_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n107 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2593 (
    .a(\u_cmsdk_mcu/HWDATA [4]),
    .b(_al_u2496_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n62 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2594 (
    .a(\u_cmsdk_mcu/HWDATA [13]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n226 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpolset [13]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2595 (
    .a(\u_cmsdk_mcu/HWDATA [13]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n181 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttypeset [13]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2596 (
    .a(\u_cmsdk_mcu/HWDATA [13]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n136 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intenset [13]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2597 (
    .a(\u_cmsdk_mcu/HWDATA [13]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n91 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_altfuncset [13]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2598 (
    .a(\u_cmsdk_mcu/HWDATA [13]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n46 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_doutenset [13]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2599 (
    .a(\u_cmsdk_mcu/HWDATA [13]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n226 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpolset [13]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2600 (
    .a(\u_cmsdk_mcu/HWDATA [13]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n181 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttypeset [13]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2601 (
    .a(\u_cmsdk_mcu/HWDATA [13]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n136 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intenset [13]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2602 (
    .a(\u_cmsdk_mcu/HWDATA [13]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n91 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_altfuncset [13]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2603 (
    .a(\u_cmsdk_mcu/HWDATA [13]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n46 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_doutenset [13]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u2604 (
    .a(\u_cmsdk_mcu/HWDATA [13]),
    .b(\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [10]),
    .c(\u_cmsdk_mcu/flash_hrdata [13]),
    .o(\u_cmsdk_mcu/u_ahb_rom/n13 [13]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2605 (
    .a(\u_cmsdk_mcu/HWDATA [13]),
    .b(\u_cmsdk_mcu/sram_hrdata [13]),
    .c(\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [10]),
    .o(\u_cmsdk_mcu/u_ahb_ram/n13 [13]));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(B*A))"),
    .INIT(8'hf8))
    _al_u2606 (
    .a(\u_cmsdk_mcu/HWDATA [5]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intclr_normal_write0 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_masked_int [5]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n281 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2607 (
    .a(\u_cmsdk_mcu/HWDATA [5]),
    .b(_al_u2476_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n244 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2608 (
    .a(\u_cmsdk_mcu/HWDATA [5]),
    .b(_al_u2478_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n199 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2609 (
    .a(\u_cmsdk_mcu/HWDATA [5]),
    .b(_al_u2480_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n154 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2610 (
    .a(\u_cmsdk_mcu/HWDATA [5]),
    .b(_al_u2482_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n109 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2611 (
    .a(\u_cmsdk_mcu/HWDATA [5]),
    .b(_al_u2484_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n64 ));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(B*A))"),
    .INIT(8'hf8))
    _al_u2612 (
    .a(\u_cmsdk_mcu/HWDATA [5]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intclr_normal_write0 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/new_masked_int [5]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n281 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2613 (
    .a(\u_cmsdk_mcu/HWDATA [5]),
    .b(_al_u2488_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n244 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2614 (
    .a(\u_cmsdk_mcu/HWDATA [5]),
    .b(_al_u2490_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n199 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2615 (
    .a(\u_cmsdk_mcu/HWDATA [5]),
    .b(_al_u2492_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n154 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2616 (
    .a(\u_cmsdk_mcu/HWDATA [5]),
    .b(_al_u2494_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n109 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2617 (
    .a(\u_cmsdk_mcu/HWDATA [5]),
    .b(_al_u2496_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n64 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2618 (
    .a(\u_cmsdk_mcu/HWDATA [14]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n226 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpolset [14]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2619 (
    .a(\u_cmsdk_mcu/HWDATA [14]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n181 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttypeset [14]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2620 (
    .a(\u_cmsdk_mcu/HWDATA [14]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n136 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intenset [14]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2621 (
    .a(\u_cmsdk_mcu/HWDATA [14]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n91 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_altfuncset [14]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2622 (
    .a(\u_cmsdk_mcu/HWDATA [14]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n46 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_doutenset [14]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2623 (
    .a(\u_cmsdk_mcu/HWDATA [14]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n226 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpolset [14]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2624 (
    .a(\u_cmsdk_mcu/HWDATA [14]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n181 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttypeset [14]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2625 (
    .a(\u_cmsdk_mcu/HWDATA [14]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n136 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intenset [14]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2626 (
    .a(\u_cmsdk_mcu/HWDATA [14]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n91 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_altfuncset [14]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2627 (
    .a(\u_cmsdk_mcu/HWDATA [14]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n46 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_doutenset [14]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u2628 (
    .a(\u_cmsdk_mcu/HWDATA [14]),
    .b(\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [10]),
    .c(\u_cmsdk_mcu/flash_hrdata [14]),
    .o(\u_cmsdk_mcu/u_ahb_rom/n13 [14]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2629 (
    .a(\u_cmsdk_mcu/HWDATA [14]),
    .b(\u_cmsdk_mcu/sram_hrdata [14]),
    .c(\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [10]),
    .o(\u_cmsdk_mcu/u_ahb_ram/n13 [14]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u263 (
    .a(\u_cmsdk_mcu/p1_out [0]),
    .b(\u_cmsdk_mcu/p1_outen [0]),
    .o(\u_cmsdk_mcu/p1_in [0]));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(B*A))"),
    .INIT(8'hf8))
    _al_u2630 (
    .a(\u_cmsdk_mcu/HWDATA [6]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intclr_normal_write0 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_masked_int [6]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n283 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2631 (
    .a(\u_cmsdk_mcu/HWDATA [6]),
    .b(_al_u2476_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n246 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2632 (
    .a(\u_cmsdk_mcu/HWDATA [6]),
    .b(_al_u2478_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n201 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2633 (
    .a(\u_cmsdk_mcu/HWDATA [6]),
    .b(_al_u2480_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n156 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2634 (
    .a(\u_cmsdk_mcu/HWDATA [6]),
    .b(_al_u2482_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n111 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2635 (
    .a(\u_cmsdk_mcu/HWDATA [6]),
    .b(_al_u2484_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n66 ));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(B*A))"),
    .INIT(8'hf8))
    _al_u2636 (
    .a(\u_cmsdk_mcu/HWDATA [6]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intclr_normal_write0 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/new_masked_int [6]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n283 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2637 (
    .a(\u_cmsdk_mcu/HWDATA [6]),
    .b(_al_u2488_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n246 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2638 (
    .a(\u_cmsdk_mcu/HWDATA [6]),
    .b(_al_u2490_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n201 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2639 (
    .a(\u_cmsdk_mcu/HWDATA [6]),
    .b(_al_u2492_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n156 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u264 (
    .a(\u_cmsdk_mcu/p1_out [10]),
    .b(\u_cmsdk_mcu/p1_outen [10]),
    .o(\u_cmsdk_mcu/p1_in [10]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2640 (
    .a(\u_cmsdk_mcu/HWDATA [6]),
    .b(_al_u2494_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n111 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2641 (
    .a(\u_cmsdk_mcu/HWDATA [6]),
    .b(_al_u2496_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n66 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u2642 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kc6ju6 ),
    .b(_al_u2399_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jckax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ubypw6 ),
    .o(_al_u2642_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*~B))"),
    .INIT(8'h8a))
    _al_u2643 (
    .a(_al_u2642_o),
    .b(_al_u1952_o),
    .c(_al_u2412_o),
    .o(_al_u2643_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*B)*~(~D*A))"),
    .INIT(16'hf351))
    _al_u2644 (
    .a(_al_u682_o),
    .b(_al_u1907_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ),
    .o(_al_u2644_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2645 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yi7ju6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(A*~(~B*~(~D*~C)))"),
    .INIT(16'h888a))
    _al_u2646 (
    .a(_al_u1658_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yi7ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 ),
    .o(_al_u2646_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u2647 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 ),
    .o(_al_u2647_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(~A*~(~C*B)))"),
    .INIT(16'hae00))
    _al_u2648 (
    .a(_al_u682_o),
    .b(_al_u2647_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 ),
    .o(_al_u2648_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~B*~(~D*~A))"),
    .INIT(16'h0302))
    _al_u2649 (
    .a(_al_u2644_o),
    .b(_al_u2646_o),
    .c(_al_u2648_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 ),
    .o(_al_u2649_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u265 (
    .a(\u_cmsdk_mcu/p1_out [11]),
    .b(\u_cmsdk_mcu/p1_outen [11]),
    .o(\u_cmsdk_mcu/p1_in [11]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*~A))"),
    .INIT(8'h23))
    _al_u2650 (
    .a(_al_u2649_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zf7ju6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vgjpw6 ),
    .o(_al_u2650_o));
  AL_MAP_LUT4 #(
    .EQN("~(B@(A*~(D*~C)))"),
    .INIT(16'h9399))
    _al_u2651 (
    .a(_al_u2643_o),
    .b(_al_u2398_o),
    .c(_al_u2650_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Umkax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E2epw6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2652 (
    .a(\u_cmsdk_mcu/HWDATA [15]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C1wpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fsdiu6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2653 (
    .a(\u_cmsdk_mcu/HWDATA [15]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n226 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpolset [15]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2654 (
    .a(\u_cmsdk_mcu/HWDATA [15]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n181 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttypeset [15]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2655 (
    .a(\u_cmsdk_mcu/HWDATA [15]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n136 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intenset [15]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2656 (
    .a(\u_cmsdk_mcu/HWDATA [15]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n91 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_altfuncset [15]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2657 (
    .a(\u_cmsdk_mcu/HWDATA [15]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n46 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_doutenset [15]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2658 (
    .a(\u_cmsdk_mcu/HWDATA [15]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n226 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpolset [15]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2659 (
    .a(\u_cmsdk_mcu/HWDATA [15]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n181 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttypeset [15]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u266 (
    .a(\u_cmsdk_mcu/p1_out [12]),
    .b(\u_cmsdk_mcu/p1_outen [12]),
    .o(\u_cmsdk_mcu/p1_in [12]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2660 (
    .a(\u_cmsdk_mcu/HWDATA [15]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n136 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intenset [15]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2661 (
    .a(\u_cmsdk_mcu/HWDATA [15]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n91 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_altfuncset [15]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2662 (
    .a(\u_cmsdk_mcu/HWDATA [15]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n46 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_doutenset [15]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u2663 (
    .a(\u_cmsdk_mcu/HWDATA [15]),
    .b(\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [10]),
    .c(\u_cmsdk_mcu/flash_hrdata [15]),
    .o(\u_cmsdk_mcu/u_ahb_rom/n13 [15]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2664 (
    .a(\u_cmsdk_mcu/HWDATA [15]),
    .b(\u_cmsdk_mcu/sram_hrdata [15]),
    .c(\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [10]),
    .o(\u_cmsdk_mcu/u_ahb_ram/n13 [15]));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(B*A))"),
    .INIT(8'hf8))
    _al_u2665 (
    .a(\u_cmsdk_mcu/HWDATA [7]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intclr_normal_write0 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_masked_int [7]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n285 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2666 (
    .a(\u_cmsdk_mcu/HWDATA [7]),
    .b(_al_u2476_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n248 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2667 (
    .a(\u_cmsdk_mcu/HWDATA [7]),
    .b(_al_u2478_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n203 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2668 (
    .a(\u_cmsdk_mcu/HWDATA [7]),
    .b(_al_u2480_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n158 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2669 (
    .a(\u_cmsdk_mcu/HWDATA [7]),
    .b(_al_u2482_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n113 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u267 (
    .a(\u_cmsdk_mcu/p1_out [13]),
    .b(\u_cmsdk_mcu/p1_outen [13]),
    .o(\u_cmsdk_mcu/p1_in [13]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2670 (
    .a(\u_cmsdk_mcu/HWDATA [7]),
    .b(_al_u2484_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n68 ));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(B*A))"),
    .INIT(8'hf8))
    _al_u2671 (
    .a(\u_cmsdk_mcu/HWDATA [7]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intclr_normal_write0 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/new_masked_int [7]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n285 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2672 (
    .a(\u_cmsdk_mcu/HWDATA [7]),
    .b(_al_u2488_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n248 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2673 (
    .a(\u_cmsdk_mcu/HWDATA [7]),
    .b(_al_u2490_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n203 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2674 (
    .a(\u_cmsdk_mcu/HWDATA [7]),
    .b(_al_u2492_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n158 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2675 (
    .a(\u_cmsdk_mcu/HWDATA [7]),
    .b(_al_u2494_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n113 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2676 (
    .a(\u_cmsdk_mcu/HWDATA [7]),
    .b(_al_u2496_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n68 ));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u2677 (
    .a(\u_cmsdk_mcu/HWDATA [17]),
    .b(\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [16]),
    .c(\u_cmsdk_mcu/flash_hrdata [17]),
    .o(\u_cmsdk_mcu/u_ahb_rom/n13 [17]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2678 (
    .a(\u_cmsdk_mcu/HWDATA [17]),
    .b(\u_cmsdk_mcu/sram_hrdata [17]),
    .c(\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [16]),
    .o(\u_cmsdk_mcu/u_ahb_ram/n13 [17]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    _al_u2679 (
    .a(\u_cmsdk_mcu/HWDATA [1]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/intr_stat_set [1]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/write_enable0c ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n117 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u268 (
    .a(\u_cmsdk_mcu/p1_out [14]),
    .b(\u_cmsdk_mcu/p1_outen [14]),
    .o(\u_cmsdk_mcu/p1_in [14]));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(B*A))"),
    .INIT(8'hf8))
    _al_u2680 (
    .a(\u_cmsdk_mcu/HWDATA [1]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intclr_normal_write0 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_masked_int [1]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n273 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2681 (
    .a(\u_cmsdk_mcu/HWDATA [1]),
    .b(_al_u2476_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n236 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2682 (
    .a(\u_cmsdk_mcu/HWDATA [1]),
    .b(_al_u2478_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n191 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2683 (
    .a(\u_cmsdk_mcu/HWDATA [1]),
    .b(_al_u2480_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n146 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2684 (
    .a(\u_cmsdk_mcu/HWDATA [1]),
    .b(_al_u2482_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n101 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2685 (
    .a(\u_cmsdk_mcu/HWDATA [1]),
    .b(_al_u2484_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n56 ));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(B*A))"),
    .INIT(8'hf8))
    _al_u2686 (
    .a(\u_cmsdk_mcu/HWDATA [1]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intclr_normal_write0 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/new_masked_int [1]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n273 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2687 (
    .a(\u_cmsdk_mcu/HWDATA [1]),
    .b(_al_u2488_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n236 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2688 (
    .a(\u_cmsdk_mcu/HWDATA [1]),
    .b(_al_u2490_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n191 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2689 (
    .a(\u_cmsdk_mcu/HWDATA [1]),
    .b(_al_u2492_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n146 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u269 (
    .a(\u_cmsdk_mcu/p1_out [15]),
    .b(\u_cmsdk_mcu/p1_outen [15]),
    .o(\u_cmsdk_mcu/p1_in [15]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2690 (
    .a(\u_cmsdk_mcu/HWDATA [1]),
    .b(_al_u2494_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n101 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2691 (
    .a(\u_cmsdk_mcu/HWDATA [1]),
    .b(_al_u2496_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n56 ));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(B*A))"),
    .INIT(8'hf8))
    _al_u2692 (
    .a(\u_cmsdk_mcu/HWDATA [9]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intclr_normal_write1 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_masked_int [9]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n289 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2693 (
    .a(\u_cmsdk_mcu/HWDATA [9]),
    .b(_al_u2500_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n252 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2694 (
    .a(\u_cmsdk_mcu/HWDATA [9]),
    .b(_al_u2502_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n207 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2695 (
    .a(\u_cmsdk_mcu/HWDATA [9]),
    .b(_al_u2504_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n162 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2696 (
    .a(\u_cmsdk_mcu/HWDATA [9]),
    .b(_al_u2506_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n117 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2697 (
    .a(\u_cmsdk_mcu/HWDATA [9]),
    .b(_al_u2508_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n72 ));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(B*A))"),
    .INIT(8'hf8))
    _al_u2698 (
    .a(\u_cmsdk_mcu/HWDATA [9]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intclr_normal_write1 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/new_masked_int [9]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n289 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2699 (
    .a(\u_cmsdk_mcu/HWDATA [9]),
    .b(_al_u2512_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n252 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u270 (
    .a(\u_cmsdk_mcu/p1_out [2]),
    .b(\u_cmsdk_mcu/p1_outen [2]),
    .o(\u_cmsdk_mcu/p1_in [2]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2700 (
    .a(\u_cmsdk_mcu/HWDATA [9]),
    .b(_al_u2514_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n207 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2701 (
    .a(\u_cmsdk_mcu/HWDATA [9]),
    .b(_al_u2516_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n162 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2702 (
    .a(\u_cmsdk_mcu/HWDATA [9]),
    .b(_al_u2518_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n117 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2703 (
    .a(\u_cmsdk_mcu/HWDATA [9]),
    .b(_al_u2520_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n72 ));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u2704 (
    .a(\u_cmsdk_mcu/HWDATA [18]),
    .b(\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [16]),
    .c(\u_cmsdk_mcu/flash_hrdata [18]),
    .o(\u_cmsdk_mcu/u_ahb_rom/n13 [18]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2705 (
    .a(\u_cmsdk_mcu/HWDATA [18]),
    .b(\u_cmsdk_mcu/sram_hrdata [18]),
    .c(\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [16]),
    .o(\u_cmsdk_mcu/u_ahb_ram/n13 [18]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u2706 (
    .a(\u_cmsdk_mcu/HWDATA [19]),
    .b(\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [16]),
    .c(\u_cmsdk_mcu/flash_hrdata [19]),
    .o(\u_cmsdk_mcu/u_ahb_rom/n13 [19]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2707 (
    .a(\u_cmsdk_mcu/HWDATA [19]),
    .b(\u_cmsdk_mcu/sram_hrdata [19]),
    .c(\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [16]),
    .o(\u_cmsdk_mcu/u_ahb_ram/n13 [19]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u2708 (
    .a(\u_cmsdk_mcu/HWDATA [20]),
    .b(\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [16]),
    .c(\u_cmsdk_mcu/flash_hrdata [20]),
    .o(\u_cmsdk_mcu/u_ahb_rom/n13 [20]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2709 (
    .a(\u_cmsdk_mcu/HWDATA [20]),
    .b(\u_cmsdk_mcu/sram_hrdata [20]),
    .c(\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [16]),
    .o(\u_cmsdk_mcu/u_ahb_ram/n13 [20]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u271 (
    .a(\u_cmsdk_mcu/p1_out [4]),
    .b(\u_cmsdk_mcu/p1_outen [4]),
    .o(\u_cmsdk_mcu/p1_in [4]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u2710 (
    .a(\u_cmsdk_mcu/HWDATA [21]),
    .b(\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [16]),
    .c(\u_cmsdk_mcu/flash_hrdata [21]),
    .o(\u_cmsdk_mcu/u_ahb_rom/n13 [21]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2711 (
    .a(\u_cmsdk_mcu/HWDATA [21]),
    .b(\u_cmsdk_mcu/sram_hrdata [21]),
    .c(\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [16]),
    .o(\u_cmsdk_mcu/u_ahb_ram/n13 [21]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u2712 (
    .a(\u_cmsdk_mcu/HWDATA [22]),
    .b(\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [16]),
    .c(\u_cmsdk_mcu/flash_hrdata [22]),
    .o(\u_cmsdk_mcu/u_ahb_rom/n13 [22]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2713 (
    .a(\u_cmsdk_mcu/HWDATA [22]),
    .b(\u_cmsdk_mcu/sram_hrdata [22]),
    .c(\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [16]),
    .o(\u_cmsdk_mcu/u_ahb_ram/n13 [22]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u2714 (
    .a(\u_cmsdk_mcu/HWDATA [23]),
    .b(\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [16]),
    .c(\u_cmsdk_mcu/flash_hrdata [23]),
    .o(\u_cmsdk_mcu/u_ahb_rom/n13 [23]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2715 (
    .a(\u_cmsdk_mcu/HWDATA [23]),
    .b(\u_cmsdk_mcu/sram_hrdata [23]),
    .c(\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [16]),
    .o(\u_cmsdk_mcu/u_ahb_ram/n13 [23]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(C*~A))"),
    .INIT(16'h8caf))
    _al_u2716 (
    .a(_al_u2439_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cz7ju6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gdqow6 ),
    .d(_al_u2272_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iexow6 ));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(D*C))"),
    .INIT(16'h0444))
    _al_u2717 (
    .a(_al_u1891_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iexow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D84iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wvgax6 ),
    .o(_al_u2717_o));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    _al_u2718 (
    .a(_al_u2717_o),
    .b(\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [24]),
    .c(\u_cmsdk_mcu/flash_hrdata [24]),
    .o(\u_cmsdk_mcu/u_ahb_rom/n13 [24]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'h5c))
    _al_u2719 (
    .a(_al_u2717_o),
    .b(\u_cmsdk_mcu/sram_hrdata [24]),
    .c(\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [24]),
    .o(\u_cmsdk_mcu/u_ahb_ram/n13 [24]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u272 (
    .a(\u_cmsdk_mcu/p1_out [6]),
    .b(\u_cmsdk_mcu/p1_outen [6]),
    .o(\u_cmsdk_mcu/p1_in [6]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*~B)*~(D*~A))"),
    .INIT(16'h8acf))
    _al_u2720 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I28ju6 ),
    .b(_al_u2261_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gdqow6 ),
    .d(_al_u2272_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Awwow6 ));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(D*C))"),
    .INIT(16'h0444))
    _al_u2721 (
    .a(_al_u1971_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Awwow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K84iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wvgax6 ),
    .o(_al_u2721_o));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    _al_u2722 (
    .a(_al_u2721_o),
    .b(\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [24]),
    .c(\u_cmsdk_mcu/flash_hrdata [25]),
    .o(\u_cmsdk_mcu/u_ahb_rom/n13 [25]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'h5c))
    _al_u2723 (
    .a(_al_u2721_o),
    .b(\u_cmsdk_mcu/sram_hrdata [25]),
    .c(\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [24]),
    .o(\u_cmsdk_mcu/u_ahb_ram/n13 [25]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*C)*~(B*~A))"),
    .INIT(16'h0bbb))
    _al_u2724 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ka8ju6 ),
    .b(_al_u2272_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R84iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wvgax6 ),
    .o(_al_u2724_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*~(D*~B))"),
    .INIT(16'h4050))
    _al_u2725 (
    .a(_al_u2032_o),
    .b(_al_u2455_o),
    .c(_al_u2724_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gdqow6 ),
    .o(_al_u2725_o));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    _al_u2726 (
    .a(_al_u2725_o),
    .b(\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [24]),
    .c(\u_cmsdk_mcu/flash_hrdata [26]),
    .o(\u_cmsdk_mcu/u_ahb_rom/n13 [26]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'h5c))
    _al_u2727 (
    .a(_al_u2725_o),
    .b(\u_cmsdk_mcu/sram_hrdata [26]),
    .c(\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [24]),
    .o(\u_cmsdk_mcu/u_ahb_ram/n13 [26]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*C)*~(B*~A))"),
    .INIT(16'h0bbb))
    _al_u2728 (
    .a(_al_u2062_o),
    .b(_al_u2272_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y84iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wvgax6 ),
    .o(_al_u2728_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*~(D*~B))"),
    .INIT(16'h4050))
    _al_u2729 (
    .a(_al_u2055_o),
    .b(_al_u2447_o),
    .c(_al_u2728_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gdqow6 ),
    .o(_al_u2729_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u273 (
    .a(\u_cmsdk_mcu/p1_out [7]),
    .b(\u_cmsdk_mcu/p1_outen [7]),
    .o(\u_cmsdk_mcu/p1_in [7]));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    _al_u2730 (
    .a(_al_u2729_o),
    .b(\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [24]),
    .c(\u_cmsdk_mcu/flash_hrdata [27]),
    .o(\u_cmsdk_mcu/u_ahb_rom/n13 [27]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'h5c))
    _al_u2731 (
    .a(_al_u2729_o),
    .b(\u_cmsdk_mcu/sram_hrdata [27]),
    .c(\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [24]),
    .o(\u_cmsdk_mcu/u_ahb_ram/n13 [27]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*C)*~(B*~A))"),
    .INIT(16'h0bbb))
    _al_u2732 (
    .a(_al_u2420_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gdqow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F94iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wvgax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W1wow6 ));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(D*~C))"),
    .INIT(16'h4044))
    _al_u2733 (
    .a(_al_u2077_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W1wow6 ),
    .c(_al_u2084_o),
    .d(_al_u2272_o),
    .o(_al_u2733_o));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    _al_u2734 (
    .a(_al_u2733_o),
    .b(\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [24]),
    .c(\u_cmsdk_mcu/flash_hrdata [28]),
    .o(\u_cmsdk_mcu/u_ahb_rom/n13 [28]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'h5c))
    _al_u2735 (
    .a(_al_u2733_o),
    .b(\u_cmsdk_mcu/sram_hrdata [28]),
    .c(\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [24]),
    .o(\u_cmsdk_mcu/u_ahb_ram/n13 [28]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u2736 (
    .a(\u_cmsdk_mcu/HWDATA [30]),
    .b(\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [24]),
    .c(\u_cmsdk_mcu/flash_hrdata [30]),
    .o(\u_cmsdk_mcu/u_ahb_rom/n13 [30]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2737 (
    .a(\u_cmsdk_mcu/HWDATA [30]),
    .b(\u_cmsdk_mcu/sram_hrdata [30]),
    .c(\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [24]),
    .o(\u_cmsdk_mcu/u_ahb_ram/n13 [30]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u2738 (
    .a(\u_cmsdk_mcu/HWDATA [31]),
    .b(\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [24]),
    .c(\u_cmsdk_mcu/flash_hrdata [31]),
    .o(\u_cmsdk_mcu/u_ahb_rom/n13 [31]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2739 (
    .a(\u_cmsdk_mcu/HWDATA [31]),
    .b(\u_cmsdk_mcu/sram_hrdata [31]),
    .c(\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [24]),
    .o(\u_cmsdk_mcu/u_ahb_ram/n13 [31]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u274 (
    .a(\u_cmsdk_mcu/p1_out [8]),
    .b(\u_cmsdk_mcu/p1_outen [8]),
    .o(\u_cmsdk_mcu/p1_in [8]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*C)*~(~B*A))"),
    .INIT(16'h0ddd))
    _al_u2740 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gdqow6 ),
    .b(_al_u2429_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M94iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wvgax6 ),
    .o(_al_u2740_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*~(D*~B))"),
    .INIT(16'h4050))
    _al_u2741 (
    .a(_al_u2099_o),
    .b(_al_u2106_o),
    .c(_al_u2740_o),
    .d(_al_u2272_o),
    .o(_al_u2741_o));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    _al_u2742 (
    .a(_al_u2741_o),
    .b(\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [24]),
    .c(\u_cmsdk_mcu/flash_hrdata [29]),
    .o(\u_cmsdk_mcu/u_ahb_rom/n13 [29]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'h5c))
    _al_u2743 (
    .a(_al_u2741_o),
    .b(\u_cmsdk_mcu/sram_hrdata [29]),
    .c(\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [24]),
    .o(\u_cmsdk_mcu/u_ahb_ram/n13 [29]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u2744 (
    .a(\u_cmsdk_mcu/HWDATA [16]),
    .b(\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [16]),
    .c(\u_cmsdk_mcu/flash_hrdata [16]),
    .o(\u_cmsdk_mcu/u_ahb_rom/n13 [16]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2745 (
    .a(\u_cmsdk_mcu/HWDATA [16]),
    .b(\u_cmsdk_mcu/sram_hrdata [16]),
    .c(\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [16]),
    .o(\u_cmsdk_mcu/u_ahb_ram/n13 [16]));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(~B*~(D*~C)))"),
    .INIT(16'h4544))
    _al_u2746 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iekax6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lgkax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oikax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rkkax6 ),
    .o(_al_u2746_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(~D*C*A))"),
    .INIT(16'h3313))
    _al_u2747 (
    .a(_al_u916_o),
    .b(_al_u2746_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fkrpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ubypw6 ),
    .o(_al_u2747_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(C*~(D*A)))"),
    .INIT(16'h8c0c))
    _al_u2748 (
    .a(_al_u1765_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L45iu6_lutinv ),
    .c(_al_u2747_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V6jax6 ),
    .o(_al_u2748_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u2749 (
    .a(_al_u696_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A95iu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iekax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wfspw6 ),
    .o(_al_u2749_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u275 (
    .a(\u_cmsdk_mcu/p1_out [9]),
    .b(\u_cmsdk_mcu/p1_outen [9]),
    .o(\u_cmsdk_mcu/p1_in [9]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u2750 (
    .a(_al_u912_o),
    .b(_al_u2749_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4jax6 ),
    .o(_al_u2750_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u2751 (
    .a(_al_u2750_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K75iu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wkipw6 ),
    .o(_al_u2751_o));
  AL_MAP_LUT3 #(
    .EQN("~(C*~B*A)"),
    .INIT(8'hdf))
    _al_u2752 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gpyiu6 ),
    .b(_al_u2748_o),
    .c(_al_u2751_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jn7ow6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u2753 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Llaow6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U98iu6 ));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u2754 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U98iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 ),
    .o(_al_u2754_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*~B*A)"),
    .INIT(16'h0020))
    _al_u2755 (
    .a(_al_u2365_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 ),
    .o(_al_u2755_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~A*~(~D*B))"),
    .INIT(16'h0501))
    _al_u2756 (
    .a(_al_u2754_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qe8iu6_lutinv ),
    .c(_al_u2755_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 ),
    .o(_al_u2756_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(~A*~(~C*B)))"),
    .INIT(16'hae00))
    _al_u2757 (
    .a(_al_u1782_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D6kiu6_lutinv ),
    .c(_al_u1271_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzjpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tc8iu6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u2758 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yljiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 ),
    .o(_al_u2758_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*A*~(D*~B))"),
    .INIT(16'h080a))
    _al_u2759 (
    .a(_al_u903_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Irmpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 ),
    .o(_al_u2759_o));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    _al_u276 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qwfax6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Utqpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n267 ));
  AL_MAP_LUT4 #(
    .EQN("(~D*~A*~(C*B))"),
    .INIT(16'h0015))
    _al_u2760 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bi0iu6 ),
    .b(_al_u681_o),
    .c(_al_u2758_o),
    .d(_al_u2759_o),
    .o(_al_u2760_o));
  AL_MAP_LUT4 #(
    .EQN("(C*A*~(D*B))"),
    .INIT(16'h20a0))
    _al_u2761 (
    .a(_al_u2756_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tc8iu6 ),
    .c(_al_u2760_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xdspw6 ),
    .o(_al_u2761_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u2762 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kxziu6_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2763 (
    .a(_al_u2365_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kxziu6_lutinv ),
    .o(_al_u2763_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2764 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P14qw6 ),
    .o(_al_u2764_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2765 (
    .a(_al_u2764_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bziiu6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(~A*~(~C*B)))"),
    .INIT(16'h00ae))
    _al_u2766 (
    .a(_al_u2763_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bziiu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9ypw6 ),
    .o(_al_u2766_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u2767 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Skjax6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9ypw6 ),
    .o(_al_u2767_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    _al_u2768 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nbkiu6_lutinv ),
    .c(_al_u2767_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M7kiu6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u2769 (
    .a(_al_u2766_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M7kiu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hd8iu6_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u277 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E8iax6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzjpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vnfpw6 [0]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2770 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P14qw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 ),
    .o(_al_u2770_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2771 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kxziu6_lutinv ),
    .b(_al_u2770_o),
    .o(_al_u2771_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u2772 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J9kiu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P14qw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Skjax6 ),
    .o(_al_u2772_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(~B*~(D*~C)))"),
    .INIT(16'h8a88))
    _al_u2773 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kxziu6_lutinv ),
    .b(_al_u2772_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujiu6 ),
    .d(_al_u2770_o),
    .o(_al_u2773_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*~A)"),
    .INIT(8'h04))
    _al_u2774 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv ),
    .b(_al_u909_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 ),
    .o(_al_u2774_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u2775 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9ypw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nyiiu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D*C*A))"),
    .INIT(16'h1333))
    _al_u2776 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ia8iu6_lutinv ),
    .b(_al_u2774_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nbkiu6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nyiiu6 ),
    .o(_al_u2776_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~B*~(~D*A))"),
    .INIT(16'h3010))
    _al_u2777 (
    .a(_al_u2771_o),
    .b(_al_u2773_o),
    .c(_al_u2776_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yb8iu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(C*~A))"),
    .INIT(16'h8caf))
    _al_u2778 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hd8iu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yb8iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4jax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wfspw6 ),
    .o(_al_u2778_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u2779 (
    .a(_al_u607_o),
    .b(_al_u1346_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 ),
    .o(_al_u2779_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u278 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzjpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W0jax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vnfpw6 [6]));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u2780 (
    .a(_al_u2779_o),
    .b(_al_u1264_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S3kiu6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u2781 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mbhow6_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u2782 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mbhow6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 ),
    .o(_al_u2782_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*~(~D*~C)))"),
    .INIT(16'h222a))
    _al_u2783 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S3kiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I6row6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yqziu6 ),
    .d(_al_u2782_o),
    .o(_al_u2783_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(~D*~C))"),
    .INIT(16'h8880))
    _al_u2784 (
    .a(_al_u2761_o),
    .b(_al_u2778_o),
    .c(_al_u2783_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sqkax6 ),
    .o(_al_u2784_o));
  AL_MAP_LUT4 #(
    .EQN("(D@C@B@A)"),
    .INIT(16'h6996))
    _al_u2785 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Irmpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S7mpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wfspw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wkipw6 ),
    .o(_al_u2785_o));
  AL_MAP_LUT3 #(
    .EQN("(C@B@A)"),
    .INIT(8'h96))
    _al_u2786 (
    .a(_al_u2785_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jckax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jgxpw6 ),
    .o(_al_u2786_o));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    _al_u2787 (
    .a(_al_u2786_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4jax6 ),
    .o(_al_u2787_o));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    _al_u2788 (
    .a(_al_u2787_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N4kax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S88iu6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*B*A)"),
    .INIT(16'h0800))
    _al_u2789 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ia8iu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J9kiu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Skjax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 ),
    .o(_al_u2789_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u279 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzjpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W2jax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vnfpw6 [7]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D*C*A))"),
    .INIT(16'h1333))
    _al_u2790 (
    .a(_al_u2771_o),
    .b(_al_u2789_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujiu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6 ),
    .o(_al_u2790_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*(A@(D*C)))"),
    .INIT(16'h1222))
    _al_u2791 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S88iu6_lutinv ),
    .b(_al_u2790_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Skjax6 ),
    .o(_al_u2791_o));
  AL_MAP_LUT2 #(
    .EQN("~(~B*A)"),
    .INIT(4'hd))
    _al_u2792 (
    .a(_al_u2784_o),
    .b(_al_u2791_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y48iu6 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*A))"),
    .INIT(8'hc4))
    _al_u2793 (
    .a(_al_u1299_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hlliu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ubypw6 ),
    .o(_al_u2793_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    _al_u2794 (
    .a(_al_u1906_o),
    .b(_al_u2793_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rskax6 ),
    .o(_al_u2794_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(~C*~B*~A))"),
    .INIT(16'h00fe))
    _al_u2795 (
    .a(_al_u2794_o),
    .b(_al_u1643_o),
    .c(_al_u1777_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fkliu6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u2796 (
    .a(_al_u1906_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rskax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jjoiu6 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u2797 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jjoiu6 ),
    .b(_al_u1299_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ubypw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ph8iu6_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2798 (
    .a(_al_u1788_o),
    .b(_al_u609_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yi8iu6_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u2799 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ph8iu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yi8iu6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ug8iu6_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u280 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzjpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wwiax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vnfpw6 [4]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D*B*~A))"),
    .INIT(16'hb0f0))
    _al_u2800 (
    .a(_al_u1336_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vo3ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 ),
    .o(_al_u2800_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u2801 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vo3ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ly2ju6 ));
  AL_MAP_LUT3 #(
    .EQN("(~C*(B@A))"),
    .INIT(8'h06))
    _al_u2802 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 ),
    .o(_al_u2802_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~(B*A))"),
    .INIT(16'h0007))
    _al_u2803 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ldoiu6_lutinv ),
    .b(_al_u1658_o),
    .c(_al_u1817_o),
    .d(_al_u2802_o),
    .o(_al_u2803_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*~(D*B))"),
    .INIT(16'h1050))
    _al_u2804 (
    .a(_al_u2800_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ly2ju6 ),
    .c(_al_u2803_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 ),
    .o(_al_u2804_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*~A))"),
    .INIT(16'h2a3f))
    _al_u2805 (
    .a(_al_u2804_o),
    .b(_al_u932_o),
    .c(_al_u2403_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fhoiu6 ));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(B*A))"),
    .INIT(8'h07))
    _al_u2806 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ug8iu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fhoiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y5liu6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2807 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sy2ju6 ));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    _al_u2808 (
    .a(_al_u1342_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sy2ju6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 ),
    .o(_al_u2808_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*~B))"),
    .INIT(8'h8a))
    _al_u2809 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vo3ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 ),
    .o(_al_u2809_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u281 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzjpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wyiax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vnfpw6 [5]));
  AL_MAP_LUT4 #(
    .EQN("(~B*A*~(~D*~C))"),
    .INIT(16'h2220))
    _al_u2810 (
    .a(_al_u2808_o),
    .b(_al_u2809_o),
    .c(_al_u1658_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ),
    .o(_al_u2810_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2811 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D31ju6 ));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u2812 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D31ju6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nz2ju6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2813 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 ),
    .o(_al_u2813_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~A*~(D*C))"),
    .INIT(16'h0111))
    _al_u2814 (
    .a(_al_u2810_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nz2ju6 ),
    .c(_al_u932_o),
    .d(_al_u2813_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Im2ju6 ));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*~(B*~A))"),
    .INIT(16'h00b0))
    _al_u2815 (
    .a(_al_u607_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 ),
    .o(_al_u2815_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(~B*~A))"),
    .INIT(8'he0))
    _al_u2816 (
    .a(_al_u2815_o),
    .b(_al_u2387_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 ),
    .o(_al_u2816_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(~A*~(~D*B)))"),
    .INIT(16'ha0e0))
    _al_u2817 (
    .a(_al_u682_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sq3ju6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 ),
    .o(_al_u2817_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u2818 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T23ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nkaju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 ),
    .o(_al_u2818_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*A)"),
    .INIT(16'h0002))
    _al_u2819 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Im2ju6 ),
    .b(_al_u2816_o),
    .c(_al_u2817_o),
    .d(_al_u2818_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ng8iu6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u282 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzjpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuiax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vnfpw6 [3]));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(B*A))"),
    .INIT(8'h07))
    _al_u2820 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ug8iu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ng8iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zf8iu6 ));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u2821 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hgrpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9ypw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dmiiu6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2822 (
    .a(_al_u2365_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dmiiu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zyoiu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~A*(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D))"),
    .INIT(16'h4450))
    _al_u2823 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hgrpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kmiiu6 ));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(B*A))"),
    .INIT(8'h07))
    _al_u2824 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kxziu6_lutinv ),
    .b(_al_u2772_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kmiiu6 ),
    .o(_al_u2824_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*A))"),
    .INIT(8'hc4))
    _al_u2825 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zyoiu6 ),
    .b(_al_u2824_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv ),
    .o(_al_u2825_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2826 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qxoiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F6ziu6 ));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*~(D*~C)))"),
    .INIT(16'h2a22))
    _al_u2827 (
    .a(_al_u2825_o),
    .b(_al_u2771_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F6ziu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Skjax6 ),
    .o(_al_u2827_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2828 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ia8iu6_lutinv ),
    .b(_al_u2772_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mldpw6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u2829 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ),
    .o(_al_u2829_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u283 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzjpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ysiax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vnfpw6 [2]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u2830 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv ),
    .b(_al_u2829_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kubow6 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u2831 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mldpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kubow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N4kax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aaiiu6 ));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u2832 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bziiu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9ypw6 ),
    .o(_al_u2832_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u2833 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aaiiu6 ),
    .b(_al_u2832_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N4kax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K8iiu6 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*~A))"),
    .INIT(8'h8c))
    _al_u2834 (
    .a(_al_u2827_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K8iiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 ),
    .o(_al_u2834_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u2835 (
    .a(_al_u2771_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Skjax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6 ),
    .o(_al_u2835_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u2836 (
    .a(_al_u2365_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9ypw6 ),
    .o(_al_u2836_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(A*~(D*~C)))"),
    .INIT(16'h4c44))
    _al_u2837 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rwjax6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Skjax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6 ),
    .o(_al_u2837_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u2838 (
    .a(_al_u2771_o),
    .b(_al_u2836_o),
    .c(_al_u2837_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljiiu6 ));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u2839 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hgrpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9ypw6 ),
    .o(_al_u2839_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u284 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzjpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zqiax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vnfpw6 [1]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*~B))"),
    .INIT(8'ha8))
    _al_u2840 (
    .a(_al_u2839_o),
    .b(_al_u2373_o),
    .c(_al_u2770_o),
    .o(_al_u2840_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*~A)"),
    .INIT(16'h0004))
    _al_u2841 (
    .a(_al_u2835_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljiiu6 ),
    .c(_al_u2763_o),
    .d(_al_u2840_o),
    .o(_al_u2841_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*~B))"),
    .INIT(8'h75))
    _al_u2842 (
    .a(_al_u2834_o),
    .b(_al_u2841_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wfspw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W7iiu6 ));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u2843 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qe8iu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D31ju6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ),
    .o(_al_u2843_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u2844 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K49ow6_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    _al_u2845 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Frziu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K49ow6_lutinv ),
    .o(_al_u2845_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(~B*~A))"),
    .INIT(8'he0))
    _al_u2846 (
    .a(_al_u2843_o),
    .b(_al_u2845_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vo3ju6_lutinv ),
    .o(_al_u2846_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2847 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yqziu6 ),
    .b(_al_u1346_o),
    .o(_al_u2847_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u2848 (
    .a(_al_u2846_o),
    .b(_al_u2847_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qa5iu6 ));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u2849 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Frziu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 ),
    .o(_al_u2849_o));
  AL_MAP_LUT2 #(
    .EQN("~(B@A)"),
    .INIT(4'h9))
    _al_u285 (
    .a(b_pad_gpio_porta_pad[7]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_int_polarity [7]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/gpio_ext_porta_int [7]));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u2850 (
    .a(_al_u2849_o),
    .b(_al_u1336_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Owoiu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ja5iu6 ));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u2851 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qa5iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ja5iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z9opw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Usaiu6_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2852 (
    .a(_al_u1342_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vo3ju6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zwcpw6_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u2853 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zwcpw6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iugiu6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2854 (
    .a(_al_u1583_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P8oiu6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(~D*~(~C*~B)))"),
    .INIT(16'h5501))
    _al_u2855 (
    .a(_al_u2847_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iugiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P8oiu6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 ),
    .o(_al_u2855_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(~B*~A))"),
    .INIT(8'he0))
    _al_u2856 (
    .a(_al_u1385_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fnnpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/SLEEPHOLDACKn ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nsaiu6_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2857 (
    .a(_al_u2855_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nsaiu6_lutinv ),
    .o(_al_u2857_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~(B*A))"),
    .INIT(16'h0007))
    _al_u2858 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ja5iu6 ),
    .b(_al_u1812_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv ),
    .o(_al_u2858_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C*~B*A))"),
    .INIT(16'hdf00))
    _al_u2859 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Usaiu6_lutinv ),
    .b(_al_u2857_o),
    .c(_al_u2858_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/SLEEPHOLDACKn ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n689 ));
  AL_MAP_LUT2 #(
    .EQN("~(B@A)"),
    .INIT(4'h9))
    _al_u286 (
    .a(b_pad_gpio_porta_pad[6]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_int_polarity [6]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/gpio_ext_porta_int [6]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u2860 (
    .a(_al_u1812_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 ),
    .o(_al_u2860_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u2861 (
    .a(_al_u1344_o),
    .b(_al_u2403_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hgrpw6 ),
    .o(_al_u2861_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u2862 (
    .a(_al_u2861_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vygax6 ),
    .o(_al_u2862_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(D*C*A))"),
    .INIT(16'h4ccc))
    _al_u2863 (
    .a(_al_u2860_o),
    .b(_al_u2862_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ldoiu6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 ),
    .o(_al_u2863_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*A)"),
    .INIT(16'h0080))
    _al_u2864 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F6ziu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujiu6 ),
    .c(_al_u2770_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dd7ow6 ));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    _al_u2865 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dd7ow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gr2qw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vygax6 ),
    .o(_al_u2865_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u2866 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mbhow6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 ),
    .o(_al_u2866_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(C*A))"),
    .INIT(16'h5f13))
    _al_u2867 (
    .a(_al_u1806_o),
    .b(_al_u2866_o),
    .c(_al_u679_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 ),
    .o(_al_u2867_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2868 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vygax6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 ),
    .o(_al_u2868_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~A*~(D*C)))"),
    .INIT(16'hc888))
    _al_u2869 (
    .a(_al_u1812_o),
    .b(_al_u2868_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hgrpw6 ),
    .o(_al_u2869_o));
  AL_MAP_LUT2 #(
    .EQN("~(B@A)"),
    .INIT(4'h9))
    _al_u287 (
    .a(b_pad_gpio_porta_pad[5]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_int_polarity [5]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/gpio_ext_porta_int [5]));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(C*A))"),
    .INIT(16'h5f13))
    _al_u2870 (
    .a(_al_u609_o),
    .b(_al_u1346_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pu1ju6_lutinv ),
    .d(_al_u1907_o),
    .o(_al_u2870_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*~(D*~C)))"),
    .INIT(16'h2a22))
    _al_u2871 (
    .a(_al_u2870_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv ),
    .c(_al_u1266_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 ),
    .o(_al_u2871_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~(~B*A))"),
    .INIT(16'h0d00))
    _al_u2872 (
    .a(_al_u1643_o),
    .b(_al_u2867_o),
    .c(_al_u2869_o),
    .d(_al_u2871_o),
    .o(_al_u2872_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~B*~(~D*~A))"),
    .INIT(16'h3020))
    _al_u2873 (
    .a(_al_u2863_o),
    .b(_al_u2865_o),
    .c(_al_u2872_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 ),
    .o(_al_u2873_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hfd11))
    _al_u2874 (
    .a(_al_u2873_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ),
    .c(_al_u1817_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oqohu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u2875 (
    .a(_al_u2399_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zf7ju6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oikax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rwjax6 ),
    .o(_al_u2875_o));
  AL_MAP_LUT4 #(
    .EQN("~(B@(D*~(C*~A)))"),
    .INIT(16'h9c33))
    _al_u2876 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ka8ju6 ),
    .b(_al_u2398_o),
    .c(_al_u2412_o),
    .d(_al_u2875_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [10]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u2877 (
    .a(_al_u2399_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zf7ju6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iekax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N4kax6 ),
    .o(_al_u2877_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u2878 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kc6ju6 ),
    .b(_al_u2877_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Umkax6 ),
    .o(_al_u2878_o));
  AL_MAP_LUT4 #(
    .EQN("~(C@(A*~(D*~B)))"),
    .INIT(16'h87a5))
    _al_u2879 (
    .a(_al_u2878_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cz7ju6 ),
    .c(_al_u2398_o),
    .d(_al_u2412_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4epw6 ));
  AL_MAP_LUT2 #(
    .EQN("~(B@A)"),
    .INIT(4'h9))
    _al_u288 (
    .a(b_pad_gpio_porta_pad[4]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_int_polarity [4]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/gpio_ext_porta_int [4]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u2880 (
    .a(_al_u2849_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vgjpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ef7ju6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u2881 (
    .a(_al_u2650_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ef7ju6 ),
    .o(_al_u2881_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(C*~A))"),
    .INIT(16'h8caf))
    _al_u2882 (
    .a(_al_u1882_o),
    .b(_al_u2881_o),
    .c(_al_u2412_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sqkax6 ),
    .o(_al_u2882_o));
  AL_MAP_LUT2 #(
    .EQN("~(B@A)"),
    .INIT(4'h9))
    _al_u2883 (
    .a(_al_u2882_o),
    .b(_al_u2398_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [0]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2884 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n24_lutinv ),
    .b(_al_u588_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_dout_normal_write0 ));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D)*~((~C*~B))+A*D*~((~C*~B))+~(A)*D*(~C*~B)+A*D*(~C*~B))"),
    .INIT(16'haba8))
    _al_u2885 (
    .a(\u_cmsdk_mcu/HWDATA [0]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_dout_normal_write0 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]),
    .d(\u_cmsdk_mcu/p1_out [0]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/nxt_dout_padded [0]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2886 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n24_lutinv ),
    .b(_al_u593_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_dout_normal_write0 ));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D)*~((~C*~B))+A*D*~((~C*~B))+~(A)*D*(~C*~B)+A*D*(~C*~B))"),
    .INIT(16'haba8))
    _al_u2887 (
    .a(\u_cmsdk_mcu/HWDATA [0]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_dout_normal_write0 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]),
    .d(\u_cmsdk_mcu/p0_out [0]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/nxt_dout_padded [0]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2888 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n24_lutinv ),
    .b(_al_u585_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_dout_normal_write1 ));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D)*~((~C*~B))+A*D*~((~C*~B))+~(A)*D*(~C*~B)+A*D*(~C*~B))"),
    .INIT(16'haba8))
    _al_u2889 (
    .a(\u_cmsdk_mcu/HWDATA [8]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_dout_normal_write1 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]),
    .d(\u_cmsdk_mcu/p1_out [8]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/nxt_dout_padded [8]));
  AL_MAP_LUT2 #(
    .EQN("~(B@A)"),
    .INIT(4'h9))
    _al_u289 (
    .a(b_pad_gpio_porta_pad[3]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_int_polarity [3]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/gpio_ext_porta_int [3]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2890 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n24_lutinv ),
    .b(_al_u591_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_dout_normal_write1 ));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D)*~((~C*~B))+A*D*~((~C*~B))+~(A)*D*(~C*~B)+A*D*(~C*~B))"),
    .INIT(16'haba8))
    _al_u2891 (
    .a(\u_cmsdk_mcu/HWDATA [8]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_dout_normal_write1 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]),
    .d(\u_cmsdk_mcu/p0_out [8]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/nxt_dout_padded [8]));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(B*A))"),
    .INIT(8'hf8))
    _al_u2892 (
    .a(\u_cmsdk_mcu/HWDATA [10]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intclr_normal_write1 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_masked_int [10]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n291 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2893 (
    .a(\u_cmsdk_mcu/HWDATA [10]),
    .b(_al_u2500_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n254 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2894 (
    .a(\u_cmsdk_mcu/HWDATA [10]),
    .b(_al_u2502_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n209 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2895 (
    .a(\u_cmsdk_mcu/HWDATA [10]),
    .b(_al_u2504_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n164 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2896 (
    .a(\u_cmsdk_mcu/HWDATA [10]),
    .b(_al_u2506_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n119 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2897 (
    .a(\u_cmsdk_mcu/HWDATA [10]),
    .b(_al_u2508_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n74 ));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(B*A))"),
    .INIT(8'hf8))
    _al_u2898 (
    .a(\u_cmsdk_mcu/HWDATA [10]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intclr_normal_write1 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/new_masked_int [10]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n291 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2899 (
    .a(\u_cmsdk_mcu/HWDATA [10]),
    .b(_al_u2512_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n254 ));
  AL_MAP_LUT2 #(
    .EQN("~(B@A)"),
    .INIT(4'h9))
    _al_u290 (
    .a(b_pad_gpio_porta_pad[2]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_int_polarity [2]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/gpio_ext_porta_int [2]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2900 (
    .a(\u_cmsdk_mcu/HWDATA [10]),
    .b(_al_u2514_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n209 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2901 (
    .a(\u_cmsdk_mcu/HWDATA [10]),
    .b(_al_u2516_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n164 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2902 (
    .a(\u_cmsdk_mcu/HWDATA [10]),
    .b(_al_u2518_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n119 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2903 (
    .a(\u_cmsdk_mcu/HWDATA [10]),
    .b(_al_u2520_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n74 ));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D)*~((~C*~B))+A*D*~((~C*~B))+~(A)*D*(~C*~B)+A*D*(~C*~B))"),
    .INIT(16'haba8))
    _al_u2904 (
    .a(\u_cmsdk_mcu/HWDATA [2]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_dout_normal_write0 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4]),
    .d(\u_cmsdk_mcu/p1_out [2]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/nxt_dout_padded [2]));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D)*~((~C*~B))+A*D*~((~C*~B))+~(A)*D*(~C*~B)+A*D*(~C*~B))"),
    .INIT(16'haba8))
    _al_u2905 (
    .a(\u_cmsdk_mcu/HWDATA [2]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_dout_normal_write0 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4]),
    .d(\u_cmsdk_mcu/p0_out [2]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/nxt_dout_padded [2]));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(B*A))"),
    .INIT(8'hf8))
    _al_u2906 (
    .a(\u_cmsdk_mcu/HWDATA [11]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intclr_normal_write1 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_masked_int [11]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n293 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2907 (
    .a(\u_cmsdk_mcu/HWDATA [11]),
    .b(_al_u2500_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n256 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2908 (
    .a(\u_cmsdk_mcu/HWDATA [11]),
    .b(_al_u2502_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n211 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2909 (
    .a(\u_cmsdk_mcu/HWDATA [11]),
    .b(_al_u2504_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n166 ));
  AL_MAP_LUT2 #(
    .EQN("~(B@A)"),
    .INIT(4'h9))
    _al_u291 (
    .a(b_pad_gpio_porta_pad[1]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_int_polarity [1]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/gpio_ext_porta_int [1]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2910 (
    .a(\u_cmsdk_mcu/HWDATA [11]),
    .b(_al_u2506_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n121 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2911 (
    .a(\u_cmsdk_mcu/HWDATA [11]),
    .b(_al_u2508_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n76 ));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(B*A))"),
    .INIT(8'hf8))
    _al_u2912 (
    .a(\u_cmsdk_mcu/HWDATA [11]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intclr_normal_write1 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/new_masked_int [11]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n293 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2913 (
    .a(\u_cmsdk_mcu/HWDATA [11]),
    .b(_al_u2512_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n256 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2914 (
    .a(\u_cmsdk_mcu/HWDATA [11]),
    .b(_al_u2514_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n211 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2915 (
    .a(\u_cmsdk_mcu/HWDATA [11]),
    .b(_al_u2516_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n166 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2916 (
    .a(\u_cmsdk_mcu/HWDATA [11]),
    .b(_al_u2518_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n121 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2917 (
    .a(\u_cmsdk_mcu/HWDATA [11]),
    .b(_al_u2520_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n76 ));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D)*~((~C*~B))+A*D*~((~C*~B))+~(A)*D*(~C*~B)+A*D*(~C*~B))"),
    .INIT(16'haba8))
    _al_u2918 (
    .a(\u_cmsdk_mcu/HWDATA [3]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_dout_normal_write0 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [5]),
    .d(\u_cmsdk_mcu/p1_out [3]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/nxt_dout_padded [3]));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D)*~((~C*~B))+A*D*~((~C*~B))+~(A)*D*(~C*~B)+A*D*(~C*~B))"),
    .INIT(16'haba8))
    _al_u2919 (
    .a(\u_cmsdk_mcu/HWDATA [3]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_dout_normal_write0 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [5]),
    .d(\u_cmsdk_mcu/p0_out [3]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/nxt_dout_padded [3]));
  AL_MAP_LUT2 #(
    .EQN("~(B@A)"),
    .INIT(4'h9))
    _al_u292 (
    .a(b_pad_gpio_porta_pad[0]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_int_polarity [0]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/gpio_ext_porta_int [0]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2920 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zf7ju6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rkkax6 ),
    .o(_al_u2920_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u2921 (
    .a(_al_u2920_o),
    .b(_al_u2399_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6 ),
    .o(_al_u2921_o));
  AL_MAP_LUT4 #(
    .EQN("~(B@(D*~(C*~A)))"),
    .INIT(16'h9c33))
    _al_u2922 (
    .a(_al_u2062_o),
    .b(_al_u2398_o),
    .c(_al_u2412_o),
    .d(_al_u2921_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C1epw6 ));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(B*A))"),
    .INIT(8'hf8))
    _al_u2923 (
    .a(\u_cmsdk_mcu/HWDATA [12]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intclr_normal_write1 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_masked_int [12]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n295 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2924 (
    .a(\u_cmsdk_mcu/HWDATA [12]),
    .b(_al_u2500_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n258 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2925 (
    .a(\u_cmsdk_mcu/HWDATA [12]),
    .b(_al_u2502_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n213 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2926 (
    .a(\u_cmsdk_mcu/HWDATA [12]),
    .b(_al_u2504_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n168 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2927 (
    .a(\u_cmsdk_mcu/HWDATA [12]),
    .b(_al_u2506_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n123 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2928 (
    .a(\u_cmsdk_mcu/HWDATA [12]),
    .b(_al_u2508_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n78 ));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(B*A))"),
    .INIT(8'hf8))
    _al_u2929 (
    .a(\u_cmsdk_mcu/HWDATA [12]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intclr_normal_write1 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/new_masked_int [12]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n295 ));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u293 (
    .a(\u_cmsdk_mcu/u_ahb_ram/buf_hwaddr [12]),
    .b(\u_cmsdk_mcu/u_ahb_rom/we ),
    .o(\u_cmsdk_mcu/u_ahb_rom/n16 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2930 (
    .a(\u_cmsdk_mcu/HWDATA [12]),
    .b(_al_u2512_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n258 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2931 (
    .a(\u_cmsdk_mcu/HWDATA [12]),
    .b(_al_u2514_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n213 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2932 (
    .a(\u_cmsdk_mcu/HWDATA [12]),
    .b(_al_u2516_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n168 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2933 (
    .a(\u_cmsdk_mcu/HWDATA [12]),
    .b(_al_u2518_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n123 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2934 (
    .a(\u_cmsdk_mcu/HWDATA [12]),
    .b(_al_u2520_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n78 ));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D)*~((~C*~B))+A*D*~((~C*~B))+~(A)*D*(~C*~B)+A*D*(~C*~B))"),
    .INIT(16'haba8))
    _al_u2935 (
    .a(\u_cmsdk_mcu/HWDATA [4]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_dout_normal_write0 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [6]),
    .d(\u_cmsdk_mcu/p1_out [4]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/nxt_dout_padded [4]));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D)*~((~C*~B))+A*D*~((~C*~B))+~(A)*D*(~C*~B)+A*D*(~C*~B))"),
    .INIT(16'haba8))
    _al_u2936 (
    .a(\u_cmsdk_mcu/HWDATA [4]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_dout_normal_write0 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [6]),
    .d(\u_cmsdk_mcu/p0_out [4]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/nxt_dout_padded [4]));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u2937 (
    .a(_al_u2920_o),
    .b(_al_u2399_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R9mpw6 ),
    .o(_al_u2937_o));
  AL_MAP_LUT4 #(
    .EQN("~(B@(D*~(C*~A)))"),
    .INIT(16'h9c33))
    _al_u2938 (
    .a(_al_u2084_o),
    .b(_al_u2398_o),
    .c(_al_u2412_o),
    .d(_al_u2937_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J1epw6 ));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(B*A))"),
    .INIT(8'hf8))
    _al_u2939 (
    .a(\u_cmsdk_mcu/HWDATA [13]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intclr_normal_write1 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_masked_int [13]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n297 ));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u294 (
    .a(\u_cmsdk_mcu/u_ahb_ram/buf_hwaddr [12]),
    .b(\u_cmsdk_mcu/u_ahb_ram/we ),
    .o(\u_cmsdk_mcu/u_ahb_ram/n16 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2940 (
    .a(\u_cmsdk_mcu/HWDATA [13]),
    .b(_al_u2500_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n260 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2941 (
    .a(\u_cmsdk_mcu/HWDATA [13]),
    .b(_al_u2502_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n215 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2942 (
    .a(\u_cmsdk_mcu/HWDATA [13]),
    .b(_al_u2504_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n170 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2943 (
    .a(\u_cmsdk_mcu/HWDATA [13]),
    .b(_al_u2506_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n125 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2944 (
    .a(\u_cmsdk_mcu/HWDATA [13]),
    .b(_al_u2508_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n80 ));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(B*A))"),
    .INIT(8'hf8))
    _al_u2945 (
    .a(\u_cmsdk_mcu/HWDATA [13]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intclr_normal_write1 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/new_masked_int [13]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n297 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2946 (
    .a(\u_cmsdk_mcu/HWDATA [13]),
    .b(_al_u2512_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n260 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2947 (
    .a(\u_cmsdk_mcu/HWDATA [13]),
    .b(_al_u2514_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n215 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2948 (
    .a(\u_cmsdk_mcu/HWDATA [13]),
    .b(_al_u2516_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n170 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2949 (
    .a(\u_cmsdk_mcu/HWDATA [13]),
    .b(_al_u2518_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n125 ));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u295 (
    .a(\u_cmsdk_mcu/p1_out [1]),
    .b(\u_cmsdk_mcu/p1_outen [1]),
    .c(\u_cmsdk_mcu/p1_altfunc [1]),
    .o(\u_cmsdk_mcu/p1_in [1]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2950 (
    .a(\u_cmsdk_mcu/HWDATA [13]),
    .b(_al_u2520_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n80 ));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D)*~((~C*~B))+A*D*~((~C*~B))+~(A)*D*(~C*~B)+A*D*(~C*~B))"),
    .INIT(16'haba8))
    _al_u2951 (
    .a(\u_cmsdk_mcu/HWDATA [5]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_dout_normal_write0 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [7]),
    .d(\u_cmsdk_mcu/p1_out [5]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/nxt_dout_padded [5]));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D)*~((~C*~B))+A*D*~((~C*~B))+~(A)*D*(~C*~B)+A*D*(~C*~B))"),
    .INIT(16'haba8))
    _al_u2952 (
    .a(\u_cmsdk_mcu/HWDATA [5]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_dout_normal_write0 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [7]),
    .d(\u_cmsdk_mcu/p0_out [5]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/nxt_dout_padded [5]));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u2953 (
    .a(_al_u2920_o),
    .b(_al_u2399_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rskax6 ),
    .o(_al_u2953_o));
  AL_MAP_LUT4 #(
    .EQN("~(B@(D*~(C*~A)))"),
    .INIT(16'h9c33))
    _al_u2954 (
    .a(_al_u2106_o),
    .b(_al_u2398_o),
    .c(_al_u2412_o),
    .d(_al_u2953_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q1epw6 ));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(B*A))"),
    .INIT(8'hf8))
    _al_u2955 (
    .a(\u_cmsdk_mcu/HWDATA [14]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intclr_normal_write1 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_masked_int [14]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n299 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2956 (
    .a(\u_cmsdk_mcu/HWDATA [14]),
    .b(_al_u2500_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n262 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2957 (
    .a(\u_cmsdk_mcu/HWDATA [14]),
    .b(_al_u2502_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n217 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2958 (
    .a(\u_cmsdk_mcu/HWDATA [14]),
    .b(_al_u2504_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n172 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2959 (
    .a(\u_cmsdk_mcu/HWDATA [14]),
    .b(_al_u2506_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n127 ));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u296 (
    .a(\u_cmsdk_mcu/p1_out [3]),
    .b(\u_cmsdk_mcu/p1_outen [3]),
    .c(\u_cmsdk_mcu/p1_altfunc [3]),
    .o(\u_cmsdk_mcu/p1_in [3]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2960 (
    .a(\u_cmsdk_mcu/HWDATA [14]),
    .b(_al_u2508_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n82 ));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(B*A))"),
    .INIT(8'hf8))
    _al_u2961 (
    .a(\u_cmsdk_mcu/HWDATA [14]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intclr_normal_write1 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/new_masked_int [14]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n299 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2962 (
    .a(\u_cmsdk_mcu/HWDATA [14]),
    .b(_al_u2512_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n262 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2963 (
    .a(\u_cmsdk_mcu/HWDATA [14]),
    .b(_al_u2514_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n217 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2964 (
    .a(\u_cmsdk_mcu/HWDATA [14]),
    .b(_al_u2516_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n172 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2965 (
    .a(\u_cmsdk_mcu/HWDATA [14]),
    .b(_al_u2518_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n127 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2966 (
    .a(\u_cmsdk_mcu/HWDATA [14]),
    .b(_al_u2520_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n82 ));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D)*~((~C*~B))+A*D*~((~C*~B))+~(A)*D*(~C*~B)+A*D*(~C*~B))"),
    .INIT(16'haba8))
    _al_u2967 (
    .a(\u_cmsdk_mcu/HWDATA [6]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_dout_normal_write0 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [8]),
    .d(\u_cmsdk_mcu/p1_out [6]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/nxt_dout_padded [6]));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D)*~((~C*~B))+A*D*~((~C*~B))+~(A)*D*(~C*~B)+A*D*(~C*~B))"),
    .INIT(16'haba8))
    _al_u2968 (
    .a(\u_cmsdk_mcu/HWDATA [6]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_dout_normal_write0 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [8]),
    .d(\u_cmsdk_mcu/p0_out [6]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/nxt_dout_padded [6]));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u2969 (
    .a(_al_u2920_o),
    .b(_al_u2399_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U1kpw6 ),
    .o(_al_u2969_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u297 (
    .a(\u_cmsdk_mcu/p1_out [5]),
    .b(\u_cmsdk_mcu/p1_outen [5]),
    .c(\u_cmsdk_mcu/p1_altfunc [5]),
    .o(\u_cmsdk_mcu/p1_in [5]));
  AL_MAP_LUT4 #(
    .EQN("~(B@(D*~(C*~A)))"),
    .INIT(16'h9c33))
    _al_u2970 (
    .a(_al_u2128_o),
    .b(_al_u2398_o),
    .c(_al_u2412_o),
    .d(_al_u2969_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X1epw6 ));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(B*A))"),
    .INIT(8'hf8))
    _al_u2971 (
    .a(\u_cmsdk_mcu/HWDATA [15]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intclr_normal_write1 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_masked_int [15]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n301 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2972 (
    .a(\u_cmsdk_mcu/HWDATA [15]),
    .b(_al_u2500_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n264 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2973 (
    .a(\u_cmsdk_mcu/HWDATA [15]),
    .b(_al_u2502_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n219 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2974 (
    .a(\u_cmsdk_mcu/HWDATA [15]),
    .b(_al_u2504_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n174 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2975 (
    .a(\u_cmsdk_mcu/HWDATA [15]),
    .b(_al_u2506_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n129 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2976 (
    .a(\u_cmsdk_mcu/HWDATA [15]),
    .b(_al_u2508_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n84 ));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(B*A))"),
    .INIT(8'hf8))
    _al_u2977 (
    .a(\u_cmsdk_mcu/HWDATA [15]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intclr_normal_write1 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/new_masked_int [15]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n301 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2978 (
    .a(\u_cmsdk_mcu/HWDATA [15]),
    .b(_al_u2512_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n264 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2979 (
    .a(\u_cmsdk_mcu/HWDATA [15]),
    .b(_al_u2514_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n219 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u298 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [4]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/apbsys_hreadyout ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2980 (
    .a(\u_cmsdk_mcu/HWDATA [15]),
    .b(_al_u2516_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n174 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2981 (
    .a(\u_cmsdk_mcu/HWDATA [15]),
    .b(_al_u2518_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n129 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2982 (
    .a(\u_cmsdk_mcu/HWDATA [15]),
    .b(_al_u2520_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n84 ));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D)*~((~C*~B))+A*D*~((~C*~B))+~(A)*D*(~C*~B)+A*D*(~C*~B))"),
    .INIT(16'haba8))
    _al_u2983 (
    .a(\u_cmsdk_mcu/HWDATA [7]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_dout_normal_write0 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [9]),
    .d(\u_cmsdk_mcu/p1_out [7]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/nxt_dout_padded [7]));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D)*~((~C*~B))+A*D*~((~C*~B))+~(A)*D*(~C*~B)+A*D*(~C*~B))"),
    .INIT(16'haba8))
    _al_u2984 (
    .a(\u_cmsdk_mcu/HWDATA [7]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_dout_normal_write0 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [9]),
    .d(\u_cmsdk_mcu/p0_out [7]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/nxt_dout_padded [7]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u2985 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kc6ju6 ),
    .b(_al_u2399_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fkrpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4jax6 ),
    .o(_al_u2985_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*~B))"),
    .INIT(8'h8a))
    _al_u2986 (
    .a(_al_u2985_o),
    .b(_al_u1961_o),
    .c(_al_u2412_o),
    .o(_al_u2986_o));
  AL_MAP_LUT4 #(
    .EQN("~(B@(A*~(D*~C)))"),
    .INIT(16'h9399))
    _al_u2987 (
    .a(_al_u2986_o),
    .b(_al_u2398_o),
    .c(_al_u2650_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V6jax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S2epw6 ));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u2988 (
    .a(_al_u2920_o),
    .b(_al_u2399_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ubypw6 ),
    .o(_al_u2988_o));
  AL_MAP_LUT4 #(
    .EQN("~(B@(D*~(C*~A)))"),
    .INIT(16'h9c33))
    _al_u2989 (
    .a(_al_u2150_o),
    .b(_al_u2398_o),
    .c(_al_u2412_o),
    .d(_al_u2988_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L2epw6 ));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~B*~A)"),
    .INIT(8'hfe))
    _al_u299 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/baud_updated ),
    .b(uart0_txen_pad),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_ctrl [1]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n38 ));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u2990 (
    .a(_al_u2920_o),
    .b(_al_u2399_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Umkax6 ),
    .o(_al_u2990_o));
  AL_MAP_LUT4 #(
    .EQN("~(B@(D*~(C*~A)))"),
    .INIT(16'h9c33))
    _al_u2991 (
    .a(_al_u2171_o),
    .b(_al_u2398_o),
    .c(_al_u2412_o),
    .d(_al_u2990_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G3epw6 ));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u2992 (
    .a(_al_u497_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [5]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [6]),
    .o(_al_u2992_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*A)"),
    .INIT(16'h0200))
    _al_u2993 (
    .a(_al_u2992_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [2]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [3]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [4]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/n34_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u2994 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/n34_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_byte_strobe [0]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_write_enable ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_resetinfo_write ));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B*A))"),
    .INIT(8'h70))
    _al_u2995 (
    .a(\u_cmsdk_mcu/HWDATA [1]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_resetinfo_write ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_resetinfo [1]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/n38 [1]));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D)*~((~C*~B))+A*D*~((~C*~B))+~(A)*D*(~C*~B)+A*D*(~C*~B))"),
    .INIT(16'haba8))
    _al_u2996 (
    .a(\u_cmsdk_mcu/HWDATA [1]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_dout_normal_write0 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .d(\u_cmsdk_mcu/p1_out [1]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/nxt_dout_padded [1]));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D)*~((~C*~B))+A*D*~((~C*~B))+~(A)*D*(~C*~B)+A*D*(~C*~B))"),
    .INIT(16'haba8))
    _al_u2997 (
    .a(\u_cmsdk_mcu/HWDATA [1]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_dout_normal_write0 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .d(\u_cmsdk_mcu/p0_out [1]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/nxt_dout_padded [1]));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D)*~((~C*~B))+A*D*~((~C*~B))+~(A)*D*(~C*~B)+A*D*(~C*~B))"),
    .INIT(16'haba8))
    _al_u2998 (
    .a(\u_cmsdk_mcu/HWDATA [9]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_dout_normal_write1 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .d(\u_cmsdk_mcu/p1_out [9]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/nxt_dout_padded [9]));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D)*~((~C*~B))+A*D*~((~C*~B))+~(A)*D*(~C*~B)+A*D*(~C*~B))"),
    .INIT(16'haba8))
    _al_u2999 (
    .a(\u_cmsdk_mcu/HWDATA [9]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_dout_normal_write1 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .d(\u_cmsdk_mcu/p0_out [9]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/nxt_dout_padded [9]));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u300 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dugax6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ksgax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E4yhu6 ));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u3000 (
    .a(_al_u2920_o),
    .b(_al_u2399_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V6jax6 ),
    .o(_al_u3000_o));
  AL_MAP_LUT4 #(
    .EQN("~(B@(D*~(C*~A)))"),
    .INIT(16'h9c33))
    _al_u3001 (
    .a(_al_u2208_o),
    .b(_al_u2398_o),
    .c(_al_u2412_o),
    .d(_al_u3000_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N3epw6 ));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u3002 (
    .a(_al_u2920_o),
    .b(_al_u2399_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iekax6 ),
    .o(_al_u3002_o));
  AL_MAP_LUT4 #(
    .EQN("~(B@(D*~(C*~A)))"),
    .INIT(16'h9c33))
    _al_u3003 (
    .a(_al_u2217_o),
    .b(_al_u2398_o),
    .c(_al_u2412_o),
    .d(_al_u3002_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U3epw6 ));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u3004 (
    .a(_al_u2920_o),
    .b(_al_u2399_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lgkax6 ),
    .o(_al_u3004_o));
  AL_MAP_LUT4 #(
    .EQN("~(B@(D*~(C*~A)))"),
    .INIT(16'h9c33))
    _al_u3005 (
    .a(_al_u2225_o),
    .b(_al_u2398_o),
    .c(_al_u2412_o),
    .d(_al_u3004_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B4epw6 ));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u3006 (
    .a(_al_u2920_o),
    .b(_al_u2399_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oikax6 ),
    .o(_al_u3006_o));
  AL_MAP_LUT4 #(
    .EQN("~(B@(D*~(C*~A)))"),
    .INIT(16'h9c33))
    _al_u3007 (
    .a(_al_u2235_o),
    .b(_al_u2398_o),
    .c(_al_u2412_o),
    .d(_al_u3006_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I4epw6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D)"),
    .INIT(16'h1f35))
    _al_u3008 (
    .a(_al_u2399_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zf7ju6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rkkax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 ),
    .o(_al_u3008_o));
  AL_MAP_LUT4 #(
    .EQN("~(B@(D*~(C*~A)))"),
    .INIT(16'h9c33))
    _al_u3009 (
    .a(_al_u2244_o),
    .b(_al_u2398_o),
    .c(_al_u2412_o),
    .d(_al_u3008_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P4epw6 ));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u301 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L5lpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pmlpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y8lpw6 ),
    .o(\u_cmsdk_mcu/dbg_swdo ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*~(B)*C*D)"),
    .INIT(16'h13f5))
    _al_u3010 (
    .a(_al_u2399_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zf7ju6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P14qw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rkkax6 ),
    .o(_al_u3010_o));
  AL_MAP_LUT4 #(
    .EQN("~(B@(D*~(C*~A)))"),
    .INIT(16'h9c33))
    _al_u3011 (
    .a(_al_u2252_o),
    .b(_al_u2398_o),
    .c(_al_u2412_o),
    .d(_al_u3010_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [23]));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u3012 (
    .a(_al_u2920_o),
    .b(_al_u2399_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fkrpw6 ),
    .o(_al_u3012_o));
  AL_MAP_LUT4 #(
    .EQN("~(B@(D*~(C*~A)))"),
    .INIT(16'h9c33))
    _al_u3013 (
    .a(_al_u2289_o),
    .b(_al_u2398_o),
    .c(_al_u2412_o),
    .d(_al_u3012_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z2epw6 ));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(B*~A))"),
    .INIT(8'h0b))
    _al_u3014 (
    .a(_al_u607_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F1jiu6_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3015 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F1jiu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ),
    .o(_al_u3015_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3016 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Difiu6 ));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'h5c))
    _al_u3017 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Difiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 ),
    .o(_al_u3017_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3018 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jf6ju6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3019 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pthiu6 ));
  AL_MAP_LUT2 #(
    .EQN("~(B*A)"),
    .INIT(4'h7))
    _al_u302 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sqfax6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uofax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n265 ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*C)*~(B*A))"),
    .INIT(16'h0777))
    _al_u3020 (
    .a(_al_u1342_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jf6ju6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pthiu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 ),
    .o(_al_u3020_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(D*~C*~A))"),
    .INIT(16'hc8cc))
    _al_u3021 (
    .a(_al_u3017_o),
    .b(_al_u3020_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 ),
    .o(_al_u3021_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C*~B*A))"),
    .INIT(16'hdf00))
    _al_u3022 (
    .a(_al_u2461_o),
    .b(_al_u3015_o),
    .c(_al_u3021_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vgjpw6 ),
    .o(_al_u3022_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*~A))"),
    .INIT(16'h23af))
    _al_u3023 (
    .a(_al_u1943_o),
    .b(_al_u3022_o),
    .c(_al_u2412_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U1kpw6 ),
    .o(_al_u3023_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*~A))"),
    .INIT(16'h23af))
    _al_u3024 (
    .a(_al_u2650_o),
    .b(_al_u2399_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fkrpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jgxpw6 ),
    .o(_al_u3024_o));
  AL_MAP_LUT3 #(
    .EQN("~(B@(C*A))"),
    .INIT(8'h93))
    _al_u3025 (
    .a(_al_u3023_o),
    .b(_al_u2398_o),
    .c(_al_u3024_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [5]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*~A))"),
    .INIT(16'h23af))
    _al_u3026 (
    .a(_al_u1925_o),
    .b(_al_u3022_o),
    .c(_al_u2412_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R9mpw6 ),
    .o(_al_u3026_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*~A))"),
    .INIT(16'h2a3f))
    _al_u3027 (
    .a(_al_u2650_o),
    .b(_al_u2399_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Irmpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U1kpw6 ),
    .o(_al_u3027_o));
  AL_MAP_LUT3 #(
    .EQN("~(B@(C*A))"),
    .INIT(8'h93))
    _al_u3028 (
    .a(_al_u3026_o),
    .b(_al_u2398_o),
    .c(_al_u3027_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [3]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*~A))"),
    .INIT(16'h23af))
    _al_u3029 (
    .a(_al_u1934_o),
    .b(_al_u3022_o),
    .c(_al_u2412_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rskax6 ),
    .o(_al_u3029_o));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    _al_u303 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qsfax6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxqpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iqzhu6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*~A))"),
    .INIT(16'h23af))
    _al_u3030 (
    .a(_al_u2650_o),
    .b(_al_u2399_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ubypw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wkipw6 ),
    .o(_al_u3030_o));
  AL_MAP_LUT3 #(
    .EQN("~(B@(C*A))"),
    .INIT(8'h93))
    _al_u3031 (
    .a(_al_u3029_o),
    .b(_al_u2398_o),
    .c(_al_u3030_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [4]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*C)*~(B*~A))"),
    .INIT(16'h0bbb))
    _al_u3032 (
    .a(_al_u1968_o),
    .b(_al_u2412_o),
    .c(_al_u2399_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wfspw6 ),
    .o(_al_u3032_o));
  AL_MAP_LUT4 #(
    .EQN("~(B@(A*~(D*~C)))"),
    .INIT(16'h9399))
    _al_u3033 (
    .a(_al_u3032_o),
    .b(_al_u2398_o),
    .c(_al_u2881_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R9mpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [1]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u3034 (
    .a(_al_u3022_o),
    .b(_al_u2399_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S7mpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sqkax6 ),
    .o(_al_u3034_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*~B))"),
    .INIT(8'h8a))
    _al_u3035 (
    .a(_al_u3034_o),
    .b(_al_u1916_o),
    .c(_al_u2412_o),
    .o(_al_u3035_o));
  AL_MAP_LUT4 #(
    .EQN("~(B@(A*~(D*~C)))"),
    .INIT(16'h9399))
    _al_u3036 (
    .a(_al_u3035_o),
    .b(_al_u2398_o),
    .c(_al_u2881_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rskax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [2]));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~(C*~(B*A)))"),
    .INIT(16'hff70))
    _al_u3037 (
    .a(\u_cmsdk_mcu/HWDATA [0]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_resetinfo_write ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_resetinfo [0]),
    .d(\u_cmsdk_mcu/SYSRESETREQ ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/nxt_resetinfo [0]));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*A)"),
    .INIT(16'h0200))
    _al_u3038 (
    .a(_al_u1048_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[4] ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[5] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[6] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n12_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3039 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n12_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n63 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u304 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iqzhu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I4rpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T24iu6 ));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*~A)"),
    .INIT(8'h04))
    _al_u3040 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_ddr [0]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/int_pre_in [0]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/ed_int_d1 [0]),
    .o(_al_u3040_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(B*A)))"),
    .INIT(16'h080f))
    _al_u3041 (
    .a(\u_cmsdk_mcu/HWDATA [0]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n63 ),
    .c(_al_u3040_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/gpio_intr_ed_pm [0]),
    .o(_al_u3041_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u3042 (
    .a(_al_u3041_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inten [0]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/n28 ));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D)*~((~C*~B))+A*D*~((~C*~B))+~(A)*D*(~C*~B)+A*D*(~C*~B))"),
    .INIT(16'haba8))
    _al_u3043 (
    .a(\u_cmsdk_mcu/HWDATA [10]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_dout_normal_write1 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4]),
    .d(\u_cmsdk_mcu/p1_out [10]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/nxt_dout_padded [10]));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D)*~((~C*~B))+A*D*~((~C*~B))+~(A)*D*(~C*~B)+A*D*(~C*~B))"),
    .INIT(16'haba8))
    _al_u3044 (
    .a(\u_cmsdk_mcu/HWDATA [10]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_dout_normal_write1 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4]),
    .d(\u_cmsdk_mcu/p0_out [10]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/nxt_dout_padded [10]));
  AL_MAP_LUT4 #(
    .EQN("~(~B*~(D*~(C*A)))"),
    .INIT(16'hdfcc))
    _al_u3045 (
    .a(\u_cmsdk_mcu/HWDATA [2]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_overrun ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n9_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_tx_overrun ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_tx_overrun ));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*~A)"),
    .INIT(8'h04))
    _al_u3046 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_ddr [2]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/int_pre_in [2]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/ed_int_d1 [2]),
    .o(_al_u3046_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(B*A)))"),
    .INIT(16'h080f))
    _al_u3047 (
    .a(\u_cmsdk_mcu/HWDATA [2]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n63 ),
    .c(_al_u3046_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/gpio_intr_ed_pm [2]),
    .o(_al_u3047_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u3048 (
    .a(_al_u3047_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inten [2]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/n44 ));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D)*~((~C*~B))+A*D*~((~C*~B))+~(A)*D*(~C*~B)+A*D*(~C*~B))"),
    .INIT(16'haba8))
    _al_u3049 (
    .a(\u_cmsdk_mcu/HWDATA [11]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_dout_normal_write1 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [5]),
    .d(\u_cmsdk_mcu/p1_out [11]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/nxt_dout_padded [11]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u305 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iqzhu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C2ypw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J44iu6 ));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D)*~((~C*~B))+A*D*~((~C*~B))+~(A)*D*(~C*~B)+A*D*(~C*~B))"),
    .INIT(16'haba8))
    _al_u3050 (
    .a(\u_cmsdk_mcu/HWDATA [11]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_dout_normal_write1 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [5]),
    .d(\u_cmsdk_mcu/p0_out [11]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/nxt_dout_padded [11]));
  AL_MAP_LUT4 #(
    .EQN("~(~B*~(D*~(C*A)))"),
    .INIT(16'hdfcc))
    _al_u3051 (
    .a(\u_cmsdk_mcu/HWDATA [3]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_overrun ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n9_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_rx_overrun ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_rx_overrun ));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*~A)"),
    .INIT(8'h04))
    _al_u3052 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_ddr [3]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/int_pre_in [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/ed_int_d1 [3]),
    .o(_al_u3052_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(B*A)))"),
    .INIT(16'h080f))
    _al_u3053 (
    .a(\u_cmsdk_mcu/HWDATA [3]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n63 ),
    .c(_al_u3052_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/gpio_intr_ed_pm [3]),
    .o(_al_u3053_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u3054 (
    .a(_al_u3053_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inten [3]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/n52 ));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D)*~((~C*~B))+A*D*~((~C*~B))+~(A)*D*(~C*~B)+A*D*(~C*~B))"),
    .INIT(16'haba8))
    _al_u3055 (
    .a(\u_cmsdk_mcu/HWDATA [12]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_dout_normal_write1 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [6]),
    .d(\u_cmsdk_mcu/p1_out [12]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/nxt_dout_padded [12]));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D)*~((~C*~B))+A*D*~((~C*~B))+~(A)*D*(~C*~B)+A*D*(~C*~B))"),
    .INIT(16'haba8))
    _al_u3056 (
    .a(\u_cmsdk_mcu/HWDATA [12]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_dout_normal_write1 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [6]),
    .d(\u_cmsdk_mcu/p0_out [12]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/nxt_dout_padded [12]));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*~A)"),
    .INIT(8'h04))
    _al_u3057 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_ddr [4]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/int_pre_in [4]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/ed_int_d1 [4]),
    .o(_al_u3057_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(B*A)))"),
    .INIT(16'h080f))
    _al_u3058 (
    .a(\u_cmsdk_mcu/HWDATA [4]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n63 ),
    .c(_al_u3057_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/gpio_intr_ed_pm [4]),
    .o(_al_u3058_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u3059 (
    .a(_al_u3058_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inten [4]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/n60 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u306 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iqzhu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xx6bx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q44iu6 ));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D)*~((~C*~B))+A*D*~((~C*~B))+~(A)*D*(~C*~B)+A*D*(~C*~B))"),
    .INIT(16'haba8))
    _al_u3060 (
    .a(\u_cmsdk_mcu/HWDATA [13]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_dout_normal_write1 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [7]),
    .d(\u_cmsdk_mcu/p1_out [13]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/nxt_dout_padded [13]));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D)*~((~C*~B))+A*D*~((~C*~B))+~(A)*D*(~C*~B)+A*D*(~C*~B))"),
    .INIT(16'haba8))
    _al_u3061 (
    .a(\u_cmsdk_mcu/HWDATA [13]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_dout_normal_write1 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [7]),
    .d(\u_cmsdk_mcu/p0_out [13]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/nxt_dout_padded [13]));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*~A)"),
    .INIT(8'h04))
    _al_u3062 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_ddr [5]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/int_pre_in [5]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/ed_int_d1 [5]),
    .o(_al_u3062_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(B*A)))"),
    .INIT(16'h080f))
    _al_u3063 (
    .a(\u_cmsdk_mcu/HWDATA [5]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n63 ),
    .c(_al_u3062_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/gpio_intr_ed_pm [5]),
    .o(_al_u3063_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u3064 (
    .a(_al_u3063_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inten [5]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/n68 ));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D)*~((~C*~B))+A*D*~((~C*~B))+~(A)*D*(~C*~B)+A*D*(~C*~B))"),
    .INIT(16'haba8))
    _al_u3065 (
    .a(\u_cmsdk_mcu/HWDATA [14]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_dout_normal_write1 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [8]),
    .d(\u_cmsdk_mcu/p1_out [14]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/nxt_dout_padded [14]));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D)*~((~C*~B))+A*D*~((~C*~B))+~(A)*D*(~C*~B)+A*D*(~C*~B))"),
    .INIT(16'haba8))
    _al_u3066 (
    .a(\u_cmsdk_mcu/HWDATA [14]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_dout_normal_write1 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [8]),
    .d(\u_cmsdk_mcu/p0_out [14]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/nxt_dout_padded [14]));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*~A)"),
    .INIT(8'h04))
    _al_u3067 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_ddr [6]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/int_pre_in [6]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/ed_int_d1 [6]),
    .o(_al_u3067_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(B*A)))"),
    .INIT(16'h080f))
    _al_u3068 (
    .a(\u_cmsdk_mcu/HWDATA [6]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n63 ),
    .c(_al_u3067_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/gpio_intr_ed_pm [6]),
    .o(_al_u3068_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u3069 (
    .a(_al_u3068_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inten [6]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/n76 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u307 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iqzhu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ns8ax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X44iu6 ));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D)*~((~C*~B))+A*D*~((~C*~B))+~(A)*D*(~C*~B)+A*D*(~C*~B))"),
    .INIT(16'haba8))
    _al_u3070 (
    .a(\u_cmsdk_mcu/HWDATA [15]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_dout_normal_write1 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [9]),
    .d(\u_cmsdk_mcu/p1_out [15]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/nxt_dout_padded [15]));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D)*~((~C*~B))+A*D*~((~C*~B))+~(A)*D*(~C*~B)+A*D*(~C*~B))"),
    .INIT(16'haba8))
    _al_u3071 (
    .a(\u_cmsdk_mcu/HWDATA [15]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_dout_normal_write1 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [9]),
    .d(\u_cmsdk_mcu/p0_out [15]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/nxt_dout_padded [15]));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*~A)"),
    .INIT(8'h04))
    _al_u3072 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_ddr [7]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/int_pre_in [7]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/ed_int_d1 [7]),
    .o(_al_u3072_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(B*A)))"),
    .INIT(16'h080f))
    _al_u3073 (
    .a(\u_cmsdk_mcu/HWDATA [7]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n63 ),
    .c(_al_u3072_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/gpio_intr_ed_pm [7]),
    .o(_al_u3073_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u3074 (
    .a(_al_u3073_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inten [7]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/n84 ));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*~A)"),
    .INIT(8'h04))
    _al_u3075 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_ddr [1]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/int_pre_in [1]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/ed_int_d1 [1]),
    .o(_al_u3075_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(B*A)))"),
    .INIT(16'h080f))
    _al_u3076 (
    .a(\u_cmsdk_mcu/HWDATA [1]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n63 ),
    .c(_al_u3075_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/gpio_intr_ed_pm [1]),
    .o(_al_u3076_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u3077 (
    .a(_al_u3076_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inten [1]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/n36 ));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*B*A)"),
    .INIT(16'h0800))
    _al_u3078 (
    .a(_al_u695_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 ),
    .o(_al_u3078_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~B*~(D*A))"),
    .INIT(16'h0103))
    _al_u3079 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hviiu6 ),
    .b(_al_u3078_o),
    .c(_al_u1264_o),
    .d(_al_u2371_o),
    .o(_al_u3079_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u308 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iqzhu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fj8ax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E54iu6 ));
  AL_MAP_LUT4 #(
    .EQN("(A*~(~D*~C*B))"),
    .INIT(16'haaa2))
    _al_u3080 (
    .a(_al_u3079_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vviiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rwjax6 ),
    .o(_al_u3080_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3081 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W0piu6_lutinv ),
    .b(_al_u2376_o),
    .o(_al_u3081_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3082 (
    .a(_al_u604_o),
    .b(_al_u2813_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 ),
    .o(_al_u3082_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*B*~A))"),
    .INIT(16'h0b0f))
    _al_u3083 (
    .a(_al_u1812_o),
    .b(_al_u1799_o),
    .c(_al_u3082_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 ),
    .o(_al_u3083_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~B*~(~D*A))"),
    .INIT(16'h3010))
    _al_u3084 (
    .a(_al_u1801_o),
    .b(_al_u3081_o),
    .c(_al_u3083_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D0jiu6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3085 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nu9ow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wkipw6 ),
    .o(_al_u3085_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*B)*~(~D*A))"),
    .INIT(16'hf351))
    _al_u3086 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wkjiu6 ),
    .b(_al_u3085_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 ),
    .o(_al_u3086_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u3087 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D0jiu6 ),
    .b(_al_u3086_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vviiu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 ),
    .o(_al_u3087_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3088 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pu1ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y0jiu6 ));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u3089 (
    .a(_al_u1802_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y0jiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Veziu6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u309 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iqzhu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Liabx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L54iu6 ));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u3090 (
    .a(_al_u2386_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qxoiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N4kax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cjiow6 ));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(D*~C*B))"),
    .INIT(16'h5155))
    _al_u3091 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cjiow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P14qw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9ypw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 ),
    .o(_al_u3091_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(A*~(D*C)))"),
    .INIT(16'hc444))
    _al_u3092 (
    .a(_al_u3091_o),
    .b(_al_u2361_o),
    .c(_al_u2365_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 ),
    .o(_al_u3092_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*A)"),
    .INIT(16'h0080))
    _al_u3093 (
    .a(_al_u3080_o),
    .b(_al_u3087_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Veziu6 ),
    .d(_al_u3092_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Epjiu6 ));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    _al_u3094 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fnnpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G0zax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[2] ),
    .o(_al_u3094_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u3095 (
    .a(_al_u1812_o),
    .b(_al_u3094_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mmjiu6_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    _al_u3096 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mmjiu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pthiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 ),
    .o(_al_u3096_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u3097 (
    .a(_al_u3096_o),
    .b(_al_u1783_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ),
    .o(_al_u3097_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3098 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uu9ow6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9ypw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ujjiu6 ));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3099 (
    .a(_al_u1812_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R9aiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wkipw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Njjiu6_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u310 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iqzhu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Va7ax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S54iu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u3100 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wkjiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ujjiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Njjiu6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6 ),
    .o(_al_u3100_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3101 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L45iu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S2ziu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 ),
    .o(_al_u3101_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u3102 (
    .a(_al_u3101_o),
    .b(_al_u2758_o),
    .c(_al_u1266_o),
    .o(_al_u3102_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3103 (
    .a(_al_u1266_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ),
    .o(_al_u3103_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u3104 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv ),
    .b(_al_u932_o),
    .c(_al_u1346_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pthiu6 ),
    .o(_al_u3104_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u3105 (
    .a(_al_u3103_o),
    .b(_al_u3104_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pu1ju6_lutinv ),
    .o(_al_u3105_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u3106 (
    .a(_al_u3097_o),
    .b(_al_u3100_o),
    .c(_al_u3102_o),
    .d(_al_u3105_o),
    .o(_al_u3106_o));
  AL_MAP_LUT4 #(
    .EQN("(A*B*~(C)*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hfee8))
    _al_u3107 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iekax6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lgkax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oikax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rkkax6 ),
    .o(_al_u3107_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*(~(A)*~(C)*~(D)+A*~(C)*~(D)+A*C*~(D)+A*~(C)*D))"),
    .INIT(16'h0223))
    _al_u3108 (
    .a(_al_u916_o),
    .b(_al_u3107_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fkrpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ubypw6 ),
    .o(_al_u3108_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(~(A)*~(C)*~(D)+A*~(C)*~(D)+A*C*~(D)+A*~(C)*D))"),
    .INIT(16'h088c))
    _al_u3109 (
    .a(_al_u1383_o),
    .b(_al_u3108_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Umkax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V6jax6 ),
    .o(_al_u3109_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u311 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iqzhu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lhbbx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G64iu6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3110 (
    .a(_al_u609_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 ),
    .o(_al_u3110_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3111 (
    .a(_al_u3109_o),
    .b(_al_u3110_o),
    .o(_al_u3111_o));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~(~C*B*A))"),
    .INIT(16'hff08))
    _al_u3112 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Epjiu6 ),
    .b(_al_u3106_o),
    .c(_al_u3111_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F58iu6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3113 (
    .a(_al_u3110_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Glaiu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(~D*~C*A))"),
    .INIT(16'h3331))
    _al_u3114 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kwuow6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Glaiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 ),
    .o(_al_u3114_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u3115 (
    .a(_al_u2868_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 ),
    .o(_al_u3115_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D*~C*B))"),
    .INIT(16'ha2aa))
    _al_u3116 (
    .a(_al_u3114_o),
    .b(_al_u3115_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yoniu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(D*~(~C*~B)))"),
    .INIT(16'h0155))
    _al_u3117 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iugiu6 ),
    .b(_al_u932_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yecpw6_lutinv ),
    .d(_al_u2813_o),
    .o(_al_u3117_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3118 (
    .a(_al_u607_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ),
    .o(_al_u3118_o));
  AL_MAP_LUT4 #(
    .EQN("~((C*B)*~(A)*~(D)+(C*B)*A*~(D)+~((C*B))*A*D+(C*B)*A*D)"),
    .INIT(16'h553f))
    _al_u3119 (
    .a(_al_u679_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 ),
    .o(_al_u3119_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u312 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iqzhu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gwwpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N64iu6 ));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D*~(C*~B)))"),
    .INIT(16'h20aa))
    _al_u3120 (
    .a(_al_u3117_o),
    .b(_al_u3118_o),
    .c(_al_u3119_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 ),
    .o(_al_u3120_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(C*~A))"),
    .INIT(16'h8caf))
    _al_u3121 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yoniu6 ),
    .b(_al_u3120_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iixpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lgkax6 ),
    .o(_al_u3121_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u3122 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vygax6 ),
    .o(_al_u3122_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(~D*B*A))"),
    .INIT(16'h0f07))
    _al_u3123 (
    .a(_al_u2866_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv ),
    .c(_al_u3122_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xiaju6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3124 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 ),
    .o(_al_u3124_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(C*~A))"),
    .INIT(16'haf23))
    _al_u3125 (
    .a(_al_u1803_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Owoiu6 ),
    .c(_al_u3124_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L0vow6 ));
  AL_MAP_LUT4 #(
    .EQN("(A*~(~D*~C*B))"),
    .INIT(16'haaa2))
    _al_u3126 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L0vow6 ),
    .b(_al_u679_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 ),
    .o(_al_u3126_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'hca00))
    _al_u3127 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yi7ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ),
    .o(_al_u3127_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3128 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Edapw6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~(~B*~A))"),
    .INIT(16'he000))
    _al_u3129 (
    .a(_al_u604_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Edapw6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 ),
    .o(_al_u3129_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u313 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iqzhu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cfvpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U64iu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    _al_u3130 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xiaju6 ),
    .b(_al_u3126_o),
    .c(_al_u3127_o),
    .d(_al_u3129_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mpniu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*B)*~(~D*A))"),
    .INIT(16'hf351))
    _al_u3131 (
    .a(_al_u1887_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Utniu6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(C*A*~(D*~B))"),
    .INIT(16'h80a0))
    _al_u3132 (
    .a(_al_u3121_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mpniu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Utniu6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wxjpw6 ),
    .o(_al_u3132_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*(~(B)*C*~(D)+B*~(C)*D+~(B)*C*D))"),
    .INIT(16'h1410))
    _al_u3133 (
    .a(_al_u1906_o),
    .b(_al_u1299_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rskax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ubypw6 ),
    .o(_al_u3133_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D*C*~A))"),
    .INIT(16'h2333))
    _al_u3134 (
    .a(_al_u3132_o),
    .b(_al_u3133_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Stuow6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cz8iu6 ));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    _al_u3135 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cz8iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n590 ));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3136 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K5eiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wjyiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C1wpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V59iu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    _al_u3137 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K5eiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C1wpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R9yax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W5ypw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O59iu6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(A*B*~(C)*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hdf88))
    _al_u3138 (
    .a(\u_cmsdk_mcu/HWDATA [0]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V59iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O59iu6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C3wpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tbvhu6 ));
  AL_MAP_LUT4 #(
    .EQN("~(~C*~(D)*~((B*A))+~C*D*~((B*A))+~(~C)*D*(B*A)+~C*D*(B*A))"),
    .INIT(16'h70f8))
    _al_u3139 (
    .a(\u_cmsdk_mcu/HWDATA [8]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O59iu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C30bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztupw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wouhu6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u314 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iqzhu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M8ipw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O34iu6 ));
  AL_MAP_LUT4 #(
    .EQN("~(~C*~(D)*~((B*A))+~C*D*~((B*A))+~(~C)*D*(B*A)+~C*D*(B*A))"),
    .INIT(16'h70f8))
    _al_u3140 (
    .a(\u_cmsdk_mcu/HWDATA [3]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O59iu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Owhbx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztupw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zmuhu6 ));
  AL_MAP_LUT4 #(
    .EQN("~(~C*~(D)*~((B*A))+~C*D*~((B*A))+~(~C)*D*(B*A)+~C*D*(B*A))"),
    .INIT(16'h70f8))
    _al_u3141 (
    .a(\u_cmsdk_mcu/HWDATA [4]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O59iu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ikhbx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztupw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gnuhu6 ));
  AL_MAP_LUT4 #(
    .EQN("~(~C*~(D)*~((B*A))+~C*D*~((B*A))+~(~C)*D*(B*A)+~C*D*(B*A))"),
    .INIT(16'h70f8))
    _al_u3142 (
    .a(\u_cmsdk_mcu/HWDATA [5]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O59iu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Czzax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztupw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nnuhu6 ));
  AL_MAP_LUT4 #(
    .EQN("~(~C*~(D)*~((B*A))+~C*D*~((B*A))+~(~C)*D*(B*A)+~C*D*(B*A))"),
    .INIT(16'h70f8))
    _al_u3143 (
    .a(\u_cmsdk_mcu/HWDATA [6]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O59iu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nt9bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztupw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bouhu6 ));
  AL_MAP_LUT4 #(
    .EQN("~(~C*~(D)*~((B*A))+~C*D*~((B*A))+~(~C)*D*(B*A)+~C*D*(B*A))"),
    .INIT(16'h70f8))
    _al_u3144 (
    .a(\u_cmsdk_mcu/HWDATA [7]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O59iu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C10bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztupw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pouhu6 ));
  AL_MAP_LUT4 #(
    .EQN("~(~C*~(D)*~((B*A))+~C*D*~((B*A))+~(~C)*D*(B*A)+~C*D*(B*A))"),
    .INIT(16'h70f8))
    _al_u3145 (
    .a(\u_cmsdk_mcu/HWDATA [9]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O59iu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tkjbx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztupw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dpuhu6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3146 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Apaiu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L45iu6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I82ju6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3147 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mmjiu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xq3pw6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u3148 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I82ju6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xq3pw6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Glaiu6 ),
    .d(_al_u1342_o),
    .o(_al_u3148_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3149 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D6kiu6_lutinv ),
    .b(_al_u1781_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Daiax6 ),
    .o(_al_u3149_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u315 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iqzhu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahdbx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B74iu6 ));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u3150 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Daiax6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 ),
    .o(_al_u3150_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(~A*~(D*B)))"),
    .INIT(16'he0a0))
    _al_u3151 (
    .a(_al_u609_o),
    .b(_al_u3150_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 ),
    .o(_al_u3151_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    _al_u3152 (
    .a(_al_u3148_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yavow6 ),
    .c(_al_u3149_o),
    .d(_al_u3151_o),
    .o(_al_u3152_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3153 (
    .a(_al_u3109_o),
    .b(_al_u1346_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vbiow6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(~B*~A)))"),
    .INIT(16'h010f))
    _al_u3154 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vbiow6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y0jiu6 ),
    .c(_al_u1264_o),
    .d(_al_u1266_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rcziu6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3155 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yljiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N3ziu6 ));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3156 (
    .a(_al_u1269_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N3ziu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 ),
    .o(_al_u3156_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(~B*~(~D*A)))"),
    .INIT(16'h0c0e))
    _al_u3157 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qe8iu6_lutinv ),
    .b(_al_u3156_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 ),
    .o(_al_u3157_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*~B))"),
    .INIT(8'ha8))
    _al_u3158 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qe8iu6_lutinv ),
    .b(_al_u606_o),
    .c(_al_u2829_o),
    .o(_al_u3158_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3159 (
    .a(_al_u1803_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vygax6 ),
    .o(_al_u3159_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u316 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iqzhu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H0ebx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I74iu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~B*~A*~(~D*C))"),
    .INIT(16'h1101))
    _al_u3160 (
    .a(_al_u3157_o),
    .b(_al_u3158_o),
    .c(_al_u3159_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ),
    .o(_al_u3160_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3161 (
    .a(_al_u3152_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rcziu6 ),
    .c(_al_u3160_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L18iu6 ));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    _al_u3162 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L18iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n1465 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3163 (
    .a(_al_u1344_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ifoiu6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*A)"),
    .INIT(16'h0080))
    _al_u3164 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ifoiu6_lutinv ),
    .b(_al_u909_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hgrpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 ),
    .o(_al_u3164_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u3165 (
    .a(_al_u3164_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F1jiu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y0jiu6 ),
    .o(_al_u3165_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(~D*C*B))"),
    .INIT(16'h5515))
    _al_u3166 (
    .a(_al_u904_o),
    .b(_al_u609_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ),
    .o(_al_u3166_o));
  AL_MAP_LUT4 #(
    .EQN("(C*A*~(D*B))"),
    .INIT(16'h20a0))
    _al_u3167 (
    .a(_al_u3165_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uyiiu6 ),
    .c(_al_u3166_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bziiu6_lutinv ),
    .o(_al_u3167_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3168 (
    .a(_al_u609_o),
    .b(_al_u903_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zzniu6_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u3169 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mmjiu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zzniu6_lutinv ),
    .o(_al_u3169_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u317 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iqzhu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ojebx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P74iu6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3170 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Us2ju6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yljiu6 ),
    .o(_al_u3170_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3171 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ldiow6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(~B*~A*~(D*C))"),
    .INIT(16'h0111))
    _al_u3172 (
    .a(_al_u3169_o),
    .b(_al_u3170_o),
    .c(_al_u1806_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ldiow6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1jiu6 ));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u3173 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gr2qw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6 ),
    .o(_al_u3173_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u3174 (
    .a(_al_u3167_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1jiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hviiu6 ),
    .d(_al_u3173_o),
    .o(_al_u3174_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~A*~(~C*~B))"),
    .INIT(16'h5400))
    _al_u3175 (
    .a(_al_u1812_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nyiiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hgrpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 ),
    .o(_al_u3175_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(~B*~(C*A)))"),
    .INIT(16'hec00))
    _al_u3176 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uyiiu6 ),
    .b(_al_u3175_o),
    .c(_al_u2373_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 ),
    .o(_al_u3176_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u3177 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N4kax6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4jax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dcziu6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3178 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dcziu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jckax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cwiiu6 ));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'h53))
    _al_u3179 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cwiiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rwjax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6 ),
    .o(_al_u3179_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u318 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iqzhu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Urgbx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W74iu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(~D*~C*A))"),
    .INIT(16'h3331))
    _al_u3180 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vviiu6 ),
    .b(_al_u3176_o),
    .c(_al_u3179_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 ),
    .o(_al_u3180_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u3181 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M1jiu6 ),
    .b(_al_u3174_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D0jiu6 ),
    .d(_al_u3180_o),
    .o(_al_u3181_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(A*~(D*B)))"),
    .INIT(16'h0d05))
    _al_u3182 (
    .a(_al_u3181_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vbiow6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ),
    .d(_al_u678_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D8iiu6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3183 (
    .a(_al_u2361_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9ypw6 ),
    .o(_al_u3183_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3184 (
    .a(_al_u1269_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nbkiu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 ),
    .o(_al_u3184_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3185 (
    .a(_al_u3183_o),
    .b(_al_u3184_o),
    .o(_al_u3185_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    _al_u3186 (
    .a(_al_u1812_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D6kiu6_lutinv ),
    .c(_al_u1813_o),
    .o(_al_u3186_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3187 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D6kiu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sy2ju6 ),
    .o(_al_u3187_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u3188 (
    .a(_al_u3186_o),
    .b(_al_u3187_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oeziu6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3189 (
    .a(_al_u3110_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 ),
    .o(_al_u3189_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u319 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iqzhu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jvkpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D84iu6 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u3190 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oeziu6 ),
    .b(_al_u3189_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 ),
    .o(_al_u3190_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3191 (
    .a(_al_u681_o),
    .b(_al_u696_o),
    .o(_al_u3191_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3192 (
    .a(_al_u606_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D6kiu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Daiax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G1aow6 ));
  AL_MAP_LUT4 #(
    .EQN("(~C*~B*~(D*A))"),
    .INIT(16'h0103))
    _al_u3193 (
    .a(_al_u604_o),
    .b(_al_u1907_o),
    .c(_al_u2392_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ),
    .o(_al_u3193_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(~C*A))"),
    .INIT(16'h31f5))
    _al_u3194 (
    .a(_al_u3191_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G1aow6 ),
    .c(_al_u3193_o),
    .d(_al_u1582_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fx9ow6 ));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B*~(~D*~A)))"),
    .INIT(16'h3070))
    _al_u3195 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rwjax6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Skjax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wv9ow6 ));
  AL_MAP_LUT4 #(
    .EQN("(C*B*~(D*A))"),
    .INIT(16'h40c0))
    _al_u3196 (
    .a(_al_u3185_o),
    .b(_al_u3190_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fx9ow6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wv9ow6 ),
    .o(_al_u3196_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u3197 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cwiiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P14qw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rwjax6 ),
    .o(_al_u3197_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u3198 (
    .a(_al_u3197_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Skjax6 ),
    .o(_al_u3198_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u3199 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vviiu6 ),
    .b(_al_u3198_o),
    .c(_al_u1269_o),
    .o(_al_u3199_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u320 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iqzhu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bp2qw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K84iu6 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u3200 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dcziu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jckax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jgxpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hbbow6 ));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u3201 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hbbow6 ),
    .b(_al_u679_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Frziu6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ya1ju6_lutinv ),
    .o(_al_u3201_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3202 (
    .a(_al_u3201_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 ),
    .o(_al_u3202_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*A*~(D*C))"),
    .INIT(16'h0222))
    _al_u3203 (
    .a(_al_u3196_o),
    .b(_al_u3199_o),
    .c(_al_u3202_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kxziu6_lutinv ),
    .o(_al_u3203_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u3204 (
    .a(_al_u1801_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ot7ow6 ));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3205 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uyiiu6 ),
    .b(_al_u3184_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hgrpw6 ),
    .o(_al_u3205_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u3206 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ot7ow6 ),
    .b(_al_u3205_o),
    .c(_al_u2767_o),
    .o(_al_u3206_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3207 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W0piu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vygax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Htyiu6 ));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*~C))"),
    .INIT(16'h8088))
    _al_u3208 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Htyiu6 ),
    .b(_al_u2771_o),
    .c(_al_u2370_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Skjax6 ),
    .o(_al_u3208_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~B*~(~D*A))"),
    .INIT(16'h0301))
    _al_u3209 (
    .a(_al_u2754_o),
    .b(_al_u1818_o),
    .c(_al_u3149_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ez1ju6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u321 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iqzhu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A6cbx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R84iu6 ));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*B*A)"),
    .INIT(16'h0800))
    _al_u3210 (
    .a(_al_u3203_o),
    .b(_al_u3206_o),
    .c(_al_u3208_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ez1ju6 ),
    .o(_al_u3210_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3211 (
    .a(_al_u3183_o),
    .b(_al_u1269_o),
    .o(_al_u3211_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    _al_u3212 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P14qw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wa0ju6 ));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3213 (
    .a(_al_u3211_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wa0ju6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Skjax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yo1ju6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3214 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N4kax6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6 ),
    .o(_al_u3214_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3215 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rwjax6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6 ),
    .o(_al_u3215_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(A*~(~D*~C)))"),
    .INIT(16'h1113))
    _al_u3216 (
    .a(_al_u3214_o),
    .b(_al_u3215_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4jax6 ),
    .o(_al_u3216_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D*~C*B))"),
    .INIT(16'ha2aa))
    _al_u3217 (
    .a(_al_u3216_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qxoiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N4kax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 ),
    .o(_al_u3217_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(~D*~C*B))"),
    .INIT(16'haaa2))
    _al_u3218 (
    .a(_al_u3217_o),
    .b(_al_u2380_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rwjax6 ),
    .o(_al_u3218_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D*~C*B))"),
    .INIT(16'ha2aa))
    _al_u3219 (
    .a(_al_u3210_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yo1ju6 ),
    .c(_al_u3218_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 ),
    .o(_al_u3219_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u322 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iqzhu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Drcbx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y84iu6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3220 (
    .a(_al_u677_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ls1ju6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u3221 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ls1ju6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pu1ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 ),
    .o(_al_u3221_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(~D*~C*B))"),
    .INIT(16'h5551))
    _al_u3222 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ujjiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mfjiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vygax6 ),
    .o(_al_u3222_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3223 (
    .a(_al_u909_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 ),
    .o(_al_u3223_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D*C*B))"),
    .INIT(16'h2aaa))
    _al_u3224 (
    .a(_al_u3222_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hs8ow6 ),
    .c(_al_u3223_o),
    .d(_al_u3124_o),
    .o(_al_u3224_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(~B*A))"),
    .INIT(8'h0d))
    _al_u3225 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qxoiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vygax6 ),
    .o(_al_u3225_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u3226 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W0piu6_lutinv ),
    .b(_al_u912_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ia8iu6_lutinv ),
    .d(_al_u3225_o),
    .o(_al_u3226_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3227 (
    .a(_al_u2364_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P14qw6 ),
    .o(_al_u3227_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(~A*~(~C*B)))"),
    .INIT(16'h00ae))
    _al_u3228 (
    .a(_al_u3227_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A95iu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xz9ow6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(D*C*B))"),
    .INIT(16'h1555))
    _al_u3229 (
    .a(_al_u3226_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W0piu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xz9ow6_lutinv ),
    .d(_al_u1269_o),
    .o(_al_u3229_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u323 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iqzhu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D2rpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F94iu6 ));
  AL_MAP_LUT4 #(
    .EQN("(C*B*~(D*~A))"),
    .INIT(16'h80c0))
    _al_u3230 (
    .a(_al_u3221_o),
    .b(_al_u3224_o),
    .c(_al_u3229_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pthiu6 ),
    .o(_al_u3230_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3231 (
    .a(_al_u2771_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F6ziu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rmiiu6 ));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u3232 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R9aiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Irmpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wkipw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wh0ju6 ));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u3233 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rmiiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Htyiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wh0ju6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 ),
    .o(_al_u3233_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~A*~(D*B))"),
    .INIT(16'h0105))
    _al_u3234 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jckax6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jgxpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N4kax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4jax6 ),
    .o(_al_u3234_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u3235 (
    .a(_al_u3219_o),
    .b(_al_u3230_o),
    .c(_al_u3233_o),
    .d(_al_u3234_o),
    .o(_al_u3235_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3236 (
    .a(_al_u609_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 ),
    .o(_al_u3236_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*B)*~(~D*A))"),
    .INIT(16'hf351))
    _al_u3237 (
    .a(_al_u1271_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D31ju6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ),
    .o(_al_u3237_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(~D*A))"),
    .INIT(16'h3f15))
    _al_u3238 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ls1ju6 ),
    .b(_al_u681_o),
    .c(_al_u3236_o),
    .d(_al_u3237_o),
    .o(_al_u3238_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    _al_u3239 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qe8iu6_lutinv ),
    .b(_al_u604_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 ),
    .o(_al_u3239_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u324 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iqzhu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bk7ax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ud4iu6 ));
  AL_MAP_LUT4 #(
    .EQN("(D*~(A*~(C*B)))"),
    .INIT(16'hd500))
    _al_u3240 (
    .a(_al_u3238_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eoyiu6_lutinv ),
    .c(_al_u3239_o),
    .d(_al_u3109_o),
    .o(_al_u3240_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*C)*~(~B*A))"),
    .INIT(16'hdd0d))
    _al_u3241 (
    .a(_al_u3235_o),
    .b(_al_u3240_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Crohu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(C*~A))"),
    .INIT(16'h8caf))
    _al_u3242 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hd8iu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yb8iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N4kax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S7mpw6 ),
    .o(_al_u3242_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*(C@B))"),
    .INIT(8'h14))
    _al_u3243 (
    .a(_al_u2783_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R9mpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sqkax6 ),
    .o(_al_u3243_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3244 (
    .a(_al_u2763_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9ypw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cbbiu6_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u3245 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cbbiu6_lutinv ),
    .b(_al_u2759_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4jax6 ),
    .o(_al_u3245_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3246 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J9kiu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 ),
    .o(_al_u3246_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    _al_u3247 (
    .a(_al_u912_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ia8iu6_lutinv ),
    .c(_al_u3246_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Habiu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u3248 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tc8iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Habiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T5mpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wfspw6 ),
    .o(_al_u3248_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u3249 (
    .a(_al_u3242_o),
    .b(_al_u3243_o),
    .c(_al_u3245_o),
    .d(_al_u3248_o),
    .o(_al_u3249_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u325 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iqzhu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ra2qw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T94iu6 ));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3250 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S88iu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Skjax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W7biu6 ));
  AL_MAP_LUT4 #(
    .EQN("(A*B*~(C)*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h7ee8))
    _al_u3251 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Irmpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S7mpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wfspw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wkipw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pyjiu6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(B@(A*C*~(D)+A*~(C)*D+~(A)*C*D+A*C*D))"),
    .INIT(16'h366c))
    _al_u3252 (
    .a(_al_u2785_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pyjiu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jckax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jgxpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ewjiu6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(B@(A*C*~(D)+A*~(C)*D+~(A)*C*D+A*C*D))"),
    .INIT(16'h366c))
    _al_u3253 (
    .a(_al_u2786_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ewjiu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N4kax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4jax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P7biu6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("~(A*~(~C*(D@B)))"),
    .INIT(16'h575d))
    _al_u3254 (
    .a(_al_u3249_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W7biu6 ),
    .c(_al_u2790_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P7biu6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S5biu6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3255 (
    .a(_al_u2467_o),
    .b(_al_u2468_o),
    .o(_al_u3255_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u3256 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U5yhu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bclpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sdlpw6 ),
    .o(_al_u3256_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*~A)"),
    .INIT(16'h0040))
    _al_u3257 (
    .a(_al_u3255_o),
    .b(_al_u3256_o),
    .c(_al_u1250_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jflpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fj1iu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~D*~A*~(C@B))"),
    .INIT(16'h0041))
    _al_u3258 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Krlpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rilpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y8lpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zslpw6 ),
    .o(_al_u3258_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3259 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fj1iu6 ),
    .b(_al_u3258_o),
    .o(_al_u3259_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u326 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iqzhu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yzqpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lm1iu6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3260 (
    .a(_al_u3259_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Golpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tezhu6 ));
  AL_MAP_LUT3 #(
    .EQN("~(C*~B*A)"),
    .INIT(8'hdf))
    _al_u3261 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tezhu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oulpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vplpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jq3iu6 ));
  AL_MAP_LUT3 #(
    .EQN("~(~C*B*A)"),
    .INIT(8'hf7))
    _al_u3262 (
    .a(_al_u3259_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Golpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vplpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W13iu6 ));
  AL_MAP_LUT4 #(
    .EQN("~(~C*~(D)*~((B*A))+~C*D*~((B*A))+~(~C)*D*(B*A)+~C*D*(B*A))"),
    .INIT(16'h70f8))
    _al_u3263 (
    .a(\u_cmsdk_mcu/HWDATA [10]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O59iu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C50bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztupw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kpuhu6 ));
  AL_MAP_LUT4 #(
    .EQN("(A*B*~(C)*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hdf88))
    _al_u3264 (
    .a(\u_cmsdk_mcu/HWDATA [2]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V59iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O59iu6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L1bbx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Smuhu6 ));
  AL_MAP_LUT4 #(
    .EQN("~(~C*~(D)*~((B*A))+~C*D*~((B*A))+~(~C)*D*(B*A)+~C*D*(B*A))"),
    .INIT(16'h70f8))
    _al_u3265 (
    .a(\u_cmsdk_mcu/HWDATA [11]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O59iu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D70bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztupw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rpuhu6 ));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3266 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wjyiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pjyiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C1wpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kwfiu6 ));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3267 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D5eiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pjyiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C1wpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K66iu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*~(B)*C*D)"),
    .INIT(16'h2077))
    _al_u3268 (
    .a(\u_cmsdk_mcu/HWDATA [3]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kwfiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K66iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Muhbx6 ),
    .o(_al_u3268_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3269 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[4] ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[5] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rmbpw6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u327 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iqzhu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L03qw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Df4iu6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3270 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M8row6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rmbpw6 ),
    .o(_al_u3270_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3271 (
    .a(_al_u3270_o),
    .b(_al_u1772_o),
    .o(_al_u3271_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u3272 (
    .a(_al_u3268_o),
    .b(_al_u1777_o),
    .c(_al_u3271_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O4phu6 ));
  AL_MAP_LUT4 #(
    .EQN("~(~C*~(D)*~((B*A))+~C*D*~((B*A))+~(~C)*D*(B*A)+~C*D*(B*A))"),
    .INIT(16'h70f8))
    _al_u3273 (
    .a(\u_cmsdk_mcu/HWDATA [12]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O59iu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E90bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztupw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ypuhu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*~(B)*C*D)"),
    .INIT(16'h2077))
    _al_u3274 (
    .a(\u_cmsdk_mcu/HWDATA [4]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kwfiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K66iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gihbx6 ),
    .o(_al_u3274_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3275 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rmbpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[2] ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[3] ),
    .o(_al_u3275_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3276 (
    .a(_al_u3275_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ukbpw6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Odfiu6_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u3277 (
    .a(_al_u3274_o),
    .b(_al_u1777_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Odfiu6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H4phu6 ));
  AL_MAP_LUT4 #(
    .EQN("~(~C*~(D)*~((B*A))+~C*D*~((B*A))+~(~C)*D*(B*A)+~C*D*(B*A))"),
    .INIT(16'h70f8))
    _al_u3278 (
    .a(\u_cmsdk_mcu/HWDATA [13]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O59iu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fb0bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztupw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fquhu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*~(B)*C*D)"),
    .INIT(16'h2077))
    _al_u3279 (
    .a(\u_cmsdk_mcu/HWDATA [5]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kwfiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K66iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mk3bx6 ),
    .o(_al_u3279_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u328 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iqzhu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P93qw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H34iu6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3280 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[0] ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[1] ),
    .o(_al_u3280_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3281 (
    .a(_al_u3275_o),
    .b(_al_u3280_o),
    .o(_al_u3281_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u3282 (
    .a(_al_u3279_o),
    .b(_al_u1777_o),
    .c(_al_u3281_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A4phu6 ));
  AL_MAP_LUT4 #(
    .EQN("~(~C*~(D)*~((B*A))+~C*D*~((B*A))+~(~C)*D*(B*A)+~C*D*(B*A))"),
    .INIT(16'h70f8))
    _al_u3283 (
    .a(\u_cmsdk_mcu/HWDATA [14]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O59iu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gd0bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztupw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tquhu6 ));
  AL_MAP_LUT4 #(
    .EQN("~(~C*~(D)*~((B*A))+~C*D*~((B*A))+~(~C)*D*(B*A)+~C*D*(B*A))"),
    .INIT(16'h70f8))
    _al_u3284 (
    .a(\u_cmsdk_mcu/HWDATA [17]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O59iu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jj0bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztupw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Csuhu6 ));
  AL_MAP_LUT4 #(
    .EQN("(A*B*~(C)*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hdf88))
    _al_u3285 (
    .a(\u_cmsdk_mcu/HWDATA [1]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V59iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O59iu6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cxzax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lmuhu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*~(B)*C*D)"),
    .INIT(16'h2077))
    _al_u3286 (
    .a(\u_cmsdk_mcu/HWDATA [9]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kwfiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K66iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rijbx6 ),
    .o(_al_u3286_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u3287 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rmbpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[2] ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[3] ),
    .o(_al_u3287_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3288 (
    .a(_al_u3287_o),
    .b(_al_u3280_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eegiu6_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u3289 (
    .a(_al_u3286_o),
    .b(_al_u1777_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eegiu6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uwdpw6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u329 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iqzhu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T3opw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oh4iu6 ));
  AL_MAP_LUT4 #(
    .EQN("~(~C*~(D)*~((B*A))+~C*D*~((B*A))+~(~C)*D*(B*A)+~C*D*(B*A))"),
    .INIT(16'h70f8))
    _al_u3290 (
    .a(\u_cmsdk_mcu/HWDATA [18]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O59iu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kl0bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztupw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qsuhu6 ));
  AL_MAP_LUT4 #(
    .EQN("~(~C*~(D)*~((B*A))+~C*D*~((B*A))+~(~C)*D*(B*A)+~C*D*(B*A))"),
    .INIT(16'h70f8))
    _al_u3291 (
    .a(\u_cmsdk_mcu/HWDATA [19]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O59iu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ln0bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztupw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Etuhu6 ));
  AL_MAP_LUT4 #(
    .EQN("~(~C*~(D)*~((B*A))+~C*D*~((B*A))+~(~C)*D*(B*A)+~C*D*(B*A))"),
    .INIT(16'h70f8))
    _al_u3292 (
    .a(\u_cmsdk_mcu/HWDATA [20]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O59iu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mp0bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztupw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Stuhu6 ));
  AL_MAP_LUT4 #(
    .EQN("~(~C*~(D)*~((B*A))+~C*D*~((B*A))+~(~C)*D*(B*A)+~C*D*(B*A))"),
    .INIT(16'h70f8))
    _al_u3293 (
    .a(\u_cmsdk_mcu/HWDATA [21]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O59iu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nr0bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztupw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Guuhu6 ));
  AL_MAP_LUT4 #(
    .EQN("~(~C*~(D)*~((B*A))+~C*D*~((B*A))+~(~C)*D*(B*A)+~C*D*(B*A))"),
    .INIT(16'h70f8))
    _al_u3294 (
    .a(\u_cmsdk_mcu/HWDATA [22]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O59iu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B3gbx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztupw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bvuhu6 ));
  AL_MAP_LUT4 #(
    .EQN("~(~C*~(D)*~((B*A))+~C*D*~((B*A))+~(~C)*D*(B*A)+~C*D*(B*A))"),
    .INIT(16'h70f8))
    _al_u3295 (
    .a(\u_cmsdk_mcu/HWDATA [23]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O59iu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ot0bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztupw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wvuhu6 ));
  AL_MAP_LUT4 #(
    .EQN("~(~C*~(D)*~((B*~A))+~C*D*~((B*~A))+~(~C)*D*(B*~A)+~C*D*(B*~A))"),
    .INIT(16'hb0f4))
    _al_u3296 (
    .a(_al_u2717_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O59iu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oxkpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztupw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dwuhu6 ));
  AL_MAP_LUT4 #(
    .EQN("~(~C*~(D)*~((B*~A))+~C*D*~((B*~A))+~(~C)*D*(B*~A)+~C*D*(B*~A))"),
    .INIT(16'hb0f4))
    _al_u3297 (
    .a(_al_u2721_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O59iu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pv0bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztupw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kwuhu6 ));
  AL_MAP_LUT4 #(
    .EQN("~(~C*~(D)*~((B*~A))+~C*D*~((B*~A))+~(~C)*D*(B*~A)+~C*D*(B*~A))"),
    .INIT(16'hb0f4))
    _al_u3298 (
    .a(_al_u2725_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O59iu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X5upw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztupw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rwuhu6 ));
  AL_MAP_LUT4 #(
    .EQN("~(~C*~(D)*~((B*~A))+~C*D*~((B*~A))+~(~C)*D*(B*~A)+~C*D*(B*~A))"),
    .INIT(16'hb0f4))
    _al_u3299 (
    .a(_al_u2729_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O59iu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qx0bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztupw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ywuhu6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u330 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iqzhu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q89bx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xi4iu6 ));
  AL_MAP_LUT4 #(
    .EQN("~(~C*~(D)*~((B*~A))+~C*D*~((B*~A))+~(~C)*D*(B*~A)+~C*D*(B*~A))"),
    .INIT(16'hb0f4))
    _al_u3300 (
    .a(_al_u2733_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O59iu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Usipw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztupw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fxuhu6 ));
  AL_MAP_LUT4 #(
    .EQN("~(~C*~(D)*~((B*A))+~C*D*~((B*A))+~(~C)*D*(B*A)+~C*D*(B*A))"),
    .INIT(16'h70f8))
    _al_u3301 (
    .a(\u_cmsdk_mcu/HWDATA [30]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O59iu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rz0bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztupw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ayuhu6 ));
  AL_MAP_LUT4 #(
    .EQN("~(~C*~(D)*~((B*A))+~C*D*~((B*A))+~(~C)*D*(B*A)+~C*D*(B*A))"),
    .INIT(16'h70f8))
    _al_u3302 (
    .a(\u_cmsdk_mcu/HWDATA [31]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O59iu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S0kbx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztupw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Acvhu6 ));
  AL_MAP_LUT4 #(
    .EQN("~(~C*~(D)*~((B*~A))+~C*D*~((B*~A))+~(~C)*D*(B*~A)+~C*D*(B*~A))"),
    .INIT(16'hb0f4))
    _al_u3303 (
    .a(_al_u2741_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O59iu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kojpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztupw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mxuhu6 ));
  AL_MAP_LUT4 #(
    .EQN("~(~C*~(D)*~((B*A))+~C*D*~((B*A))+~(~C)*D*(B*A)+~C*D*(B*A))"),
    .INIT(16'h70f8))
    _al_u3304 (
    .a(\u_cmsdk_mcu/HWDATA [16]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O59iu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ih0bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztupw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oruhu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*~B)*~(D*~A))"),
    .INIT(16'h8acf))
    _al_u3305 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hd8iu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yb8iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Irmpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 ),
    .o(_al_u3305_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*(C@(D*B)))"),
    .INIT(16'h1450))
    _al_u3306 (
    .a(_al_u2783_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R9mpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rskax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sqkax6 ),
    .o(_al_u3306_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u3307 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cbbiu6_lutinv ),
    .b(_al_u2759_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N4kax6 ),
    .o(_al_u3307_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u3308 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tc8iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Habiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jpmpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S7mpw6 ),
    .o(_al_u3308_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u3309 (
    .a(_al_u3305_o),
    .b(_al_u3306_o),
    .c(_al_u3307_o),
    .d(_al_u3308_o),
    .o(_al_u3309_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u331 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iqzhu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O1mpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gk4iu6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3310 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W7biu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P7biu6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zbjiu6 ));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3311 (
    .a(_al_u2787_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ewjiu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N4kax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ncjiu6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u3312 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Irmpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S7mpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wfspw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wkipw6 ),
    .o(_al_u3312_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u3313 (
    .a(_al_u3312_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pyjiu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ewjiu6_lutinv ),
    .o(_al_u3313_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D*C*B))"),
    .INIT(16'h2aaa))
    _al_u3314 (
    .a(_al_u3313_o),
    .b(_al_u2786_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ewjiu6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4jax6 ),
    .o(_al_u3314_o));
  AL_MAP_LUT2 #(
    .EQN("~(B@A)"),
    .INIT(4'h9))
    _al_u3315 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ncjiu6_lutinv ),
    .b(_al_u3314_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gcjiu6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("~(A*~(~D*(C@B)))"),
    .INIT(16'h557d))
    _al_u3316 (
    .a(_al_u3309_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zbjiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gcjiu6_lutinv ),
    .d(_al_u2790_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Agjiu6 ));
  AL_MAP_LUT3 #(
    .EQN("(~A*(C@B))"),
    .INIT(8'h14))
    _al_u3317 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Krlpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rilpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y8lpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yi1iu6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u3318 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fj1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yi1iu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P13iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zslpw6 ),
    .o(_al_u3318_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u3319 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cjqpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ehqpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T0ipw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/cpu0cdbgpwrupreq ),
    .o(_al_u3319_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u332 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iqzhu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gc1qw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pl4iu6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3320 (
    .a(_al_u3318_o),
    .b(_al_u3319_o),
    .o(_al_u3320_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(D*C*~B))"),
    .INIT(16'h4555))
    _al_u3321 (
    .a(_al_u3320_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cjqpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qwfax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Utqpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C53iu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u3322 (
    .a(_al_u3255_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mmyhu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Agyhu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A1zhu6_lutinv ),
    .o(_al_u3322_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(~D*C*~B))"),
    .INIT(16'haa8a))
    _al_u3323 (
    .a(_al_u3322_o),
    .b(_al_u3255_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T0zhu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y8lpw6 ),
    .o(_al_u3323_o));
  AL_MAP_LUT4 #(
    .EQN("~(D*~(A)*~((C*B))+D*A*~((C*B))+~(D)*A*(C*B)+D*A*(C*B))"),
    .INIT(16'h407f))
    _al_u3324 (
    .a(\u_cmsdk_mcu/dbg_swdo ),
    .b(_al_u1676_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Krlpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rilpw6 ),
    .o(_al_u3324_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u3325 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U03iu6 ),
    .b(_al_u3324_o),
    .c(_al_u1676_o),
    .o(_al_u3325_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u3326 (
    .a(_al_u529_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kalpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yklpw6 ),
    .o(_al_u3326_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u3327 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Agyhu6 ),
    .b(_al_u3326_o),
    .c(_al_u1757_o),
    .o(_al_u3327_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*A)"),
    .INIT(16'h0200))
    _al_u3328 (
    .a(_al_u1251_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jflpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kalpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yklpw6 ),
    .o(_al_u3328_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~B*~(~C*A))"),
    .INIT(16'h3100))
    _al_u3329 (
    .a(_al_u3327_o),
    .b(_al_u530_o),
    .c(_al_u3328_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U5yhu6 ),
    .o(_al_u3329_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u333 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iqzhu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gl1qw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ym4iu6 ));
  AL_MAP_LUT3 #(
    .EQN("(~(A)*~(B)*~(C)+~(A)*B*~(C)+A*~(B)*C+~(A)*B*C+A*B*C)"),
    .INIT(8'he5))
    _al_u3330 (
    .a(_al_u3325_o),
    .b(_al_u3329_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y8lpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/It3iu6_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C*~A))"),
    .INIT(8'h73))
    _al_u3331 (
    .a(_al_u3323_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/It3iu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U5yhu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rfxhu6 ));
  AL_MAP_LUT3 #(
    .EQN("(A*(C@B))"),
    .INIT(8'h28))
    _al_u3332 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/state_reg [0]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/state_reg [1]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/state_reg [2]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/next_state [2]));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*C)*~(B*A))"),
    .INIT(16'h7707))
    _al_u3333 (
    .a(\u_cmsdk_mcu/HWDATA [0]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kwfiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/apbsubsys_interrupt [0]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S11bx6 ),
    .o(_al_u3333_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D*~(C*B)))"),
    .INIT(16'h80aa))
    _al_u3334 (
    .a(_al_u3333_o),
    .b(\u_cmsdk_mcu/HWDATA [0]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K66iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U31bx6 ),
    .o(_al_u3334_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3335 (
    .a(_al_u3270_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ukbpw6_lutinv ),
    .o(_al_u3335_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u3336 (
    .a(_al_u3334_o),
    .b(_al_u1777_o),
    .c(_al_u3335_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J5phu6 ));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u3337 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/uart0_txovrint ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_ctrl [5]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_rx_overrun ),
    .o(_al_u3337_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*~C)*~(B*A))"),
    .INIT(16'h7770))
    _al_u3338 (
    .a(\u_cmsdk_mcu/HWDATA [8]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kwfiu6 ),
    .c(_al_u3337_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sq3bx6 ),
    .o(_al_u3338_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D*~(C*B)))"),
    .INIT(16'h80aa))
    _al_u3339 (
    .a(_al_u3338_o),
    .b(\u_cmsdk_mcu/HWDATA [8]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K66iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Us3bx6 ),
    .o(_al_u3339_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u334 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iqzhu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nv3qw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M94iu6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3340 (
    .a(_al_u3287_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ukbpw6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bggiu6_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u3341 (
    .a(_al_u3339_o),
    .b(_al_u1777_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bggiu6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bxdpw6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*~(B)*C*D)"),
    .INIT(16'h2077))
    _al_u3342 (
    .a(\u_cmsdk_mcu/HWDATA [2]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kwfiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K66iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5bbx6 ),
    .o(_al_u3342_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3343 (
    .a(_al_u3270_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A9row6_lutinv ),
    .o(_al_u3343_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u3344 (
    .a(_al_u3342_o),
    .b(_al_u1777_o),
    .c(_al_u3343_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V4phu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*~(B)*C*D)"),
    .INIT(16'h2077))
    _al_u3345 (
    .a(\u_cmsdk_mcu/HWDATA [11]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kwfiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K66iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lg1bx6 ),
    .o(_al_u3345_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3346 (
    .a(_al_u3287_o),
    .b(_al_u1772_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dagiu6_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u3347 (
    .a(_al_u3345_o),
    .b(_al_u1777_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dagiu6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y2phu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*~(B)*C*D)"),
    .INIT(16'h2077))
    _al_u3348 (
    .a(\u_cmsdk_mcu/HWDATA [13]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kwfiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K66iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rk1bx6 ),
    .o(_al_u3348_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3349 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[2] ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[3] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljbpw6_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u335 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iqzhu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ymwpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z54iu6 ));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3350 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rmbpw6 ),
    .b(_al_u3280_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljbpw6_lutinv ),
    .o(_al_u3350_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u3351 (
    .a(_al_u3348_o),
    .b(_al_u1777_o),
    .c(_al_u3350_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K2phu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*~(B)*C*D)"),
    .INIT(16'h2077))
    _al_u3352 (
    .a(\u_cmsdk_mcu/HWDATA [14]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kwfiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K66iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xo1bx6 ),
    .o(_al_u3352_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3353 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A9row6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rmbpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljbpw6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3giu6 ));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u3354 (
    .a(_al_u3352_o),
    .b(_al_u1777_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3giu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D2phu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u3355 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [12]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [13]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [14]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [15]),
    .o(_al_u3355_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u3356 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [0]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [1]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [10]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [11]),
    .o(_al_u3356_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u3357 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [6]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [7]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [8]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [9]),
    .o(_al_u3357_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u3358 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [2]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [4]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [5]),
    .o(_al_u3358_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u3359 (
    .a(_al_u3355_o),
    .b(_al_u3356_o),
    .c(_al_u3357_o),
    .d(_al_u3358_o),
    .o(_al_u3359_o));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~B*~A)"),
    .INIT(8'hfe))
    _al_u336 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D2opw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yzlpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgfax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T33iu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*~C)*~(B*A))"),
    .INIT(16'h7770))
    _al_u3360 (
    .a(\u_cmsdk_mcu/HWDATA [6]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kwfiu6 ),
    .c(_al_u3359_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jp9bx6 ),
    .o(_al_u3360_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D*~(C*B)))"),
    .INIT(16'h80aa))
    _al_u3361 (
    .a(_al_u3360_o),
    .b(\u_cmsdk_mcu/HWDATA [6]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K66iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lr9bx6 ),
    .o(_al_u3361_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3362 (
    .a(_al_u3275_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A9row6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G9fiu6_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u3363 (
    .a(_al_u3361_o),
    .b(_al_u1777_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G9fiu6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T3phu6 ));
  AL_MAP_LUT4 #(
    .EQN("(A*B*~(C)*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hdf88))
    _al_u3364 (
    .a(\u_cmsdk_mcu/HWDATA [15]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V59iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O59iu6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hf0bx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hruhu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u3365 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[12] ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[13] ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[14] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[15] ),
    .o(_al_u3365_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u3366 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[0] ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[1] ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[10] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[11] ),
    .o(_al_u3366_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u3367 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[6] ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[7] ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[8] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[9] ),
    .o(_al_u3367_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u3368 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[2] ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[3] ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[4] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[5] ),
    .o(_al_u3368_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u3369 (
    .a(_al_u3365_o),
    .b(_al_u3366_o),
    .c(_al_u3367_o),
    .d(_al_u3368_o),
    .o(_al_u3369_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u337 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inten_padded [0]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttype_padded [0]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpol_padded [0]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/new_masked_int [0]));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*~C)*~(B*A))"),
    .INIT(16'h7770))
    _al_u3370 (
    .a(\u_cmsdk_mcu/HWDATA [7]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kwfiu6 ),
    .c(_al_u3369_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Om3bx6 ),
    .o(_al_u3370_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D*~(C*B)))"),
    .INIT(16'h80aa))
    _al_u3371 (
    .a(_al_u3370_o),
    .b(\u_cmsdk_mcu/HWDATA [7]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K66iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qo3bx6 ),
    .o(_al_u3371_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3372 (
    .a(_al_u3275_o),
    .b(_al_u1772_o),
    .o(_al_u3372_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u3373 (
    .a(_al_u3371_o),
    .b(_al_u1777_o),
    .c(_al_u3372_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M3phu6 ));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3374 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K5eiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dtjow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C1wpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ch5iu6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*~A))"),
    .INIT(16'h23af))
    _al_u3375 (
    .a(_al_u2725_o),
    .b(_al_u1301_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ch5iu6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Avzax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ag5iu6 ));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u3376 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljbpw6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[4] ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[5] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ejbpw6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3377 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ejbpw6 ),
    .b(_al_u1772_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ajgiu6 ));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B*A))"),
    .INIT(8'h70))
    _al_u3378 (
    .a(_al_u1777_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ajgiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zdtpw6 ),
    .o(_al_u3378_o));
  AL_MAP_LUT4 #(
    .EQN("~(A*~(C*~(D*~B)))"),
    .INIT(16'hd5f5))
    _al_u3379 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ag5iu6 ),
    .b(_al_u2721_o),
    .c(_al_u3378_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ch5iu6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qmthu6 ));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u338 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inten_padded [1]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttype_padded [1]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpol_padded [1]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/new_masked_int [1]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3380 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ejbpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A9row6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rhgiu6 ));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B*A))"),
    .INIT(8'h70))
    _al_u3381 (
    .a(_al_u1777_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rhgiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mnmpw6 ),
    .o(_al_u3381_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+A*B*C*D)"),
    .INIT(16'hb3f0))
    _al_u3382 (
    .a(_al_u2729_o),
    .b(_al_u2733_o),
    .c(_al_u3381_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ch5iu6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xmthu6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u3383 (
    .a(_al_u2293_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M7zhu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lbyhu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u3384 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lbyhu6 ),
    .b(_al_u2299_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Krlpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y8lpw6 ),
    .o(_al_u3384_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    _al_u3385 (
    .a(_al_u3384_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pyyhu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rilpw6 ),
    .o(_al_u3385_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*~A)"),
    .INIT(8'h04))
    _al_u3386 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jflpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kalpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yklpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Swyhu6 ));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u3387 (
    .a(_al_u2296_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Swyhu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sdlpw6 ),
    .o(_al_u3387_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D*C*B))"),
    .INIT(16'h2aaa))
    _al_u3388 (
    .a(_al_u3387_o),
    .b(_al_u1308_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bclpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rilpw6 ),
    .o(_al_u3388_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3389 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Epyhu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kalpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sdlpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rkzhu6 ));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u339 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inten_padded [10]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttype_padded [10]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpol_padded [10]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/new_masked_int [10]));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3390 (
    .a(_al_u529_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Epyhu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kalpw6 ),
    .o(_al_u3390_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf513))
    _al_u3391 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rkzhu6 ),
    .b(_al_u3390_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bclpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rilpw6 ),
    .o(_al_u3391_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*A)"),
    .INIT(16'h0080))
    _al_u3392 (
    .a(_al_u3388_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I6yhu6_lutinv ),
    .c(_al_u3391_o),
    .d(_al_u2305_o),
    .o(_al_u3392_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*(C@B))"),
    .INIT(8'h14))
    _al_u3393 (
    .a(_al_u1761_o),
    .b(_al_u529_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kalpw6 ),
    .o(_al_u3393_o));
  AL_MAP_LUT4 #(
    .EQN("~(~C*~(D*~(B*~A)))"),
    .INIT(16'hfbf0))
    _al_u3394 (
    .a(_al_u3385_o),
    .b(_al_u3392_o),
    .c(_al_u3393_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U5yhu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zehpw6 [2]));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3395 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pthiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ),
    .o(_al_u3395_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u3396 (
    .a(_al_u1775_o),
    .b(_al_u3395_o),
    .c(_al_u1266_o),
    .o(_al_u3396_o));
  AL_MAP_LUT4 #(
    .EQN("(C*A*~(~D*B))"),
    .INIT(16'ha020))
    _al_u3397 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1jiu6 ),
    .b(_al_u1783_o),
    .c(_al_u3396_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 ),
    .o(_al_u3397_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(~D*C))"),
    .INIT(16'h8808))
    _al_u3398 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Epjiu6 ),
    .b(_al_u3397_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hviiu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P14qw6 ),
    .o(_al_u3398_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(A*~(D*B)))"),
    .INIT(16'h0d05))
    _al_u3399 (
    .a(_al_u3398_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vbiow6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ),
    .d(_al_u609_o),
    .o(_al_u3399_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u340 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inten_padded [11]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttype_padded [11]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpol_padded [11]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/new_masked_int [11]));
  AL_MAP_LUT4 #(
    .EQN("(~C*~B*~(D*A))"),
    .INIT(16'h0103))
    _al_u3400 (
    .a(_al_u2771_o),
    .b(_al_u2773_o),
    .c(_al_u2836_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6 ),
    .o(_al_u3400_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3401 (
    .a(_al_u2365_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 ),
    .o(_al_u3401_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(~C*~(~D*~B)))"),
    .INIT(16'ha0a2))
    _al_u3402 (
    .a(_al_u3400_o),
    .b(_al_u3401_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv ),
    .d(_al_u909_o),
    .o(_al_u3402_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3403 (
    .a(_al_u3402_o),
    .b(_al_u2771_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hm7ow6_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u3404 (
    .a(_al_u2832_o),
    .b(_al_u912_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ia8iu6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cn7ow6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*~B)*~(D*~A))"),
    .INIT(16'h8acf))
    _al_u3405 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hm7ow6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cn7ow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jckax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4jax6 ),
    .o(_al_u3405_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3406 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L45iu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dr7ow6 ));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C))"),
    .INIT(16'h02a2))
    _al_u3407 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S3kiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dr7ow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dk7ow6 ));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    _al_u3408 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dk7ow6 ),
    .b(_al_u1383_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Umkax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z6iow6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("~(~C*(~D*~(B)*~(A)+~D*B*~(A)+~(~D)*B*A+~D*B*A))"),
    .INIT(16'hf7f2))
    _al_u3409 (
    .a(_al_u3399_o),
    .b(_al_u3405_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z6iow6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Umkax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Leohu6 ));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u341 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inten_padded [12]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttype_padded [12]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpol_padded [12]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/new_masked_int [12]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(C*~A))"),
    .INIT(16'h8caf))
    _al_u3410 (
    .a(_al_u3402_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cn7ow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N4kax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4jax6 ),
    .o(_al_u3410_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    _al_u3411 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dk7ow6 ),
    .b(_al_u1765_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V6jax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jkhow6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("~(~C*(~D*~(B)*~(A)+~D*B*~(A)+~(~D)*B*A+~D*B*A))"),
    .INIT(16'hf7f2))
    _al_u3412 (
    .a(_al_u3399_o),
    .b(_al_u3410_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jkhow6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V6jax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Miohu6 ));
  AL_MAP_LUT4 #(
    .EQN("(D*~(~C*~B*~A))"),
    .INIT(16'hfe00))
    _al_u3413 (
    .a(_al_u906_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mfjiu6 ),
    .c(_al_u1359_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzjpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Am7ow6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u3414 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cbbiu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Am7ow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F4iax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6 ),
    .o(_al_u3414_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*~B))"),
    .INIT(8'h8a))
    _al_u3415 (
    .a(_al_u3414_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cn7ow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jgxpw6 ),
    .o(_al_u3415_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*~A))"),
    .INIT(8'h8c))
    _al_u3416 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hm7ow6_lutinv ),
    .b(_al_u3415_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jckax6 ),
    .o(_al_u3416_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*~(~D*B))"),
    .INIT(16'h5010))
    _al_u3417 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dk7ow6 ),
    .b(_al_u916_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fkrpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ubypw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pj7ow6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("~(~C*(~D*~(B)*~(A)+~D*B*~(A)+~(~D)*B*A+~D*B*A))"),
    .INIT(16'hf7f2))
    _al_u3418 (
    .a(_al_u3399_o),
    .b(_al_u3416_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pj7ow6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fkrpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssohu6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3419 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Skjax6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 ),
    .o(_al_u3419_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u342 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inten_padded [13]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttype_padded [13]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpol_padded [13]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/new_masked_int [13]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u3420 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rmiiu6 ),
    .b(_al_u2832_o),
    .c(_al_u3419_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6 ),
    .o(_al_u3420_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u3421 (
    .a(_al_u3420_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aaiiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kmiiu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 ),
    .o(_al_u3421_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*~B))"),
    .INIT(8'h8a))
    _al_u3422 (
    .a(_al_u3421_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljiiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wkipw6 ),
    .o(_al_u3422_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u3423 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I6row6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 ),
    .o(_al_u3423_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(~C*~B*~A))"),
    .INIT(16'hfe00))
    _al_u3424 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iekax6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lgkax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oikax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rkkax6 ),
    .o(_al_u3424_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u3425 (
    .a(_al_u3423_o),
    .b(_al_u3424_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hoiiu6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("~(~C*(~D*~(B)*~(A)+~D*B*~(A)+~(~D)*B*A+~D*B*A))"),
    .INIT(16'hf7f2))
    _al_u3426 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D8iiu6 ),
    .b(_al_u3422_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hoiiu6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rkkax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cfthu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(D@C)*~(B*A))"),
    .INIT(16'h7007))
    _al_u3427 (
    .a(_al_u1255_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Krlpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qwfax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Utqpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S63iu6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("~(~A*~(D*~(C*B)))"),
    .INIT(16'hbfaa))
    _al_u3428 (
    .a(_al_u3320_o),
    .b(_al_u1253_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S63iu6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ryfax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rtxhu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~C*B*~(D*~A))"),
    .INIT(16'h080c))
    _al_u3429 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I6yhu6_lutinv ),
    .b(_al_u3391_o),
    .c(_al_u3328_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yklpw6 ),
    .o(_al_u3429_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u343 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inten_padded [14]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttype_padded [14]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpol_padded [14]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/new_masked_int [14]));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(~B*(D@A)))"),
    .INIT(16'h0e0d))
    _al_u3430 (
    .a(_al_u1756_o),
    .b(_al_u1761_o),
    .c(_al_u1763_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yklpw6 ),
    .o(_al_u3430_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*~A))"),
    .INIT(8'h8c))
    _al_u3431 (
    .a(_al_u3429_o),
    .b(_al_u3430_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U5yhu6 ),
    .o(_al_u3431_o));
  AL_MAP_LUT4 #(
    .EQN("~(B*~(~D*C*~A))"),
    .INIT(16'h3373))
    _al_u3432 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mmyhu6 ),
    .b(_al_u3431_o),
    .c(_al_u1253_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kwlpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zehpw6 [4]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3433 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_raw_intstatus [0]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_intmask [0]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/apbsubsys_interrupt [10]));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(C*A))"),
    .INIT(16'h5f13))
    _al_u3434 (
    .a(\u_cmsdk_mcu/HWDATA [10]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/apbsubsys_interrupt [10]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kwfiu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ca1bx6 ),
    .o(_al_u3434_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D*~(C*B)))"),
    .INIT(16'h80aa))
    _al_u3435 (
    .a(_al_u3434_o),
    .b(\u_cmsdk_mcu/HWDATA [10]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K66iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fc1bx6 ),
    .o(_al_u3435_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3436 (
    .a(_al_u3287_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A9row6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hcgiu6_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u3437 (
    .a(_al_u3435_o),
    .b(_al_u1777_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hcgiu6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F3phu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*B)*~(~D*A))"),
    .INIT(16'hf351))
    _al_u3438 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_raw_intstatus [4]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_raw_intstatus [2]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_intmask [2]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_intmask [4]),
    .o(_al_u3438_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*B)*~(~D*A))"),
    .INIT(16'hf351))
    _al_u3439 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_raw_intstatus [5]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_raw_intstatus [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_intmask [3]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_intmask [5]),
    .o(_al_u3439_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u344 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inten_padded [15]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttype_padded [15]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpol_padded [15]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/new_masked_int [15]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3440 (
    .a(_al_u3438_o),
    .b(_al_u3439_o),
    .o(_al_u3440_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*~B)*~(C*A))"),
    .INIT(16'h5f4c))
    _al_u3441 (
    .a(\u_cmsdk_mcu/HWDATA [12]),
    .b(_al_u3440_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kwfiu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W51bx6 ),
    .o(_al_u3441_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D*~(C*B)))"),
    .INIT(16'h80aa))
    _al_u3442 (
    .a(_al_u3441_o),
    .b(\u_cmsdk_mcu/HWDATA [12]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K66iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z71bx6 ),
    .o(_al_u3442_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3443 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ukbpw6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rmbpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljbpw6_lutinv ),
    .o(_al_u3443_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u3444 (
    .a(_al_u3442_o),
    .b(_al_u1777_o),
    .c(_al_u3443_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R2phu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*~(B)*C*D)"),
    .INIT(16'h2077))
    _al_u3445 (
    .a(\u_cmsdk_mcu/HWDATA [15]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kwfiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K66iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yxrpw6 ),
    .o(_al_u3445_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3446 (
    .a(_al_u1772_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rmbpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljbpw6_lutinv ),
    .o(_al_u3446_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u3447 (
    .a(_al_u3445_o),
    .b(_al_u1777_o),
    .c(_al_u3446_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W1phu6 ));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B*A))"),
    .INIT(8'h70))
    _al_u3448 (
    .a(\u_cmsdk_mcu/HWDATA [17]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K66iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dt1bx6 ),
    .o(_al_u3448_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3449 (
    .a(\u_cmsdk_mcu/HWDATA [17]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kwfiu6 ),
    .o(_al_u3449_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u345 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inten_padded [2]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttype_padded [2]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpol_padded [2]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/new_masked_int [2]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u3450 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_raw_intstatus [7]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [1]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_intmask [7]),
    .o(_al_u3450_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~A*~(~D*~C))"),
    .INIT(16'h1110))
    _al_u3451 (
    .a(_al_u3448_o),
    .b(_al_u3449_o),
    .c(_al_u3450_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ar1bx6 ),
    .o(_al_u3451_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u3452 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[4] ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[5] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uybpw6_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3453 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M8row6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uybpw6_lutinv ),
    .o(_al_u3453_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3454 (
    .a(_al_u3453_o),
    .b(_al_u3280_o),
    .o(_al_u3454_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u3455 (
    .a(_al_u3451_o),
    .b(_al_u1777_o),
    .c(_al_u3454_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I1phu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*C)*~(B*A))"),
    .INIT(16'h7707))
    _al_u3456 (
    .a(\u_cmsdk_mcu/HWDATA [1]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kwfiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/apbsubsys_interrupt [1]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y72bx6 ),
    .o(_al_u3456_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D*~(C*B)))"),
    .INIT(16'h80aa))
    _al_u3457 (
    .a(_al_u3456_o),
    .b(\u_cmsdk_mcu/HWDATA [1]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K66iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aa2bx6 ),
    .o(_al_u3457_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3458 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M8row6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rmbpw6 ),
    .c(_al_u3280_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yogiu6_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u3459 (
    .a(_al_u3457_o),
    .b(_al_u1777_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yogiu6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C5phu6 ));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u346 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inten_padded [3]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttype_padded [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpol_padded [3]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/new_masked_int [3]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B*A))"),
    .INIT(8'h70))
    _al_u3460 (
    .a(\u_cmsdk_mcu/HWDATA [18]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K66iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P12bx6 ),
    .o(_al_u3460_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3461 (
    .a(\u_cmsdk_mcu/HWDATA [18]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kwfiu6 ),
    .o(_al_u3461_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~A*~(~D*C))"),
    .INIT(16'h1101))
    _al_u3462 (
    .a(_al_u3460_o),
    .b(_al_u3461_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [2]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mz1bx6 ),
    .o(_al_u3462_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3463 (
    .a(_al_u3453_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A9row6_lutinv ),
    .o(_al_u3463_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u3464 (
    .a(_al_u3462_o),
    .b(_al_u1777_o),
    .c(_al_u3463_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B1phu6 ));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B*A))"),
    .INIT(8'h70))
    _al_u3465 (
    .a(\u_cmsdk_mcu/HWDATA [19]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K66iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V52bx6 ),
    .o(_al_u3465_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3466 (
    .a(\u_cmsdk_mcu/HWDATA [19]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kwfiu6 ),
    .o(_al_u3466_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~A*~(~D*C))"),
    .INIT(16'h1101))
    _al_u3467 (
    .a(_al_u3465_o),
    .b(_al_u3466_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [3]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S32bx6 ),
    .o(_al_u3467_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3468 (
    .a(_al_u3453_o),
    .b(_al_u1772_o),
    .o(_al_u3468_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u3469 (
    .a(_al_u3467_o),
    .b(_al_u1777_o),
    .c(_al_u3468_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U0phu6 ));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u347 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inten_padded [4]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttype_padded [4]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpol_padded [4]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/new_masked_int [4]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B*A))"),
    .INIT(8'h70))
    _al_u3470 (
    .a(\u_cmsdk_mcu/HWDATA [20]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K66iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fe2bx6 ),
    .o(_al_u3470_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3471 (
    .a(\u_cmsdk_mcu/HWDATA [20]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kwfiu6 ),
    .o(_al_u3471_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~A*~(~D*C))"),
    .INIT(16'h1101))
    _al_u3472 (
    .a(_al_u3470_o),
    .b(_al_u3471_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [4]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cc2bx6 ),
    .o(_al_u3472_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3473 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uybpw6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[2] ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[3] ),
    .o(_al_u3473_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3474 (
    .a(_al_u3473_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ukbpw6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lhdiu6_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u3475 (
    .a(_al_u3472_o),
    .b(_al_u1777_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lhdiu6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N0phu6 ));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B*A))"),
    .INIT(8'h70))
    _al_u3476 (
    .a(\u_cmsdk_mcu/HWDATA [21]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K66iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Li2bx6 ),
    .o(_al_u3476_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3477 (
    .a(\u_cmsdk_mcu/HWDATA [21]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kwfiu6 ),
    .o(_al_u3477_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~A*~(~D*C))"),
    .INIT(16'h1101))
    _al_u3478 (
    .a(_al_u3476_o),
    .b(_al_u3477_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [5]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ig2bx6 ),
    .o(_al_u3478_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3479 (
    .a(_al_u3473_o),
    .b(_al_u3280_o),
    .o(_al_u3479_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u348 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inten_padded [5]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttype_padded [5]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpol_padded [5]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/new_masked_int [5]));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u3480 (
    .a(_al_u3478_o),
    .b(_al_u1777_o),
    .c(_al_u3479_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G0phu6 ));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B*A))"),
    .INIT(8'h70))
    _al_u3481 (
    .a(\u_cmsdk_mcu/HWDATA [22]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K66iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y0gbx6 ),
    .o(_al_u3481_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3482 (
    .a(\u_cmsdk_mcu/HWDATA [22]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kwfiu6 ),
    .o(_al_u3482_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~A*~(~D*C))"),
    .INIT(16'h1101))
    _al_u3483 (
    .a(_al_u3481_o),
    .b(_al_u3482_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [6]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vyfbx6 ),
    .o(_al_u3483_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3484 (
    .a(_al_u3473_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A9row6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nbdiu6_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u3485 (
    .a(_al_u3483_o),
    .b(_al_u1777_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nbdiu6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zzohu6 ));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B*A))"),
    .INIT(8'h70))
    _al_u3486 (
    .a(\u_cmsdk_mcu/HWDATA [23]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K66iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xq2bx6 ),
    .o(_al_u3486_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3487 (
    .a(\u_cmsdk_mcu/HWDATA [23]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kwfiu6 ),
    .o(_al_u3487_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~A*~(~D*C))"),
    .INIT(16'h1101))
    _al_u3488 (
    .a(_al_u3486_o),
    .b(_al_u3487_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [7]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uo2bx6 ),
    .o(_al_u3488_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3489 (
    .a(_al_u3473_o),
    .b(_al_u1772_o),
    .o(_al_u3489_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u349 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inten_padded [6]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttype_padded [6]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpol_padded [6]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/new_masked_int [6]));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u3490 (
    .a(_al_u3488_o),
    .b(_al_u1777_o),
    .c(_al_u3489_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Szohu6 ));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B*~A))"),
    .INIT(8'hb0))
    _al_u3491 (
    .a(_al_u2717_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K66iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dv2bx6 ),
    .o(_al_u3491_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u3492 (
    .a(_al_u2717_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kwfiu6 ),
    .o(_al_u3492_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~A*~(~D*C))"),
    .INIT(16'h1101))
    _al_u3493 (
    .a(_al_u3491_o),
    .b(_al_u3492_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [8]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/At2bx6 ),
    .o(_al_u3493_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u3494 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uybpw6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[2] ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[3] ),
    .o(_al_u3494_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3495 (
    .a(_al_u3494_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ukbpw6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jzfiu6_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u3496 (
    .a(_al_u3493_o),
    .b(_al_u1777_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jzfiu6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nwdpw6 ));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B*~A))"),
    .INIT(8'hb0))
    _al_u3497 (
    .a(_al_u2721_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K66iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rm2bx6 ),
    .o(_al_u3497_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u3498 (
    .a(_al_u2721_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kwfiu6 ),
    .o(_al_u3498_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~A*~(~D*C))"),
    .INIT(16'h1101))
    _al_u3499 (
    .a(_al_u3497_o),
    .b(_al_u3498_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [9]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ok2bx6 ),
    .o(_al_u3499_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u350 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inten_padded [7]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttype_padded [7]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpol_padded [7]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/new_masked_int [7]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3500 (
    .a(_al_u3494_o),
    .b(_al_u3280_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mxfiu6_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u3501 (
    .a(_al_u3499_o),
    .b(_al_u1777_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mxfiu6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gwdpw6 ));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B*~A))"),
    .INIT(8'hb0))
    _al_u3502 (
    .a(_al_u2725_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K66iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jz2bx6 ),
    .o(_al_u3502_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u3503 (
    .a(_al_u2725_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kwfiu6 ),
    .o(_al_u3503_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~A*~(~D*C))"),
    .INIT(16'h1101))
    _al_u3504 (
    .a(_al_u3502_o),
    .b(_al_u3503_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [10]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gx2bx6 ),
    .o(_al_u3504_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3505 (
    .a(_al_u3494_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A9row6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ivfiu6_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u3506 (
    .a(_al_u3504_o),
    .b(_al_u1777_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ivfiu6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lzohu6 ));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B*~A))"),
    .INIT(8'hb0))
    _al_u3507 (
    .a(_al_u2729_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K66iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P33bx6 ),
    .o(_al_u3507_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u3508 (
    .a(_al_u2729_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kwfiu6 ),
    .o(_al_u3508_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~A*~(~D*C))"),
    .INIT(16'h1101))
    _al_u3509 (
    .a(_al_u3507_o),
    .b(_al_u3508_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [11]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M13bx6 ),
    .o(_al_u3509_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u351 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inten_padded [8]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttype_padded [8]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpol_padded [8]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/new_masked_int [8]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3510 (
    .a(_al_u3494_o),
    .b(_al_u1772_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Etfiu6_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u3511 (
    .a(_al_u3509_o),
    .b(_al_u1777_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Etfiu6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ezohu6 ));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B*~A))"),
    .INIT(8'hb0))
    _al_u3512 (
    .a(_al_u2733_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K66iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V73bx6 ),
    .o(_al_u3512_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u3513 (
    .a(_al_u2733_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kwfiu6 ),
    .o(_al_u3513_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~A*~(~D*C))"),
    .INIT(16'h1101))
    _al_u3514 (
    .a(_al_u3512_o),
    .b(_al_u3513_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [12]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S53bx6 ),
    .o(_al_u3514_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3515 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ukbpw6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljbpw6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uybpw6_lutinv ),
    .o(_al_u3515_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u3516 (
    .a(_al_u3514_o),
    .b(_al_u1777_o),
    .c(_al_u3515_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xyohu6 ));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B*A))"),
    .INIT(8'h70))
    _al_u3517 (
    .a(\u_cmsdk_mcu/HWDATA [30]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K66iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tcipw6 ),
    .o(_al_u3517_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3518 (
    .a(\u_cmsdk_mcu/HWDATA [30]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kwfiu6 ),
    .o(_al_u3518_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~A*~(~D*C))"),
    .INIT(16'h1101))
    _al_u3519 (
    .a(_al_u3517_o),
    .b(_al_u3518_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [14]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qaipw6 ),
    .o(_al_u3519_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u352 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inten_padded [9]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttype_padded [9]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpol_padded [9]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/new_masked_int [9]));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3520 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A9row6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljbpw6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uybpw6_lutinv ),
    .o(_al_u3520_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u3521 (
    .a(_al_u3519_o),
    .b(_al_u1777_o),
    .c(_al_u3520_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jyohu6 ));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B*A))"),
    .INIT(8'h70))
    _al_u3522 (
    .a(\u_cmsdk_mcu/HWDATA [31]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K66iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hg3bx6 ),
    .o(_al_u3522_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3523 (
    .a(\u_cmsdk_mcu/HWDATA [31]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kwfiu6 ),
    .o(_al_u3523_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~A*~(~D*C))"),
    .INIT(16'h1101))
    _al_u3524 (
    .a(_al_u3522_o),
    .b(_al_u3523_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [15]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ee3bx6 ),
    .o(_al_u3524_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3525 (
    .a(_al_u1772_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljbpw6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uybpw6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Webiu6 ));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u3526 (
    .a(_al_u3524_o),
    .b(_al_u1777_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Webiu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cyohu6 ));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B*~A))"),
    .INIT(8'hb0))
    _al_u3527 (
    .a(_al_u2741_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K66iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bc3bx6 ),
    .o(_al_u3527_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u3528 (
    .a(_al_u2741_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kwfiu6 ),
    .o(_al_u3528_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~A*~(~D*C))"),
    .INIT(16'h1101))
    _al_u3529 (
    .a(_al_u3527_o),
    .b(_al_u3528_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [13]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y93bx6 ),
    .o(_al_u3529_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u353 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .o(\u_cmsdk_mcu/u_ahb_ram/mux3_b0_sel_is_2_o ));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3530 (
    .a(_al_u3280_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljbpw6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uybpw6_lutinv ),
    .o(_al_u3530_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u3531 (
    .a(_al_u3529_o),
    .b(_al_u1777_o),
    .c(_al_u3530_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qyohu6 ));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B*A))"),
    .INIT(8'h70))
    _al_u3532 (
    .a(\u_cmsdk_mcu/HWDATA [16]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K66iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jx1bx6 ),
    .o(_al_u3532_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3533 (
    .a(\u_cmsdk_mcu/HWDATA [16]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kwfiu6 ),
    .o(_al_u3533_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u3534 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_raw_intstatus [6]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [0]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_intmask [6]),
    .o(_al_u3534_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~A*~(~D*~C))"),
    .INIT(16'h1110))
    _al_u3535 (
    .a(_al_u3532_o),
    .b(_al_u3533_o),
    .c(_al_u3534_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gv1bx6 ),
    .o(_al_u3535_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3536 (
    .a(_al_u3453_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ukbpw6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hwhiu6_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u3537 (
    .a(_al_u3535_o),
    .b(_al_u1777_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hwhiu6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P1phu6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3538 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cbbiu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rwjax6 ),
    .o(_al_u3538_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B@A))"),
    .INIT(8'h90))
    _al_u3539 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P14qw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 ),
    .o(_al_u3539_o));
  AL_MAP_LUT3 #(
    .EQN("(A*B*~(C)+A*~(B)*C+~(A)*B*C+A*B*C)"),
    .INIT(8'he8))
    _al_u354 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rxd_lpf [0]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rxd_lpf [1]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rxd_lpf [2]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_shift_in ));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*~A)"),
    .INIT(16'h0040))
    _al_u3540 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv ),
    .b(_al_u3539_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9ypw6 ),
    .o(_al_u3540_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*B*~(D*A))"),
    .INIT(16'h040c))
    _al_u3541 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Am7ow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kubow6 ),
    .c(_al_u3540_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G2iax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wtbow6 ));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*~(D*~B))"),
    .INIT(16'h4050))
    _al_u3542 (
    .a(_al_u3538_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cn7ow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wtbow6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wkipw6 ),
    .o(_al_u3542_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*~A))"),
    .INIT(8'h8c))
    _al_u3543 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hm7ow6_lutinv ),
    .b(_al_u3542_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jgxpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Itbow6 ));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    _al_u3544 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dk7ow6 ),
    .b(_al_u916_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ubypw6 ),
    .o(_al_u3544_o));
  AL_MAP_LUT4 #(
    .EQN("~(~C*(~D*~(B)*~(A)+~D*B*~(A)+~(~D)*B*A+~D*B*A))"),
    .INIT(16'hf7f2))
    _al_u3545 (
    .a(_al_u3399_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Itbow6 ),
    .c(_al_u3544_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ubypw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tpohu6 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u3546 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aaiiu6 ),
    .b(_al_u2832_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eciiu6 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*~A))"),
    .INIT(8'h8c))
    _al_u3547 (
    .a(_al_u2827_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eciiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rwjax6 ),
    .o(_al_u3547_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*~B))"),
    .INIT(8'h8a))
    _al_u3548 (
    .a(_al_u3547_o),
    .b(_al_u2841_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S7mpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xbiiu6 ));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    _al_u3549 (
    .a(_al_u3423_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iekax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lgkax6 ),
    .o(_al_u3549_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u355 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_tick_cnt [2]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_tick_cnt [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/BAUDTICK ),
    .o(_al_u355_o));
  AL_MAP_LUT4 #(
    .EQN("~(~C*(~D*~(B)*~(A)+~D*B*~(A)+~(~D)*B*A+~D*B*A))"),
    .INIT(16'hf7f2))
    _al_u3550 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D8iiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xbiiu6 ),
    .c(_al_u3549_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lgkax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qfthu6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3551 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cwiiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujiu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yy7ow6 ));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*A)"),
    .INIT(16'h0080))
    _al_u3552 (
    .a(_al_u2771_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yy7ow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qxoiu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 ),
    .o(_al_u3552_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(D*C*~B))"),
    .INIT(16'h4555))
    _al_u3553 (
    .a(_al_u3552_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nbkiu6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dmiiu6 ),
    .o(_al_u3553_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*~A)"),
    .INIT(8'h04))
    _al_u3554 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jckax6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N4kax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4jax6 ),
    .o(_al_u3554_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u3555 (
    .a(_al_u2369_o),
    .b(_al_u3554_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Skjax6 ),
    .o(_al_u3555_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(A*~(D*C)))"),
    .INIT(16'hc444))
    _al_u3556 (
    .a(_al_u3553_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uyiiu6 ),
    .c(_al_u2832_o),
    .d(_al_u3555_o),
    .o(_al_u3556_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3557 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ot7ow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wkipw6 ),
    .o(_al_u3557_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3558 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dr7ow6 ),
    .b(_al_u604_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ),
    .o(_al_u3558_o));
  AL_MAP_LUT4 #(
    .EQN("(A*(~C*~(B)*~(D)+~C*B*~(D)+~(~C)*B*D+~C*B*D))"),
    .INIT(16'h880a))
    _al_u3559 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U98iu6 ),
    .b(_al_u1266_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 ),
    .o(_al_u3559_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u356 (
    .a(_al_u355_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_tick_cnt [0]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_tick_cnt [1]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_state_inc ));
  AL_MAP_LUT4 #(
    .EQN("(~C*B*~(~D*~A))"),
    .INIT(16'h0c08))
    _al_u3560 (
    .a(_al_u682_o),
    .b(_al_u1346_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ),
    .o(_al_u3560_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u3561 (
    .a(_al_u3169_o),
    .b(_al_u3558_o),
    .c(_al_u3559_o),
    .d(_al_u3560_o),
    .o(_al_u3561_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(~B*~(~D*C)))"),
    .INIT(16'h88a8))
    _al_u3562 (
    .a(_al_u2361_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6 ),
    .o(_al_u3562_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~A*~(D*C))"),
    .INIT(16'h0111))
    _al_u3563 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ujjiu6 ),
    .b(_al_u3186_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zzniu6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv ),
    .o(_al_u3563_o));
  AL_MAP_LUT4 #(
    .EQN("(C*A*~(D*B))"),
    .INIT(16'h20a0))
    _al_u3564 (
    .a(_al_u3561_o),
    .b(_al_u3562_o),
    .c(_al_u3563_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M7kiu6 ),
    .o(_al_u3564_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*~A)"),
    .INIT(16'h1000))
    _al_u3565 (
    .a(_al_u3556_o),
    .b(_al_u3557_o),
    .c(_al_u3564_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lv7ow6 ),
    .o(_al_u3565_o));
  AL_MAP_LUT4 #(
    .EQN("~(~C*~(A*~(D*B)))"),
    .INIT(16'hf2fa))
    _al_u3566 (
    .a(_al_u3565_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vbiow6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ),
    .d(_al_u678_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O25iu6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3567 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N98iu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vxniu6_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3568 (
    .a(_al_u1266_o),
    .b(_al_u1271_o),
    .c(_al_u1342_o),
    .o(_al_u3568_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D*~C*A))"),
    .INIT(16'h3133))
    _al_u3569 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vxniu6_lutinv ),
    .b(_al_u3568_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ),
    .o(_al_u3569_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u357 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [12]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [13]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [14]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [15]),
    .o(_al_u357_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u3570 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P8oiu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 ),
    .o(_al_u3570_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*A*~(D*C))"),
    .INIT(16'h0222))
    _al_u3571 (
    .a(_al_u3569_o),
    .b(_al_u3570_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y0jiu6 ),
    .d(_al_u604_o),
    .o(_al_u3571_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u3572 (
    .a(_al_u906_o),
    .b(_al_u932_o),
    .c(_al_u2403_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rvniu6 ));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u3573 (
    .a(_al_u3571_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rvniu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mfjiu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pthiu6 ),
    .o(_al_u3573_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3574 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Llaow6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ldoiu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 ),
    .o(_al_u3574_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3575 (
    .a(_al_u1296_o),
    .b(_al_u1344_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vo3ju6_lutinv ),
    .o(_al_u3575_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u3576 (
    .a(_al_u3575_o),
    .b(_al_u1781_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pthiu6 ),
    .o(_al_u3576_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(C*~(~D*~A)))"),
    .INIT(16'h0c4c))
    _al_u3577 (
    .a(_al_u3574_o),
    .b(_al_u3576_o),
    .c(_al_u607_o),
    .d(_al_u1329_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Faoiu6 ));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3578 (
    .a(_al_u1781_o),
    .b(_al_u3122_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 ),
    .o(_al_u3578_o));
  AL_MAP_LUT4 #(
    .EQN("(C*A*~(D*~B))"),
    .INIT(16'h80a0))
    _al_u3579 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qyniu6_lutinv ),
    .b(_al_u2403_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 ),
    .o(_al_u3579_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u358 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [0]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [1]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [10]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [11]),
    .o(_al_u358_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~B*~(D*A))"),
    .INIT(16'h0103))
    _al_u3580 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zzniu6_lutinv ),
    .b(_al_u3578_o),
    .c(_al_u3579_o),
    .d(_al_u607_o),
    .o(_al_u3580_o));
  AL_MAP_LUT4 #(
    .EQN("(C*A*~(D*~B))"),
    .INIT(16'h80a0))
    _al_u3581 (
    .a(_al_u3573_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Faoiu6 ),
    .c(_al_u3580_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ),
    .o(_al_u3581_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3582 (
    .a(_al_u1635_o),
    .b(_al_u678_o),
    .c(_al_u679_o),
    .o(_al_u3582_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3583 (
    .a(_al_u3118_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Edapw6_lutinv ),
    .o(_al_u3583_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u3584 (
    .a(_al_u678_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 ),
    .o(_al_u3584_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(~C*~B*~A))"),
    .INIT(16'h00fe))
    _al_u3585 (
    .a(_al_u3582_o),
    .b(_al_u3583_o),
    .c(_al_u3584_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vygax6 ),
    .o(_al_u3585_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3586 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pthiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 ),
    .o(_al_u3586_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*(~(B)*~(C)*~(D)+B*~(C)*~(D)+~(B)*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'h5015))
    _al_u3587 (
    .a(_al_u3586_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 ),
    .o(_al_u3587_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(~B*~(A)*~(D)+~B*A*~(D)+~(~B)*A*D+~B*A*D))"),
    .INIT(16'h050c))
    _al_u3588 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 ),
    .o(_al_u3588_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(C*~(~D*B)))"),
    .INIT(16'h0545))
    _al_u3589 (
    .a(_al_u3585_o),
    .b(_al_u3587_o),
    .c(_al_u2868_o),
    .d(_al_u3588_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U0oiu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u359 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [6]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [7]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [8]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [9]),
    .o(_al_u359_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(~D*A))"),
    .INIT(16'h3f15))
    _al_u3590 (
    .a(_al_u1659_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ifoiu6_lutinv ),
    .c(_al_u932_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sdoiu6 ));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    _al_u3591 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 ),
    .o(_al_u3591_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(A*~(C*B)))"),
    .INIT(16'h00d5))
    _al_u3592 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sdoiu6 ),
    .b(_al_u3591_o),
    .c(_al_u1582_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ),
    .o(_al_u3592_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(~C*B*A))"),
    .INIT(16'h00f7))
    _al_u3593 (
    .a(_al_u3581_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U0oiu6 ),
    .c(_al_u3592_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ),
    .o(_al_u3593_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3594 (
    .a(_al_u3593_o),
    .b(_al_u1806_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Crniu6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3595 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Crniu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Utniu6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Umniu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*~B)*~(D*~A))"),
    .INIT(16'h8acf))
    _al_u3596 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yoniu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mpniu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6kax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vmipw6 ),
    .o(_al_u3596_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*~C))"),
    .INIT(16'h8088))
    _al_u3597 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Umniu6 ),
    .b(_al_u3596_o),
    .c(_al_u3120_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rkkax6 ),
    .o(_al_u3597_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3598 (
    .a(_al_u3132_o),
    .b(_al_u3593_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qkniu6_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3599 (
    .a(_al_u3597_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qkniu6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dhniu6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u360 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [2]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [4]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [5]),
    .o(_al_u360_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*~B)*~(D*~A))"),
    .INIT(16'h8acf))
    _al_u3600 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yoniu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mpniu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dzvpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Htmpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Inniu6 ));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*~C))"),
    .INIT(16'h8088))
    _al_u3601 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Umniu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Inniu6 ),
    .c(_al_u3120_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oikax6 ),
    .o(_al_u3601_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(C*~A))"),
    .INIT(16'h8caf))
    _al_u3602 (
    .a(_al_u3120_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mpniu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iekax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Shopw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aqniu6 ));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*~C))"),
    .INIT(16'h8088))
    _al_u3603 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Crniu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aqniu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yoniu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vhspw6 ),
    .o(_al_u3603_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3604 (
    .a(_al_u3601_o),
    .b(_al_u3603_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ckniu6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3605 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dhniu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ckniu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Etmiu6 ));
  AL_MAP_LUT2 #(
    .EQN("~(B@A)"),
    .INIT(4'h9))
    _al_u3606 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C53iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Utqpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fuxhu6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3607 (
    .a(_al_u3211_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yv1ju6 ));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*B*A)"),
    .INIT(16'h0800))
    _al_u3608 (
    .a(_al_u2835_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Htyiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rwjax6 ),
    .o(_al_u3608_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(~D*C*B))"),
    .INIT(16'haa2a))
    _al_u3609 (
    .a(_al_u3608_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N4kax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4jax6 ),
    .o(_al_u3609_o));
  AL_MAP_LUT4 #(
    .EQN("~(D*C*B*A)"),
    .INIT(16'h7fff))
    _al_u361 (
    .a(_al_u357_o),
    .b(_al_u358_o),
    .c(_al_u359_o),
    .d(_al_u360_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n304 ));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u3610 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yv1ju6 ),
    .b(_al_u3609_o),
    .c(_al_u2365_o),
    .o(_al_u3610_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*A)"),
    .INIT(16'h0002))
    _al_u3611 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pu1ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Daiax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ),
    .o(_al_u3611_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(~B*~(~D*A)))"),
    .INIT(16'hc0e0))
    _al_u3612 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qe8iu6_lutinv ),
    .b(_al_u3611_o),
    .c(_al_u1582_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ),
    .o(_al_u3612_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*A*~(~D*B))"),
    .INIT(16'h0a02))
    _al_u3613 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ez1ju6 ),
    .b(_al_u3185_o),
    .c(_al_u3612_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 ),
    .o(_al_u3613_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D*C*A))"),
    .INIT(16'h1333))
    _al_u3614 (
    .a(_al_u3110_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ),
    .c(_al_u2829_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 ),
    .o(_al_u3614_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*~(D*B))"),
    .INIT(16'h1050))
    _al_u3615 (
    .a(_al_u3157_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U98iu6 ),
    .c(_al_u3614_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vxniu6_lutinv ),
    .o(_al_u3615_o));
  AL_MAP_LUT4 #(
    .EQN("(A*(B@(~D*C)))"),
    .INIT(16'h8828))
    _al_u3616 (
    .a(_al_u3215_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N4kax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4jax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ro1ju6 ));
  AL_MAP_LUT4 #(
    .EQN("(C*B*~(D*A))"),
    .INIT(16'h40c0))
    _al_u3617 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yo1ju6 ),
    .b(_al_u3613_o),
    .c(_al_u3615_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ro1ju6 ),
    .o(_al_u3617_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3618 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Apaiu6_lutinv ),
    .b(_al_u607_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 ),
    .o(_al_u3618_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(~A*~(C*B)))"),
    .INIT(16'h00ea))
    _al_u3619 (
    .a(_al_u3618_o),
    .b(_al_u681_o),
    .c(_al_u2829_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jr1ju6_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("~(B*~A)"),
    .INIT(4'hb))
    _al_u362 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n3685 ));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u3620 (
    .a(_al_u3610_o),
    .b(_al_u3617_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jr1ju6_lutinv ),
    .d(_al_u1342_o),
    .o(_al_u3620_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u3621 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xq3pw6_lutinv ),
    .b(_al_u3109_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ),
    .o(_al_u3621_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    _al_u3622 (
    .a(_al_u3621_o),
    .b(_al_u3110_o),
    .c(_al_u607_o),
    .o(_al_u3622_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*C)*~(~B*A))"),
    .INIT(16'hdd0d))
    _al_u3623 (
    .a(_al_u3620_o),
    .b(_al_u3622_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fpnpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iuohu6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3624 (
    .a(_al_u909_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ),
    .o(_al_u3624_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u3625 (
    .a(_al_u2364_o),
    .b(_al_u930_o),
    .c(_al_u2764_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yljiu6 ),
    .o(_al_u3625_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(~D*C))"),
    .INIT(16'h4404))
    _al_u3626 (
    .a(_al_u3624_o),
    .b(_al_u3625_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J9kiu6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Skjax6 ),
    .o(_al_u3626_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(~D*~(~C*~B)))"),
    .INIT(16'haa02))
    _al_u3627 (
    .a(_al_u3626_o),
    .b(_al_u3110_o),
    .c(_al_u903_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 ),
    .o(_al_u3627_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~A*~(D*C))"),
    .INIT(16'h0111))
    _al_u3628 (
    .a(_al_u2758_o),
    .b(_al_u1583_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hgrpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 ),
    .o(_al_u3628_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3629 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D6kiu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ),
    .o(_al_u3629_o));
  AL_MAP_LUT2 #(
    .EQN("~(B*~A)"),
    .INIT(4'hb))
    _al_u363 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U8jax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qqhiu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u3630 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y0jiu6 ),
    .b(_al_u3629_o),
    .c(_al_u1266_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D31ju6 ),
    .o(_al_u3630_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u3631 (
    .a(_al_u3627_o),
    .b(_al_u3189_o),
    .c(_al_u3628_o),
    .d(_al_u3630_o),
    .o(_al_u3631_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3632 (
    .a(_al_u606_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yljiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 ),
    .o(_al_u3632_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u3633 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bziiu6_lutinv ),
    .b(_al_u3632_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 ),
    .o(_al_u3633_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3634 (
    .a(_al_u696_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S2ziu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 ),
    .o(_al_u3634_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*A*~(D*B))"),
    .INIT(16'h020a))
    _al_u3635 (
    .a(_al_u3633_o),
    .b(_al_u1812_o),
    .c(_al_u3634_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 ),
    .o(_al_u3635_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*~C))"),
    .INIT(16'h8088))
    _al_u3636 (
    .a(_al_u3631_o),
    .b(_al_u3635_o),
    .c(_al_u1643_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N3ziu6 ),
    .o(_al_u3636_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    _al_u3637 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F6ziu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wh0ju6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jgxpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4jax6 ),
    .o(_al_u3637_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(~D*~C*B))"),
    .INIT(16'h5551))
    _al_u3638 (
    .a(_al_u3637_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qxoiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 ),
    .o(_al_u3638_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*B*~A)"),
    .INIT(16'h0400))
    _al_u3639 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jckax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N4kax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P14qw6 ),
    .o(_al_u3639_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~((~C*~B))*~(D)+A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D)"),
    .INIT(16'h03fe))
    _al_u364 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_state [0]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_state [1]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_state [2]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_state [3]),
    .o(_al_u364_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(~D*~C))"),
    .INIT(16'h4440))
    _al_u3640 (
    .a(_al_u3638_o),
    .b(_al_u3639_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4jax6 ),
    .o(_al_u3640_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~C)*~(~B*A))"),
    .INIT(16'hd0dd))
    _al_u3641 (
    .a(_al_u1342_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 ),
    .o(_al_u3641_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~A*~(D*~B))"),
    .INIT(16'h0405))
    _al_u3642 (
    .a(_al_u1802_o),
    .b(_al_u3641_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vygax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T41ju6 ));
  AL_MAP_LUT4 #(
    .EQN("(C*A*~(D*~B))"),
    .INIT(16'h80a0))
    _al_u3643 (
    .a(_al_u3636_o),
    .b(_al_u3640_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T41ju6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J9kiu6_lutinv ),
    .o(_al_u3643_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u3644 (
    .a(_al_u3109_o),
    .b(_al_u903_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I30ju6_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3645 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nsaiu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wxyiu6 ));
  AL_MAP_LUT4 #(
    .EQN("(A*~(~D*~C*B))"),
    .INIT(16'haaa2))
    _al_u3646 (
    .a(_al_u3643_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I30ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wxyiu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 ),
    .o(_al_u3646_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u3647 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nbkiu6_lutinv ),
    .b(_al_u2364_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qxoiu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 ),
    .o(_al_u3647_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D*~C*B))"),
    .INIT(16'ha2aa))
    _al_u3648 (
    .a(_al_u3647_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 ),
    .o(_al_u3648_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u3649 (
    .a(_al_u3648_o),
    .b(_al_u912_o),
    .c(_al_u3215_o),
    .o(_al_u3649_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u365 (
    .a(_al_u364_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n102 [2]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_rx_state [2]));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u3650 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N4kax6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rwjax6 ),
    .o(_al_u3650_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D*~(~C*~A)))"),
    .INIT(16'h0133))
    _al_u3651 (
    .a(_al_u2380_o),
    .b(_al_u3650_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qz0ju6 ));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*A)"),
    .INIT(16'h0002))
    _al_u3652 (
    .a(_al_u3215_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N4kax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4jax6 ),
    .o(_al_u3652_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(A*~(C)*~(D)+~(A)*C*D))"),
    .INIT(16'h4008))
    _al_u3653 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N4kax6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rwjax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4jax6 ),
    .o(_al_u3653_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(~D*~B*A))"),
    .INIT(16'hf0d0))
    _al_u3654 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qz0ju6 ),
    .b(_al_u3652_o),
    .c(_al_u2364_o),
    .d(_al_u3653_o),
    .o(_al_u3654_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D*~(~C*B)))"),
    .INIT(16'h08aa))
    _al_u3655 (
    .a(_al_u3646_o),
    .b(_al_u3649_o),
    .c(_al_u3654_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 ),
    .o(_al_u3655_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3656 (
    .a(_al_u1346_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Daiax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z37ow6_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3657 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z37ow6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 ),
    .o(_al_u3657_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(~B*~(C*A)))"),
    .INIT(16'h00ec))
    _al_u3658 (
    .a(_al_u607_o),
    .b(_al_u2813_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 ),
    .o(_al_u3658_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~B*~(~D*A))"),
    .INIT(16'h0301))
    _al_u3659 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I30ju6_lutinv ),
    .b(_al_u3657_o),
    .c(_al_u3658_o),
    .d(_al_u3094_o),
    .o(_al_u3659_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u366 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T24iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M8ipw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F24iu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h7705))
    _al_u3660 (
    .a(_al_u3655_o),
    .b(_al_u3659_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Twohu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*~A)"),
    .INIT(16'h0004))
    _al_u3661 (
    .a(_al_u1643_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K49ow6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 ),
    .o(_al_u3661_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(D*~C*B))"),
    .INIT(16'h5155))
    _al_u3662 (
    .a(_al_u2365_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 ),
    .o(_al_u3662_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(D*~C*B))"),
    .INIT(16'h5155))
    _al_u3663 (
    .a(_al_u3661_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W0piu6_lutinv ),
    .c(_al_u3662_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 ),
    .o(_al_u3663_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u3664 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ujjiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R9aiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wkipw6 ),
    .o(_al_u3664_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*A*~(~D*C))"),
    .INIT(16'h2202))
    _al_u3665 (
    .a(_al_u3663_o),
    .b(_al_u3664_o),
    .c(_al_u2847_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wxyiu6 ),
    .o(_al_u3665_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3666 (
    .a(_al_u3629_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yecpw6_lutinv ),
    .o(_al_u3666_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3667 (
    .a(_al_u3236_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 ),
    .o(_al_u3667_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(~C*A))"),
    .INIT(16'hf531))
    _al_u3668 (
    .a(_al_u3666_o),
    .b(_al_u3667_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U99ow6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(~D*A))"),
    .INIT(16'h3f15))
    _al_u3669 (
    .a(_al_u3187_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T23ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K49ow6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 ),
    .o(_al_u3669_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u367 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S2cbx6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Stkpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wt3qw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zwnpw6 ),
    .o(_al_u367_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*A*~(~D*C))"),
    .INIT(16'h2202))
    _al_u3670 (
    .a(_al_u909_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ),
    .o(_al_u3670_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u3671 (
    .a(_al_u1813_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hwaiu6_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u3672 (
    .a(_al_u3670_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hwaiu6_lutinv ),
    .c(_al_u1662_o),
    .o(_al_u3672_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u3673 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T41ju6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U99ow6 ),
    .c(_al_u3669_o),
    .d(_al_u3672_o),
    .o(_al_u3673_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*~B*A)"),
    .INIT(16'h0020))
    _al_u3674 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D31ju6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 ),
    .o(_al_u3674_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(~C*~(D*B)))"),
    .INIT(16'ha8a0))
    _al_u3675 (
    .a(_al_u3109_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N3ziu6 ),
    .c(_al_u3674_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jf6ju6 ),
    .o(_al_u3675_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(A*~(C*~B)))"),
    .INIT(16'h7500))
    _al_u3676 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P14qw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kb9ow6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(A*~(~B*~(~D*C)))"),
    .INIT(16'h88a8))
    _al_u3677 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uyiiu6 ),
    .b(_al_u2772_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kb9ow6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9ypw6 ),
    .o(_al_u3677_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    _al_u3678 (
    .a(_al_u3665_o),
    .b(_al_u3673_o),
    .c(_al_u3675_o),
    .d(_al_u3677_o),
    .o(_al_u3678_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(~D*~C))"),
    .INIT(16'h8880))
    _al_u3679 (
    .a(_al_u3214_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jckax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jgxpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4jax6 ),
    .o(_al_u3679_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u368 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C72qw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J4cbx6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kn2qw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nfqpw6 ),
    .o(_al_u368_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3680 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujiu6 ),
    .b(_al_u2369_o),
    .o(_al_u3680_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*(~(A)*C*~(D)+A*C*~(D)+~(A)*~(C)*D+A*~(C)*D+A*C*D))"),
    .INIT(16'h2330))
    _al_u3681 (
    .a(_al_u3679_o),
    .b(_al_u3680_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9ypw6 ),
    .o(_al_u3681_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u3682 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Skjax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y40ju6 ));
  AL_MAP_LUT4 #(
    .EQN("(~B*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))"),
    .INIT(16'h2203))
    _al_u3683 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N4kax6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4jax6 ),
    .o(_al_u3683_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(A*~(~D*C)))"),
    .INIT(16'h44c4))
    _al_u3684 (
    .a(_al_u3681_o),
    .b(_al_u2770_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y40ju6 ),
    .d(_al_u3683_o),
    .o(_al_u3684_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+A*B*C*D)"),
    .INIT(16'h8dfb))
    _al_u3685 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N4kax6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rwjax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4jax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wh9ow6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(A*~(~B*~(~D*C)))"),
    .INIT(16'h88a8))
    _al_u3686 (
    .a(_al_u2386_o),
    .b(_al_u2764_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wh9ow6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9ypw6 ),
    .o(_al_u3686_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(~C*~B*A))"),
    .INIT(16'h00fd))
    _al_u3687 (
    .a(_al_u2767_o),
    .b(_al_u2369_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hgrpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Io9ow6 ));
  AL_MAP_LUT4 #(
    .EQN("(D*~(A*~(~C*B)))"),
    .INIT(16'h5d00))
    _al_u3688 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Io9ow6 ),
    .b(_al_u1367_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 ),
    .o(_al_u3688_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3689 (
    .a(_al_u2371_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fm6ow6_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u369 (
    .a(_al_u367_o),
    .b(_al_u368_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I13iu6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3690 (
    .a(_al_u1344_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ),
    .o(_al_u3690_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*C)*~(B*A))"),
    .INIT(16'h0777))
    _al_u3691 (
    .a(_al_u912_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fm6ow6_lutinv ),
    .c(_al_u3690_o),
    .d(_al_u696_o),
    .o(_al_u3691_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*~A)"),
    .INIT(16'h0100))
    _al_u3692 (
    .a(_al_u3684_o),
    .b(_al_u3686_o),
    .c(_al_u3688_o),
    .d(_al_u3691_o),
    .o(_al_u3692_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0cf5))
    _al_u3693 (
    .a(_al_u1643_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 ),
    .o(_al_u3693_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(~B*~(D*~A)))"),
    .INIT(16'hd0c0))
    _al_u3694 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eoyiu6_lutinv ),
    .b(_al_u3693_o),
    .c(_al_u1806_o),
    .d(_al_u1266_o),
    .o(_al_u3694_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*A*~(~D*~B))"),
    .INIT(16'h0a08))
    _al_u3695 (
    .a(_al_u3678_o),
    .b(_al_u3692_o),
    .c(_al_u3694_o),
    .d(_al_u1812_o),
    .o(_al_u3695_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D*C*~A))"),
    .INIT(16'h2333))
    _al_u3696 (
    .a(_al_u3109_o),
    .b(_al_u696_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yljiu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 ),
    .o(_al_u3696_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~A*~(~C*~B))"),
    .INIT(16'h5400))
    _al_u3697 (
    .a(_al_u3696_o),
    .b(_al_u607_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Difiu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ),
    .o(_al_u3697_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*C)*~(~B*A))"),
    .INIT(16'hdd0d))
    _al_u3698 (
    .a(_al_u3695_o),
    .b(_al_u3697_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jrohu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u3699 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bggiu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yogiu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xozax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z9abx6 ),
    .o(_al_u3699_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u370 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_state [2]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_state [3]),
    .o(_al_u370_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u3700 (
    .a(_al_u3271_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Webiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aw4bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uizax6 ),
    .o(_al_u3700_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u3701 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nbdiu6_lutinv ),
    .b(_al_u3446_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lfgbx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M85bx6 ),
    .o(_al_u3701_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u3702 (
    .a(_al_u3454_o),
    .b(_al_u3463_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J6zax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nhgbx6 ),
    .o(_al_u3702_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u3703 (
    .a(_al_u3699_o),
    .b(_al_u3700_o),
    .c(_al_u3701_o),
    .d(_al_u3702_o),
    .o(_al_u3703_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u3704 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Etfiu6_lutinv ),
    .b(_al_u3520_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E34bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hbgbx6 ),
    .o(_al_u3704_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u3705 (
    .a(_al_u3703_o),
    .b(_al_u3704_o),
    .c(_al_u3530_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Up4bx6 ),
    .o(_al_u3705_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u3706 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Odfiu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ivfiu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bcabx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jdgbx6 ),
    .o(_al_u3706_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u3707 (
    .a(_al_u3281_o),
    .b(_al_u3479_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ohyax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vbspw6 ),
    .o(_al_u3707_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u3708 (
    .a(_al_u3372_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3giu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cwyax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pjgbx6 ),
    .o(_al_u3708_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u3709 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eegiu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lhdiu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K94bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T3abx6 ),
    .o(_al_u3709_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*A)"),
    .INIT(16'h0080))
    _al_u371 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_state_inc ),
    .b(_al_u370_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_state [0]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_state [1]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rxbuf_sample ));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u3710 (
    .a(_al_u3706_o),
    .b(_al_u3707_o),
    .c(_al_u3708_o),
    .d(_al_u3709_o),
    .o(_al_u3710_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u3711 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dagiu6_lutinv ),
    .b(_al_u3443_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qf4bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X7abx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Isbpw6 ));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u3712 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F8row6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[2] ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[3] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qrgiu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u3713 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rhgiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qrgiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tl4bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vpgbx6 ),
    .o(_al_u3713_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u3714 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jzfiu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mxfiu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R1abx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yw3bx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A2cpw6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u3715 (
    .a(_al_u3468_o),
    .b(_al_u3350_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G25bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pczax6 ),
    .o(_al_u3715_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u3716 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Isbpw6 ),
    .b(_al_u3713_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A2cpw6 ),
    .d(_al_u3715_o),
    .o(_al_u3716_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u3717 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ajgiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hwhiu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V5abx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wgipw6 ),
    .o(_al_u3717_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u3718 (
    .a(_al_u3335_o),
    .b(_al_u3343_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C5gbx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nv9bx6 ),
    .o(_al_u3718_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u3719 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G9fiu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hcgiu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rlgbx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tngbx6 ),
    .o(_al_u3719_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(D*C*~B))"),
    .INIT(16'h4555))
    _al_u372 (
    .a(XTAL1_wire),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bciax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cokbx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I2zax6 ),
    .o(XTAL2_pad));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u3720 (
    .a(_al_u3489_o),
    .b(_al_u3515_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pz9bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Unyax6 ),
    .o(_al_u3720_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u3721 (
    .a(_al_u3717_o),
    .b(_al_u3718_o),
    .c(_al_u3719_o),
    .d(_al_u3720_o),
    .o(_al_u3721_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u3722 (
    .a(_al_u3705_o),
    .b(_al_u3710_o),
    .c(_al_u3716_o),
    .d(_al_u3721_o),
    .o(_al_u3722_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3723 (
    .a(_al_u3722_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tl4bx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vwapw6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u3724 (
    .a(_al_u3343_o),
    .b(_al_u3350_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I45bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vkzax6 ),
    .o(_al_u3724_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u3725 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hwhiu6_lutinv ),
    .b(_al_u3446_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H4zax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oa5bx6 ),
    .o(_al_u3725_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u3726 (
    .a(_al_u3463_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nbdiu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nazax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Slyax6 ),
    .o(_al_u3726_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u3727 (
    .a(_al_u3443_o),
    .b(_al_u3520_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E05bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yt4bx6 ),
    .o(_al_u3727_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u3728 (
    .a(_al_u3724_o),
    .b(_al_u3725_o),
    .c(_al_u3726_o),
    .d(_al_u3727_o),
    .o(_al_u3728_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u3729 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ivfiu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Webiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C14bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cy4bx6 ),
    .o(_al_u3729_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(D*C*~A))"),
    .INIT(16'h8ccc))
    _al_u373 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cjqpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Okfax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qwfax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Utqpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qq3iu6 ));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u3730 (
    .a(_al_u3728_o),
    .b(_al_u3729_o),
    .c(_al_u3530_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wr4bx6 ),
    .o(_al_u3730_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u3731 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bggiu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Etfiu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G54bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I74bx6 ),
    .o(_al_u3731_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u3732 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dagiu6_lutinv ),
    .b(_al_u3468_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rezax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sh4bx6 ),
    .o(_al_u3732_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u3733 (
    .a(_al_u3271_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qrgiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgzax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uj4bx6 ),
    .o(_al_u3733_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u3734 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Odfiu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lhdiu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mfyax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S3mpw6 ),
    .o(_al_u3734_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u3735 (
    .a(_al_u3731_o),
    .b(_al_u3732_o),
    .c(_al_u3733_o),
    .d(_al_u3734_o),
    .o(_al_u3735_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u3736 (
    .a(_al_u3335_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ajgiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Elnpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yqzax6 ),
    .o(_al_u3736_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u3737 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eegiu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hcgiu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mb4bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Od4bx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H3bpw6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u3738 (
    .a(_al_u3489_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mxfiu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Az3bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wpyax6 ),
    .o(_al_u3738_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u3739 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rhgiu6 ),
    .b(_al_u3479_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gz6ax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qjyax6 ),
    .o(_al_u3739_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u374 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D43qw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pe7ax6 ),
    .o(_al_u374_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u3740 (
    .a(_al_u3736_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H3bpw6 ),
    .c(_al_u3738_o),
    .d(_al_u3739_o),
    .o(_al_u3740_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u3741 (
    .a(_al_u3372_o),
    .b(_al_u3454_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eyyax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L8zax6 ),
    .o(_al_u3741_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u3742 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G9fiu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3giu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Auyax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K65bx6 ),
    .o(_al_u3742_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u3743 (
    .a(_al_u3281_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yogiu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wmzax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yryax6 ),
    .o(_al_u3743_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u3744 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jzfiu6_lutinv ),
    .b(_al_u3515_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sn4bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wu3bx6 ),
    .o(_al_u3744_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u3745 (
    .a(_al_u3741_o),
    .b(_al_u3742_o),
    .c(_al_u3743_o),
    .d(_al_u3744_o),
    .o(_al_u3745_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u3746 (
    .a(_al_u3730_o),
    .b(_al_u3735_o),
    .c(_al_u3740_o),
    .d(_al_u3745_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sbrow6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3747 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qrgiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rmbpw6 ),
    .o(_al_u3747_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3748 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ejbpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[1] ),
    .o(_al_u3748_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u3749 (
    .a(_al_u3747_o),
    .b(_al_u3748_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uybpw6_lutinv ),
    .o(_al_u3749_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u375 (
    .a(_al_u374_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Di3qw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Le2qw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vowiu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~C*(~(A)*B*~(D)+~(A)*~(B)*D+~(A)*B*D+A*B*D))"),
    .INIT(16'h0d04))
    _al_u3750 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vwapw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sbrow6 ),
    .c(_al_u3749_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uj4bx6 ),
    .o(_al_u3750_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u3751 (
    .a(_al_u3750_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B0biu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_primask_o ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0biu6 ));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3752 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zwcpw6_lutinv ),
    .b(_al_u607_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Utgiu6 ));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u3753 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Utgiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 ),
    .o(_al_u3753_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3754 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yljiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pthiu6 ),
    .o(_al_u3754_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(~B*~(D*C)))"),
    .INIT(16'ha888))
    _al_u3755 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0biu6 ),
    .b(_al_u3753_o),
    .c(_al_u3754_o),
    .d(_al_u3124_o),
    .o(_al_u3755_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u3756 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K5eiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R9yax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W5ypw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztupw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xrgiu6 ));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u3757 (
    .a(_al_u3755_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fsdiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xrgiu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qh5iu6 ));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B*A))"),
    .INIT(8'h70))
    _al_u3758 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xrgiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C1wpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F17ax6 ),
    .o(_al_u3758_o));
  AL_MAP_LUT4 #(
    .EQN("~(A*~(D*~(C*B)))"),
    .INIT(16'h7f55))
    _al_u3759 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qh5iu6 ),
    .b(_al_u1777_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qrgiu6 ),
    .d(_al_u3758_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rjthu6 ));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*A)"),
    .INIT(16'h0200))
    _al_u376 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vowiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hw8ax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sqwpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zm8ax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ve7iu6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3760 (
    .a(_al_u3597_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qkniu6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Miniu6_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3761 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ckniu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Miniu6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztmiu6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3762 (
    .a(_al_u3601_o),
    .b(_al_u3603_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Finiu6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3763 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Miniu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Finiu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jsmiu6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3764 (
    .a(_al_u3597_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qkniu6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vjniu6_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3765 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Finiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vjniu6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qsmiu6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3766 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ckniu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vjniu6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gumiu6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u3767 (
    .a(_al_u3597_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qkniu6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rhniu6_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3768 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ckniu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rhniu6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ltmiu6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3769 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Finiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rhniu6_lutinv ),
    .o(_al_u3769_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u377 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ve7iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dg2qw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oe7iu6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3770 (
    .a(_al_u3769_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jrypw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydkiu6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u3771 (
    .a(_al_u3601_o),
    .b(_al_u3603_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Khniu6_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3772 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vjniu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Khniu6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xsmiu6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3773 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rhniu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Khniu6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Csmiu6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3774 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tezhu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vplpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Di1iu6 ));
  AL_MAP_LUT4 #(
    .EQN("(D*~(~B*~(C*A)))"),
    .INIT(16'hec00))
    _al_u3775 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Di1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B7lpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L5lpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ryfax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fwohu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*~A)"),
    .INIT(16'h0040))
    _al_u3776 (
    .a(_al_u3255_o),
    .b(_al_u1757_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Krlpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yklpw6 ),
    .o(_al_u3776_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u3777 (
    .a(_al_u1253_o),
    .b(_al_u1676_o),
    .c(\u_cmsdk_mcu/dbg_swdo_en ),
    .o(_al_u3777_o));
  AL_MAP_LUT4 #(
    .EQN("~(B*~(D*~(C*~A)))"),
    .INIT(16'hbf33))
    _al_u3778 (
    .a(_al_u3776_o),
    .b(_al_u3777_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I6yhu6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U5yhu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I5nhu6 ));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*B*A)"),
    .INIT(16'h0800))
    _al_u3779 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K5eiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R9yax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W5ypw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztupw6 ),
    .o(_al_u3779_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u378 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rxbuf_sample ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_ctrl [3]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/intr_stat_set [1]));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*B*~A)"),
    .INIT(16'h0400))
    _al_u3780 (
    .a(\u_cmsdk_mcu/HWDATA [30]),
    .b(\u_cmsdk_mcu/HWDATA [17]),
    .c(\u_cmsdk_mcu/HWDATA [16]),
    .d(_al_u3779_o),
    .o(_al_u3780_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u3781 (
    .a(_al_u3780_o),
    .b(\u_cmsdk_mcu/HWDATA [31]),
    .c(_al_u2725_o),
    .o(_al_u3781_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3782 (
    .a(_al_u2729_o),
    .b(_al_u2733_o),
    .c(_al_u2741_o),
    .o(_al_u3782_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*B*A)"),
    .INIT(16'h0800))
    _al_u3783 (
    .a(\u_cmsdk_mcu/HWDATA [22]),
    .b(\u_cmsdk_mcu/HWDATA [23]),
    .c(_al_u2717_o),
    .d(_al_u2721_o),
    .o(_al_u3783_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*~A)"),
    .INIT(16'h4000))
    _al_u3784 (
    .a(\u_cmsdk_mcu/HWDATA [18]),
    .b(\u_cmsdk_mcu/HWDATA [19]),
    .c(\u_cmsdk_mcu/HWDATA [20]),
    .d(\u_cmsdk_mcu/HWDATA [21]),
    .o(_al_u3784_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u3785 (
    .a(_al_u3781_o),
    .b(_al_u3782_o),
    .c(_al_u3783_o),
    .d(_al_u3784_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T9qow6 ));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(B*A))"),
    .INIT(8'hf8))
    _al_u3786 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T9qow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G3eiu6 ),
    .c(\u_cmsdk_mcu/SYSRESETREQ ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yaohu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(D*C*B))"),
    .INIT(16'h1555))
    _al_u3787 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G1aow6 ),
    .b(_al_u607_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vo3ju6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 ),
    .o(_al_u3787_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B*~A))"),
    .INIT(8'hb0))
    _al_u3788 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I82ju6 ),
    .b(_al_u3787_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 ),
    .o(_al_u3788_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u3789 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qe8iu6_lutinv ),
    .b(_al_u3156_o),
    .c(_al_u2392_o),
    .o(_al_u3789_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u379 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_state [2]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_state [3]),
    .o(_al_u379_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u3790 (
    .a(_al_u3789_o),
    .b(_al_u1297_o),
    .c(_al_u606_o),
    .o(_al_u3790_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~A*~(D*C))"),
    .INIT(16'h0111))
    _al_u3791 (
    .a(_al_u697_o),
    .b(_al_u3159_o),
    .c(_al_u609_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ),
    .o(_al_u3791_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u3792 (
    .a(_al_u1269_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yljiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ),
    .o(_al_u3792_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u3793 (
    .a(_al_u696_o),
    .b(_al_u2392_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mbhow6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ),
    .o(_al_u3793_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u3794 (
    .a(_al_u3624_o),
    .b(_al_u3793_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 ),
    .o(_al_u3794_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*~A)"),
    .INIT(16'h0040))
    _al_u3795 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv ),
    .b(_al_u1266_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 ),
    .o(_al_u3795_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*~B*A)"),
    .INIT(16'h0020))
    _al_u3796 (
    .a(_al_u3791_o),
    .b(_al_u3792_o),
    .c(_al_u3794_o),
    .d(_al_u3795_o),
    .o(_al_u3796_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u3797 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rcziu6 ),
    .b(_al_u3788_o),
    .c(_al_u3790_o),
    .d(_al_u3796_o),
    .o(_al_u3797_o));
  AL_MAP_LUT4 #(
    .EQN("~(A*~((D*B))*~(C)+A*(D*B)*~(C)+~(A)*(D*B)*C+A*(D*B)*C)"),
    .INIT(16'h35f5))
    _al_u3798 (
    .a(_al_u682_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 ),
    .o(_al_u3798_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf53f))
    _al_u3799 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Edapw6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 ),
    .o(_al_u3799_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*B*A)"),
    .INIT(16'h0800))
    _al_u380 (
    .a(_al_u379_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_state [0]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_state [1]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/BAUDTICK ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n53 ));
  AL_MAP_LUT4 #(
    .EQN("(A*~(~B*~(D*C)))"),
    .INIT(16'ha888))
    _al_u3800 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 ),
    .o(_al_u3800_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*~A)"),
    .INIT(16'h0100))
    _al_u3801 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jf6ju6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pthiu6 ),
    .c(_al_u3800_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 ),
    .o(_al_u3801_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(D*C*B))"),
    .INIT(16'h1555))
    _al_u3802 (
    .a(_al_u3797_o),
    .b(_al_u3798_o),
    .c(_al_u3799_o),
    .d(_al_u3801_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A3iiu6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3803 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ly2ju6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Np7ow6_lutinv ),
    .o(_al_u3803_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3804 (
    .a(_al_u604_o),
    .b(_al_u2813_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ),
    .o(_al_u3804_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~A*~(D*B))"),
    .INIT(16'h0105))
    _al_u3805 (
    .a(_al_u3803_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vxniu6_lutinv ),
    .c(_al_u3804_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ),
    .o(_al_u3805_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*C)*~(B*A))"),
    .INIT(16'h0777))
    _al_u3806 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Btoiu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vo3ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Owoiu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 ),
    .o(_al_u3806_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*A)"),
    .INIT(16'h0002))
    _al_u3807 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ),
    .o(_al_u3807_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(~D*C*B))"),
    .INIT(16'h5515))
    _al_u3808 (
    .a(_al_u3797_o),
    .b(_al_u3805_o),
    .c(_al_u3806_o),
    .d(_al_u3807_o),
    .o(_al_u3808_o));
  AL_MAP_LUT4 #(
    .EQN("~(~(C*B)*~(D*A))"),
    .INIT(16'heac0))
    _al_u3809 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A3iiu6 ),
    .b(_al_u3808_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Go0iu6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [1]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ay8iu6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u381 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n53 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n55 [3]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_tx_tick_cnt [3]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3810 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U98iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 ),
    .o(_al_u3810_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3811 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M8fax6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wkipw6 ),
    .o(_al_u3811_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u3812 (
    .a(_al_u1812_o),
    .b(_al_u2380_o),
    .c(_al_u3811_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9ypw6 ),
    .o(_al_u3812_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*~B)*~(D*A))"),
    .INIT(16'h45cf))
    _al_u3813 (
    .a(_al_u3810_o),
    .b(_al_u3812_o),
    .c(_al_u903_o),
    .d(_al_u1342_o),
    .o(_al_u3813_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u3814 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Llaow6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vygax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 ),
    .o(_al_u3814_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u3815 (
    .a(_al_u3814_o),
    .b(_al_u1782_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 ),
    .o(_al_u3815_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~B*~(C*A))"),
    .INIT(16'h0013))
    _al_u3816 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qe8iu6_lutinv ),
    .b(_al_u1783_o),
    .c(_al_u2849_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ),
    .o(_al_u3816_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u3817 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9ypw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 ),
    .o(_al_u3817_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u3818 (
    .a(_al_u3815_o),
    .b(_al_u3816_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kxziu6_lutinv ),
    .d(_al_u3817_o),
    .o(_al_u3818_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(~D*C))"),
    .INIT(16'h8808))
    _al_u3819 (
    .a(_al_u903_o),
    .b(_al_u2392_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vygax6 ),
    .o(_al_u3819_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u382 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n53 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n55 [2]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_tx_tick_cnt [2]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(~D*~C*A))"),
    .INIT(16'h3331))
    _al_u3820 (
    .a(_al_u3629_o),
    .b(_al_u3819_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Np7ow6_lutinv ),
    .d(_al_u3150_o),
    .o(_al_u3820_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(D*~C*A))"),
    .INIT(16'hc4cc))
    _al_u3821 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U98iu6 ),
    .b(_al_u3820_o),
    .c(_al_u1266_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Btoiu6_lutinv ),
    .o(_al_u3821_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*~(D*~A))"),
    .INIT(16'h80c0))
    _al_u3822 (
    .a(_al_u3813_o),
    .b(_al_u3818_o),
    .c(_al_u3821_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 ),
    .o(_al_u3822_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D*C*B))"),
    .INIT(16'h2aaa))
    _al_u3823 (
    .a(_al_u3822_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eoyiu6_lutinv ),
    .c(_al_u2754_o),
    .d(_al_u1266_o),
    .o(_al_u3823_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3824 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I30ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 ),
    .o(_al_u3824_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u3825 (
    .a(_al_u3823_o),
    .b(_al_u3824_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qyniu6_lutinv ),
    .o(_al_u3825_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3826 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 ),
    .o(_al_u3826_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    _al_u3827 (
    .a(_al_u1643_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N3ziu6 ),
    .c(_al_u3826_o),
    .o(_al_u3827_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(B*~(~D*~C)))"),
    .INIT(16'h1115))
    _al_u3828 (
    .a(_al_u2772_o),
    .b(_al_u2364_o),
    .c(_al_u2764_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nyiiu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gc6ow6 ));
  AL_MAP_LUT4 #(
    .EQN("(~D*A*~(C*~B))"),
    .INIT(16'h008a))
    _al_u3829 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vo3ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D31ju6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 ),
    .o(_al_u3829_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u383 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n53 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n55 [1]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_tx_tick_cnt [1]));
  AL_MAP_LUT4 #(
    .EQN("(~C*A*~(D*B))"),
    .INIT(16'h020a))
    _al_u3830 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gc6ow6 ),
    .b(_al_u1799_o),
    .c(_al_u3829_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 ),
    .o(_al_u3830_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u3831 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rwjax6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 ),
    .o(_al_u3831_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(~C*A))"),
    .INIT(16'h31f5))
    _al_u3832 (
    .a(_al_u3754_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A95iu6_lutinv ),
    .c(_al_u1813_o),
    .d(_al_u3831_o),
    .o(_al_u3832_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3833 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wa0ju6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Skjax6 ),
    .o(_al_u3833_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*~A)"),
    .INIT(16'h0040))
    _al_u3834 (
    .a(_al_u3827_o),
    .b(_al_u3830_o),
    .c(_al_u3832_o),
    .d(_al_u3833_o),
    .o(_al_u3834_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(~A*~(D*B)))"),
    .INIT(16'h0e0a))
    _al_u3835 (
    .a(_al_u604_o),
    .b(_al_u2647_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 ),
    .o(_al_u3835_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D*C*B))"),
    .INIT(16'h2aaa))
    _al_u3836 (
    .a(_al_u3834_o),
    .b(_al_u3109_o),
    .c(_al_u3835_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Frziu6_lutinv ),
    .o(_al_u3836_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*~A)"),
    .INIT(16'h0004))
    _al_u3837 (
    .a(_al_u1643_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 ),
    .o(_al_u3837_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3838 (
    .a(_al_u3837_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 ),
    .o(_al_u3838_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+~(A)*B*~(C)+A*B*~(C)+~(A)*~(B)*C+~(A)*B*C)"),
    .INIT(8'h5e))
    _al_u3839 (
    .a(_al_u2767_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P14qw6 ),
    .o(_al_u3839_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u384 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n53 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n55 [0]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_tx_tick_cnt [0]));
  AL_MAP_LUT4 #(
    .EQN("(C*A*~(D*B))"),
    .INIT(16'h20a0))
    _al_u3840 (
    .a(_al_u3839_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qxoiu6 ),
    .c(_al_u2868_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Skjax6 ),
    .o(_al_u3840_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C@A))"),
    .INIT(8'h84))
    _al_u3841 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jckax6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N4kax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4jax6 ),
    .o(_al_u3841_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3842 (
    .a(_al_u3841_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rwjax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuyiu6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*~C))"),
    .INIT(16'h8088))
    _al_u3843 (
    .a(_al_u2361_o),
    .b(_al_u3840_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuyiu6_lutinv ),
    .d(_al_u2764_o),
    .o(_al_u3843_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(~D*~(C*B)))"),
    .INIT(16'h5540))
    _al_u3844 (
    .a(_al_u2369_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N4kax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 ),
    .o(_al_u3844_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(~A*~(~C*~B)))"),
    .INIT(16'h00ab))
    _al_u3845 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fm6ow6_lutinv ),
    .b(_al_u3844_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P14qw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9ypw6 ),
    .o(_al_u3845_o));
  AL_MAP_LUT4 #(
    .EQN("(C*(~(A)*~(B)*~(D)+A*~(B)*~(D)+~(A)*B*D))"),
    .INIT(16'h4030))
    _al_u3846 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N4kax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Skjax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4jax6 ),
    .o(_al_u3846_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(D*C*B))"),
    .INIT(16'h1555))
    _al_u3847 (
    .a(_al_u3846_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N4kax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P14qw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 ),
    .o(_al_u3847_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*A*~(D*~C))"),
    .INIT(16'h2022))
    _al_u3848 (
    .a(_al_u3843_o),
    .b(_al_u3845_o),
    .c(_al_u3847_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rwjax6 ),
    .o(_al_u3848_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(A*~(~C*~B)))"),
    .INIT(16'h0057))
    _al_u3849 (
    .a(_al_u3836_o),
    .b(_al_u3838_o),
    .c(_al_u3848_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv ),
    .o(_al_u3849_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u385 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_shift_in ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_ctrl [1]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n100 ));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*C)*~(~B*A))"),
    .INIT(16'hdd0d))
    _al_u3850 (
    .a(_al_u3825_o),
    .b(_al_u3849_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Utohu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~B*(A*~(C)*~(D)+~(A)*C*~(D)+A*C*~(D)+A*C*D))"),
    .INIT(16'h2032))
    _al_u3851 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zbjiu6 ),
    .b(_al_u2790_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ncjiu6_lutinv ),
    .d(_al_u3314_o),
    .o(_al_u3851_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3852 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R9mpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rskax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sqkax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jajiu6 ));
  AL_MAP_LUT3 #(
    .EQN("(~A*(C@B))"),
    .INIT(8'h14))
    _al_u3853 (
    .a(_al_u2783_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jajiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U1kpw6 ),
    .o(_al_u3853_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3854 (
    .a(_al_u2763_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9ypw6 ),
    .o(_al_u3854_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u3855 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv ),
    .b(_al_u1803_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 ),
    .o(_al_u3855_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*~(D*B))"),
    .INIT(16'h1050))
    _al_u3856 (
    .a(_al_u3854_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tc8iu6 ),
    .c(_al_u3855_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xiipw6 ),
    .o(_al_u3856_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(D*C))"),
    .INIT(16'h0444))
    _al_u3857 (
    .a(_al_u3853_o),
    .b(_al_u3856_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Habiu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Irmpw6 ),
    .o(_al_u3857_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(~A*~(~D*B)))"),
    .INIT(16'ha0e0))
    _al_u3858 (
    .a(_al_u2766_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M7kiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rwjax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 ),
    .o(_al_u3858_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*A*~(D*~C))"),
    .INIT(16'h2022))
    _al_u3859 (
    .a(_al_u3857_o),
    .b(_al_u3858_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yb8iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wkipw6 ),
    .o(_al_u3859_o));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    _al_u386 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_state_inc ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n100 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_state_update ));
  AL_MAP_LUT2 #(
    .EQN("~(B*~A)"),
    .INIT(4'hb))
    _al_u3860 (
    .a(_al_u3851_o),
    .b(_al_u3859_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y7jiu6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3861 (
    .a(_al_u3601_o),
    .b(_al_u3603_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jkniu6_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3862 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vjniu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jkniu6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Numiu6 ));
  AL_MAP_LUT2 #(
    .EQN("~(B*A)"),
    .INIT(4'h7))
    _al_u3863 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Miniu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jkniu6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ickiu6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3864 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rhniu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jkniu6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Stmiu6 ));
  AL_MAP_LUT2 #(
    .EQN("~(B*A)"),
    .INIT(4'h7))
    _al_u3865 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dhniu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jkniu6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hfkiu6 ));
  AL_MAP_LUT2 #(
    .EQN("~(~B*A)"),
    .INIT(4'hd))
    _al_u3866 (
    .a(_al_u3769_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jrypw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n1552 ));
  AL_MAP_LUT2 #(
    .EQN("~(B*A)"),
    .INIT(4'h7))
    _al_u3867 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Miniu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Khniu6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kdkiu6 ));
  AL_MAP_LUT2 #(
    .EQN("~(B*A)"),
    .INIT(4'h7))
    _al_u3868 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dhniu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Khniu6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mekiu6 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    _al_u3869 (
    .a(_al_u3255_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A1zhu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y8lpw6 ),
    .o(_al_u3869_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u387 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_state [0]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_state [1]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_state [2]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_state [3]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n88_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(C*~(~B*~(~D*A)))"),
    .INIT(16'hc0e0))
    _al_u3870 (
    .a(_al_u3869_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahlpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kwlpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pmlpw6 ),
    .o(_al_u3870_o));
  AL_MAP_LUT4 #(
    .EQN("~(~B*~(C*~(D*A)))"),
    .INIT(16'hdcfc))
    _al_u3871 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Di1iu6 ),
    .b(_al_u3870_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A5ipw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z73qw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nrxhu6 ));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B*A))"),
    .INIT(8'h70))
    _al_u3872 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Di1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bx2qw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ry2qw6 ),
    .o(_al_u3872_o));
  AL_MAP_LUT3 #(
    .EQN("~(~A*~(C*B))"),
    .INIT(8'hea))
    _al_u3873 (
    .a(_al_u3872_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fj1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yi1iu6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J3yhu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    _al_u3874 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T9qow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I4eiu6 ),
    .c(_al_u1299_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ur4iu6 ),
    .o(_al_u3874_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*~A))"),
    .INIT(16'h2a3f))
    _al_u3875 (
    .a(_al_u3874_o),
    .b(\u_cmsdk_mcu/HWDATA [31]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ch5iu6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pdyax6 ),
    .o(_al_u3875_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u3876 (
    .a(_al_u3875_o),
    .b(_al_u1777_o),
    .c(_al_u1791_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Npghu6 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u3877 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aaiiu6 ),
    .b(_al_u2832_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rwjax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yfiiu6 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*~A))"),
    .INIT(8'h8c))
    _al_u3878 (
    .a(_al_u2827_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yfiiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6 ),
    .o(_al_u3878_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*~B))"),
    .INIT(8'h8a))
    _al_u3879 (
    .a(_al_u3878_o),
    .b(_al_u2841_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Irmpw6 ),
    .o(_al_u3879_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u388 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_shift_in ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n88_lutinv ),
    .o(_al_u388_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*~B))"),
    .INIT(8'h54))
    _al_u3880 (
    .a(_al_u3423_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iekax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lgkax6 ),
    .o(_al_u3880_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B)*~(C)*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf722))
    _al_u3881 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D8iiu6 ),
    .b(_al_u3879_o),
    .c(_al_u3880_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oikax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jfthu6 ));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u3882 (
    .a(_al_u3318_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ph1iu6 ),
    .c(_al_u3319_o),
    .o(_al_u3882_o));
  AL_MAP_LUT4 #(
    .EQN("~(B*~(C*~(D*A)))"),
    .INIT(16'h73f3))
    _al_u3883 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Di1iu6 ),
    .b(_al_u3882_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I0opw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Li7ax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q3yhu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*C)*~(B*A))"),
    .INIT(16'h0777))
    _al_u3884 (
    .a(_al_u3808_o),
    .b(_al_u1533_o),
    .c(_al_u3797_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [28]),
    .o(_al_u3884_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u3885 (
    .a(_al_u3884_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A3iiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [30]),
    .o(_al_u3885_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u3886 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A3iiu6 ),
    .b(_al_u3797_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [30]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [32]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/If3pw6 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u3887 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/If3pw6 ),
    .b(_al_u3808_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/To2ju6_lutinv ),
    .o(_al_u3887_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u3888 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A3iiu6 ),
    .b(_al_u3797_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [29]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [31]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gd4pw6 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u3889 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gd4pw6 ),
    .b(_al_u3808_o),
    .c(_al_u1541_o),
    .o(_al_u3889_o));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    _al_u389 (
    .a(_al_u388_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/BAUDTICK ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/update_rx_tick_cnt ));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u3890 (
    .a(_al_u3885_o),
    .b(_al_u3887_o),
    .c(_al_u3889_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I7cow6 ));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3891 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hs8ow6 ),
    .b(_al_u3624_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 ),
    .o(_al_u3891_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(~D*C*A))"),
    .INIT(16'h3313))
    _al_u3892 (
    .a(_al_u696_o),
    .b(_al_u909_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pthiu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 ),
    .o(_al_u3892_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(~A*~(~D*B)))"),
    .INIT(16'h0a0e))
    _al_u3893 (
    .a(_al_u3891_o),
    .b(_al_u681_o),
    .c(_al_u3892_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ),
    .o(_al_u3893_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~A*~(D*C))"),
    .INIT(16'h0111))
    _al_u3894 (
    .a(_al_u2846_o),
    .b(_al_u3893_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P8oiu6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 ),
    .o(_al_u3894_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u3895 (
    .a(_al_u2771_o),
    .b(_al_u2832_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6 ),
    .o(_al_u3895_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3896 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qe8iu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vs0iu6 ),
    .c(_al_u1266_o),
    .o(_al_u3896_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D*~C*~A))"),
    .INIT(16'h3233))
    _al_u3897 (
    .a(_al_u3895_o),
    .b(_al_u3896_o),
    .c(_al_u1812_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 ),
    .o(_al_u3897_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u3898 (
    .a(_al_u1269_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N3ziu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Difiu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 ),
    .o(_al_u3898_o));
  AL_MAP_LUT4 #(
    .EQN("~(B*~((D*C))*~(A)+B*(D*C)*~(A)+~(B)*(D*C)*A+B*(D*C)*A)"),
    .INIT(16'h1bbb))
    _al_u3899 (
    .a(_al_u3109_o),
    .b(_al_u3898_o),
    .c(_al_u2779_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S2ziu6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fy8ow6_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    _al_u390 (
    .a(_al_u388_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n92 [3]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_rx_tick_cnt [3]));
  AL_MAP_LUT4 #(
    .EQN("(C*A*~(~D*~B))"),
    .INIT(16'ha080))
    _al_u3900 (
    .a(_al_u3894_o),
    .b(_al_u3897_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fy8ow6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vygax6 ),
    .o(_al_u3900_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3901 (
    .a(_al_u2371_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 ),
    .o(_al_u3901_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(~D*~C))"),
    .INIT(16'h4440))
    _al_u3902 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N4kax6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4jax6 ),
    .o(_al_u3902_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(~D*~C*B))"),
    .INIT(16'h5551))
    _al_u3903 (
    .a(_al_u3902_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rwjax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4jax6 ),
    .o(_al_u3903_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*~A)"),
    .INIT(16'h0004))
    _al_u3904 (
    .a(_al_u3901_o),
    .b(_al_u3903_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P14qw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 ),
    .o(_al_u3904_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(~D*C))"),
    .INIT(16'h8808))
    _al_u3905 (
    .a(_al_u2369_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N4kax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4jax6 ),
    .o(_al_u3905_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~(~B*A))"),
    .INIT(16'hd000))
    _al_u3906 (
    .a(_al_u3904_o),
    .b(_al_u3905_o),
    .c(_al_u2364_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 ),
    .o(_al_u3906_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(~A*~(C*B)))"),
    .INIT(16'h00ea))
    _al_u3907 (
    .a(_al_u3906_o),
    .b(_al_u2373_o),
    .c(_al_u3831_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hgrpw6 ),
    .o(_al_u3907_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3908 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nyiiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 ),
    .o(_al_u3908_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u3909 (
    .a(_al_u3908_o),
    .b(_al_u2367_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y40ju6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hgrpw6 ),
    .o(_al_u3909_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u391 (
    .a(_al_u388_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n92 [2]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_rx_tick_cnt [2]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u3910 (
    .a(_al_u2364_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P14qw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 ),
    .o(_al_u3910_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*A*~(D*C))"),
    .INIT(16'h0222))
    _al_u3911 (
    .a(_al_u3909_o),
    .b(_al_u3910_o),
    .c(_al_u2373_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dmiiu6 ),
    .o(_al_u3911_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u3912 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gr2qw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 ),
    .o(_al_u3912_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u3913 (
    .a(_al_u3912_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yj8ow6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D)"),
    .INIT(16'h035f))
    _al_u3914 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P14qw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 ),
    .o(_al_u3914_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(C*~(~D*B)))"),
    .INIT(16'h0a8a))
    _al_u3915 (
    .a(_al_u3911_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yj8ow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J9kiu6_lutinv ),
    .d(_al_u3914_o),
    .o(_al_u3915_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~(B*~A))"),
    .INIT(16'h000b))
    _al_u3916 (
    .a(_al_u3907_o),
    .b(_al_u3915_o),
    .c(_al_u1812_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vygax6 ),
    .o(_al_u3916_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u3917 (
    .a(_al_u678_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 ),
    .o(_al_u3917_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(D*C*~B))"),
    .INIT(16'h4555))
    _al_u3918 (
    .a(_al_u3666_o),
    .b(_al_u3917_o),
    .c(_al_u909_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ),
    .o(_al_u3918_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(~B*~(~D*C)))"),
    .INIT(16'h88a8))
    _al_u3919 (
    .a(_al_u1806_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ly2ju6 ),
    .c(_al_u604_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 ),
    .o(_al_u3919_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u392 (
    .a(_al_u388_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n92 [1]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_rx_tick_cnt [1]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*~A)"),
    .INIT(16'h0004))
    _al_u3920 (
    .a(_al_u3827_o),
    .b(_al_u3918_o),
    .c(_al_u697_o),
    .d(_al_u3919_o),
    .o(_al_u3920_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~(B*~A))"),
    .INIT(16'h000b))
    _al_u3921 (
    .a(_al_u3916_o),
    .b(_al_u3920_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv ),
    .o(_al_u3921_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(~A*~(C*~B)))"),
    .INIT(16'hba00))
    _al_u3922 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 ),
    .o(_al_u3922_o));
  AL_MAP_LUT4 #(
    .EQN("~(~C*~B*~(~D*~A))"),
    .INIT(16'hfcfd))
    _al_u3923 (
    .a(_al_u3900_o),
    .b(_al_u3921_o),
    .c(_al_u3922_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qrohu6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3924 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 ),
    .o(_al_u3924_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3925 (
    .a(_al_u1346_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Difiu6 ),
    .c(_al_u3924_o),
    .o(_al_u3925_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B*A))"),
    .INIT(8'h70))
    _al_u3926 (
    .a(_al_u3520_o),
    .b(_al_u3925_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [14]),
    .o(_al_u3926_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~D*~(C*A)))"),
    .INIT(16'hcc80))
    _al_u3927 (
    .a(_al_u1777_o),
    .b(_al_u3926_o),
    .c(_al_u3520_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qaipw6 ),
    .o(_al_u3927_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    _al_u3928 (
    .a(_al_u3874_o),
    .b(_al_u3518_o),
    .c(_al_u3927_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sgthu6 ));
  AL_MAP_LUT4 #(
    .EQN("(A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h3f08))
    _al_u3929 (
    .a(_al_u1777_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hwhiu6_lutinv ),
    .c(_al_u3925_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gv1bx6 ),
    .o(_al_u3929_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u393 (
    .a(_al_u388_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n92 [0]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_rx_tick_cnt [0]));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*~A)"),
    .INIT(16'h0100))
    _al_u3930 (
    .a(_al_u3874_o),
    .b(_al_u3533_o),
    .c(_al_u3534_o),
    .d(_al_u3929_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgthu6 ));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B*A))"),
    .INIT(8'h70))
    _al_u3931 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yogiu6_lutinv ),
    .b(_al_u3925_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/apbsubsys_interrupt [1]),
    .o(_al_u3931_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~D*~(C*A)))"),
    .INIT(16'hcc80))
    _al_u3932 (
    .a(_al_u1777_o),
    .b(_al_u3931_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yogiu6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y72bx6 ),
    .o(_al_u3932_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*~(D*B))"),
    .INIT(16'h1050))
    _al_u3933 (
    .a(_al_u3874_o),
    .b(\u_cmsdk_mcu/HWDATA [1]),
    .c(_al_u3932_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kwfiu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cmthu6 ));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u3934 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bggiu6_lutinv ),
    .b(_al_u3337_o),
    .c(_al_u3925_o),
    .o(_al_u3934_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(~D*~(C*B)))"),
    .INIT(16'haa80))
    _al_u3935 (
    .a(_al_u3934_o),
    .b(_al_u1777_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bggiu6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sq3bx6 ),
    .o(_al_u3935_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*~(D*B))"),
    .INIT(16'h1050))
    _al_u3936 (
    .a(_al_u3874_o),
    .b(\u_cmsdk_mcu/HWDATA [8]),
    .c(_al_u3935_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kwfiu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Enthu6 ));
  AL_MAP_LUT4 #(
    .EQN("(A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h3f08))
    _al_u3937 (
    .a(_al_u1777_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hcgiu6_lutinv ),
    .c(_al_u3925_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ca1bx6 ),
    .o(_al_u3937_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*~(D*A))"),
    .INIT(16'h40c0))
    _al_u3938 (
    .a(\u_cmsdk_mcu/HWDATA [10]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/apbsubsys_interrupt [10]),
    .c(_al_u3937_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kwfiu6 ),
    .o(_al_u3938_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u3939 (
    .a(_al_u3874_o),
    .b(_al_u3938_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Snthu6 ));
  AL_MAP_LUT4 #(
    .EQN("~(~B*~(D*C*~A))"),
    .INIT(16'hdccc))
    _al_u394 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cjqpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pifax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qwfax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Utqpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H43iu6 ));
  AL_MAP_LUT4 #(
    .EQN("(A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h3f08))
    _al_u3940 (
    .a(_al_u1777_o),
    .b(_al_u3443_o),
    .c(_al_u3925_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W51bx6 ),
    .o(_al_u3940_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~B*~(D*A))"),
    .INIT(16'h1030))
    _al_u3941 (
    .a(\u_cmsdk_mcu/HWDATA [12]),
    .b(_al_u3440_o),
    .c(_al_u3940_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kwfiu6 ),
    .o(_al_u3941_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u3942 (
    .a(_al_u3874_o),
    .b(_al_u3941_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gothu6 ));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B*A))"),
    .INIT(8'h70))
    _al_u3943 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jzfiu6_lutinv ),
    .b(_al_u3925_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [8]),
    .o(_al_u3943_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(~D*~(C*B)))"),
    .INIT(16'haa80))
    _al_u3944 (
    .a(_al_u3943_o),
    .b(_al_u1777_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jzfiu6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/At2bx6 ),
    .o(_al_u3944_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    _al_u3945 (
    .a(_al_u3874_o),
    .b(_al_u3492_o),
    .c(_al_u3944_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ipthu6 ));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B*A))"),
    .INIT(8'h70))
    _al_u3946 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mxfiu6_lutinv ),
    .b(_al_u3925_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [9]),
    .o(_al_u3946_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(~D*~(C*B)))"),
    .INIT(16'haa80))
    _al_u3947 (
    .a(_al_u3946_o),
    .b(_al_u1777_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mxfiu6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ok2bx6 ),
    .o(_al_u3947_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    _al_u3948 (
    .a(_al_u3874_o),
    .b(_al_u3498_o),
    .c(_al_u3947_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ppthu6 ));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B*A))"),
    .INIT(8'h70))
    _al_u3949 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ivfiu6_lutinv ),
    .b(_al_u3925_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [10]),
    .o(_al_u3949_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u395 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I5xax6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yzspw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K5eiu6 ));
  AL_MAP_LUT4 #(
    .EQN("(A*~(~D*~(C*B)))"),
    .INIT(16'haa80))
    _al_u3950 (
    .a(_al_u3949_o),
    .b(_al_u1777_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ivfiu6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gx2bx6 ),
    .o(_al_u3950_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    _al_u3951 (
    .a(_al_u3874_o),
    .b(_al_u3503_o),
    .c(_al_u3950_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wpthu6 ));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B*A))"),
    .INIT(8'h70))
    _al_u3952 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Etfiu6_lutinv ),
    .b(_al_u3925_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [11]),
    .o(_al_u3952_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(~D*~(C*B)))"),
    .INIT(16'haa80))
    _al_u3953 (
    .a(_al_u3952_o),
    .b(_al_u1777_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Etfiu6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M13bx6 ),
    .o(_al_u3953_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    _al_u3954 (
    .a(_al_u3874_o),
    .b(_al_u3508_o),
    .c(_al_u3953_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dqthu6 ));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B*A))"),
    .INIT(8'h70))
    _al_u3955 (
    .a(_al_u3515_o),
    .b(_al_u3925_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [12]),
    .o(_al_u3955_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~D*~(C*A)))"),
    .INIT(16'hcc80))
    _al_u3956 (
    .a(_al_u1777_o),
    .b(_al_u3955_o),
    .c(_al_u3515_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S53bx6 ),
    .o(_al_u3956_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    _al_u3957 (
    .a(_al_u3874_o),
    .b(_al_u3513_o),
    .c(_al_u3956_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kqthu6 ));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u3958 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G9fiu6_lutinv ),
    .b(_al_u3359_o),
    .c(_al_u3925_o),
    .o(_al_u3958_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(~D*~(C*B)))"),
    .INIT(16'haa80))
    _al_u3959 (
    .a(_al_u3958_o),
    .b(_al_u1777_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G9fiu6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jp9bx6 ),
    .o(_al_u3959_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u396 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R9yax6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W5ypw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztupw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jcpow6 ));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*~(D*B))"),
    .INIT(16'h1050))
    _al_u3960 (
    .a(_al_u3874_o),
    .b(\u_cmsdk_mcu/HWDATA [6]),
    .c(_al_u3959_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kwfiu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Osthu6 ));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u3961 (
    .a(_al_u3372_o),
    .b(_al_u3369_o),
    .c(_al_u3925_o),
    .o(_al_u3961_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(~D*~(C*B)))"),
    .INIT(16'haa80))
    _al_u3962 (
    .a(_al_u3961_o),
    .b(_al_u1777_o),
    .c(_al_u3372_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Om3bx6 ),
    .o(_al_u3962_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*~(D*B))"),
    .INIT(16'h1050))
    _al_u3963 (
    .a(_al_u3874_o),
    .b(\u_cmsdk_mcu/HWDATA [7]),
    .c(_al_u3962_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kwfiu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vsthu6 ));
  AL_MAP_LUT4 #(
    .EQN("(A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h3f08))
    _al_u3964 (
    .a(_al_u1777_o),
    .b(_al_u3454_o),
    .c(_al_u3925_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ar1bx6 ),
    .o(_al_u3964_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*~A)"),
    .INIT(16'h0100))
    _al_u3965 (
    .a(_al_u3874_o),
    .b(_al_u3449_o),
    .c(_al_u3450_o),
    .d(_al_u3964_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vruhu6 ));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B*A))"),
    .INIT(8'h70))
    _al_u3966 (
    .a(_al_u3463_o),
    .b(_al_u3925_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [2]),
    .o(_al_u3966_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(~D*~(C*B)))"),
    .INIT(16'haa80))
    _al_u3967 (
    .a(_al_u3966_o),
    .b(_al_u1777_o),
    .c(_al_u3463_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mz1bx6 ),
    .o(_al_u3967_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    _al_u3968 (
    .a(_al_u3874_o),
    .b(_al_u3461_o),
    .c(_al_u3967_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jsuhu6 ));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B*A))"),
    .INIT(8'h70))
    _al_u3969 (
    .a(_al_u3468_o),
    .b(_al_u3925_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [3]),
    .o(_al_u3969_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u397 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K5eiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jcpow6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hqgiu6 ));
  AL_MAP_LUT4 #(
    .EQN("(A*~(~D*~(C*B)))"),
    .INIT(16'haa80))
    _al_u3970 (
    .a(_al_u3969_o),
    .b(_al_u1777_o),
    .c(_al_u3468_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S32bx6 ),
    .o(_al_u3970_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    _al_u3971 (
    .a(_al_u3874_o),
    .b(_al_u3466_o),
    .c(_al_u3970_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xsuhu6 ));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B*A))"),
    .INIT(8'h70))
    _al_u3972 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lhdiu6_lutinv ),
    .b(_al_u3925_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [4]),
    .o(_al_u3972_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(~D*~(C*B)))"),
    .INIT(16'haa80))
    _al_u3973 (
    .a(_al_u3972_o),
    .b(_al_u1777_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lhdiu6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cc2bx6 ),
    .o(_al_u3973_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    _al_u3974 (
    .a(_al_u3874_o),
    .b(_al_u3471_o),
    .c(_al_u3973_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ltuhu6 ));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B*A))"),
    .INIT(8'h70))
    _al_u3975 (
    .a(_al_u3479_o),
    .b(_al_u3925_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [5]),
    .o(_al_u3975_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(~D*~(C*B)))"),
    .INIT(16'haa80))
    _al_u3976 (
    .a(_al_u3975_o),
    .b(_al_u1777_o),
    .c(_al_u3479_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ig2bx6 ),
    .o(_al_u3976_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    _al_u3977 (
    .a(_al_u3874_o),
    .b(_al_u3477_o),
    .c(_al_u3976_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztuhu6 ));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B*A))"),
    .INIT(8'h70))
    _al_u3978 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nbdiu6_lutinv ),
    .b(_al_u3925_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [6]),
    .o(_al_u3978_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(~D*~(C*B)))"),
    .INIT(16'haa80))
    _al_u3979 (
    .a(_al_u3978_o),
    .b(_al_u1777_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nbdiu6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vyfbx6 ),
    .o(_al_u3979_o));
  AL_MAP_LUT2 #(
    .EQN("~(B*A)"),
    .INIT(4'h7))
    _al_u398 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hqgiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C1wpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aqgiu6 ));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    _al_u3980 (
    .a(_al_u3874_o),
    .b(_al_u3482_o),
    .c(_al_u3979_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uuuhu6 ));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B*A))"),
    .INIT(8'h70))
    _al_u3981 (
    .a(_al_u3489_o),
    .b(_al_u3925_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [7]),
    .o(_al_u3981_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(~D*~(C*B)))"),
    .INIT(16'haa80))
    _al_u3982 (
    .a(_al_u3981_o),
    .b(_al_u1777_o),
    .c(_al_u3489_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uo2bx6 ),
    .o(_al_u3982_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    _al_u3983 (
    .a(_al_u3874_o),
    .b(_al_u3487_o),
    .c(_al_u3982_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pvuhu6 ));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B*A))"),
    .INIT(8'h70))
    _al_u3984 (
    .a(_al_u3530_o),
    .b(_al_u3925_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [13]),
    .o(_al_u3984_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~D*~(C*A)))"),
    .INIT(16'hcc80))
    _al_u3985 (
    .a(_al_u1777_o),
    .b(_al_u3984_o),
    .c(_al_u3530_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y93bx6 ),
    .o(_al_u3985_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    _al_u3986 (
    .a(_al_u3874_o),
    .b(_al_u3528_o),
    .c(_al_u3985_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J6vhu6 ));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B*A))"),
    .INIT(8'h70))
    _al_u3987 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Webiu6 ),
    .b(_al_u3925_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [15]),
    .o(_al_u3987_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~D*~(C*A)))"),
    .INIT(16'hcc80))
    _al_u3988 (
    .a(_al_u1777_o),
    .b(_al_u3987_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Webiu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ee3bx6 ),
    .o(_al_u3988_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    _al_u3989 (
    .a(_al_u3874_o),
    .b(_al_u3523_o),
    .c(_al_u3988_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q6vhu6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u399 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I5xax6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yzspw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vynow6_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B*A))"),
    .INIT(8'h70))
    _al_u3990 (
    .a(_al_u3335_o),
    .b(_al_u3925_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/apbsubsys_interrupt [0]),
    .o(_al_u3990_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(~D*~(C*B)))"),
    .INIT(16'haa80))
    _al_u3991 (
    .a(_al_u3990_o),
    .b(_al_u1777_o),
    .c(_al_u3335_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S11bx6 ),
    .o(_al_u3991_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*~(D*B))"),
    .INIT(16'h1050))
    _al_u3992 (
    .a(_al_u3874_o),
    .b(\u_cmsdk_mcu/HWDATA [0]),
    .c(_al_u3991_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kwfiu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mivhu6 ));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3993 (
    .a(_al_u909_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ),
    .o(_al_u3993_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3994 (
    .a(_al_u3993_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ),
    .o(_al_u3994_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3995 (
    .a(_al_u679_o),
    .b(_al_u1582_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 ),
    .o(_al_u3995_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~B*~(C*A))"),
    .INIT(16'h0013))
    _al_u3996 (
    .a(_al_u3183_o),
    .b(_al_u3994_o),
    .c(_al_u3910_o),
    .d(_al_u3995_o),
    .o(_al_u3996_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*~A)"),
    .INIT(8'h04))
    _al_u3997 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N4kax6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4jax6 ),
    .o(_al_u3997_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3998 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wh0ju6 ),
    .b(_al_u3997_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jckax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J8ziu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D*A)))"),
    .INIT(16'h2303))
    _al_u3999 (
    .a(_al_u2371_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P14qw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Skjax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ea7ow6_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    _al_u400 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R9yax6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W5ypw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztupw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D5eiu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*C)*~(B*A))"),
    .INIT(16'h0777))
    _al_u4000 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dd7ow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J8ziu6 ),
    .c(_al_u3246_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ea7ow6_lutinv ),
    .o(_al_u4000_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u4001 (
    .a(_al_u2373_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dmiiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P14qw6 ),
    .o(_al_u4001_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*~A)"),
    .INIT(16'h4000))
    _al_u4002 (
    .a(_al_u1812_o),
    .b(_al_u4001_o),
    .c(_al_u2369_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 ),
    .o(_al_u4002_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*A*~(~D*~B))"),
    .INIT(16'h0a08))
    _al_u4003 (
    .a(_al_u3996_o),
    .b(_al_u4000_o),
    .c(_al_u4002_o),
    .d(_al_u1812_o),
    .o(_al_u4003_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D*C*~B))"),
    .INIT(16'h8aaa))
    _al_u4004 (
    .a(_al_u4003_o),
    .b(_al_u3109_o),
    .c(_al_u1806_o),
    .d(_al_u1266_o),
    .o(_al_u4004_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u4005 (
    .a(_al_u3227_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nbkiu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qxoiu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sh7ow6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(C*~A))"),
    .INIT(16'haf23))
    _al_u4006 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sh7ow6 ),
    .b(_al_u4001_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dmiiu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rwjax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yd7ow6_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u4007 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N4kax6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rwjax6 ),
    .o(_al_u4007_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~(B*~A))"),
    .INIT(16'h000b))
    _al_u4008 (
    .a(_al_u4007_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4jax6 ),
    .o(_al_u4008_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(C*~B*A))"),
    .INIT(16'h00df))
    _al_u4009 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qz0ju6 ),
    .b(_al_u4008_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hgrpw6 ),
    .o(_al_u4009_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u401 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vynow6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D5eiu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6eiu6 ));
  AL_MAP_LUT4 #(
    .EQN("(A*~(C*~(~D*~B)))"),
    .INIT(16'h0a2a))
    _al_u4010 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yd7ow6_lutinv ),
    .b(_al_u4009_o),
    .c(_al_u2365_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9ypw6 ),
    .o(_al_u4010_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(A*~(C*~B)))"),
    .INIT(16'h0075))
    _al_u4011 (
    .a(_al_u4004_o),
    .b(_al_u4010_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uyiiu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vygax6 ),
    .o(_al_u4011_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u4012 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pu1ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yi7ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ),
    .o(_al_u4012_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~A*~(D*B))"),
    .INIT(16'h0105))
    _al_u4013 (
    .a(_al_u3189_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z37ow6_lutinv ),
    .c(_al_u4012_o),
    .d(_al_u1582_o),
    .o(_al_u4013_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~A*~(D*C))"),
    .INIT(16'h0111))
    _al_u4014 (
    .a(_al_u904_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pu1ju6_lutinv ),
    .d(_al_u2392_o),
    .o(_al_u4014_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*~B*A)"),
    .INIT(16'h0020))
    _al_u4015 (
    .a(_al_u4013_o),
    .b(_al_u3186_o),
    .c(_al_u4014_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uu9ow6_lutinv ),
    .o(_al_u4015_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u4016 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nu9ow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ),
    .o(_al_u4016_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(~B*~(C*A)))"),
    .INIT(16'hec00))
    _al_u4017 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv ),
    .b(_al_u903_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D6kiu6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yecpw6_lutinv ),
    .o(_al_u4017_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*A)"),
    .INIT(16'h0002))
    _al_u4018 (
    .a(_al_u4015_o),
    .b(_al_u1784_o),
    .c(_al_u4016_o),
    .d(_al_u4017_o),
    .o(_al_u4018_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u4019 (
    .a(_al_u1802_o),
    .b(_al_u1268_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 ),
    .o(_al_u4019_o));
  AL_MAP_LUT2 #(
    .EQN("~(B*A)"),
    .INIT(4'h7))
    _al_u402 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6eiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C1wpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F6eiu6 ));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*~A)"),
    .INIT(16'h0100))
    _al_u4020 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P14qw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Skjax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V17ow6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u4021 (
    .a(_al_u4018_o),
    .b(_al_u4019_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Htyiu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V17ow6_lutinv ),
    .o(_al_u4021_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*C)*~(B*A))"),
    .INIT(16'h0777))
    _al_u4022 (
    .a(_al_u908_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nsaiu6_lutinv ),
    .c(_al_u932_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 ),
    .o(_al_u4022_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(~D*~(C*~B)))"),
    .INIT(16'haa20))
    _al_u4023 (
    .a(_al_u4021_o),
    .b(_al_u3824_o),
    .c(_al_u4022_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 ),
    .o(_al_u4023_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*C)*~(B*~A))"),
    .INIT(16'hbb0b))
    _al_u4024 (
    .a(_al_u4011_o),
    .b(_al_u4023_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsohu6 ));
  AL_MAP_LUT4 #(
    .EQN("(D*A*~(~C*~B))"),
    .INIT(16'ha800))
    _al_u4025 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oulpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qa1qw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qj1qw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vplpw6 ),
    .o(_al_u4025_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u4026 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tezhu6 ),
    .b(_al_u4025_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sbyhu6 ));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u4027 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rkzhu6 ),
    .b(_al_u3390_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bclpw6 ),
    .o(_al_u4027_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B*A))"),
    .INIT(8'h70))
    _al_u4028 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ffyhu6 ),
    .b(_al_u4027_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rilpw6 ),
    .o(_al_u4028_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(~A*~(~C*B)))"),
    .INIT(16'h00ae))
    _al_u4029 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Agyhu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rkzhu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bclpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rilpw6 ),
    .o(_al_u4029_o));
  AL_MAP_LUT4 #(
    .EQN("(C*(~(A)*~(B)*~(D)+A*B*D))"),
    .INIT(16'h8010))
    _al_u403 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D2opw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yzlpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z73qw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgfax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ne3iu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D)"),
    .INIT(16'h1bf0))
    _al_u4030 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bclpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jflpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kalpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sdlpw6 ),
    .o(_al_u4030_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~A*~(D*~C))"),
    .INIT(16'h1011))
    _al_u4031 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lbyhu6 ),
    .b(_al_u4029_o),
    .c(_al_u4030_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yklpw6 ),
    .o(_al_u4031_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C*~B*~A))"),
    .INIT(16'hef00))
    _al_u4032 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sbyhu6 ),
    .b(_al_u4028_o),
    .c(_al_u4031_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U5yhu6 ),
    .o(_al_u4032_o));
  AL_MAP_LUT4 #(
    .EQN("~(~A*~(C*~(~D*B)))"),
    .INIT(16'hfaba))
    _al_u4033 (
    .a(_al_u4032_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cayhu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahlpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rilpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zehpw6 [6]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*C)*~(B*A))"),
    .INIT(16'h0777))
    _al_u4034 (
    .a(_al_u3808_o),
    .b(_al_u1397_o),
    .c(_al_u3797_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [11]),
    .o(_al_u4034_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u4035 (
    .a(_al_u4034_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A3iiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [13]),
    .o(_al_u4035_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~(~B*~A))"),
    .INIT(16'he000))
    _al_u4036 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vviiu6 ),
    .b(_al_u3081_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Skjax6 ),
    .o(_al_u4036_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u4037 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W0piu6_lutinv ),
    .b(_al_u3227_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 ),
    .o(_al_u4037_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*A*~(~D*~C))"),
    .INIT(16'h2220))
    _al_u4038 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zyoiu6 ),
    .b(_al_u1812_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6 ),
    .o(_al_u4038_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u4039 (
    .a(_al_u4037_o),
    .b(_al_u4038_o),
    .c(_al_u697_o),
    .d(_al_u3667_o),
    .o(_al_u4039_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u404 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R9yax6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W5ypw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztupw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wjyiu6 ));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(B*~A))"),
    .INIT(8'h0b))
    _al_u4040 (
    .a(_al_u4036_o),
    .b(_al_u4039_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv ),
    .o(_al_u4040_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u4041 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qe8iu6_lutinv ),
    .b(_al_u604_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 ),
    .o(_al_u4041_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u4042 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F85iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y0jiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Owoiu6 ),
    .o(_al_u4042_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(D*C))"),
    .INIT(16'h0444))
    _al_u4043 (
    .a(_al_u4041_o),
    .b(_al_u4042_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L0niu6 ),
    .d(_al_u3110_o),
    .o(_al_u4043_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*B*~(D*~A))"),
    .INIT(16'h080c))
    _al_u4044 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R9aiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M8fax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9ypw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wkipw6 ),
    .o(_al_u4044_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~(~B*A))"),
    .INIT(16'hd000))
    _al_u4045 (
    .a(_al_u1812_o),
    .b(_al_u4044_o),
    .c(_al_u930_o),
    .d(_al_u1359_o),
    .o(_al_u4045_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*A*~(~D*B))"),
    .INIT(16'h0a02))
    _al_u4046 (
    .a(_al_u4043_o),
    .b(_al_u2754_o),
    .c(_al_u4045_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 ),
    .o(_al_u4046_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u4047 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D5eiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rzciu6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ar1iu6 ));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u4048 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/HALTED ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ar1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C1wpw6 ),
    .o(_al_u4048_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(~D*~(B*~A)))"),
    .INIT(16'h0f04))
    _al_u4049 (
    .a(_al_u4040_o),
    .b(_al_u4046_o),
    .c(_al_u4048_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ),
    .o(_al_u4049_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u405 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vynow6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wjyiu6 ),
    .o(_al_u405_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*~(~D*B))"),
    .INIT(16'h5010))
    _al_u4050 (
    .a(_al_u4049_o),
    .b(_al_u2860_o),
    .c(_al_u903_o),
    .d(_al_u3811_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ok8iu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4051 (
    .a(_al_u4049_o),
    .b(_al_u4048_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X44iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dm6bx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Emmiu6 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u4052 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ok8iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Emmiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[11] ),
    .o(_al_u4052_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u4053 (
    .a(_al_u4049_o),
    .b(_al_u903_o),
    .c(_al_u1264_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jl8iu6 ));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C*~A))"),
    .INIT(8'h73))
    _al_u4054 (
    .a(_al_u4035_o),
    .b(_al_u4052_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jl8iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K8qhu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*C)*~(B*A))"),
    .INIT(16'h0777))
    _al_u4055 (
    .a(_al_u3808_o),
    .b(_al_u1429_o),
    .c(_al_u3797_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [15]),
    .o(_al_u4055_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u4056 (
    .a(_al_u4055_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A3iiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [17]),
    .o(_al_u4056_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4057 (
    .a(_al_u4049_o),
    .b(_al_u4048_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z54iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Chwpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dbmiu6 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u4058 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ok8iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dbmiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[15] ),
    .o(_al_u4058_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C*~A))"),
    .INIT(8'h73))
    _al_u4059 (
    .a(_al_u4056_o),
    .b(_al_u4058_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jl8iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sqqhu6 ));
  AL_MAP_LUT2 #(
    .EQN("~(B*A)"),
    .INIT(4'h7))
    _al_u406 (
    .a(_al_u405_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C1wpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R5eiu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*C)*~(B*A))"),
    .INIT(16'h0777))
    _al_u4060 (
    .a(_al_u3808_o),
    .b(_al_u1437_o),
    .c(_al_u3797_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [16]),
    .o(_al_u4060_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u4061 (
    .a(_al_u4060_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A3iiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [18]),
    .o(_al_u4061_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4062 (
    .a(_al_u4049_o),
    .b(_al_u4048_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G64iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pbbbx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E8miu6 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u4063 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ok8iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E8miu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[16] ),
    .o(_al_u4063_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C*~A))"),
    .INIT(8'h73))
    _al_u4064 (
    .a(_al_u4061_o),
    .b(_al_u4063_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jl8iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hvqhu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*C)*~(B*A))"),
    .INIT(16'h0777))
    _al_u4065 (
    .a(_al_u3808_o),
    .b(_al_u1445_o),
    .c(_al_u3797_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [17]),
    .o(_al_u4065_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u4066 (
    .a(_al_u4065_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A3iiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [19]),
    .o(_al_u4066_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4067 (
    .a(_al_u4049_o),
    .b(_al_u4048_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N64iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Syjbx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F5miu6 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u4068 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ok8iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F5miu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[17] ),
    .o(_al_u4068_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C*~A))"),
    .INIT(8'h73))
    _al_u4069 (
    .a(_al_u4066_o),
    .b(_al_u4068_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jl8iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wzqhu6 ));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*~A)"),
    .INIT(8'h04))
    _al_u407 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R9yax6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W5ypw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztupw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xznow6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*C)*~(B*A))"),
    .INIT(16'h0777))
    _al_u4070 (
    .a(_al_u3808_o),
    .b(_al_u1453_o),
    .c(_al_u3797_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [18]),
    .o(_al_u4070_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u4071 (
    .a(_al_u4070_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A3iiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [20]),
    .o(_al_u4071_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4072 (
    .a(_al_u4049_o),
    .b(_al_u4048_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U64iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T6kbx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G2miu6 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u4073 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ok8iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G2miu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[18] ),
    .o(_al_u4073_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C*~A))"),
    .INIT(8'h73))
    _al_u4074 (
    .a(_al_u4071_o),
    .b(_al_u4073_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jl8iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L4rhu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*C)*~(B*A))"),
    .INIT(16'h0777))
    _al_u4075 (
    .a(_al_u3808_o),
    .b(_al_u1461_o),
    .c(_al_u3797_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [19]),
    .o(_al_u4075_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u4076 (
    .a(_al_u4075_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A3iiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [21]),
    .o(_al_u4076_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4077 (
    .a(_al_u4049_o),
    .b(_al_u4048_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B74iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fjdbx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hzliu6 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u4078 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ok8iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hzliu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[19] ),
    .o(_al_u4078_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C*~A))"),
    .INIT(8'h73))
    _al_u4079 (
    .a(_al_u4076_o),
    .b(_al_u4078_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jl8iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A9rhu6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u408 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I5xax6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yzspw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rzciu6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*C)*~(B*A))"),
    .INIT(16'h0777))
    _al_u4080 (
    .a(_al_u3808_o),
    .b(_al_u1469_o),
    .c(_al_u3797_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [20]),
    .o(_al_u4080_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u4081 (
    .a(_al_u4080_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A3iiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [22]),
    .o(_al_u4081_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4082 (
    .a(_al_u4049_o),
    .b(_al_u4048_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I74iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M2ebx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bwliu6 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u4083 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ok8iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bwliu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[20] ),
    .o(_al_u4083_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C*~A))"),
    .INIT(8'h73))
    _al_u4084 (
    .a(_al_u4081_o),
    .b(_al_u4083_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jl8iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pdrhu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*C)*~(B*A))"),
    .INIT(16'h0777))
    _al_u4085 (
    .a(_al_u3808_o),
    .b(_al_u1477_o),
    .c(_al_u3797_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [21]),
    .o(_al_u4085_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u4086 (
    .a(_al_u4085_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A3iiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [23]),
    .o(_al_u4086_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4087 (
    .a(_al_u4049_o),
    .b(_al_u4048_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P74iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tlebx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ctliu6 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u4088 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ok8iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ctliu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[21] ),
    .o(_al_u4088_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C*~A))"),
    .INIT(8'h73))
    _al_u4089 (
    .a(_al_u4086_o),
    .b(_al_u4088_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jl8iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eirhu6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u409 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xznow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rzciu6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fpgiu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*C)*~(B*A))"),
    .INIT(16'h0777))
    _al_u4090 (
    .a(_al_u3808_o),
    .b(_al_u1485_o),
    .c(_al_u3797_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [22]),
    .o(_al_u4090_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u4091 (
    .a(_al_u4090_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A3iiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [24]),
    .o(_al_u4091_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4092 (
    .a(_al_u4049_o),
    .b(_al_u4048_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W74iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztgbx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kv9iu6 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u4093 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ok8iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kv9iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[22] ),
    .o(_al_u4093_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C*~A))"),
    .INIT(8'h73))
    _al_u4094 (
    .a(_al_u4091_o),
    .b(_al_u4093_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jl8iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kavhu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*C)*~(~B*A))"),
    .INIT(16'h0ddd))
    _al_u4095 (
    .a(_al_u3808_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E17ju6_lutinv ),
    .c(_al_u3797_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [25]),
    .o(_al_u4095_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u4096 (
    .a(_al_u4095_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A3iiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [27]),
    .o(_al_u4096_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4097 (
    .a(_al_u4049_o),
    .b(_al_u4048_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R84iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F8cbx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mzkiu6 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u4098 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ok8iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mzkiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[25] ),
    .o(_al_u4098_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C*~A))"),
    .INIT(8'h73))
    _al_u4099 (
    .a(_al_u4096_o),
    .b(_al_u4098_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jl8iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W5shu6 ));
  AL_MAP_LUT2 #(
    .EQN("~(B*A)"),
    .INIT(4'h7))
    _al_u410 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fpgiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C1wpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P3fiu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*C)*~(~B*A))"),
    .INIT(16'h0ddd))
    _al_u4100 (
    .a(_al_u3808_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F57ju6_lutinv ),
    .c(_al_u3797_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [26]),
    .o(_al_u4100_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u4101 (
    .a(_al_u4100_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A3iiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [28]),
    .o(_al_u4101_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4102 (
    .a(_al_u4049_o),
    .b(_al_u4048_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y84iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nybbx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E2liu6 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u4103 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ok8iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E2liu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[26] ),
    .o(_al_u4103_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C*~A))"),
    .INIT(8'h73))
    _al_u4104 (
    .a(_al_u4101_o),
    .b(_al_u4103_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jl8iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H1shu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*C)*~(B*A))"),
    .INIT(16'h0777))
    _al_u4105 (
    .a(_al_u3808_o),
    .b(_al_u1608_o),
    .c(_al_u3797_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [7]),
    .o(_al_u4105_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u4106 (
    .a(_al_u4105_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A3iiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [9]),
    .o(_al_u4106_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4107 (
    .a(_al_u4049_o),
    .b(_al_u4048_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pl4iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N61qw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y3niu6 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u4108 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ok8iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y3niu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[7] ),
    .o(_al_u4108_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C*~A))"),
    .INIT(8'h73))
    _al_u4109 (
    .a(_al_u4106_o),
    .b(_al_u4108_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jl8iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vpphu6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u411 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I5xax6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yzspw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pjyiu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*C)*~(B*A))"),
    .INIT(16'h0777))
    _al_u4110 (
    .a(_al_u3808_o),
    .b(_al_u1624_o),
    .c(_al_u3797_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [9]),
    .o(_al_u4110_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u4111 (
    .a(_al_u4110_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A3iiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [11]),
    .o(_al_u4111_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4112 (
    .a(_al_u4049_o),
    .b(_al_u4048_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J44iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gwxpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ivmiu6 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u4113 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ok8iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ivmiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[9] ),
    .o(_al_u4113_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C*~A))"),
    .INIT(8'h73))
    _al_u4114 (
    .a(_al_u4111_o),
    .b(_al_u4113_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jl8iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gzphu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4115 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A3iiu6 ),
    .b(_al_u3797_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [10]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [12]),
    .o(_al_u4115_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u4116 (
    .a(_al_u4115_o),
    .b(_al_u3808_o),
    .c(_al_u1632_o),
    .o(_al_u4116_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4117 (
    .a(_al_u4049_o),
    .b(_al_u4048_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q44iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C07bx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Womiu6 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u4118 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ok8iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Womiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[10] ),
    .o(_al_u4118_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C*~A))"),
    .INIT(8'h73))
    _al_u4119 (
    .a(_al_u4116_o),
    .b(_al_u4118_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jl8iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V3qhu6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u412 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xznow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pjyiu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tzdiu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*C)*~(B*A))"),
    .INIT(16'h0777))
    _al_u4120 (
    .a(_al_u3808_o),
    .b(_al_u1616_o),
    .c(_al_u3797_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [6]),
    .o(_al_u4120_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u4121 (
    .a(_al_u4120_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A3iiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [8]),
    .o(_al_u4121_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4122 (
    .a(_al_u4049_o),
    .b(_al_u4048_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gk4iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Asupw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Krkiu6 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u4123 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ok8iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Krkiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[6] ),
    .o(_al_u4123_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C*~A))"),
    .INIT(8'h73))
    _al_u4124 (
    .a(_al_u4121_o),
    .b(_al_u4123_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jl8iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hfshu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4125 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A3iiu6 ),
    .b(_al_u3797_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [12]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [14]),
    .o(_al_u4125_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u4126 (
    .a(_al_u4125_o),
    .b(_al_u3808_o),
    .c(_al_u1405_o),
    .o(_al_u4126_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4127 (
    .a(_al_u4049_o),
    .b(_al_u4048_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E54iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xpxax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mjmiu6 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u4128 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ok8iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mjmiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[12] ),
    .o(_al_u4128_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C*~A))"),
    .INIT(8'h73))
    _al_u4129 (
    .a(_al_u4126_o),
    .b(_al_u4128_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jl8iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zcqhu6 ));
  AL_MAP_LUT2 #(
    .EQN("~(B*A)"),
    .INIT(4'h7))
    _al_u413 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tzdiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C1wpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dv9iu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4130 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A3iiu6 ),
    .b(_al_u3797_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [13]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [15]),
    .o(_al_u4130_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u4131 (
    .a(_al_u4130_o),
    .b(_al_u3808_o),
    .c(_al_u1413_o),
    .o(_al_u4131_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4132 (
    .a(_al_u4049_o),
    .b(_al_u4048_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L54iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sb8ax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ugmiu6 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u4133 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ok8iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ugmiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[13] ),
    .o(_al_u4133_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C*~A))"),
    .INIT(8'h73))
    _al_u4134 (
    .a(_al_u4131_o),
    .b(_al_u4133_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jl8iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ohqhu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4135 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A3iiu6 ),
    .b(_al_u3797_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [14]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [16]),
    .o(_al_u4135_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u4136 (
    .a(_al_u4135_o),
    .b(_al_u3808_o),
    .c(_al_u1421_o),
    .o(_al_u4136_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4137 (
    .a(_al_u4049_o),
    .b(_al_u4048_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S54iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z47ax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cemiu6 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u4138 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ok8iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cemiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[14] ),
    .o(_al_u4138_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C*~A))"),
    .INIT(8'h73))
    _al_u4139 (
    .a(_al_u4136_o),
    .b(_al_u4138_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jl8iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dmqhu6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u414 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vynow6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xznow6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S1fiu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*C)*~(~B*A))"),
    .INIT(16'h0ddd))
    _al_u4140 (
    .a(_al_u3808_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mk6ju6_lutinv ),
    .c(_al_u3797_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [5]),
    .o(_al_u4140_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u4141 (
    .a(_al_u4140_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A3iiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [7]),
    .o(_al_u4141_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4142 (
    .a(_al_u4049_o),
    .b(_al_u4048_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xi4iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ua9bx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zokiu6 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u4143 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ok8iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zokiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[5] ),
    .o(_al_u4143_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C*~A))"),
    .INIT(8'h73))
    _al_u4144 (
    .a(_al_u4141_o),
    .b(_al_u4143_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jl8iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wjshu6 ));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u4145 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nz2ju6 ),
    .b(_al_u2868_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 ),
    .o(_al_u4145_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u4146 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qyniu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yljiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Owoiu6 ),
    .o(_al_u4146_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*A*~(D*C))"),
    .INIT(16'h0222))
    _al_u4147 (
    .a(_al_u4145_o),
    .b(_al_u4146_o),
    .c(_al_u682_o),
    .d(_al_u1329_o),
    .o(_al_u4147_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(~C*~B*~A))"),
    .INIT(16'hfe00))
    _al_u4148 (
    .a(_al_u604_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sq3ju6 ),
    .c(_al_u1336_o),
    .d(_al_u2868_o),
    .o(_al_u4148_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(A*~(C*~B)))"),
    .INIT(16'h0075))
    _al_u4149 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wrcpw6 ));
  AL_MAP_LUT2 #(
    .EQN("~(B*A)"),
    .INIT(4'h7))
    _al_u415 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S1fiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C1wpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L1fiu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~C*A*~(D*B))"),
    .INIT(16'h020a))
    _al_u4150 (
    .a(_al_u4147_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Obbow6_lutinv ),
    .c(_al_u4148_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wrcpw6 ),
    .o(_al_u4150_o));
  AL_MAP_LUT4 #(
    .EQN("(A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .INIT(16'ha280))
    _al_u4151 (
    .a(_al_u3122_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 ),
    .o(_al_u4151_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D*~C*A))"),
    .INIT(16'h3133))
    _al_u4152 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zwcpw6_lutinv ),
    .b(_al_u4151_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 ),
    .o(_al_u4152_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u4153 (
    .a(_al_u1813_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N98iu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ),
    .o(_al_u4153_o));
  AL_MAP_LUT4 #(
    .EQN("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'hc0a0))
    _al_u4154 (
    .a(_al_u2849_o),
    .b(_al_u4153_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 ),
    .o(_al_u4154_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*A*~(D*~B))"),
    .INIT(16'h080a))
    _al_u4155 (
    .a(_al_u4150_o),
    .b(_al_u4152_o),
    .c(_al_u4154_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F9vpw6 ),
    .o(_al_u4155_o));
  AL_MAP_LUT4 #(
    .EQN("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'ha088))
    _al_u4156 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hgrpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Skjax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9ypw6 ),
    .o(_al_u4156_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u4157 (
    .a(_al_u1799_o),
    .b(_al_u4156_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ),
    .o(_al_u4157_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~A*~(~D*C)))"),
    .INIT(16'h88c8))
    _al_u4158 (
    .a(_al_u4157_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Llaow6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vo3ju6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 ),
    .o(_al_u4158_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u4159 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kxziu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hbbow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 ),
    .o(_al_u4159_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    _al_u416 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pjyiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R9yax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W5ypw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztupw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U2fiu6 ));
  AL_MAP_LUT4 #(
    .EQN("(C*~(~A*~(~D*B)))"),
    .INIT(16'ha0e0))
    _al_u4160 (
    .a(_al_u4158_o),
    .b(_al_u4159_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F9vpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ),
    .o(_al_u4160_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u4161 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D6kiu6_lutinv ),
    .b(_al_u1582_o),
    .o(_al_u4161_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*~A)"),
    .INIT(16'h1000))
    _al_u4162 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vygax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 ),
    .o(_al_u4162_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~A*~(D*B))"),
    .INIT(16'h0105))
    _al_u4163 (
    .a(_al_u4161_o),
    .b(_al_u903_o),
    .c(_al_u4162_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vygax6 ),
    .o(_al_u4163_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~A*~(D*C))"),
    .INIT(16'h0111))
    _al_u4164 (
    .a(_al_u908_o),
    .b(_al_u3591_o),
    .c(_al_u607_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vo3ju6_lutinv ),
    .o(_al_u4164_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u4165 (
    .a(_al_u4163_o),
    .b(_al_u4164_o),
    .c(_al_u1269_o),
    .d(_al_u678_o),
    .o(_al_u4165_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D*~(C*~B)))"),
    .INIT(16'h20aa))
    _al_u4166 (
    .a(_al_u4155_o),
    .b(_al_u4160_o),
    .c(_al_u4165_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 ),
    .o(_al_u4166_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*~A)"),
    .INIT(8'h04))
    _al_u4167 (
    .a(_al_u1336_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Et8iu6_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u4168 (
    .a(_al_u4166_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Et8iu6_lutinv ),
    .o(_al_u4168_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u4169 (
    .a(_al_u4168_o),
    .b(_al_u1299_o),
    .o(_al_u4169_o));
  AL_MAP_LUT2 #(
    .EQN("~(B*A)"),
    .INIT(4'h7))
    _al_u417 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U2fiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C1wpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N2fiu6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u4170 (
    .a(_al_u4169_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6lax6 ),
    .o(_al_u4170_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u4171 (
    .a(_al_u4170_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J0iax6 ),
    .o(_al_u4171_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u4172 (
    .a(_al_u3993_o),
    .b(_al_u679_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 ),
    .o(_al_u4172_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u4173 (
    .a(_al_u4166_o),
    .b(_al_u4172_o),
    .o(_al_u4173_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u4174 (
    .a(_al_u4171_o),
    .b(_al_u4173_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qqiow6 ));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u4175 (
    .a(_al_u2860_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M8fax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wkipw6 ),
    .o(_al_u4175_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*~B))"),
    .INIT(8'h54))
    _al_u4176 (
    .a(_al_u4049_o),
    .b(_al_u4175_o),
    .c(_al_u906_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vpoiu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(D*C*B))"),
    .INIT(16'h1555))
    _al_u4177 (
    .a(_al_u2373_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wa0ju6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rwjax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cqoiu6 ));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D*B*A))"),
    .INIT(16'h70f0))
    _al_u4178 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xqoiu6_lutinv ),
    .b(_al_u1812_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cqoiu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Irmpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U19iu6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u4179 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vpoiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U19iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ql8iu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    _al_u418 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vynow6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R9yax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W5ypw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztupw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q0fiu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4180 (
    .a(_al_u4049_o),
    .b(_al_u4048_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D84iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgkbx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gwkiu6 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u4181 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ok8iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gwkiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[23] ),
    .o(_al_u4181_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u4182 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ql8iu6 ),
    .b(_al_u4181_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_tbit_o ),
    .o(_al_u4182_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*C)*~(B*A))"),
    .INIT(16'h0777))
    _al_u4183 (
    .a(_al_u3808_o),
    .b(_al_u1493_o),
    .c(_al_u3797_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [23]),
    .o(_al_u4183_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u4184 (
    .a(_al_u4183_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A3iiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [25]),
    .o(_al_u4184_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*~B))"),
    .INIT(8'h75))
    _al_u4185 (
    .a(_al_u4182_o),
    .b(_al_u4184_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jl8iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lashu6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u4186 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vpoiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U19iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B29iu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4187 (
    .a(_al_u4049_o),
    .b(_al_u4048_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K84iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nwbbx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ipliu6 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u4188 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ok8iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ipliu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[24] ),
    .o(_al_u4188_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u4189 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B29iu6 ),
    .b(_al_u4188_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_control_o ),
    .o(_al_u4189_o));
  AL_MAP_LUT2 #(
    .EQN("~(B*A)"),
    .INIT(4'h7))
    _al_u419 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q0fiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C1wpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J0fiu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*C)*~(~B*A))"),
    .INIT(16'h0ddd))
    _al_u4190 (
    .a(_al_u3808_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mi8ju6_lutinv ),
    .c(_al_u3797_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [24]),
    .o(_al_u4190_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u4191 (
    .a(_al_u4190_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A3iiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [26]),
    .o(_al_u4191_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*~B))"),
    .INIT(8'h75))
    _al_u4192 (
    .a(_al_u4189_o),
    .b(_al_u4191_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jl8iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Anrhu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4193 (
    .a(_al_u4049_o),
    .b(_al_u4048_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F94iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ibqpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ocniu6 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u4194 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ok8iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ocniu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[27] ),
    .o(_al_u4194_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u4195 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ql8iu6 ),
    .b(_al_u4194_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_apsr_o[0] ),
    .o(_al_u4195_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*C)*~(B*A))"),
    .INIT(16'h0777))
    _al_u4196 (
    .a(_al_u3808_o),
    .b(_al_u1525_o),
    .c(_al_u3797_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [27]),
    .o(_al_u4196_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u4197 (
    .a(_al_u4196_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A3iiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [29]),
    .o(_al_u4197_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*~B))"),
    .INIT(8'h75))
    _al_u4198 (
    .a(_al_u4195_o),
    .b(_al_u4197_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jl8iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zkphu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4199 (
    .a(_al_u4049_o),
    .b(_al_u4048_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M94iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sx3qw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mj8iu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*~(B)*C*D)"),
    .INIT(16'h25a1))
    _al_u420 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [0]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [0]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpol_padded [0]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_last_datain [0]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_raw_int [0]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u4200 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ok8iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mj8iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[28] ),
    .o(_al_u4200_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u4201 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ql8iu6 ),
    .b(_al_u4200_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_apsr_o[1] ),
    .o(_al_u4201_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*~B))"),
    .INIT(8'h75))
    _al_u4202 (
    .a(_al_u4201_o),
    .b(_al_u3885_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jl8iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufvhu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4203 (
    .a(_al_u4049_o),
    .b(_al_u4048_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T94iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F6dbx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C8liu6 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u4204 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ok8iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C8liu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[29] ),
    .o(_al_u4204_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u4205 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ql8iu6 ),
    .b(_al_u4204_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_apsr_o[2] ),
    .o(_al_u4205_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*~B))"),
    .INIT(8'h75))
    _al_u4206 (
    .a(_al_u4205_o),
    .b(_al_u3889_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jl8iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dsrhu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4207 (
    .a(_al_u4049_o),
    .b(_al_u4048_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lm1iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Usnpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pmoiu6 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u4208 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ok8iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pmoiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[30] ),
    .o(_al_u4208_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u4209 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ql8iu6 ),
    .b(_al_u4208_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_apsr_o[3] ),
    .o(_al_u4209_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u421 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_raw_int [0]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inten_padded [0]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_masked_int [0]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*~B))"),
    .INIT(8'h75))
    _al_u4210 (
    .a(_al_u4209_o),
    .b(_al_u3887_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jl8iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dgphu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4211 (
    .a(_al_u4049_o),
    .b(_al_u4048_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T24iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I1lpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jz8iu6 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u4212 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B29iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jz8iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_primask_o ),
    .o(_al_u4212_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~A*~(D*~C)))"),
    .INIT(16'h8c88))
    _al_u4213 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ay8iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jl8iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U19iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_tbit_o ),
    .o(_al_u4213_o));
  AL_MAP_LUT4 #(
    .EQN("~(~C*A*~(D*B))"),
    .INIT(16'hfdf5))
    _al_u4214 (
    .a(_al_u4212_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ql8iu6 ),
    .c(_al_u4213_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[0] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qdvhu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4215 (
    .a(_al_u4049_o),
    .b(_al_u4048_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oh4iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qc5bx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ykkiu6 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u4216 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ok8iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ykkiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[4] ),
    .o(_al_u4216_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u4217 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ql8iu6 ),
    .b(_al_u4216_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[5] ),
    .o(_al_u4217_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4218 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A3iiu6 ),
    .b(_al_u3797_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [4]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [6]),
    .o(_al_u4218_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u4219 (
    .a(_al_u4218_o),
    .b(_al_u3808_o),
    .c(_al_u1600_o),
    .o(_al_u4219_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*~(B)*C*D)"),
    .INIT(16'h25a1))
    _al_u422 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [1]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [1]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpol_padded [1]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_last_datain [1]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_raw_int [1]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*~B))"),
    .INIT(8'h75))
    _al_u4220 (
    .a(_al_u4217_o),
    .b(_al_u4219_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jl8iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Loshu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4221 (
    .a(_al_u4049_o),
    .b(_al_u4048_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Df4iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T5yax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qgkiu6 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u4222 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ok8iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qgkiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[2] ),
    .o(_al_u4222_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u4223 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ql8iu6 ),
    .b(_al_u4222_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[3] ),
    .o(_al_u4223_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4224 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A3iiu6 ),
    .b(_al_u3797_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [2]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [4]),
    .o(_al_u4224_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u4225 (
    .a(_al_u4224_o),
    .b(_al_u3808_o),
    .c(_al_u1592_o),
    .o(_al_u4225_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*~B))"),
    .INIT(8'h75))
    _al_u4226 (
    .a(_al_u4223_o),
    .b(_al_u4225_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jl8iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Htshu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4227 (
    .a(_al_u4049_o),
    .b(_al_u4048_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H34iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wtxax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B0iiu6 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u4228 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ok8iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B0iiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[3] ),
    .o(_al_u4228_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u4229 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ql8iu6 ),
    .b(_al_u4228_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[4] ),
    .o(_al_u4229_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u423 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_raw_int [1]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inten_padded [1]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_masked_int [1]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4230 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A3iiu6 ),
    .b(_al_u3797_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [3]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [5]),
    .o(_al_u4230_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u4231 (
    .a(_al_u4230_o),
    .b(_al_u3808_o),
    .c(_al_u1573_o),
    .o(_al_u4231_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*~B))"),
    .INIT(8'h75))
    _al_u4232 (
    .a(_al_u4229_o),
    .b(_al_u4231_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jl8iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lgthu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4233 (
    .a(_al_u4049_o),
    .b(_al_u4048_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ym4iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kn1qw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z0niu6 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u4234 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ok8iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z0niu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[8] ),
    .o(_al_u4234_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(D*C*A))"),
    .INIT(16'h4ccc))
    _al_u4235 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ql8iu6 ),
    .b(_al_u4234_o),
    .c(_al_u1299_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F26bx6 ),
    .o(_al_u4235_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4236 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A3iiu6 ),
    .b(_al_u3797_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [8]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [10]),
    .o(_al_u4236_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*B))"),
    .INIT(8'ha2))
    _al_u4237 (
    .a(_al_u4236_o),
    .b(_al_u3808_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N18ju6_lutinv ),
    .o(_al_u4237_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*~B))"),
    .INIT(8'h75))
    _al_u4238 (
    .a(_al_u4235_o),
    .b(_al_u4237_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jl8iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kuphu6 ));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*~A)"),
    .INIT(8'h04))
    _al_u4239 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sbyhu6 ),
    .b(_al_u1250_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jflpw6 ),
    .o(_al_u4239_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*~(B)*C*D)"),
    .INIT(16'h25a1))
    _al_u424 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [10]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [10]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpol_padded [10]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_last_datain [10]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_raw_int [10]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u4240 (
    .a(_al_u1308_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bclpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rilpw6 ),
    .o(_al_u4240_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~A*~(D*B))"),
    .INIT(16'h0105))
    _al_u4241 (
    .a(_al_u4240_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Agyhu6 ),
    .c(_al_u2296_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rilpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J9zhu6 ));
  AL_MAP_LUT4 #(
    .EQN("~(A*~((D*B))*~(C)+A*(D*B)*~(C)+~(A)*(D*B)*C+A*(D*B)*C)"),
    .INIT(16'h35f5))
    _al_u4242 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Swyhu6 ),
    .b(_al_u1757_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bclpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yklpw6 ),
    .o(_al_u4242_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*A)"),
    .INIT(16'h0200))
    _al_u4243 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J9zhu6 ),
    .b(_al_u2295_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A1zhu6_lutinv ),
    .d(_al_u4242_o),
    .o(_al_u4243_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*~B))"),
    .INIT(8'h8a))
    _al_u4244 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Golpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Krlpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vplpw6 ),
    .o(_al_u4244_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*~B))"),
    .INIT(8'h8a))
    _al_u4245 (
    .a(_al_u2299_o),
    .b(_al_u4244_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y8lpw6 ),
    .o(_al_u4245_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u4246 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M7zhu6 ),
    .b(_al_u4244_o),
    .o(_al_u4246_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(D*~C*B))"),
    .INIT(16'h5155))
    _al_u4247 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rkzhu6 ),
    .b(_al_u1251_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jflpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yklpw6 ),
    .o(_al_u4247_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C*~B*~A))"),
    .INIT(16'hef00))
    _al_u4248 (
    .a(_al_u4245_o),
    .b(_al_u4246_o),
    .c(_al_u4247_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rilpw6 ),
    .o(_al_u4248_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*B*~(~D*A))"),
    .INIT(16'h0c04))
    _al_u4249 (
    .a(_al_u4239_o),
    .b(_al_u4243_o),
    .c(_al_u4248_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bclpw6 ),
    .o(_al_u4249_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u425 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_raw_int [10]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inten_padded [10]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_masked_int [10]));
  AL_MAP_LUT4 #(
    .EQN("~(~(~D*~B)*~(C*~A))"),
    .INIT(16'h5073))
    _al_u4250 (
    .a(_al_u4249_o),
    .b(_al_u1761_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U5yhu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bclpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zehpw6 [0]));
  AL_MAP_LUT4 #(
    .EQN("(D*~A*~(C*B))"),
    .INIT(16'h1500))
    _al_u4251 (
    .a(_al_u3874_o),
    .b(_al_u1774_o),
    .c(_al_u1777_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T8kbx6 ),
    .o(_al_u4251_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*A)"),
    .INIT(16'h0080))
    _al_u4252 (
    .a(_al_u4159_o),
    .b(_al_u679_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Frziu6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 ),
    .o(_al_u4252_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u4253 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ya1ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hgrpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fpaow6_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u4254 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fpaow6_lutinv ),
    .b(_al_u1367_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y7cpw6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*~A)"),
    .INIT(16'h4000))
    _al_u4255 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv ),
    .b(_al_u1296_o),
    .c(_al_u1344_o),
    .d(_al_u2403_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jxaiu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~C*~A*~(D*B))"),
    .INIT(16'h0105))
    _al_u4256 (
    .a(_al_u4252_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y7cpw6_lutinv ),
    .c(_al_u4151_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jxaiu6 ),
    .o(_al_u4256_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(D*C*~A))"),
    .INIT(16'h8ccc))
    _al_u4257 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0biu6 ),
    .b(_al_u4256_o),
    .c(_al_u3754_o),
    .d(_al_u3124_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxaiu6 ));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u4258 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jxaiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vo3ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 ),
    .o(_al_u4258_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u4259 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I8lax6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vygax6 ),
    .o(_al_u4259_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*~(B)*C*D)"),
    .INIT(16'h25a1))
    _al_u426 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [11]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [11]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpol_padded [11]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_last_datain [11]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_raw_int [11]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(C*B*A))"),
    .INIT(16'h007f))
    _al_u4260 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hwaiu6_lutinv ),
    .b(_al_u604_o),
    .c(_al_u1336_o),
    .d(_al_u4259_o),
    .o(_al_u4260_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(C*~B*A))"),
    .INIT(16'h00df))
    _al_u4261 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxaiu6 ),
    .b(_al_u4258_o),
    .c(_al_u4260_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F9vpw6 ),
    .o(_al_u4261_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    _al_u4262 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I8lax6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vygax6 ),
    .o(_al_u4262_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B*A))"),
    .INIT(8'h70))
    _al_u4263 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uzaiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B0biu6 ),
    .c(_al_u4262_o),
    .o(_al_u4263_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~A*~(D*~B))"),
    .INIT(16'h0405))
    _al_u4264 (
    .a(_al_u4261_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0biu6 ),
    .c(_al_u4263_o),
    .d(_al_u3753_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Li5iu6 ));
  AL_MAP_LUT2 #(
    .EQN("~(B*~A)"),
    .INIT(4'hb))
    _al_u4265 (
    .a(_al_u4251_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Li5iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G8vhu6 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u4266 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pyyhu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Krlpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zslpw6 ),
    .o(_al_u4266_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u4267 (
    .a(_al_u2299_o),
    .b(_al_u4266_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y8lpw6 ),
    .o(_al_u4267_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(~D*~C*B))"),
    .INIT(16'h5551))
    _al_u4268 (
    .a(_al_u2305_o),
    .b(_al_u2298_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jflpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yklpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X2zhu6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*~B*A)"),
    .INIT(16'h0020))
    _al_u4269 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J9zhu6 ),
    .b(_al_u4267_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X2zhu6_lutinv ),
    .d(_al_u3328_o),
    .o(_al_u4269_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u427 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_raw_int [11]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inten_padded [11]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_masked_int [11]));
  AL_MAP_LUT4 #(
    .EQN("(A*~(~D*C*B))"),
    .INIT(16'haa2a))
    _al_u4270 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Golpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Krlpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vplpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zslpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F7zhu6 ));
  AL_MAP_LUT4 #(
    .EQN("(D*~B*~(C*A))"),
    .INIT(16'h1300))
    _al_u4271 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lbyhu6 ),
    .b(_al_u3390_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F7zhu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rilpw6 ),
    .o(_al_u4271_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~A*~(C*B))"),
    .INIT(16'h0015))
    _al_u4272 (
    .a(_al_u2299_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rkzhu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bclpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rilpw6 ),
    .o(_al_u4272_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*~B))"),
    .INIT(8'ha8))
    _al_u4273 (
    .a(_al_u4269_o),
    .b(_al_u4271_o),
    .c(_al_u4272_o),
    .o(_al_u4273_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~D*~C*A))"),
    .INIT(16'hccc4))
    _al_u4274 (
    .a(_al_u4239_o),
    .b(_al_u4273_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bclpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Krlpw6 ),
    .o(_al_u4274_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(~A*(D@C)))"),
    .INIT(16'h3223))
    _al_u4275 (
    .a(_al_u1761_o),
    .b(_al_u1763_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bclpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sdlpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H1zhu6 ));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C*~A))"),
    .INIT(8'h73))
    _al_u4276 (
    .a(_al_u4274_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H1zhu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U5yhu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zehpw6 [1]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u4277 (
    .a(_al_u4170_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[0] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vtzhu6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u4278 (
    .a(_al_u4169_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J0iax6 ),
    .o(_al_u4278_o));
  AL_MAP_LUT3 #(
    .EQN("(A*B*~(C)+A*~(B)*C+~(A)*B*C+A*B*C)"),
    .INIT(8'he8))
    _al_u4279 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vtzhu6 ),
    .b(_al_u4278_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[1] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R0ghu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*~(B)*C*D)"),
    .INIT(16'h25a1))
    _al_u428 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [12]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [12]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpol_padded [12]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_last_datain [12]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_raw_int [12]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u4280 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kxziu6_lutinv ),
    .b(_al_u3690_o),
    .c(_al_u604_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F9vpw6 ),
    .o(_al_u4280_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(~A*~(D*B)))"),
    .INIT(16'he0a0))
    _al_u4281 (
    .a(_al_u4280_o),
    .b(_al_u2782_o),
    .c(_al_u696_o),
    .d(_al_u3924_o),
    .o(_al_u4281_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(D*C*B))"),
    .INIT(16'h1555))
    _al_u4282 (
    .a(_al_u4281_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mfjiu6 ),
    .c(_al_u1296_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vygax6 ),
    .o(_al_u4282_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u4283 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ldoiu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vo3ju6_lutinv ),
    .c(_al_u3924_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 ),
    .o(_al_u4283_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(D*~(~C*A)))"),
    .INIT(16'h08cc))
    _al_u4284 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxaiu6 ),
    .b(_al_u4282_o),
    .c(_al_u4283_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F9vpw6 ),
    .o(_al_u4284_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u4285 (
    .a(_al_u4284_o),
    .b(\u_cmsdk_mcu/LOCKUPRESET ),
    .o(\u_cmsdk_mcu/n1 ));
  AL_MAP_LUT4 #(
    .EQN("~(~A*~(D*~(C*B)))"),
    .INIT(16'hbfaa))
    _al_u4286 (
    .a(\u_cmsdk_mcu/n1 ),
    .b(\u_cmsdk_mcu/HWDATA [2]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_resetinfo_write ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_resetinfo [2]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/nxt_resetinfo [2]));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u4287 (
    .a(\u_cmsdk_mcu/n1 ),
    .b(\u_cmsdk_mcu/SYSRESETREQ ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/nxt_hrst ));
  AL_MAP_LUT2 #(
    .EQN("~(~B*A)"),
    .INIT(4'hd))
    _al_u4288 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/nxt_hrst ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_resetinfo_write ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_resetinfo_en ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u4289 (
    .a(_al_u4166_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ),
    .o(_al_u4289_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u429 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_raw_int [12]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inten_padded [12]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_masked_int [12]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u4290 (
    .a(_al_u4172_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Et8iu6_lutinv ),
    .o(_al_u4290_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(~C*~A))"),
    .INIT(16'hfa32))
    _al_u4291 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ),
    .o(_al_u4291_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*~(~D*C)))"),
    .INIT(16'h22a2))
    _al_u4292 (
    .a(_al_u4291_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 ),
    .o(_al_u4292_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    _al_u4293 (
    .a(_al_u4284_o),
    .b(_al_u4289_o),
    .c(_al_u4290_o),
    .d(_al_u4292_o),
    .o(_al_u4293_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u4294 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jjoiu6 ),
    .b(_al_u1299_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ),
    .o(_al_u4294_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    _al_u4295 (
    .a(_al_u1788_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ),
    .c(_al_u609_o),
    .o(_al_u4295_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u4296 (
    .a(_al_u4293_o),
    .b(_al_u4294_o),
    .c(_al_u4295_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nn8iu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(~B*~(~D*A)))"),
    .INIT(16'h0c0e))
    _al_u4297 (
    .a(_al_u4170_o),
    .b(_al_u4278_o),
    .c(_al_u4173_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ),
    .o(_al_u4297_o));
  AL_MAP_LUT3 #(
    .EQN("~(~A*~(C*B))"),
    .INIT(8'hea))
    _al_u4298 (
    .a(_al_u4297_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J0iax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hjohu6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u4299 (
    .a(_al_u4284_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zrhiu6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*~(B)*C*D)"),
    .INIT(16'h25a1))
    _al_u430 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [13]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [13]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpol_padded [13]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_last_datain [13]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_raw_int [13]));
  AL_MAP_LUT4 #(
    .EQN("(D*~B*~(~C*A))"),
    .INIT(16'h3100))
    _al_u4300 (
    .a(_al_u927_o),
    .b(_al_u933_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dg2qw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uh2qw6 ),
    .o(_al_u4300_o));
  AL_MAP_LUT2 #(
    .EQN("~(~B*A)"),
    .INIT(4'hd))
    _al_u4301 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zrhiu6_lutinv ),
    .b(_al_u4300_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ghthu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4302 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A3iiu6 ),
    .b(_al_u3808_o),
    .c(_al_u1354_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [2]),
    .o(_al_u4302_o));
  AL_MAP_LUT4 #(
    .EQN("~(B*~(C*(D@A)))"),
    .INIT(16'h73b3))
    _al_u4303 (
    .a(_al_u4170_o),
    .b(_al_u4302_o),
    .c(_al_u3797_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[0] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iiliu6 ));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    _al_u4304 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0biu6 ),
    .b(_al_u678_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 ),
    .o(_al_u4304_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u4305 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kxziu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sy2ju6 ),
    .o(_al_u4305_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(~A*~(C*B)))"),
    .INIT(16'h00ea))
    _al_u4306 (
    .a(_al_u4305_o),
    .b(_al_u681_o),
    .c(_al_u1342_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F9vpw6 ),
    .o(_al_u4306_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(D*~C*B))"),
    .INIT(16'h5155))
    _al_u4307 (
    .a(_al_u4306_o),
    .b(_al_u607_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B8bow6 ));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~C*~(~D*~A)))"),
    .INIT(16'hc0c4))
    _al_u4308 (
    .a(_al_u1643_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Obbow6_lutinv ),
    .c(_al_u604_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 ),
    .o(_al_u4308_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*A*~(D*C))"),
    .INIT(16'h0222))
    _al_u4309 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B8bow6 ),
    .b(_al_u4308_o),
    .c(_al_u3201_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kxziu6_lutinv ),
    .o(_al_u4309_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u431 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_raw_int [13]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inten_padded [13]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_masked_int [13]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u4310 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Apaiu6_lutinv ),
    .b(_al_u3917_o),
    .o(_al_u4310_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(B*~(C*~A)))"),
    .INIT(16'h7300))
    _al_u4311 (
    .a(_al_u4304_o),
    .b(_al_u4309_o),
    .c(_al_u4310_o),
    .d(_al_u696_o),
    .o(_al_u4311_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u4312 (
    .a(_al_u3211_o),
    .b(_al_u2770_o),
    .o(_al_u4312_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(~A*~(C*~B)))"),
    .INIT(16'hba00))
    _al_u4313 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qe8iu6_lutinv ),
    .b(_al_u1643_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U98iu6 ),
    .d(_al_u1817_o),
    .o(_al_u4313_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(~D*C*A))"),
    .INIT(16'h3313))
    _al_u4314 (
    .a(_al_u4312_o),
    .b(_al_u4313_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 ),
    .o(_al_u4314_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D*C*B))"),
    .INIT(16'h2aaa))
    _al_u4315 (
    .a(_al_u4314_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yv1ju6 ),
    .c(_al_u2364_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 ),
    .o(_al_u4315_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hd3df))
    _al_u4316 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cwiiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rwjax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6 ),
    .o(_al_u4316_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*~B*A)"),
    .INIT(16'h0020))
    _al_u4317 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vviiu6 ),
    .b(_al_u4316_o),
    .c(_al_u1269_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 ),
    .o(_al_u4317_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    _al_u4318 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jckax6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jgxpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N4kax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4jax6 ),
    .o(_al_u4318_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~A*~(D*B))"),
    .INIT(16'h0105))
    _al_u4319 (
    .a(_al_u4312_o),
    .b(_al_u3233_o),
    .c(_al_u4317_o),
    .d(_al_u4318_o),
    .o(_al_u4319_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*~(B)*C*D)"),
    .INIT(16'h25a1))
    _al_u432 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [14]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [14]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpol_padded [14]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_last_datain [14]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_raw_int [14]));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u4320 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Htyiu6 ),
    .b(_al_u2365_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv ),
    .o(_al_u4320_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D*C*A))"),
    .INIT(16'h1333))
    _al_u4321 (
    .a(_al_u3211_o),
    .b(_al_u4320_o),
    .c(_al_u2367_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rwjax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O4bow6 ));
  AL_MAP_LUT4 #(
    .EQN("(C*~(A*~(D*B)))"),
    .INIT(16'hd050))
    _al_u4322 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O4bow6 ),
    .b(_al_u3608_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4jax6 ),
    .o(_al_u4322_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*A*~(D*~B))"),
    .INIT(16'h080a))
    _al_u4323 (
    .a(_al_u4315_o),
    .b(_al_u4319_o),
    .c(_al_u4322_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Skjax6 ),
    .o(_al_u4323_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u4324 (
    .a(_al_u2371_o),
    .b(_al_u2380_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 ),
    .o(_al_u4324_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(~B*~(D*C)))"),
    .INIT(16'ha888))
    _al_u4325 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yo1ju6 ),
    .b(_al_u4324_o),
    .c(_al_u3902_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rwjax6 ),
    .o(_al_u4325_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(B*A))"),
    .INIT(8'h07))
    _al_u4326 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Frziu6_lutinv ),
    .b(_al_u1582_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D31ju6 ),
    .o(_al_u4326_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*~(D*C)))"),
    .INIT(16'ha222))
    _al_u4327 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qe8iu6_lutinv ),
    .b(_al_u4326_o),
    .c(_al_u1342_o),
    .d(_al_u2829_o),
    .o(_al_u4327_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(~D*~(C*~B)))"),
    .INIT(16'h5510))
    _al_u4328 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 ),
    .o(_al_u4328_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D*C*A))"),
    .INIT(16'h1333))
    _al_u4329 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ia8iu6_lutinv ),
    .b(_al_u4328_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Frziu6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujiu6 ),
    .o(_al_u4329_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u433 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_raw_int [14]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inten_padded [14]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_masked_int [14]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~A*~(D*~C))"),
    .INIT(16'h1011))
    _al_u4330 (
    .a(_al_u3205_o),
    .b(_al_u4327_o),
    .c(_al_u4329_o),
    .d(_al_u909_o),
    .o(_al_u4330_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(~A*~(D*B)))"),
    .INIT(16'h0e0a))
    _al_u4331 (
    .a(_al_u4016_o),
    .b(_al_u1806_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv ),
    .d(_al_u3124_o),
    .o(_al_u4331_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~A*~(D*C))"),
    .INIT(16'h0111))
    _al_u4332 (
    .a(_al_u3186_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ),
    .c(_al_u932_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pu1ju6_lutinv ),
    .o(_al_u4332_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(~D*C*B))"),
    .INIT(16'haa2a))
    _al_u4333 (
    .a(_al_u4332_o),
    .b(_al_u1346_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D31ju6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 ),
    .o(_al_u4333_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u4334 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L45iu6_lutinv ),
    .b(_al_u1269_o),
    .c(_al_u1342_o),
    .d(_al_u1344_o),
    .o(_al_u4334_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u4335 (
    .a(_al_u903_o),
    .b(_al_u1266_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gebow6_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u4336 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gebow6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pu1ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yi7ju6_lutinv ),
    .o(_al_u4336_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(D*C))"),
    .INIT(16'h0444))
    _al_u4337 (
    .a(_al_u4334_o),
    .b(_al_u4336_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nkaju6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 ),
    .o(_al_u4337_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u4338 (
    .a(_al_u4330_o),
    .b(_al_u4331_o),
    .c(_al_u4333_o),
    .d(_al_u4337_o),
    .o(_al_u4338_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(~D*C))"),
    .INIT(16'h4404))
    _al_u4339 (
    .a(_al_u4325_o),
    .b(_al_u4338_o),
    .c(_al_u3608_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N4kax6 ),
    .o(_al_u4339_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*~(B)*C*D)"),
    .INIT(16'h25a1))
    _al_u434 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [15]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [15]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpol_padded [15]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_last_datain [15]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_raw_int [15]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*C)*~(B*A))"),
    .INIT(16'h0777))
    _al_u4340 (
    .a(_al_u607_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D6kiu6_lutinv ),
    .c(_al_u1346_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jf6ju6 ),
    .o(_al_u4340_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C*~(~B*A)))"),
    .INIT(16'h2f00))
    _al_u4341 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I82ju6 ),
    .b(_al_u3109_o),
    .c(_al_u4340_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 ),
    .o(_al_u4341_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(~A*~(D*~B)))"),
    .INIT(16'hb0a0))
    _al_u4342 (
    .a(_al_u930_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vygax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 ),
    .o(_al_u4342_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u4343 (
    .a(_al_u4342_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yi7ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 ),
    .o(_al_u4343_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u4344 (
    .a(_al_u4343_o),
    .b(_al_u3624_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fpaow6_lutinv ),
    .o(_al_u4344_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(~A*~(~D*~B)))"),
    .INIT(16'ha0b0))
    _al_u4345 (
    .a(_al_u3085_o),
    .b(_al_u4344_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Llaow6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F9vpw6 ),
    .o(_al_u4345_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    _al_u4346 (
    .a(_al_u4323_o),
    .b(_al_u4339_o),
    .c(_al_u4341_o),
    .d(_al_u4345_o),
    .o(_al_u4346_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*C)*~(B*~A))"),
    .INIT(16'hbb0b))
    _al_u4347 (
    .a(_al_u4311_o),
    .b(_al_u4346_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vqohu6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u4348 (
    .a(_al_u4284_o),
    .b(_al_u1809_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aphiu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~C)*~(~B*~A))"),
    .INIT(16'he0ee))
    _al_u4349 (
    .a(_al_u4278_o),
    .b(_al_u4173_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U8jax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dgapw6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u435 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_raw_int [15]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inten_padded [15]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_masked_int [15]));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(~D*~B*~A))"),
    .INIT(16'h0f0e))
    _al_u4350 (
    .a(_al_u4170_o),
    .b(_al_u4173_o),
    .c(_al_u4168_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[0] ),
    .o(_al_u4350_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u4351 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N3ziu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv ),
    .o(_al_u4351_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*~B))"),
    .INIT(8'h8a))
    _al_u4352 (
    .a(_al_u4351_o),
    .b(_al_u678_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 ),
    .o(_al_u4352_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(~A*~(~D*B)))"),
    .INIT(16'ha0e0))
    _al_u4353 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bi0iu6 ),
    .b(_al_u903_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 ),
    .o(_al_u4353_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u4354 (
    .a(_al_u1784_o),
    .b(_al_u4352_o),
    .c(_al_u697_o),
    .d(_al_u4353_o),
    .o(_al_u4354_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*~A)"),
    .INIT(16'h4000))
    _al_u4355 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vygax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 ),
    .o(_al_u4355_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*A)"),
    .INIT(16'h0002))
    _al_u4356 (
    .a(_al_u4354_o),
    .b(_al_u4012_o),
    .c(_al_u4283_o),
    .d(_al_u4355_o),
    .o(_al_u4356_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*~A)"),
    .INIT(16'h0040))
    _al_u4357 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xq3pw6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I30ju6_lutinv ),
    .c(_al_u1271_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 ),
    .o(_al_u4357_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*~A))"),
    .INIT(8'h32))
    _al_u4358 (
    .a(_al_u1643_o),
    .b(_al_u1336_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ),
    .o(_al_u4358_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(C*A))"),
    .INIT(16'h5f13))
    _al_u4359 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L45iu6_lutinv ),
    .b(_al_u682_o),
    .c(_al_u1342_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 ),
    .o(_al_u4359_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*~(B)*C*D)"),
    .INIT(16'h25a1))
    _al_u436 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [2]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [2]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpol_padded [2]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_last_datain [2]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_raw_int [2]));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u4360 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N98iu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 ),
    .o(_al_u4360_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~A*~(~D*~B))"),
    .INIT(16'h0504))
    _al_u4361 (
    .a(_al_u3666_o),
    .b(_al_u4359_o),
    .c(_al_u4360_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 ),
    .o(_al_u4361_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(B*~(C*~A)))"),
    .INIT(16'h7300))
    _al_u4362 (
    .a(_al_u4358_o),
    .b(_al_u4361_o),
    .c(_al_u1806_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv ),
    .o(_al_u4362_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*C)*~(B*A))"),
    .INIT(16'h0777))
    _al_u4363 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zwcpw6_lutinv ),
    .b(_al_u607_o),
    .c(_al_u903_o),
    .d(_al_u2829_o),
    .o(_al_u4363_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(A*~(C*B)))"),
    .INIT(16'h00d5))
    _al_u4364 (
    .a(_al_u4363_o),
    .b(_al_u4161_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Daiax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 ),
    .o(_al_u4364_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*A)"),
    .INIT(16'h0002))
    _al_u4365 (
    .a(_al_u4356_o),
    .b(_al_u4357_o),
    .c(_al_u4362_o),
    .d(_al_u4364_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lrhiu6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u4366 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lrhiu6 ),
    .b(_al_u4151_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ueapw6 ));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B*~(D*~A)))"),
    .INIT(16'h7030))
    _al_u4367 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dgapw6 ),
    .b(_al_u4350_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ueapw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[0] ),
    .o(_al_u4367_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u4368 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aphiu6 ),
    .b(_al_u4367_o),
    .o(_al_u4368_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u4369 (
    .a(_al_u4368_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L18iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W7cow6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u437 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_raw_int [2]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inten_padded [2]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_masked_int [2]));
  AL_MAP_LUT2 #(
    .EQN("~(~B*A)"),
    .INIT(4'hd))
    _al_u4370 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W7cow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n3436 ));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u4371 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y40ju6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 ),
    .o(_al_u4371_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(D*~C*~A))"),
    .INIT(16'hc8cc))
    _al_u4372 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0biu6 ),
    .b(_al_u4371_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F9vpw6 ),
    .o(_al_u4372_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u4373 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N4kax6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4jax6 ),
    .o(_al_u4373_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u4374 (
    .a(_al_u3831_o),
    .b(_al_u4373_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6 ),
    .o(_al_u4374_o));
  AL_MAP_LUT4 #(
    .EQN("(A*(~(B)*~(C)*~(D)+~(B)*C*~(D)+B*C*~(D)+B*~(C)*D+B*C*D))"),
    .INIT(16'h88a2))
    _al_u4375 (
    .a(_al_u4374_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qxoiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gr2qw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 ),
    .o(_al_u4375_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u4376 (
    .a(_al_u3997_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jgxpw6 ),
    .o(_al_u4376_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(~B*~(C*~A)))"),
    .INIT(16'hdc00))
    _al_u4377 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wh0ju6 ),
    .b(_al_u4376_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P14qw6 ),
    .o(_al_u4377_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(~B*~(D*~A)))"),
    .INIT(16'hd0c0))
    _al_u4378 (
    .a(_al_u4375_o),
    .b(_al_u4377_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J9kiu6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Skjax6 ),
    .o(_al_u4378_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u4379 (
    .a(_al_u3246_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Skjax6 ),
    .o(_al_u4379_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*~(B)*C*D)"),
    .INIT(16'h25a1))
    _al_u438 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [3]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpol_padded [3]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_last_datain [3]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_raw_int [3]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    _al_u4380 (
    .a(_al_u604_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 ),
    .o(_al_u4380_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~A*~(~D*B))"),
    .INIT(16'h0501))
    _al_u4381 (
    .a(_al_u4379_o),
    .b(_al_u2772_o),
    .c(_al_u4380_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 ),
    .o(_al_u4381_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u4382 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yljiu6 ),
    .b(_al_u3122_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 ),
    .o(_al_u4382_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u4383 (
    .a(_al_u4382_o),
    .b(_al_u682_o),
    .c(_al_u696_o),
    .o(_al_u4383_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u4384 (
    .a(_al_u696_o),
    .b(_al_u2392_o),
    .c(_al_u2647_o),
    .o(_al_u4384_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*A*~(D*B))"),
    .INIT(16'h020a))
    _al_u4385 (
    .a(_al_u4383_o),
    .b(_al_u1812_o),
    .c(_al_u4384_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 ),
    .o(_al_u4385_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(~D*~(C@B)))"),
    .INIT(16'haa28))
    _al_u4386 (
    .a(_al_u3246_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N4kax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rwjax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6 ),
    .o(_al_u4386_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(D*~C*B))"),
    .INIT(16'h5155))
    _al_u4387 (
    .a(_al_u4386_o),
    .b(_al_u908_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nsaiu6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 ),
    .o(_al_u4387_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*~A)"),
    .INIT(16'h4000))
    _al_u4388 (
    .a(_al_u4378_o),
    .b(_al_u4381_o),
    .c(_al_u4385_o),
    .d(_al_u4387_o),
    .o(_al_u4388_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~B*~(~D*A))"),
    .INIT(16'h0301))
    _al_u4389 (
    .a(_al_u2369_o),
    .b(_al_u4007_o),
    .c(_al_u4373_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 ),
    .o(_al_u4389_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u439 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_raw_int [3]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inten_padded [3]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_masked_int [3]));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D*~(~C*B)))"),
    .INIT(16'h08aa))
    _al_u4390 (
    .a(_al_u4389_o),
    .b(_al_u2369_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dcziu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 ),
    .o(_al_u4390_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(A*~(D*~C)))"),
    .INIT(16'h4c44))
    _al_u4391 (
    .a(_al_u4390_o),
    .b(_al_u2386_o),
    .c(_al_u2380_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6 ),
    .o(_al_u4391_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u4392 (
    .a(_al_u912_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6 ),
    .o(_al_u4392_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u4393 (
    .a(_al_u2770_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 ),
    .o(_al_u4393_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u4394 (
    .a(_al_u4393_o),
    .b(_al_u2364_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nyiiu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ia0ju6 ));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(D*C))"),
    .INIT(16'h0444))
    _al_u4395 (
    .a(_al_u4392_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ia0ju6 ),
    .c(_al_u2371_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wa0ju6 ),
    .o(_al_u4395_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(~D*~(C*~B)))"),
    .INIT(16'haa20))
    _al_u4396 (
    .a(_al_u4388_o),
    .b(_al_u4391_o),
    .c(_al_u4395_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hgrpw6 ),
    .o(_al_u4396_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D*C*~B))"),
    .INIT(16'h8aaa))
    _al_u4397 (
    .a(_al_u4396_o),
    .b(_al_u3109_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mmjiu6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gebow6_lutinv ),
    .o(_al_u4397_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D*C*~B))"),
    .INIT(16'h8aaa))
    _al_u4398 (
    .a(_al_u4397_o),
    .b(_al_u3109_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ldoiu6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yljiu6 ),
    .o(_al_u4398_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(B*~(D*~A)))"),
    .INIT(16'h0703))
    _al_u4399 (
    .a(_al_u4372_o),
    .b(_al_u4398_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv ),
    .d(_al_u909_o),
    .o(_al_u4399_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*~(B)*C*D)"),
    .INIT(16'h25a1))
    _al_u440 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [4]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [4]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpol_padded [4]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_last_datain [4]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_raw_int [4]));
  AL_MAP_LUT4 #(
    .EQN("~((C*B)*~(A)*~(D)+(C*B)*A*~(D)+~((C*B))*A*D+(C*B)*A*D)"),
    .INIT(16'h553f))
    _al_u4400 (
    .a(_al_u3810_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ia8iu6_lutinv ),
    .c(_al_u909_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 ),
    .o(_al_u4400_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u4401 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yqziu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 ),
    .o(_al_u4401_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~D*~C*~A))"),
    .INIT(16'hccc8))
    _al_u4402 (
    .a(_al_u4401_o),
    .b(_al_u681_o),
    .c(_al_u3754_o),
    .d(_al_u909_o),
    .o(_al_u4402_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(D*~(~C*~B)))"),
    .INIT(16'h0155))
    _al_u4403 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ),
    .b(_al_u604_o),
    .c(_al_u679_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 ),
    .o(_al_u4403_o));
  AL_MAP_LUT4 #(
    .EQN("(C*A*~(D*B))"),
    .INIT(16'h20a0))
    _al_u4404 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F85iu6 ),
    .b(_al_u4161_o),
    .c(_al_u4403_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ),
    .o(_al_u4404_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(D*C))"),
    .INIT(16'h0444))
    _al_u4405 (
    .a(_al_u4402_o),
    .b(_al_u4404_o),
    .c(_al_u1643_o),
    .d(_al_u1635_o),
    .o(_al_u4405_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~A*~(D*C))"),
    .INIT(16'h0111))
    _al_u4406 (
    .a(_al_u912_o),
    .b(_al_u2386_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hgrpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 ),
    .o(_al_u4406_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u4407 (
    .a(_al_u909_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wkipw6 ),
    .o(_al_u4407_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u4408 (
    .a(_al_u3223_o),
    .b(_al_u4407_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9ypw6 ),
    .o(_al_u4408_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B*A))"),
    .INIT(8'h70))
    _al_u4409 (
    .a(_al_u4406_o),
    .b(_al_u4408_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kxziu6_lutinv ),
    .o(_al_u4409_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u441 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_raw_int [4]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inten_padded [4]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_masked_int [4]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u4410 (
    .a(_al_u2771_o),
    .b(_al_u2832_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Skjax6 ),
    .o(_al_u4410_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(~D*C))"),
    .INIT(16'h4404))
    _al_u4411 (
    .a(_al_u4409_o),
    .b(_al_u4410_o),
    .c(_al_u3574_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 ),
    .o(_al_u4411_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*~(~D*~A))"),
    .INIT(16'hc080))
    _al_u4412 (
    .a(_al_u4400_o),
    .b(_al_u4405_o),
    .c(_al_u4411_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hgrpw6 ),
    .o(_al_u4412_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D*~C*B))"),
    .INIT(16'ha2aa))
    _al_u4413 (
    .a(_al_u4412_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qe8iu6_lutinv ),
    .c(_al_u3109_o),
    .d(_al_u1266_o),
    .o(_al_u4413_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u4414 (
    .a(_al_u3109_o),
    .b(_al_u1775_o),
    .o(_al_u4414_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~(~B*~A))"),
    .INIT(16'he000))
    _al_u4415 (
    .a(_al_u1812_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 ),
    .o(_al_u4415_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D*~(~C*~B)))"),
    .INIT(16'h02aa))
    _al_u4416 (
    .a(_al_u4413_o),
    .b(_al_u4414_o),
    .c(_al_u4415_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 ),
    .o(_al_u4416_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*C)*~(B*~A))"),
    .INIT(16'hbb0b))
    _al_u4417 (
    .a(_al_u4399_o),
    .b(_al_u4416_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Axohu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*A)"),
    .INIT(16'h0002))
    _al_u4418 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lrhiu6 ),
    .b(_al_u3797_o),
    .c(_al_u1809_o),
    .d(_al_u3122_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S18iu6 ));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u4419 (
    .a(_al_u4368_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S18iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jxgax6 ),
    .o(_al_u4419_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*~(B)*C*D)"),
    .INIT(16'h25a1))
    _al_u442 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [5]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [5]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpol_padded [5]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_last_datain [5]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_raw_int [5]));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u4420 (
    .a(_al_u4419_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sqfax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uofax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xg6iu6 ));
  AL_MAP_LUT4 #(
    .EQN("(C*(D@B@A))"),
    .INIT(16'h9060))
    _al_u4421 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vtzhu6 ),
    .b(_al_u4278_o),
    .c(_al_u3797_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[1] ),
    .o(_al_u4421_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*B)*~(D*A))"),
    .INIT(16'h51f3))
    _al_u4422 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A3iiu6 ),
    .b(_al_u3808_o),
    .c(_al_u1581_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [3]),
    .o(_al_u4422_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u4423 (
    .a(_al_u4421_o),
    .b(_al_u4422_o),
    .o(_al_u4423_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4424 (
    .a(_al_u4049_o),
    .b(_al_u4048_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ud4iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xrxax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C4iiu6 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u4425 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ok8iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C4iiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[1] ),
    .o(_al_u4425_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u4426 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ql8iu6 ),
    .b(_al_u4425_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[2] ),
    .o(_al_u4426_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C*~A))"),
    .INIT(8'h73))
    _al_u4427 (
    .a(_al_u4423_o),
    .b(_al_u4426_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jl8iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Egthu6 ));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u4428 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xg6iu6 ),
    .b(_al_u4111_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H4ypw6 ),
    .o(\u_cmsdk_mcu/HADDR [10]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u4429 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xg6iu6 ),
    .b(_al_u4237_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yf1qw6 ),
    .o(\u_cmsdk_mcu/HADDR [9]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u443 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_raw_int [5]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inten_padded [5]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_masked_int [5]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u4430 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xg6iu6 ),
    .b(_al_u4106_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ke1qw6 ),
    .o(\u_cmsdk_mcu/HADDR [8]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u4431 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xg6iu6 ),
    .b(_al_u4121_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nd3qw6 ),
    .o(\u_cmsdk_mcu/HADDR [7]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u4432 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xg6iu6 ),
    .b(_al_u4141_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vn9bx6 ),
    .o(\u_cmsdk_mcu/HADDR [6]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u4433 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xg6iu6 ),
    .b(_al_u4219_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bf3qw6 ),
    .o(\u_cmsdk_mcu/HADDR [5]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u4434 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xg6iu6 ),
    .b(_al_u4231_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pg3qw6 ),
    .o(\u_cmsdk_mcu/HADDR [4]));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u4435 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iqzhu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J0gax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nmfax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wqzhu6 ));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    _al_u4436 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wqzhu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nrqpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P23qw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Am6iu6_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u4437 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xg6iu6 ),
    .b(_al_u4225_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Am6iu6_lutinv ),
    .o(\u_cmsdk_mcu/HADDR [3]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u4438 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wqzhu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gpqpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xn7ax6 ),
    .o(_al_u4438_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u4439 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xg6iu6 ),
    .b(_al_u4423_o),
    .c(_al_u4438_o),
    .o(\u_cmsdk_mcu/HADDR [2]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*~(B)*C*D)"),
    .INIT(16'h25a1))
    _al_u444 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [6]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [6]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpol_padded [6]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_last_datain [6]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_raw_int [6]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u4440 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xg6iu6 ),
    .b(_al_u4136_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ad7ax6 ),
    .o(\u_cmsdk_mcu/HADDR [15]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u4441 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xg6iu6 ),
    .b(_al_u4131_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvabx6 ),
    .o(\u_cmsdk_mcu/HADDR [14]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u4442 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xg6iu6 ),
    .b(_al_u4126_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kl8ax6 ),
    .o(\u_cmsdk_mcu/HADDR [13]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u4443 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xg6iu6 ),
    .b(_al_u4035_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Su8ax6 ),
    .o(\u_cmsdk_mcu/HADDR [12]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u4444 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xg6iu6 ),
    .b(_al_u4116_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B79bx6 ),
    .o(\u_cmsdk_mcu/HADDR [11]));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*~B))"),
    .INIT(8'h54))
    _al_u4445 (
    .a(_al_u4368_o),
    .b(_al_u3797_o),
    .c(_al_u1888_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jc3pw6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u4446 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wqzhu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dugax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qc3pw6_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u4447 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xg6iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jc3pw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qc3pw6_lutinv ),
    .o(\u_cmsdk_mcu/HSIZE [1]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u4448 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iqzhu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gnqpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sq4iu6 ));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'h4e))
    _al_u4449 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xg6iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fnpiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sq4iu6 ),
    .o(\u_cmsdk_mcu/HWRITE ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u445 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_raw_int [6]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inten_padded [6]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_masked_int [6]));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*~A)"),
    .INIT(16'h0040))
    _al_u4450 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fm7ax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gr2qw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Isjpw6 ),
    .o(_al_u4450_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(~C*~B*A))"),
    .INIT(16'hfd00))
    _al_u4451 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zrhiu6_lutinv ),
    .b(_al_u1777_o),
    .c(_al_u3925_o),
    .d(_al_u4450_o),
    .o(_al_u4451_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(D*C*B))"),
    .INIT(16'h1555))
    _al_u4452 (
    .a(_al_u4451_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tu4iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O34iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I4rpw6 ),
    .o(_al_u4452_o));
  AL_MAP_LUT4 #(
    .EQN("~(A*~(D*~(C*B)))"),
    .INIT(16'h7f55))
    _al_u4453 (
    .a(_al_u4452_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Scbiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T24iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lmkbx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pfphu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4454 (
    .a(_al_u4049_o),
    .b(_al_u4048_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O34iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nu5bx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xfliu6 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u4455 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ok8iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xfliu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[0] ),
    .o(_al_u4455_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u4456 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ql8iu6 ),
    .b(_al_u4455_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[1] ),
    .o(_al_u4456_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u4457 (
    .a(_al_u2364_o),
    .b(_al_u2367_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 ),
    .o(_al_u4457_o));
  AL_MAP_LUT4 #(
    .EQN("~(B*~(D*C*A))"),
    .INIT(16'hb333))
    _al_u4458 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iiliu6 ),
    .b(_al_u4456_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jl8iu6 ),
    .d(_al_u4457_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Irrhu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*B)*~(~D*A))"),
    .INIT(16'hf351))
    _al_u4459 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R2phu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bxdpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Us3bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z71bx6 ),
    .o(_al_u4459_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*~(B)*C*D)"),
    .INIT(16'h25a1))
    _al_u446 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [7]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [7]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpol_padded [7]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_last_datain [7]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_raw_int [7]));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*B)*~(~D*A))"),
    .INIT(16'hf351))
    _al_u4460 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W1phu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U0phu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V52bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yxrpw6 ),
    .o(_al_u4460_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*B)*~(~D*A))"),
    .INIT(16'hf351))
    _al_u4461 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Szohu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gwdpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rm2bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xq2bx6 ),
    .o(_al_u4461_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*B)*~(~D*A))"),
    .INIT(16'hf351))
    _al_u4462 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B1phu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nwdpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dv2bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P12bx6 ),
    .o(_al_u4462_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u4463 (
    .a(_al_u4459_o),
    .b(_al_u4460_o),
    .c(_al_u4461_o),
    .d(_al_u4462_o),
    .o(_al_u4463_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(~C*A))"),
    .INIT(16'hf531))
    _al_u4464 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F3phu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zzohu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fc1bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y0gbx6 ),
    .o(_al_u4464_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(~C*A))"),
    .INIT(16'hf531))
    _al_u4465 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N0phu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G0phu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fe2bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Li2bx6 ),
    .o(_al_u4465_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u4466 (
    .a(_al_u4463_o),
    .b(_al_u4464_o),
    .c(_al_u4465_o),
    .o(_al_u4466_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*~B))"),
    .INIT(8'ha8))
    _al_u4467 (
    .a(_al_u4466_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Li5iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T8kbx6 ),
    .o(_al_u4467_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*~B)*~(~D*A))"),
    .INIT(16'hfc54))
    _al_u4468 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jyohu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qh5iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F17ax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tcipw6 ),
    .o(_al_u4468_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(~C*A))"),
    .INIT(16'hf531))
    _al_u4469 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H4phu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A4phu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gihbx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mk3bx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ux5iu6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u447 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_raw_int [7]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inten_padded [7]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_masked_int [7]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*A))"),
    .INIT(8'hc4))
    _al_u4470 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M3phu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ux5iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qo3bx6 ),
    .o(_al_u4470_o));
  AL_MAP_LUT4 #(
    .EQN("(C*A*~(~D*B))"),
    .INIT(16'ha020))
    _al_u4471 (
    .a(_al_u4468_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cyohu6 ),
    .c(_al_u4470_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hg3bx6 ),
    .o(_al_u4471_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*B)*~(~D*A))"),
    .INIT(16'hf351))
    _al_u4472 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T3phu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I1phu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dt1bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lr9bx6 ),
    .o(_al_u4472_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*~A)"),
    .INIT(8'h04))
    _al_u4473 (
    .a(_al_u2733_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ch5iu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mnmpw6 ),
    .o(_al_u4473_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u4474 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J5phu6 ),
    .b(_al_u4473_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U31bx6 ),
    .o(_al_u4474_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*B)*~(~D*~A))"),
    .INIT(16'hf3a2))
    _al_u4475 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ag5iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P1phu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jx1bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zdtpw6 ),
    .o(_al_u4475_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(~D*C))"),
    .INIT(16'h8808))
    _al_u4476 (
    .a(_al_u4474_o),
    .b(_al_u4475_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C5phu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aa2bx6 ),
    .o(_al_u4476_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(~C*A))"),
    .INIT(16'hf531))
    _al_u4477 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O4phu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V4phu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Muhbx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5bbx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O16iu6 ));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u4478 (
    .a(_al_u4472_o),
    .b(_al_u4476_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O16iu6 ),
    .o(_al_u4478_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(~C*A))"),
    .INIT(16'hf531))
    _al_u4479 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K2phu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D2phu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rk1bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xo1bx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vu5iu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*~(B)*C*D)"),
    .INIT(16'h25a1))
    _al_u448 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [8]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [8]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpol_padded [8]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_last_datain [8]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_raw_int [8]));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(~C*A))"),
    .INIT(16'hf531))
    _al_u4480 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y2phu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uwdpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lg1bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rijbx6 ),
    .o(_al_u4480_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u4481 (
    .a(_al_u4471_o),
    .b(_al_u4478_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vu5iu6 ),
    .d(_al_u4480_o),
    .o(_al_u4481_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(~C*A))"),
    .INIT(16'hf531))
    _al_u4482 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lzohu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ezohu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jz2bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P33bx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zi5iu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*B)*~(~D*A))"),
    .INIT(16'hf351))
    _al_u4483 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xyohu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qyohu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bc3bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V73bx6 ),
    .o(_al_u4483_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u4484 (
    .a(_al_u4467_o),
    .b(_al_u4481_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zi5iu6 ),
    .d(_al_u4483_o),
    .o(_al_u4484_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(A*~(~D*B)))"),
    .INIT(16'h50d0))
    _al_u4485 (
    .a(_al_u4484_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Npghu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kqhbx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pdyax6 ),
    .o(_al_u4485_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u4486 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N98iu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 ),
    .o(_al_u4486_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~B*~(C*A))"),
    .INIT(16'h0013))
    _al_u4487 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zwcpw6_lutinv ),
    .b(_al_u3925_o),
    .c(_al_u4486_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z9opw6 ),
    .o(_al_u4487_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*B*~A)"),
    .INIT(16'h0400))
    _al_u4488 (
    .a(_al_u4485_o),
    .b(_al_u1299_o),
    .c(_al_u1777_o),
    .d(_al_u4487_o),
    .o(_al_u4488_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(D*C*B))"),
    .INIT(16'h1555))
    _al_u4489 (
    .a(_al_u4488_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qa5iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ja5iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z9opw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J4xhu6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u449 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_raw_int [8]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inten_padded [8]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_masked_int [8]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*~A))"),
    .INIT(8'h32))
    _al_u4490 (
    .a(_al_u4419_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wvgax6 ),
    .o(_al_u4490_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u4491 (
    .a(_al_u4490_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sqfax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uofax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tszhu6 ));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u4492 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iqzhu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gpqpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nrqpw6 ),
    .o(_al_u4492_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u4493 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wqzhu6 ),
    .b(_al_u4492_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J0gax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bqzhu6_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u4494 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tszhu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bqzhu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n265 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sf1iu6 ));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u4495 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cq3qw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vqgax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wc2qw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydgax6 ),
    .o(_al_u4495_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u4496 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xg6iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ),
    .c(_al_u4495_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nr4iu6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*B)*~(C)*~(A)+~(D*B)*C*~(A)+~(~(D*B))*C*A+~(D*B)*C*A)"),
    .INIT(16'h4e0a))
    _al_u4497 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nr4iu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ur4iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sq4iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dg2qw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G6xhu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(~D*~(C*A)))"),
    .INIT(16'h3320))
    _al_u4498 (
    .a(_al_u4171_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U8jax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hphiu6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*A)"),
    .INIT(16'h0200))
    _al_u4499 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hphiu6_lutinv ),
    .b(_al_u4173_o),
    .c(_al_u4168_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ueapw6 ),
    .o(_al_u4499_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*~(B)*C*D)"),
    .INIT(16'h25a1))
    _al_u450 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [9]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [9]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpol_padded [9]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_last_datain [9]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_raw_int [9]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u4500 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aphiu6 ),
    .b(_al_u4499_o),
    .o(_al_u4500_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u4501 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/HALTED ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jcpow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rzciu6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C1wpw6 ),
    .o(_al_u4501_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u4502 (
    .a(_al_u4500_o),
    .b(_al_u4501_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R05iu6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u4503 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R05iu6 ),
    .b(_al_u1299_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vihiu6_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u4504 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vihiu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X7ypw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A25iu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4505 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A25iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R05iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E6iax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uu8iu6 ));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u4506 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vihiu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[0] ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pz4iu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(A*~(~D*B)))"),
    .INIT(16'h050d))
    _al_u4507 (
    .a(_al_u4170_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[0] ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U8jax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X7ypw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ekhiu6_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u4508 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vihiu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ekhiu6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uy4iu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u4509 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pz4iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uy4iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rw8iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Swjbx6 ),
    .o(_al_u4509_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u451 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_raw_int [9]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inten_padded [9]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_masked_int [9]));
  AL_MAP_LUT4 #(
    .EQN("(C*A*~(~D*B))"),
    .INIT(16'ha020))
    _al_u4510 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vihiu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[0] ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U8jax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M15iu6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u4511 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/mux4_b10_sel_is_4_o ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [5]),
    .o(_al_u4511_o));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u4512 (
    .a(_al_u1986_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inten_padded [14]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttype_padded [14]),
    .o(_al_u4512_o));
  AL_MAP_LUT4 #(
    .EQN("~(C*~((D*~A))*~(B)+C*(D*~A)*~(B)+~(C)*(D*~A)*B+C*(D*~A)*B)"),
    .INIT(16'h8bcf))
    _al_u4513 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpol_padded [14]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [14]),
    .o(_al_u4513_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u4514 (
    .a(_al_u4512_o),
    .b(_al_u1982_o),
    .c(_al_u4513_o),
    .o(_al_u4514_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u4515 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .o(_al_u4515_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u4516 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4]),
    .c(\u_cmsdk_mcu/p0_outen [14]),
    .d(\u_cmsdk_mcu/p0_altfunc [14]),
    .o(_al_u4516_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D*~C*A))"),
    .INIT(16'h3133))
    _al_u4517 (
    .a(_al_u4515_o),
    .b(_al_u4516_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4]),
    .d(\u_cmsdk_mcu/p0_out [14]),
    .o(_al_u4517_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*~(~D*~C)))"),
    .INIT(16'h222a))
    _al_u4518 (
    .a(_al_u4511_o),
    .b(_al_u4514_o),
    .c(_al_u4517_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [5]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n31 [14]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u4519 (
    .a(_al_u1986_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inten_padded [14]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [14]),
    .o(_al_u4519_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u452 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_tick_cnt [2]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_tick_cnt [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/BAUDTICK ),
    .o(_al_u452_o));
  AL_MAP_LUT4 #(
    .EQN("~(C*~((D*~A))*~(B)+C*(D*~A)*~(B)+~(C)*(D*~A)*B+C*(D*~A)*B)"),
    .INIT(16'h8bcf))
    _al_u4520 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpol_padded [14]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[14] ),
    .o(_al_u4520_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u4521 (
    .a(_al_u4519_o),
    .b(_al_u1982_o),
    .c(_al_u4520_o),
    .o(_al_u4521_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h3210))
    _al_u4522 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [14]),
    .d(\u_cmsdk_mcu/p1_out [14]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/mux0_b14/B1_0 ));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u4523 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4]),
    .c(\u_cmsdk_mcu/p1_outen [14]),
    .d(\u_cmsdk_mcu/p1_altfunc [14]),
    .o(_al_u4523_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(~B*~(~C*A)))"),
    .INIT(16'h00ce))
    _al_u4524 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/mux0_b14/B1_0 ),
    .b(_al_u4523_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [5]),
    .o(_al_u4524_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*~A)"),
    .INIT(16'h4000))
    _al_u4525 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [10]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [11]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [8]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [14]),
    .o(_al_u4525_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(A*~(~C*B)))"),
    .INIT(16'h005d))
    _al_u4526 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/mux4_b10_sel_is_4_o ),
    .b(_al_u4521_o),
    .c(_al_u4524_o),
    .d(_al_u4525_o),
    .o(_al_u4526_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4527 (
    .a(\u_cmsdk_mcu/sram_hrdata [14]),
    .b(\u_cmsdk_mcu/flash_hrdata [14]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [0]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [1]),
    .o(_al_u4527_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(D*C))"),
    .INIT(16'h0444))
    _al_u4528 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n37 [14]),
    .b(_al_u4527_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [4]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/rwdata_reg [14]),
    .o(_al_u4528_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*~(D*~B))"),
    .INIT(16'h4050))
    _al_u4529 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n31 [14]),
    .b(_al_u4526_o),
    .c(_al_u4528_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [6]),
    .o(_al_u4529_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u453 (
    .a(_al_u452_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_tick_cnt [0]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_tick_cnt [1]),
    .o(_al_u453_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(B*~A))"),
    .INIT(8'h0b))
    _al_u4530 (
    .a(_al_u4529_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vobiu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jvvpw6 ),
    .o(_al_u4530_o));
  AL_MAP_LUT4 #(
    .EQN("~(B*A*~(~D*C))"),
    .INIT(16'h77f7))
    _al_u4531 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uu8iu6 ),
    .b(_al_u4509_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M15iu6 ),
    .d(_al_u4530_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gfvhu6 ));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*~A))"),
    .INIT(8'h23))
    _al_u4532 (
    .a(_al_u4500_o),
    .b(_al_u4501_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hgrpw6 ),
    .o(_al_u4532_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u4533 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vobiu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jvvpw6 ),
    .o(_al_u4533_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*A))"),
    .INIT(8'hc4))
    _al_u4534 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M15iu6 ),
    .b(_al_u4532_o),
    .c(_al_u4533_o),
    .o(_al_u4534_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u4535 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pz4iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uy4iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wz4iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tajax6 ),
    .o(_al_u4535_o));
  AL_MAP_LUT4 #(
    .EQN("~(B*A*~(D*C))"),
    .INIT(16'hf777))
    _al_u4536 (
    .a(_al_u4534_o),
    .b(_al_u4535_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A25iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L4lax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X4xhu6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u4537 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bqzhu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iqzhu6_lutinv ),
    .o(_al_u4537_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u4538 (
    .a(_al_u4490_o),
    .b(_al_u4537_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sqfax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uofax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pkhpw6 [1]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u4539 (
    .a(_al_u4368_o),
    .b(_al_u1888_o),
    .o(_al_u4539_o));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~B*~A)"),
    .INIT(8'hfe))
    _al_u454 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n53 ),
    .b(_al_u453_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_ctrl [6]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_state_inc ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u4540 (
    .a(_al_u4539_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iiliu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hz0iu6 ));
  AL_MAP_LUT4 #(
    .EQN("(B*~((D*C))*~(A)+B*(D*C)*~(A)+~(B)*(D*C)*A+B*(D*C)*A)"),
    .INIT(16'he444))
    _al_u4541 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xg6iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hz0iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qc3pw6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vj3qw6 ),
    .o(\u_cmsdk_mcu/HADDR [1]));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u4542 (
    .a(_al_u4539_o),
    .b(_al_u3797_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qk9pw6_lutinv ),
    .o(_al_u4542_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~((D*~C))*~(A)+B*(D*~C)*~(A)+~(B)*(D*~C)*A+B*(D*~C)*A)"),
    .INIT(16'h4e44))
    _al_u4543 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xg6iu6 ),
    .b(_al_u4542_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wqzhu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ksgax6 ),
    .o(\u_cmsdk_mcu/HSIZE [0]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u4544 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xg6iu6 ),
    .b(_al_u3887_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydgax6 ),
    .o(_al_u4544_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u4545 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xg6iu6 ),
    .b(_al_u4197_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vqgax6 ),
    .o(_al_u4545_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u4546 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xg6iu6 ),
    .b(_al_u3885_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cq3qw6 ),
    .o(_al_u4546_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u4547 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xg6iu6 ),
    .b(_al_u4101_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q4dbx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/HADDR[27]_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u4548 (
    .a(_al_u4544_o),
    .b(_al_u4545_o),
    .c(_al_u4546_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/HADDR[27]_lutinv ),
    .o(_al_u4548_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u4549 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nlcbx6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/No3qw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q2ibx6 ),
    .o(_al_u4549_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B)*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hdf0a))
    _al_u455 (
    .a(_al_u379_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_state [0]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_state [1]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_shift_buf [0]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_txd ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*B))"),
    .INIT(8'ha2))
    _al_u4550 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xg6iu6 ),
    .b(_al_u4549_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H7hbx6 ),
    .o(_al_u4550_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u4551 (
    .a(_al_u4096_o),
    .b(_al_u4184_o),
    .c(_al_u4191_o),
    .o(_al_u4551_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(~B*~(D*C)))"),
    .INIT(16'h5444))
    _al_u4552 (
    .a(_al_u4550_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xg6iu6 ),
    .c(_al_u4551_o),
    .d(_al_u4091_o),
    .o(_al_u4552_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u4553 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xg6iu6 ),
    .b(_al_u3889_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wc2qw6 ),
    .o(_al_u4553_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u4554 (
    .a(_al_u4548_o),
    .b(_al_u4552_o),
    .c(_al_u4553_o),
    .o(\u_cmsdk_mcu/flash_hsel ));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u4555 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pz4iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wz4iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kq7iu6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u4556 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M15iu6 ),
    .b(_al_u4533_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pp7iu6 ));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u4557 (
    .a(_al_u1986_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inten_padded [1]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttype_padded [1]),
    .o(_al_u4557_o));
  AL_MAP_LUT4 #(
    .EQN("~(C*~((D*~A))*~(B)+C*(D*~A)*~(B)+~(C)*(D*~A)*B+C*(D*~A)*B)"),
    .INIT(16'h8bcf))
    _al_u4558 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpol_padded [1]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [1]),
    .o(_al_u4558_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u4559 (
    .a(_al_u4557_o),
    .b(_al_u1982_o),
    .c(_al_u4558_o),
    .o(_al_u4559_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u456 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/state_reg [1]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/state_reg [2]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/i_paddr [15]),
    .o(_al_u456_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u4560 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4]),
    .c(\u_cmsdk_mcu/p0_outen [1]),
    .d(\u_cmsdk_mcu/p0_altfunc [1]),
    .o(_al_u4560_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D*~C*A))"),
    .INIT(16'h3133))
    _al_u4561 (
    .a(_al_u4515_o),
    .b(_al_u4560_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4]),
    .d(\u_cmsdk_mcu/p0_out [1]),
    .o(_al_u4561_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*~(~D*~C)))"),
    .INIT(16'h222a))
    _al_u4562 (
    .a(_al_u4511_o),
    .b(_al_u4559_o),
    .c(_al_u4561_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [5]),
    .o(_al_u4562_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4563 (
    .a(\u_cmsdk_mcu/sram_hrdata [1]),
    .b(\u_cmsdk_mcu/flash_hrdata [1]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [0]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [1]),
    .o(_al_u4563_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(D*C))"),
    .INIT(16'h0444))
    _al_u4564 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n37 [1]),
    .b(_al_u4563_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [4]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/rwdata_reg [1]),
    .o(_al_u4564_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u4565 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [6]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [7]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [8]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [9]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n12_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u4566 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [10]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [11]),
    .o(_al_u4566_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u4567 (
    .a(_al_u1988_o),
    .b(_al_u1986_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n12_lutinv ),
    .d(_al_u4566_o),
    .o(_al_u4567_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(D*C))"),
    .INIT(16'h0444))
    _al_u4568 (
    .a(_al_u4562_o),
    .b(_al_u4564_o),
    .c(_al_u4567_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [5]),
    .o(_al_u4568_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u4569 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [8]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [9]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [10]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [11]),
    .o(_al_u4569_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*A)"),
    .INIT(16'h0200))
    _al_u457 (
    .a(_al_u456_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/i_paddr [12]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/i_paddr [13]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/i_paddr [14]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_apb_slave_mux/n4 ));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u4570 (
    .a(_al_u4569_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [6]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [7]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/mux6_b3_sel_is_2_o ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4571 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/n34_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/mux6_b3_sel_is_2_o ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/n19 [1]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_resetinfo [1]),
    .o(_al_u4571_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h3210))
    _al_u4572 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [1]),
    .d(\u_cmsdk_mcu/p1_out [1]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/mux0_b1/B1_0 ));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u4573 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4]),
    .c(\u_cmsdk_mcu/p1_outen [1]),
    .d(\u_cmsdk_mcu/p1_altfunc [1]),
    .o(_al_u4573_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(~B*~(~C*A)))"),
    .INIT(16'h00ce))
    _al_u4574 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/mux0_b1/B1_0 ),
    .b(_al_u4573_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [5]),
    .o(_al_u4574_o));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u4575 (
    .a(_al_u1986_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inten_padded [1]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [1]),
    .o(_al_u4575_o));
  AL_MAP_LUT4 #(
    .EQN("~(C*~((D*~A))*~(B)+C*(D*~A)*~(B)+~(C)*(D*~A)*B+C*(D*~A)*B)"),
    .INIT(16'h8bcf))
    _al_u4576 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpol_padded [1]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[1] ),
    .o(_al_u4576_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~A*~(~D*C))"),
    .INIT(16'h1101))
    _al_u4577 (
    .a(_al_u4574_o),
    .b(_al_u4575_o),
    .c(_al_u1982_o),
    .d(_al_u4576_o),
    .o(_al_u4577_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(D*C*B))"),
    .INIT(16'h1555))
    _al_u4578 (
    .a(_al_u4567_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n26_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [1]),
    .o(_al_u4578_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C*~(~B*A)))"),
    .INIT(16'h2f00))
    _al_u4579 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/mux4_b10_sel_is_4_o ),
    .b(_al_u4577_o),
    .c(_al_u4578_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [6]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n33 [1]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u458 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_apb_slave_mux/n4 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PWRITE ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/read_enable ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u4580 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [7]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_read_enable ),
    .o(_al_u4580_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*A*~(D*~B))"),
    .INIT(16'h080a))
    _al_u4581 (
    .a(_al_u4568_o),
    .b(_al_u4571_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n33 [1]),
    .d(_al_u4580_o),
    .o(_al_u4581_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*B)*~(~D*A))"),
    .INIT(16'hf351))
    _al_u4582 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kq7iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pp7iu6 ),
    .c(_al_u4581_o),
    .d(_al_u1833_o),
    .o(_al_u4582_o));
  AL_MAP_LUT4 #(
    .EQN("~((D*~A)*~(C)*~(B)+(D*~A)*C*~(B)+~((D*~A))*C*B+(D*~A)*C*B)"),
    .INIT(16'h2e3f))
    _al_u4583 (
    .a(_al_u4500_o),
    .b(_al_u4501_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O34iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S7mpw6 ),
    .o(_al_u4583_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u4584 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uy4iu6 ),
    .b(_al_u4583_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tujbx6 ),
    .o(_al_u4584_o));
  AL_MAP_LUT4 #(
    .EQN("~(B*A*~(D*C))"),
    .INIT(16'hf777))
    _al_u4585 (
    .a(_al_u4582_o),
    .b(_al_u4584_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A25iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T5mpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nhthu6 ));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u4586 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n12_lutinv ),
    .b(_al_u4566_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n13 [2]),
    .o(_al_u4586_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u4587 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n26_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [2]),
    .o(_al_u4587_o));
  AL_MAP_LUT4 #(
    .EQN("~(C*~((D*~A))*~(B)+C*(D*~A)*~(B)+~(C)*(D*~A)*B+C*(D*~A)*B)"),
    .INIT(16'h8bcf))
    _al_u4588 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpol_padded [2]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[2] ),
    .o(_al_u4588_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~B*~(~D*A))"),
    .INIT(16'h0301))
    _al_u4589 (
    .a(_al_u1983_o),
    .b(_al_u4586_o),
    .c(_al_u4587_o),
    .d(_al_u4588_o),
    .o(_al_u4589_o));
  AL_MAP_LUT4 #(
    .EQN("(D*A*(C@B))"),
    .INIT(16'h2800))
    _al_u459 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [4]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/state_reg [0]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/state_reg [1]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/state_reg [2]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n43 ));
  AL_MAP_LUT4 #(
    .EQN("(~B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h3210))
    _al_u4590 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [2]),
    .d(\u_cmsdk_mcu/p1_out [2]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/mux0_b2/B1_0 ));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u4591 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4]),
    .c(\u_cmsdk_mcu/p1_outen [2]),
    .d(\u_cmsdk_mcu/p1_altfunc [2]),
    .o(_al_u4591_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(~B*~(~C*A)))"),
    .INIT(16'h00ce))
    _al_u4592 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/mux0_b2/B1_0 ),
    .b(_al_u4591_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [5]),
    .o(_al_u4592_o));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u4593 (
    .a(_al_u1986_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inten_padded [2]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [2]),
    .o(_al_u4593_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*~(~D*~C)))"),
    .INIT(16'h222a))
    _al_u4594 (
    .a(_al_u4589_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/mux4_b10_sel_is_4_o ),
    .c(_al_u4592_o),
    .d(_al_u4593_o),
    .o(_al_u4594_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4595 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/n34_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/mux6_b3_sel_is_2_o ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/n19 [2]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_resetinfo [2]),
    .o(_al_u4595_o));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u4596 (
    .a(_al_u1986_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inten_padded [2]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttype_padded [2]),
    .o(_al_u4596_o));
  AL_MAP_LUT4 #(
    .EQN("~(C*~((D*~A))*~(B)+C*(D*~A)*~(B)+~(C)*(D*~A)*B+C*(D*~A)*B)"),
    .INIT(16'h8bcf))
    _al_u4597 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpol_padded [2]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [2]),
    .o(_al_u4597_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u4598 (
    .a(_al_u4596_o),
    .b(_al_u1982_o),
    .c(_al_u4597_o),
    .o(_al_u4598_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u4599 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4]),
    .c(\u_cmsdk_mcu/p0_outen [2]),
    .d(\u_cmsdk_mcu/p0_altfunc [2]),
    .o(_al_u4599_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u460 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n43 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wvgax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lf1iu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D*~C*A))"),
    .INIT(16'h3133))
    _al_u4600 (
    .a(_al_u4515_o),
    .b(_al_u4599_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4]),
    .d(\u_cmsdk_mcu/p0_out [2]),
    .o(_al_u4600_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*~(~D*~C)))"),
    .INIT(16'h222a))
    _al_u4601 (
    .a(_al_u4511_o),
    .b(_al_u4598_o),
    .c(_al_u4600_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [5]),
    .o(_al_u4601_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u4602 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/haddr_reg [7]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/haddr_reg [8]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/haddr_reg [9]),
    .o(_al_u4602_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u4603 (
    .a(_al_u4602_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/haddr_reg [5]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/haddr_reg [6]),
    .o(_al_u4603_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u4604 (
    .a(_al_u4603_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/haddr_reg [0]),
    .o(_al_u4604_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u4605 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [8]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/haddr_reg [2]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/haddr_reg [3]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/haddr_reg [4]),
    .o(_al_u4605_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u4606 (
    .a(_al_u4604_o),
    .b(_al_u4605_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n37 [2]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*C)*~(B*A))"),
    .INIT(16'h0777))
    _al_u4607 (
    .a(\u_cmsdk_mcu/sram_hrdata [2]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [1]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [4]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/rwdata_reg [2]),
    .o(_al_u4607_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u4608 (
    .a(_al_u4607_o),
    .b(\u_cmsdk_mcu/flash_hrdata [2]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [0]),
    .o(_al_u4608_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*~(D*B))"),
    .INIT(16'h1050))
    _al_u4609 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n37 [2]),
    .b(_al_u4586_o),
    .c(_al_u4608_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [5]),
    .o(_al_u4609_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u461 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n43 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wvgax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V3xhu6 ));
  AL_MAP_LUT4 #(
    .EQN("(C*~B*~(D*~A))"),
    .INIT(16'h2030))
    _al_u4610 (
    .a(_al_u4595_o),
    .b(_al_u4601_o),
    .c(_al_u4609_o),
    .d(_al_u4580_o),
    .o(_al_u4610_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*~A))"),
    .INIT(8'h8c))
    _al_u4611 (
    .a(_al_u4594_o),
    .b(_al_u4610_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [6]),
    .o(_al_u4611_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*B)*~(~D*A))"),
    .INIT(16'hf351))
    _al_u4612 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kq7iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pp7iu6 ),
    .c(_al_u4611_o),
    .d(_al_u1836_o),
    .o(_al_u4612_o));
  AL_MAP_LUT4 #(
    .EQN("~((D*~A)*~(C)*~(B)+(D*~A)*C*~(B)+~((D*~A))*C*B+(D*~A)*C*B)"),
    .INIT(16'h2e3f))
    _al_u4613 (
    .a(_al_u4500_o),
    .b(_al_u4501_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ud4iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Irmpw6 ),
    .o(_al_u4613_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u4614 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A25iu6 ),
    .b(_al_u4613_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jpmpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uehiu6 ));
  AL_MAP_LUT4 #(
    .EQN("~(B*A*~(D*C))"),
    .INIT(16'hf777))
    _al_u4615 (
    .a(_al_u4612_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uehiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uy4iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Usjbx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uhthu6 ));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u4616 (
    .a(_al_u1986_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inten_padded [3]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttype_padded [3]),
    .o(_al_u4616_o));
  AL_MAP_LUT4 #(
    .EQN("~(C*~((D*~A))*~(B)+C*(D*~A)*~(B)+~(C)*(D*~A)*B+C*(D*~A)*B)"),
    .INIT(16'h8bcf))
    _al_u4617 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpol_padded [3]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [3]),
    .o(_al_u4617_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u4618 (
    .a(_al_u4616_o),
    .b(_al_u1982_o),
    .c(_al_u4617_o),
    .o(_al_u4618_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u4619 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4]),
    .c(\u_cmsdk_mcu/p0_outen [3]),
    .d(\u_cmsdk_mcu/p0_altfunc [3]),
    .o(_al_u4619_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u462 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[9] ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[10] ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[11] ),
    .o(_al_u462_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D*~C*A))"),
    .INIT(16'h3133))
    _al_u4620 (
    .a(_al_u4515_o),
    .b(_al_u4619_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4]),
    .d(\u_cmsdk_mcu/p0_out [3]),
    .o(_al_u4620_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*~(~D*~C)))"),
    .INIT(16'h222a))
    _al_u4621 (
    .a(_al_u4511_o),
    .b(_al_u4618_o),
    .c(_al_u4620_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [5]),
    .o(_al_u4621_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h3210))
    _al_u4622 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [3]),
    .d(\u_cmsdk_mcu/p1_out [3]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/mux0_b3/B1_0 ));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u4623 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4]),
    .c(\u_cmsdk_mcu/p1_outen [3]),
    .d(\u_cmsdk_mcu/p1_altfunc [3]),
    .o(_al_u4623_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(~B*~(~C*A)))"),
    .INIT(16'h00ce))
    _al_u4624 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/mux0_b3/B1_0 ),
    .b(_al_u4623_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [5]),
    .o(_al_u4624_o));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u4625 (
    .a(_al_u1986_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inten_padded [3]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [3]),
    .o(_al_u4625_o));
  AL_MAP_LUT4 #(
    .EQN("~(C*~((D*~A))*~(B)+C*(D*~A)*~(B)+~(C)*(D*~A)*B+C*(D*~A)*B)"),
    .INIT(16'h8bcf))
    _al_u4626 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpol_padded [3]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[3] ),
    .o(_al_u4626_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~A*~(~D*C))"),
    .INIT(16'h1101))
    _al_u4627 (
    .a(_al_u4624_o),
    .b(_al_u4625_o),
    .c(_al_u1982_o),
    .d(_al_u4626_o),
    .o(_al_u4627_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u4628 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n26_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [5]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [3]),
    .o(_al_u4628_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(D*C*B))"),
    .INIT(16'h1555))
    _al_u4629 (
    .a(_al_u4628_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n12_lutinv ),
    .c(_al_u4566_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n13 [3]),
    .o(_al_u4629_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u463 (
    .a(_al_u462_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[7] ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[8] ),
    .o(_al_u463_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C*~(~B*A)))"),
    .INIT(16'h2f00))
    _al_u4630 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/mux4_b10_sel_is_4_o ),
    .b(_al_u4627_o),
    .c(_al_u4629_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [6]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n33 [3]));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u4631 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [8]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/haddr_reg [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/haddr_reg [4]),
    .o(_al_u4631_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*(D@C))"),
    .INIT(16'h0880))
    _al_u4632 (
    .a(_al_u4604_o),
    .b(_al_u4631_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/haddr_reg [1]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/haddr_reg [2]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n37 [3]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u4633 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n12_lutinv ),
    .b(_al_u4566_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n13 [3]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [5]),
    .o(_al_u4633_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*C)*~(B*A))"),
    .INIT(16'h0777))
    _al_u4634 (
    .a(\u_cmsdk_mcu/flash_hrdata [3]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [0]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [4]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/rwdata_reg [3]),
    .o(_al_u4634_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(D*C))"),
    .INIT(16'h0444))
    _al_u4635 (
    .a(_al_u4633_o),
    .b(_al_u4634_o),
    .c(\u_cmsdk_mcu/sram_hrdata [3]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [1]),
    .o(_al_u4635_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D*C*B))"),
    .INIT(16'h2aaa))
    _al_u4636 (
    .a(_al_u4635_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/mux6_b3_sel_is_2_o ),
    .c(_al_u4580_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/n19 [3]),
    .o(_al_u4636_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*~A)"),
    .INIT(16'h0100))
    _al_u4637 (
    .a(_al_u4621_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n33 [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n37 [3]),
    .d(_al_u4636_o),
    .o(_al_u4637_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*B)*~(~D*A))"),
    .INIT(16'hf351))
    _al_u4638 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kq7iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pp7iu6 ),
    .c(_al_u4637_o),
    .d(_al_u1839_o),
    .o(_al_u4638_o));
  AL_MAP_LUT4 #(
    .EQN("~((D*~A)*~(C)*~(B)+(D*~A)*C*~(B)+~((D*~A))*C*B+(D*~A)*C*B)"),
    .INIT(16'h2e3f))
    _al_u4639 (
    .a(_al_u4500_o),
    .b(_al_u4501_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H34iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wkipw6 ),
    .o(_al_u4639_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u464 (
    .a(_al_u463_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[5] ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[6] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n25_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u4640 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A25iu6 ),
    .b(_al_u4639_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xiipw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cchiu6 ));
  AL_MAP_LUT4 #(
    .EQN("~(B*A*~(D*C))"),
    .INIT(16'hf777))
    _al_u4641 (
    .a(_al_u4638_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cchiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uy4iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vqjbx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bithu6 ));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u4642 (
    .a(_al_u1986_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inten_padded [4]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttype_padded [4]),
    .o(_al_u4642_o));
  AL_MAP_LUT4 #(
    .EQN("~(C*~((D*~A))*~(B)+C*(D*~A)*~(B)+~(C)*(D*~A)*B+C*(D*~A)*B)"),
    .INIT(16'h8bcf))
    _al_u4643 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpol_padded [4]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [4]),
    .o(_al_u4643_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u4644 (
    .a(_al_u4642_o),
    .b(_al_u1982_o),
    .c(_al_u4643_o),
    .o(_al_u4644_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u4645 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4]),
    .c(\u_cmsdk_mcu/p0_outen [4]),
    .d(\u_cmsdk_mcu/p0_altfunc [4]),
    .o(_al_u4645_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D*~C*A))"),
    .INIT(16'h3133))
    _al_u4646 (
    .a(_al_u4515_o),
    .b(_al_u4645_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4]),
    .d(\u_cmsdk_mcu/p0_out [4]),
    .o(_al_u4646_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*~(~D*~C)))"),
    .INIT(16'h222a))
    _al_u4647 (
    .a(_al_u4511_o),
    .b(_al_u4644_o),
    .c(_al_u4646_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [5]),
    .o(_al_u4647_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h3210))
    _al_u4648 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [4]),
    .d(\u_cmsdk_mcu/p1_out [4]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/mux0_b4/B1_0 ));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u4649 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4]),
    .c(\u_cmsdk_mcu/p1_outen [4]),
    .d(\u_cmsdk_mcu/p1_altfunc [4]),
    .o(_al_u4649_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u465 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[8] ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[9] ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[10] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[11] ),
    .o(_al_u465_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(~B*~(~C*A)))"),
    .INIT(16'h00ce))
    _al_u4650 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/mux0_b4/B1_0 ),
    .b(_al_u4649_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [5]),
    .o(_al_u4650_o));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u4651 (
    .a(_al_u1986_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inten_padded [4]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [4]),
    .o(_al_u4651_o));
  AL_MAP_LUT4 #(
    .EQN("~(C*~((D*~A))*~(B)+C*(D*~A)*~(B)+~(C)*(D*~A)*B+C*(D*~A)*B)"),
    .INIT(16'h8bcf))
    _al_u4652 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpol_padded [4]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[4] ),
    .o(_al_u4652_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~A*~(~D*C))"),
    .INIT(16'h1101))
    _al_u4653 (
    .a(_al_u4650_o),
    .b(_al_u4651_o),
    .c(_al_u1982_o),
    .d(_al_u4652_o),
    .o(_al_u4653_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u4654 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n26_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [6]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [4]),
    .o(_al_u4654_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(D*C*B))"),
    .INIT(16'h1555))
    _al_u4655 (
    .a(_al_u4654_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n12_lutinv ),
    .c(_al_u4566_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n13 [4]),
    .o(_al_u4655_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C*~(~B*A)))"),
    .INIT(16'h2f00))
    _al_u4656 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/mux4_b10_sel_is_4_o ),
    .b(_al_u4653_o),
    .c(_al_u4655_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [6]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n33 [4]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u4657 (
    .a(_al_u4603_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/haddr_reg [0]),
    .o(_al_u4657_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u4658 (
    .a(_al_u4657_o),
    .b(_al_u4605_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n37 [4]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u4659 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n12_lutinv ),
    .b(_al_u4566_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n13 [4]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [5]),
    .o(_al_u4659_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u466 (
    .a(_al_u465_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[6] ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[7] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n27_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*C)*~(B*A))"),
    .INIT(16'h0777))
    _al_u4660 (
    .a(\u_cmsdk_mcu/sram_hrdata [4]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [1]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [4]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/rwdata_reg [4]),
    .o(_al_u4660_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(D*C))"),
    .INIT(16'h0444))
    _al_u4661 (
    .a(_al_u4659_o),
    .b(_al_u4660_o),
    .c(\u_cmsdk_mcu/flash_hrdata [4]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [0]),
    .o(_al_u4661_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D*C*B))"),
    .INIT(16'h2aaa))
    _al_u4662 (
    .a(_al_u4661_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/mux6_b3_sel_is_2_o ),
    .c(_al_u4580_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/n19 [4]),
    .o(_al_u4662_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*~A)"),
    .INIT(16'h0100))
    _al_u4663 (
    .a(_al_u4647_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n33 [4]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n37 [4]),
    .d(_al_u4662_o),
    .o(_al_u4663_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*B)*~(~D*A))"),
    .INIT(16'hf351))
    _al_u4664 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kq7iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pp7iu6 ),
    .c(_al_u4663_o),
    .d(_al_u1841_o),
    .o(_al_u4664_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4665 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uy4iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R05iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jgxpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tokax6 ),
    .o(_al_u4665_o));
  AL_MAP_LUT4 #(
    .EQN("~(B*A*~(D*C))"),
    .INIT(16'hf777))
    _al_u4666 (
    .a(_al_u4664_o),
    .b(_al_u4665_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A25iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G2iax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iithu6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u4667 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n37 [4]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/haddr_reg [1]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n37 [5]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u4668 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/mux6_b3_sel_is_2_o ),
    .b(_al_u4580_o),
    .o(_al_u4668_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u4669 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n12_lutinv ),
    .b(_al_u4566_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n13 [5]),
    .o(_al_u4669_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u467 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] ),
    .o(_al_u467_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*C)*~(B*A))"),
    .INIT(16'h0777))
    _al_u4670 (
    .a(\u_cmsdk_mcu/sram_hrdata [5]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [1]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [4]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/rwdata_reg [5]),
    .o(_al_u4670_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u4671 (
    .a(_al_u4670_o),
    .b(\u_cmsdk_mcu/flash_hrdata [5]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [0]),
    .o(_al_u4671_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u4672 (
    .a(_al_u4669_o),
    .b(_al_u4671_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [5]),
    .o(_al_u4672_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*~(D*B))"),
    .INIT(16'h1050))
    _al_u4673 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n37 [5]),
    .b(_al_u4668_o),
    .c(_al_u4672_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/n19 [5]),
    .o(_al_u4673_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h3210))
    _al_u4674 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [5]),
    .d(\u_cmsdk_mcu/p1_out [5]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/mux0_b5/B1_0 ));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u4675 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4]),
    .c(\u_cmsdk_mcu/p1_outen [5]),
    .d(\u_cmsdk_mcu/p1_altfunc [5]),
    .o(_al_u4675_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(~B*~(~C*A)))"),
    .INIT(16'h00ce))
    _al_u4676 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/mux0_b5/B1_0 ),
    .b(_al_u4675_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [5]),
    .o(_al_u4676_o));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u4677 (
    .a(_al_u1986_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inten_padded [5]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [5]),
    .o(_al_u4677_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*~B))"),
    .INIT(8'ha8))
    _al_u4678 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/mux4_b10_sel_is_4_o ),
    .b(_al_u4676_o),
    .c(_al_u4677_o),
    .o(_al_u4678_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(D*C*B))"),
    .INIT(16'h1555))
    _al_u4679 (
    .a(_al_u4669_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n26_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [7]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [5]),
    .o(_al_u4679_o));
  AL_MAP_LUT4 #(
    .EQN("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'ha088))
    _al_u468 (
    .a(_al_u467_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_rx_buf [7]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [7]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[4] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n26 [7]));
  AL_MAP_LUT4 #(
    .EQN("~(C*~((D*~A))*~(B)+C*(D*~A)*~(B)+~(C)*(D*~A)*B+C*(D*~A)*B)"),
    .INIT(16'h8bcf))
    _al_u4680 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpol_padded [5]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[5] ),
    .o(_al_u4680_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~B*~(~D*A))"),
    .INIT(16'h3010))
    _al_u4681 (
    .a(_al_u1983_o),
    .b(_al_u4678_o),
    .c(_al_u4679_o),
    .d(_al_u4680_o),
    .o(_al_u4681_o));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u4682 (
    .a(_al_u1986_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inten_padded [5]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttype_padded [5]),
    .o(_al_u4682_o));
  AL_MAP_LUT4 #(
    .EQN("~(C*~((D*~A))*~(B)+C*(D*~A)*~(B)+~(C)*(D*~A)*B+C*(D*~A)*B)"),
    .INIT(16'h8bcf))
    _al_u4683 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpol_padded [5]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [5]),
    .o(_al_u4683_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u4684 (
    .a(_al_u4682_o),
    .b(_al_u1982_o),
    .c(_al_u4683_o),
    .o(_al_u4684_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u4685 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4]),
    .c(\u_cmsdk_mcu/p0_outen [5]),
    .d(\u_cmsdk_mcu/p0_altfunc [5]),
    .o(_al_u4685_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D*~C*A))"),
    .INIT(16'h3133))
    _al_u4686 (
    .a(_al_u4515_o),
    .b(_al_u4685_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4]),
    .d(\u_cmsdk_mcu/p0_out [5]),
    .o(_al_u4686_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*~(~D*~C)))"),
    .INIT(16'h222a))
    _al_u4687 (
    .a(_al_u4511_o),
    .b(_al_u4684_o),
    .c(_al_u4686_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [5]),
    .o(_al_u4687_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*A*~(D*~B))"),
    .INIT(16'h080a))
    _al_u4688 (
    .a(_al_u4673_o),
    .b(_al_u4681_o),
    .c(_al_u4687_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [6]),
    .o(_al_u4688_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*B)*~(~D*A))"),
    .INIT(16'hf351))
    _al_u4689 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kq7iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pp7iu6 ),
    .c(_al_u4688_o),
    .d(_al_u1844_o),
    .o(_al_u4689_o));
  AL_MAP_LUT4 #(
    .EQN("((D*B)*~(C)*~(A)+(D*B)*C*~(A)+~((D*B))*C*A+(D*B)*C*A)"),
    .INIT(16'he4a0))
    _al_u469 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n25_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n27_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n26 [7]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n28 [7]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/read_mux_byte0 [7]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4690 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uy4iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R05iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jckax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kakax6 ),
    .o(_al_u4690_o));
  AL_MAP_LUT4 #(
    .EQN("~(B*A*~(D*C))"),
    .INIT(16'hf777))
    _al_u4691 (
    .a(_al_u4689_o),
    .b(_al_u4690_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A25iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F4iax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pithu6 ));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u4692 (
    .a(_al_u1982_o),
    .b(_al_u4515_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n12_lutinv ),
    .d(_al_u4566_o),
    .o(_al_u4692_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u4693 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n26_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [8]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [6]),
    .o(_al_u4693_o));
  AL_MAP_LUT4 #(
    .EQN("~(C*~((D*~A))*~(B)+C*(D*~A)*~(B)+~(C)*(D*~A)*B+C*(D*~A)*B)"),
    .INIT(16'h8bcf))
    _al_u4694 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpol_padded [6]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[6] ),
    .o(_al_u4694_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~B*~(~D*A))"),
    .INIT(16'h0301))
    _al_u4695 (
    .a(_al_u1983_o),
    .b(_al_u4692_o),
    .c(_al_u4693_o),
    .d(_al_u4694_o),
    .o(_al_u4695_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h3210))
    _al_u4696 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [6]),
    .d(\u_cmsdk_mcu/p1_out [6]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/mux0_b6/B1_0 ));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u4697 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4]),
    .c(\u_cmsdk_mcu/p1_outen [6]),
    .d(\u_cmsdk_mcu/p1_altfunc [6]),
    .o(_al_u4697_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(~B*~(~C*A)))"),
    .INIT(16'h00ce))
    _al_u4698 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/mux0_b6/B1_0 ),
    .b(_al_u4697_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [5]),
    .o(_al_u4698_o));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u4699 (
    .a(_al_u1986_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inten_padded [6]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [6]),
    .o(_al_u4699_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u470 (
    .a(_al_u467_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[4] ),
    .o(_al_u470_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*~(~D*~C)))"),
    .INIT(16'h222a))
    _al_u4700 (
    .a(_al_u4695_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/mux4_b10_sel_is_4_o ),
    .c(_al_u4698_o),
    .d(_al_u4699_o),
    .o(_al_u4700_o));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u4701 (
    .a(_al_u1986_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inten_padded [6]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttype_padded [6]),
    .o(_al_u4701_o));
  AL_MAP_LUT4 #(
    .EQN("~(C*~((D*~A))*~(B)+C*(D*~A)*~(B)+~(C)*(D*~A)*B+C*(D*~A)*B)"),
    .INIT(16'h8bcf))
    _al_u4702 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpol_padded [6]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [6]),
    .o(_al_u4702_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u4703 (
    .a(_al_u4701_o),
    .b(_al_u1982_o),
    .c(_al_u4702_o),
    .o(_al_u4703_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u4704 (
    .a(_al_u4515_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4]),
    .c(\u_cmsdk_mcu/p0_out [6]),
    .o(_al_u4704_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u4705 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4]),
    .c(\u_cmsdk_mcu/p0_outen [6]),
    .d(\u_cmsdk_mcu/p0_altfunc [6]),
    .o(_al_u4705_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(~D*~(~C*~B)))"),
    .INIT(16'haa02))
    _al_u4706 (
    .a(_al_u4703_o),
    .b(_al_u4704_o),
    .c(_al_u4705_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [5]),
    .o(_al_u4706_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(~C*~(B*~A)))"),
    .INIT(16'hf400))
    _al_u4707 (
    .a(_al_u4706_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/mux4_b10_sel_is_4_o ),
    .c(_al_u4692_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [5]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n31 [6]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4708 (
    .a(\u_cmsdk_mcu/sram_hrdata [6]),
    .b(\u_cmsdk_mcu/flash_hrdata [6]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [0]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [1]),
    .o(_al_u4708_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u4709 (
    .a(_al_u4708_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [4]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/rwdata_reg [6]),
    .o(_al_u4709_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u471 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n25_lutinv ),
    .b(_al_u470_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n7_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u4710 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [2]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [4]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [5]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/mux4_b6_sel_is_13_o ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u4711 (
    .a(_al_u4668_o),
    .b(_al_u4709_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/mux4_b6_sel_is_13_o ),
    .o(_al_u4711_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~B*~(D*~A))"),
    .INIT(16'h2030))
    _al_u4712 (
    .a(_al_u4700_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n31 [6]),
    .c(_al_u4711_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [6]),
    .o(_al_u4712_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*B)*~(~D*A))"),
    .INIT(16'hf351))
    _al_u4713 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kq7iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pp7iu6 ),
    .c(_al_u4712_o),
    .d(_al_u1846_o),
    .o(_al_u4713_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u4714 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A25iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R05iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E8iax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4jax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q5hiu6 ));
  AL_MAP_LUT4 #(
    .EQN("~(B*A*~(D*C))"),
    .INIT(16'hf777))
    _al_u4715 (
    .a(_al_u4713_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q5hiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uy4iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L8kax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Withu6 ));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u4716 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n12_lutinv ),
    .b(_al_u4566_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n13 [7]),
    .o(_al_u4716_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*C)*~(B*A))"),
    .INIT(16'h0777))
    _al_u4717 (
    .a(\u_cmsdk_mcu/sram_hrdata [7]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [1]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [4]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/rwdata_reg [7]),
    .o(_al_u4717_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u4718 (
    .a(_al_u4717_o),
    .b(\u_cmsdk_mcu/flash_hrdata [7]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [0]),
    .o(_al_u4718_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u4719 (
    .a(_al_u4716_o),
    .b(_al_u4718_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [5]),
    .o(_al_u4719_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u472 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[4] ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[5] ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[6] ),
    .o(_al_u472_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*~(D*B))"),
    .INIT(16'h1050))
    _al_u4720 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n37 [5]),
    .b(_al_u4668_o),
    .c(_al_u4719_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/n19 [7]),
    .o(_al_u4720_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h3210))
    _al_u4721 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [7]),
    .d(\u_cmsdk_mcu/p1_out [7]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/mux0_b7/B1_0 ));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u4722 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4]),
    .c(\u_cmsdk_mcu/p1_outen [7]),
    .d(\u_cmsdk_mcu/p1_altfunc [7]),
    .o(_al_u4722_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(~B*~(~C*A)))"),
    .INIT(16'h00ce))
    _al_u4723 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/mux0_b7/B1_0 ),
    .b(_al_u4722_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [5]),
    .o(_al_u4723_o));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u4724 (
    .a(_al_u1986_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inten_padded [7]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [7]),
    .o(_al_u4724_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*~B))"),
    .INIT(8'ha8))
    _al_u4725 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/mux4_b10_sel_is_4_o ),
    .b(_al_u4723_o),
    .c(_al_u4724_o),
    .o(_al_u4725_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(D*C*B))"),
    .INIT(16'h1555))
    _al_u4726 (
    .a(_al_u4716_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n26_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [9]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [7]),
    .o(_al_u4726_o));
  AL_MAP_LUT4 #(
    .EQN("~(C*~((D*~A))*~(B)+C*(D*~A)*~(B)+~(C)*(D*~A)*B+C*(D*~A)*B)"),
    .INIT(16'h8bcf))
    _al_u4727 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpol_padded [7]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[7] ),
    .o(_al_u4727_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~B*~(~D*A))"),
    .INIT(16'h3010))
    _al_u4728 (
    .a(_al_u1983_o),
    .b(_al_u4725_o),
    .c(_al_u4726_o),
    .d(_al_u4727_o),
    .o(_al_u4728_o));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u4729 (
    .a(_al_u1986_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inten_padded [7]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttype_padded [7]),
    .o(_al_u4729_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u473 (
    .a(_al_u463_o),
    .b(_al_u472_o),
    .o(_al_u473_o));
  AL_MAP_LUT4 #(
    .EQN("~(C*~((D*~A))*~(B)+C*(D*~A)*~(B)+~(C)*(D*~A)*B+C*(D*~A)*B)"),
    .INIT(16'h8bcf))
    _al_u4730 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpol_padded [7]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [7]),
    .o(_al_u4730_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u4731 (
    .a(_al_u4729_o),
    .b(_al_u1982_o),
    .c(_al_u4730_o),
    .o(_al_u4731_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u4732 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4]),
    .c(\u_cmsdk_mcu/p0_outen [7]),
    .d(\u_cmsdk_mcu/p0_altfunc [7]),
    .o(_al_u4732_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D*~C*A))"),
    .INIT(16'h3133))
    _al_u4733 (
    .a(_al_u4515_o),
    .b(_al_u4732_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4]),
    .d(\u_cmsdk_mcu/p0_out [7]),
    .o(_al_u4733_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*~(~D*~C)))"),
    .INIT(16'h222a))
    _al_u4734 (
    .a(_al_u4511_o),
    .b(_al_u4731_o),
    .c(_al_u4733_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [5]),
    .o(_al_u4734_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*A*~(D*~B))"),
    .INIT(16'h080a))
    _al_u4735 (
    .a(_al_u4720_o),
    .b(_al_u4728_o),
    .c(_al_u4734_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [6]),
    .o(_al_u4735_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*B)*~(~D*A))"),
    .INIT(16'hf351))
    _al_u4736 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kq7iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pp7iu6 ),
    .c(_al_u4735_o),
    .d(_al_u1848_o),
    .o(_al_u4736_o));
  AL_MAP_LUT4 #(
    .EQN("~((D*~A)*~(C)*~(B)+(D*~A)*C*~(B)+~((D*~A))*C*B+(D*~A)*C*B)"),
    .INIT(16'h2e3f))
    _al_u4737 (
    .a(_al_u4500_o),
    .b(_al_u4501_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Df4iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N4kax6 ),
    .o(_al_u4737_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u4738 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A25iu6 ),
    .b(_al_u4737_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zqiax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y2hiu6 ));
  AL_MAP_LUT4 #(
    .EQN("~(B*A*~(D*C))"),
    .INIT(16'hf777))
    _al_u4739 (
    .a(_al_u4736_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y2hiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uy4iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O2kax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Djthu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'h0a0c))
    _al_u474 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_ctrl [5]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_rx_buf [5]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/mux3_b5/B1_0 ));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u4740 (
    .a(_al_u1986_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inten_padded [9]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttype_padded [9]),
    .o(_al_u4740_o));
  AL_MAP_LUT4 #(
    .EQN("~(C*~((D*~A))*~(B)+C*(D*~A)*~(B)+~(C)*(D*~A)*B+C*(D*~A)*B)"),
    .INIT(16'h8bcf))
    _al_u4741 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpol_padded [9]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [9]),
    .o(_al_u4741_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u4742 (
    .a(_al_u4740_o),
    .b(_al_u1982_o),
    .c(_al_u4741_o),
    .o(_al_u4742_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u4743 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4]),
    .c(\u_cmsdk_mcu/p0_outen [9]),
    .d(\u_cmsdk_mcu/p0_altfunc [9]),
    .o(_al_u4743_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D*~C*A))"),
    .INIT(16'h3133))
    _al_u4744 (
    .a(_al_u4515_o),
    .b(_al_u4743_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4]),
    .d(\u_cmsdk_mcu/p0_out [9]),
    .o(_al_u4744_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*~(~D*~C)))"),
    .INIT(16'h222a))
    _al_u4745 (
    .a(_al_u4511_o),
    .b(_al_u4742_o),
    .c(_al_u4744_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [5]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n31 [9]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*C)*~(B*A))"),
    .INIT(16'h0777))
    _al_u4746 (
    .a(\u_cmsdk_mcu/sram_hrdata [9]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [1]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [4]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/rwdata_reg [9]),
    .o(_al_u4746_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(D*C))"),
    .INIT(16'h0444))
    _al_u4747 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n31 [9]),
    .b(_al_u4746_o),
    .c(\u_cmsdk_mcu/flash_hrdata [9]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [0]),
    .o(_al_u4747_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h3210))
    _al_u4748 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [9]),
    .d(\u_cmsdk_mcu/p1_out [9]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/mux0_b9/B1_0 ));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u4749 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4]),
    .c(\u_cmsdk_mcu/p1_outen [9]),
    .d(\u_cmsdk_mcu/p1_altfunc [9]),
    .o(_al_u4749_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u475 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n7_lutinv ),
    .b(_al_u473_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/mux3_b5/B1_0 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [5]),
    .o(_al_u475_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(~B*~(~C*A)))"),
    .INIT(16'h00ce))
    _al_u4750 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/mux0_b9/B1_0 ),
    .b(_al_u4749_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [5]),
    .o(_al_u4750_o));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u4751 (
    .a(_al_u1986_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inten_padded [9]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [9]),
    .o(_al_u4751_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*~B))"),
    .INIT(8'ha8))
    _al_u4752 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/mux4_b10_sel_is_4_o ),
    .b(_al_u4750_o),
    .c(_al_u4751_o),
    .o(_al_u4752_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*~A)"),
    .INIT(16'h4000))
    _al_u4753 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [10]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [11]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [9]),
    .o(_al_u4753_o));
  AL_MAP_LUT4 #(
    .EQN("~(C*~((D*~A))*~(B)+C*(D*~A)*~(B)+~(C)*(D*~A)*B+C*(D*~A)*B)"),
    .INIT(16'h8bcf))
    _al_u4754 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpol_padded [9]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[9] ),
    .o(_al_u4754_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~B*~(~D*A))"),
    .INIT(16'h0301))
    _al_u4755 (
    .a(_al_u1983_o),
    .b(_al_u4752_o),
    .c(_al_u4753_o),
    .d(_al_u4754_o),
    .o(_al_u4755_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*~B))"),
    .INIT(8'h8a))
    _al_u4756 (
    .a(_al_u4747_o),
    .b(_al_u4755_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [6]),
    .o(_al_u4756_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*B)*~(~D*A))"),
    .INIT(16'hf351))
    _al_u4757 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kq7iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pp7iu6 ),
    .c(_al_u4756_o),
    .d(_al_u1852_o),
    .o(_al_u4757_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4758 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uy4iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R05iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rwjax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sujax6 ),
    .o(_al_u4758_o));
  AL_MAP_LUT4 #(
    .EQN("~(B*A*~(D*C))"),
    .INIT(16'hf777))
    _al_u4759 (
    .a(_al_u4757_o),
    .b(_al_u4758_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A25iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuiax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jzuhu6 ));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*B))"),
    .INIT(8'hd5))
    _al_u476 (
    .a(_al_u475_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n27_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n28 [5]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/read_mux_byte0 [5]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u4760 (
    .a(_al_u1986_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inten_padded [10]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttype_padded [10]),
    .o(_al_u4760_o));
  AL_MAP_LUT4 #(
    .EQN("~(C*~((D*~A))*~(B)+C*(D*~A)*~(B)+~(C)*(D*~A)*B+C*(D*~A)*B)"),
    .INIT(16'h8bcf))
    _al_u4761 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpol_padded [10]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [10]),
    .o(_al_u4761_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u4762 (
    .a(_al_u4760_o),
    .b(_al_u1982_o),
    .c(_al_u4761_o),
    .o(_al_u4762_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u4763 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4]),
    .c(\u_cmsdk_mcu/p0_outen [10]),
    .d(\u_cmsdk_mcu/p0_altfunc [10]),
    .o(_al_u4763_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D*~C*A))"),
    .INIT(16'h3133))
    _al_u4764 (
    .a(_al_u4515_o),
    .b(_al_u4763_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4]),
    .d(\u_cmsdk_mcu/p0_out [10]),
    .o(_al_u4764_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*~(~D*~C)))"),
    .INIT(16'h222a))
    _al_u4765 (
    .a(_al_u4511_o),
    .b(_al_u4762_o),
    .c(_al_u4764_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [5]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n31 [10]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*C)*~(B*A))"),
    .INIT(16'h0777))
    _al_u4766 (
    .a(\u_cmsdk_mcu/sram_hrdata [10]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [1]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [4]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/rwdata_reg [10]),
    .o(_al_u4766_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(D*C))"),
    .INIT(16'h0444))
    _al_u4767 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n31 [10]),
    .b(_al_u4766_o),
    .c(\u_cmsdk_mcu/flash_hrdata [10]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [0]),
    .o(_al_u4767_o));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u4768 (
    .a(_al_u1986_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inten_padded [10]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [10]),
    .o(_al_u4768_o));
  AL_MAP_LUT4 #(
    .EQN("~(C*~((D*~A))*~(B)+C*(D*~A)*~(B)+~(C)*(D*~A)*B+C*(D*~A)*B)"),
    .INIT(16'h8bcf))
    _al_u4769 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpol_padded [10]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[10] ),
    .o(_al_u4769_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'h0a0c))
    _al_u477 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_ctrl [4]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_rx_buf [4]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/mux3_b4/B1_0 ));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u4770 (
    .a(_al_u4768_o),
    .b(_al_u1982_o),
    .c(_al_u4769_o),
    .o(_al_u4770_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h3210))
    _al_u4771 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [10]),
    .d(\u_cmsdk_mcu/p1_out [10]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/mux0_b10/B1_0 ));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u4772 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4]),
    .c(\u_cmsdk_mcu/p1_outen [10]),
    .d(\u_cmsdk_mcu/p1_altfunc [10]),
    .o(_al_u4772_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(~B*~(~C*A)))"),
    .INIT(16'h00ce))
    _al_u4773 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/mux0_b10/B1_0 ),
    .b(_al_u4772_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [5]),
    .o(_al_u4773_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*~A)"),
    .INIT(16'h4000))
    _al_u4774 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [10]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [11]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [10]),
    .o(_al_u4774_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(A*~(~C*B)))"),
    .INIT(16'h005d))
    _al_u4775 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/mux4_b10_sel_is_4_o ),
    .b(_al_u4770_o),
    .c(_al_u4773_o),
    .d(_al_u4774_o),
    .o(_al_u4775_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*~B))"),
    .INIT(8'h8a))
    _al_u4776 (
    .a(_al_u4767_o),
    .b(_al_u4775_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [6]),
    .o(_al_u4776_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*B)*~(~D*A))"),
    .INIT(16'hf351))
    _al_u4777 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kq7iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pp7iu6 ),
    .c(_al_u4776_o),
    .d(_al_u1854_o),
    .o(_al_u4777_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4778 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A25iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R05iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wwiax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Epciu6 ));
  AL_MAP_LUT4 #(
    .EQN("~(B*A*~(D*C))"),
    .INIT(16'hf777))
    _al_u4779 (
    .a(_al_u4777_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Epciu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uy4iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sqjax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qzuhu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u478 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n7_lutinv ),
    .b(_al_u473_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/mux3_b4/B1_0 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [4]),
    .o(_al_u478_o));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u4780 (
    .a(_al_u1986_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inten_padded [11]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttype_padded [11]),
    .o(_al_u4780_o));
  AL_MAP_LUT4 #(
    .EQN("~(C*~((D*~A))*~(B)+C*(D*~A)*~(B)+~(C)*(D*~A)*B+C*(D*~A)*B)"),
    .INIT(16'h8bcf))
    _al_u4781 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpol_padded [11]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [11]),
    .o(_al_u4781_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u4782 (
    .a(_al_u4780_o),
    .b(_al_u1982_o),
    .c(_al_u4781_o),
    .o(_al_u4782_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u4783 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4]),
    .c(\u_cmsdk_mcu/p0_outen [11]),
    .d(\u_cmsdk_mcu/p0_altfunc [11]),
    .o(_al_u4783_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D*~C*A))"),
    .INIT(16'h3133))
    _al_u4784 (
    .a(_al_u4515_o),
    .b(_al_u4783_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4]),
    .d(\u_cmsdk_mcu/p0_out [11]),
    .o(_al_u4784_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*~(~D*~C)))"),
    .INIT(16'h222a))
    _al_u4785 (
    .a(_al_u4511_o),
    .b(_al_u4782_o),
    .c(_al_u4784_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [5]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n31 [11]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4786 (
    .a(\u_cmsdk_mcu/sram_hrdata [11]),
    .b(\u_cmsdk_mcu/flash_hrdata [11]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [0]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [1]),
    .o(_al_u4786_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(D*C))"),
    .INIT(16'h0444))
    _al_u4787 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n31 [11]),
    .b(_al_u4786_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [4]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/rwdata_reg [11]),
    .o(_al_u4787_o));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u4788 (
    .a(_al_u1986_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inten_padded [11]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [11]),
    .o(_al_u4788_o));
  AL_MAP_LUT4 #(
    .EQN("~(C*~((D*~A))*~(B)+C*(D*~A)*~(B)+~(C)*(D*~A)*B+C*(D*~A)*B)"),
    .INIT(16'h8bcf))
    _al_u4789 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpol_padded [11]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[11] ),
    .o(_al_u4789_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*B))"),
    .INIT(8'hd5))
    _al_u479 (
    .a(_al_u478_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n27_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n28 [4]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/read_mux_byte0 [4]));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u4790 (
    .a(_al_u4788_o),
    .b(_al_u1982_o),
    .c(_al_u4789_o),
    .o(_al_u4790_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h3210))
    _al_u4791 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [11]),
    .d(\u_cmsdk_mcu/p1_out [11]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/mux0_b11/B1_0 ));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u4792 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4]),
    .c(\u_cmsdk_mcu/p1_outen [11]),
    .d(\u_cmsdk_mcu/p1_altfunc [11]),
    .o(_al_u4792_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(~B*~(~C*A)))"),
    .INIT(16'h00ce))
    _al_u4793 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/mux0_b11/B1_0 ),
    .b(_al_u4792_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [5]),
    .o(_al_u4793_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*~A)"),
    .INIT(16'h4000))
    _al_u4794 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [10]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [11]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [5]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [11]),
    .o(_al_u4794_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(A*~(~C*B)))"),
    .INIT(16'h005d))
    _al_u4795 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/mux4_b10_sel_is_4_o ),
    .b(_al_u4790_o),
    .c(_al_u4793_o),
    .d(_al_u4794_o),
    .o(_al_u4795_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*~B))"),
    .INIT(8'h8a))
    _al_u4796 (
    .a(_al_u4787_o),
    .b(_al_u4795_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [6]),
    .o(_al_u4796_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*B)*~(~D*A))"),
    .INIT(16'hf351))
    _al_u4797 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kq7iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pp7iu6 ),
    .c(_al_u4796_o),
    .d(_al_u1856_o),
    .o(_al_u4797_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4798 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A25iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R05iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wyiax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Anciu6 ));
  AL_MAP_LUT4 #(
    .EQN("~(B*A*~(D*C))"),
    .INIT(16'hf777))
    _al_u4799 (
    .a(_al_u4797_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Anciu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uy4iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Smjax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xzuhu6 ));
  AL_MAP_LUT4 #(
    .EQN("(C*B*~(D*~A))"),
    .INIT(16'h80c0))
    _al_u480 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_ctrl [5]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_rx_overrun ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] ),
    .o(_al_u480_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h3210))
    _al_u4800 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [12]),
    .d(\u_cmsdk_mcu/p1_out [12]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/mux0_b12/B1_0 ));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u4801 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4]),
    .c(\u_cmsdk_mcu/p1_outen [12]),
    .d(\u_cmsdk_mcu/p1_altfunc [12]),
    .o(_al_u4801_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(~B*~(~C*A)))"),
    .INIT(16'h00ce))
    _al_u4802 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/mux0_b12/B1_0 ),
    .b(_al_u4801_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [5]),
    .o(_al_u4802_o));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u4803 (
    .a(_al_u1986_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inten_padded [12]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [12]),
    .o(_al_u4803_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*~B))"),
    .INIT(8'ha8))
    _al_u4804 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/mux4_b10_sel_is_4_o ),
    .b(_al_u4802_o),
    .c(_al_u4803_o),
    .o(_al_u4804_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*~A)"),
    .INIT(16'h4000))
    _al_u4805 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [10]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [11]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [6]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [12]),
    .o(_al_u4805_o));
  AL_MAP_LUT4 #(
    .EQN("~(C*~((D*~A))*~(B)+C*(D*~A)*~(B)+~(C)*(D*~A)*B+C*(D*~A)*B)"),
    .INIT(16'h8bcf))
    _al_u4806 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpol_padded [12]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[12] ),
    .o(_al_u4806_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~B*~(~D*A))"),
    .INIT(16'h0301))
    _al_u4807 (
    .a(_al_u1983_o),
    .b(_al_u4804_o),
    .c(_al_u4805_o),
    .d(_al_u4806_o),
    .o(_al_u4807_o));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u4808 (
    .a(_al_u1986_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inten_padded [12]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttype_padded [12]),
    .o(_al_u4808_o));
  AL_MAP_LUT4 #(
    .EQN("~(C*~((D*~A))*~(B)+C*(D*~A)*~(B)+~(C)*(D*~A)*B+C*(D*~A)*B)"),
    .INIT(16'h8bcf))
    _al_u4809 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpol_padded [12]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [12]),
    .o(_al_u4809_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'h0a0c))
    _al_u481 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_ctrl [3]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_rx_buf [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] ),
    .o(_al_u481_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u4810 (
    .a(_al_u4808_o),
    .b(_al_u1982_o),
    .c(_al_u4809_o),
    .o(_al_u4810_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u4811 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4]),
    .c(\u_cmsdk_mcu/p0_outen [12]),
    .d(\u_cmsdk_mcu/p0_altfunc [12]),
    .o(_al_u4811_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D*~C*A))"),
    .INIT(16'h3133))
    _al_u4812 (
    .a(_al_u4515_o),
    .b(_al_u4811_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4]),
    .d(\u_cmsdk_mcu/p0_out [12]),
    .o(_al_u4812_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*~(~D*~C)))"),
    .INIT(16'h222a))
    _al_u4813 (
    .a(_al_u4511_o),
    .b(_al_u4810_o),
    .c(_al_u4812_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [5]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n31 [12]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4814 (
    .a(\u_cmsdk_mcu/sram_hrdata [12]),
    .b(\u_cmsdk_mcu/flash_hrdata [12]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [0]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [1]),
    .o(_al_u4814_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(D*C))"),
    .INIT(16'h0444))
    _al_u4815 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n37 [14]),
    .b(_al_u4814_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [4]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/rwdata_reg [12]),
    .o(_al_u4815_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~B*~(D*~A))"),
    .INIT(16'h2030))
    _al_u4816 (
    .a(_al_u4807_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n31 [12]),
    .c(_al_u4815_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [6]),
    .o(_al_u4816_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*B)*~(~D*A))"),
    .INIT(16'hf351))
    _al_u4817 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kq7iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pp7iu6 ),
    .c(_al_u4816_o),
    .d(_al_u1859_o),
    .o(_al_u4817_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4818 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A25iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R05iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Skjax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W0jax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wkciu6 ));
  AL_MAP_LUT4 #(
    .EQN("~(B*A*~(D*C))"),
    .INIT(16'hf777))
    _al_u4819 (
    .a(_al_u4817_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wkciu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uy4iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sijax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E0vhu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~D*A*~(~C*~B))"),
    .INIT(16'h00a8))
    _al_u482 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n25_lutinv ),
    .b(_al_u480_o),
    .c(_al_u481_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[4] ),
    .o(_al_u482_o));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u4820 (
    .a(_al_u1986_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inten_padded [8]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttype_padded [8]),
    .o(_al_u4820_o));
  AL_MAP_LUT4 #(
    .EQN("~(C*~((D*~A))*~(B)+C*(D*~A)*~(B)+~(C)*(D*~A)*B+C*(D*~A)*B)"),
    .INIT(16'h8bcf))
    _al_u4821 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpol_padded [8]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [8]),
    .o(_al_u4821_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u4822 (
    .a(_al_u4820_o),
    .b(_al_u1982_o),
    .c(_al_u4821_o),
    .o(_al_u4822_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u4823 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4]),
    .c(\u_cmsdk_mcu/p0_outen [8]),
    .d(\u_cmsdk_mcu/p0_altfunc [8]),
    .o(_al_u4823_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D*~C*A))"),
    .INIT(16'h3133))
    _al_u4824 (
    .a(_al_u4515_o),
    .b(_al_u4823_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4]),
    .d(\u_cmsdk_mcu/p0_out [8]),
    .o(_al_u4824_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*~(~D*~C)))"),
    .INIT(16'h222a))
    _al_u4825 (
    .a(_al_u4511_o),
    .b(_al_u4822_o),
    .c(_al_u4824_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [5]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n31 [8]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4826 (
    .a(\u_cmsdk_mcu/sram_hrdata [8]),
    .b(\u_cmsdk_mcu/flash_hrdata [8]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [0]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [1]),
    .o(_al_u4826_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(D*C))"),
    .INIT(16'h0444))
    _al_u4827 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n31 [8]),
    .b(_al_u4826_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [4]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/rwdata_reg [8]),
    .o(_al_u4827_o));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u4828 (
    .a(_al_u1986_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inten_padded [8]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [8]),
    .o(_al_u4828_o));
  AL_MAP_LUT4 #(
    .EQN("~(C*~((D*~A))*~(B)+C*(D*~A)*~(B)+~(C)*(D*~A)*B+C*(D*~A)*B)"),
    .INIT(16'h8bcf))
    _al_u4829 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpol_padded [8]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[8] ),
    .o(_al_u4829_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u483 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n27_lutinv ),
    .b(_al_u482_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n28 [3]),
    .o(_al_u483_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u4830 (
    .a(_al_u4828_o),
    .b(_al_u1982_o),
    .c(_al_u4829_o),
    .o(_al_u4830_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h3210))
    _al_u4831 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [8]),
    .d(\u_cmsdk_mcu/p1_out [8]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/mux0_b8/B1_0 ));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u4832 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4]),
    .c(\u_cmsdk_mcu/p1_outen [8]),
    .d(\u_cmsdk_mcu/p1_altfunc [8]),
    .o(_al_u4832_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(~B*~(~C*A)))"),
    .INIT(16'h00ce))
    _al_u4833 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/mux0_b8/B1_0 ),
    .b(_al_u4832_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [5]),
    .o(_al_u4833_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*~A)"),
    .INIT(16'h4000))
    _al_u4834 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [10]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [11]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [8]),
    .o(_al_u4834_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(A*~(~C*B)))"),
    .INIT(16'h005d))
    _al_u4835 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/mux4_b10_sel_is_4_o ),
    .b(_al_u4830_o),
    .c(_al_u4833_o),
    .d(_al_u4834_o),
    .o(_al_u4835_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*~B))"),
    .INIT(8'h8a))
    _al_u4836 (
    .a(_al_u4827_o),
    .b(_al_u4835_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [6]),
    .o(_al_u4836_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*B)*~(~D*A))"),
    .INIT(16'hf351))
    _al_u4837 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kq7iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pp7iu6 ),
    .c(_al_u4836_o),
    .d(_al_u1850_o),
    .o(_al_u4837_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4838 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uy4iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R05iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qyjax6 ),
    .o(_al_u4838_o));
  AL_MAP_LUT4 #(
    .EQN("~(B*A*~(D*C))"),
    .INIT(16'hf777))
    _al_u4839 (
    .a(_al_u4837_o),
    .b(_al_u4838_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A25iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ysiax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V5vhu6 ));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*B))"),
    .INIT(8'hd5))
    _al_u484 (
    .a(_al_u483_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n7_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [3]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/read_mux_byte0 [3]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .INIT(16'h5140))
    _al_u4840 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [2]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [3]),
    .c(\u_cmsdk_mcu/LOCKUPRESET ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/remap_ctrl ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/mux3_b0/B1_0 ));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u4841 (
    .a(_al_u2992_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/mux3_b0/B1_0 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [4]),
    .o(_al_u4841_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u4842 (
    .a(_al_u4841_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/mux6_b3_sel_is_2_o ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/n19 [0]),
    .o(_al_u4842_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(A*~(D*B)))"),
    .INIT(16'hd050))
    _al_u4843 (
    .a(_al_u4842_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/n34_lutinv ),
    .c(_al_u4580_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_resetinfo [0]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n35 [0]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u4844 (
    .a(_al_u1986_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inten_padded [0]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttype_padded [0]),
    .o(_al_u4844_o));
  AL_MAP_LUT4 #(
    .EQN("~(C*~((D*~A))*~(B)+C*(D*~A)*~(B)+~(C)*(D*~A)*B+C*(D*~A)*B)"),
    .INIT(16'h8bcf))
    _al_u4845 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpol_padded [0]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [0]),
    .o(_al_u4845_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u4846 (
    .a(_al_u4844_o),
    .b(_al_u1982_o),
    .c(_al_u4845_o),
    .o(_al_u4846_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u4847 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4]),
    .c(\u_cmsdk_mcu/p0_outen [0]),
    .d(\u_cmsdk_mcu/p0_altfunc [0]),
    .o(_al_u4847_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D*~C*A))"),
    .INIT(16'h3133))
    _al_u4848 (
    .a(_al_u4515_o),
    .b(_al_u4847_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4]),
    .d(\u_cmsdk_mcu/p0_out [0]),
    .o(_al_u4848_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*~(~D*~C)))"),
    .INIT(16'h222a))
    _al_u4849 (
    .a(_al_u4511_o),
    .b(_al_u4846_o),
    .c(_al_u4848_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [5]),
    .o(_al_u4849_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u485 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_ctrl [4]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_tx_overrun ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/uart0_txovrint ));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B@A))"),
    .INIT(8'h90))
    _al_u4850 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/haddr_reg [2]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/haddr_reg [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/haddr_reg [4]),
    .o(_al_u4850_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u4851 (
    .a(_al_u4657_o),
    .b(_al_u4850_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [8]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/haddr_reg [1]),
    .o(_al_u4851_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u4852 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n12_lutinv ),
    .b(_al_u4566_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n13 [0]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [5]),
    .o(_al_u4852_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*C)*~(B*A))"),
    .INIT(16'h0777))
    _al_u4853 (
    .a(\u_cmsdk_mcu/flash_hrdata [0]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [0]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [4]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/rwdata_reg [0]),
    .o(_al_u4853_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(D*C))"),
    .INIT(16'h0444))
    _al_u4854 (
    .a(_al_u4852_o),
    .b(_al_u4853_o),
    .c(\u_cmsdk_mcu/sram_hrdata [0]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [1]),
    .o(_al_u4854_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*~A)"),
    .INIT(16'h0100))
    _al_u4855 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n37 [2]),
    .b(_al_u4851_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n37 [14]),
    .d(_al_u4854_o),
    .o(_al_u4855_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h3210))
    _al_u4856 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [0]),
    .d(\u_cmsdk_mcu/p1_out [0]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/mux0_b0/B1_0 ));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u4857 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4]),
    .c(\u_cmsdk_mcu/p1_outen [0]),
    .d(\u_cmsdk_mcu/p1_altfunc [0]),
    .o(_al_u4857_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(~B*~(~C*A)))"),
    .INIT(16'h00ce))
    _al_u4858 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/mux0_b0/B1_0 ),
    .b(_al_u4857_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [5]),
    .o(_al_u4858_o));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u4859 (
    .a(_al_u1986_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inten_padded [0]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [0]),
    .o(_al_u4859_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h5ff3))
    _al_u486 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/uart0_txovrint ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_rx_buf [2]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] ),
    .o(_al_u486_o));
  AL_MAP_LUT4 #(
    .EQN("~(C*~((D*~A))*~(B)+C*(D*~A)*~(B)+~(C)*(D*~A)*B+C*(D*~A)*B)"),
    .INIT(16'h8bcf))
    _al_u4860 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpol_padded [0]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[0] ),
    .o(_al_u4860_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~A*~(~D*C))"),
    .INIT(16'h1101))
    _al_u4861 (
    .a(_al_u4858_o),
    .b(_al_u4859_o),
    .c(_al_u1982_o),
    .d(_al_u4860_o),
    .o(_al_u4861_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u4862 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n26_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [0]),
    .o(_al_u4862_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(D*C*B))"),
    .INIT(16'h1555))
    _al_u4863 (
    .a(_al_u4862_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n12_lutinv ),
    .c(_al_u4566_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n13 [0]),
    .o(_al_u4863_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C*~(~B*A)))"),
    .INIT(16'h2f00))
    _al_u4864 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/mux4_b10_sel_is_4_o ),
    .b(_al_u4861_o),
    .c(_al_u4863_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [6]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n33 [0]));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*~B*~A)"),
    .INIT(16'h0010))
    _al_u4865 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n35 [0]),
    .b(_al_u4849_o),
    .c(_al_u4855_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n33 [0]),
    .o(_al_u4865_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*B)*~(~D*A))"),
    .INIT(16'hf351))
    _al_u4866 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kq7iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pp7iu6 ),
    .c(_al_u4865_o),
    .d(_al_u1868_o),
    .o(_al_u4866_o));
  AL_MAP_LUT4 #(
    .EQN("~((D*~A)*~(C)*~(B)+(D*~A)*C*~(B)+~((D*~A))*C*B+(D*~A)*C*B)"),
    .INIT(16'h2e3f))
    _al_u4867 (
    .a(_al_u4500_o),
    .b(_al_u4501_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T24iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wfspw6 ),
    .o(_al_u4867_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u4868 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A25iu6 ),
    .b(_al_u4867_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xdspw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A3biu6 ));
  AL_MAP_LUT4 #(
    .EQN("~(B*A*~(D*C))"),
    .INIT(16'hf777))
    _al_u4869 (
    .a(_al_u4866_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A3biu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uy4iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tcjax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S7vhu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf53f))
    _al_u487 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_ctrl [2]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_tx_overrun ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] ),
    .o(_al_u487_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h3210))
    _al_u4870 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [13]),
    .d(\u_cmsdk_mcu/p1_out [13]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/mux0_b13/B1_0 ));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u4871 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4]),
    .c(\u_cmsdk_mcu/p1_outen [13]),
    .d(\u_cmsdk_mcu/p1_altfunc [13]),
    .o(_al_u4871_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(~B*~(~C*A)))"),
    .INIT(16'h00ce))
    _al_u4872 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/mux0_b13/B1_0 ),
    .b(_al_u4871_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [5]),
    .o(_al_u4872_o));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u4873 (
    .a(_al_u1986_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inten_padded [13]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [13]),
    .o(_al_u4873_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*~B))"),
    .INIT(8'ha8))
    _al_u4874 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/mux4_b10_sel_is_4_o ),
    .b(_al_u4872_o),
    .c(_al_u4873_o),
    .o(_al_u4874_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*~A)"),
    .INIT(16'h4000))
    _al_u4875 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [10]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [11]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [7]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [13]),
    .o(_al_u4875_o));
  AL_MAP_LUT4 #(
    .EQN("~(C*~((D*~A))*~(B)+C*(D*~A)*~(B)+~(C)*(D*~A)*B+C*(D*~A)*B)"),
    .INIT(16'h8bcf))
    _al_u4876 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpol_padded [13]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[13] ),
    .o(_al_u4876_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~B*~(~D*A))"),
    .INIT(16'h0301))
    _al_u4877 (
    .a(_al_u1983_o),
    .b(_al_u4874_o),
    .c(_al_u4875_o),
    .d(_al_u4876_o),
    .o(_al_u4877_o));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u4878 (
    .a(_al_u1986_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inten_padded [13]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttype_padded [13]),
    .o(_al_u4878_o));
  AL_MAP_LUT4 #(
    .EQN("~(C*~((D*~A))*~(B)+C*(D*~A)*~(B)+~(C)*(D*~A)*B+C*(D*~A)*B)"),
    .INIT(16'h8bcf))
    _al_u4879 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpol_padded [13]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [13]),
    .o(_al_u4879_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*A*~(C*B))"),
    .INIT(16'h002a))
    _al_u488 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n25_lutinv ),
    .b(_al_u486_o),
    .c(_al_u487_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[4] ),
    .o(_al_u488_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u4880 (
    .a(_al_u4878_o),
    .b(_al_u1982_o),
    .c(_al_u4879_o),
    .o(_al_u4880_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u4881 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4]),
    .c(\u_cmsdk_mcu/p0_outen [13]),
    .d(\u_cmsdk_mcu/p0_altfunc [13]),
    .o(_al_u4881_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D*~C*A))"),
    .INIT(16'h3133))
    _al_u4882 (
    .a(_al_u4515_o),
    .b(_al_u4881_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4]),
    .d(\u_cmsdk_mcu/p0_out [13]),
    .o(_al_u4882_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*~(~D*~C)))"),
    .INIT(16'h222a))
    _al_u4883 (
    .a(_al_u4511_o),
    .b(_al_u4880_o),
    .c(_al_u4882_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [5]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n31 [13]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4884 (
    .a(\u_cmsdk_mcu/sram_hrdata [13]),
    .b(\u_cmsdk_mcu/flash_hrdata [13]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [0]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [1]),
    .o(_al_u4884_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(D*C))"),
    .INIT(16'h0444))
    _al_u4885 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n37 [14]),
    .b(_al_u4884_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [4]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/rwdata_reg [13]),
    .o(_al_u4885_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~B*~(D*~A))"),
    .INIT(16'h2030))
    _al_u4886 (
    .a(_al_u4877_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n31 [13]),
    .c(_al_u4885_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [6]),
    .o(_al_u4886_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*B)*~(~D*A))"),
    .INIT(16'hf351))
    _al_u4887 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kq7iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pp7iu6 ),
    .c(_al_u4886_o),
    .d(_al_u1862_o),
    .o(_al_u4887_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4888 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A25iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R05iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P14qw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W2jax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U28iu6 ));
  AL_MAP_LUT4 #(
    .EQN("~(B*A*~(D*C))"),
    .INIT(16'hf777))
    _al_u4889 (
    .a(_al_u4887_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U28iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uy4iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sgjax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wgvhu6 ));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u489 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n27_lutinv ),
    .b(_al_u488_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n28 [2]),
    .o(_al_u489_o));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u4890 (
    .a(_al_u1986_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inten_padded [15]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttype_padded [15]),
    .o(_al_u4890_o));
  AL_MAP_LUT4 #(
    .EQN("~(C*~((D*~A))*~(B)+C*(D*~A)*~(B)+~(C)*(D*~A)*B+C*(D*~A)*B)"),
    .INIT(16'h8bcf))
    _al_u4891 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpol_padded [15]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [15]),
    .o(_al_u4891_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u4892 (
    .a(_al_u4890_o),
    .b(_al_u1982_o),
    .c(_al_u4891_o),
    .o(_al_u4892_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u4893 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4]),
    .c(\u_cmsdk_mcu/p0_outen [15]),
    .d(\u_cmsdk_mcu/p0_altfunc [15]),
    .o(_al_u4893_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D*~C*A))"),
    .INIT(16'h3133))
    _al_u4894 (
    .a(_al_u4515_o),
    .b(_al_u4893_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4]),
    .d(\u_cmsdk_mcu/p0_out [15]),
    .o(_al_u4894_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*~(~D*~C)))"),
    .INIT(16'h222a))
    _al_u4895 (
    .a(_al_u4511_o),
    .b(_al_u4892_o),
    .c(_al_u4894_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [5]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n31 [15]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u4896 (
    .a(_al_u1986_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inten_padded [15]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [15]),
    .o(_al_u4896_o));
  AL_MAP_LUT4 #(
    .EQN("~(C*~((D*~A))*~(B)+C*(D*~A)*~(B)+~(C)*(D*~A)*B+C*(D*~A)*B)"),
    .INIT(16'h8bcf))
    _al_u4897 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpol_padded [15]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[15] ),
    .o(_al_u4897_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u4898 (
    .a(_al_u4896_o),
    .b(_al_u1982_o),
    .c(_al_u4897_o),
    .o(_al_u4898_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h3210))
    _al_u4899 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [15]),
    .d(\u_cmsdk_mcu/p1_out [15]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/mux0_b15/B1_0 ));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*B))"),
    .INIT(8'hd5))
    _al_u490 (
    .a(_al_u489_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n7_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [2]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/read_mux_byte0 [2]));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u4900 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4]),
    .c(\u_cmsdk_mcu/p1_outen [15]),
    .d(\u_cmsdk_mcu/p1_altfunc [15]),
    .o(_al_u4900_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(~B*~(~C*A)))"),
    .INIT(16'h00ce))
    _al_u4901 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/mux0_b15/B1_0 ),
    .b(_al_u4900_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [5]),
    .o(_al_u4901_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*~A)"),
    .INIT(16'h4000))
    _al_u4902 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [10]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [11]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [9]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [15]),
    .o(_al_u4902_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(A*~(~C*B)))"),
    .INIT(16'h005d))
    _al_u4903 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/mux4_b10_sel_is_4_o ),
    .b(_al_u4898_o),
    .c(_al_u4901_o),
    .d(_al_u4902_o),
    .o(_al_u4903_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4904 (
    .a(\u_cmsdk_mcu/sram_hrdata [15]),
    .b(\u_cmsdk_mcu/flash_hrdata [15]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [0]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [1]),
    .o(_al_u4904_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(D*C))"),
    .INIT(16'h0444))
    _al_u4905 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n37 [14]),
    .b(_al_u4904_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [4]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/rwdata_reg [15]),
    .o(_al_u4905_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*~(D*~B))"),
    .INIT(16'h4050))
    _al_u4906 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n31 [15]),
    .b(_al_u4903_o),
    .c(_al_u4905_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [6]),
    .o(_al_u4906_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u4907 (
    .a(_al_u4906_o),
    .b(_al_u4533_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sn7iu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u4908 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M15iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uy4iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sn7iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sejax6 ),
    .o(_al_u4908_o));
  AL_MAP_LUT4 #(
    .EQN("~((D*~A)*~(C)*~(B)+(D*~A)*C*~(B)+~((D*~A))*C*B+(D*~A)*C*B)"),
    .INIT(16'h2e3f))
    _al_u4909 (
    .a(_al_u4500_o),
    .b(_al_u4501_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z54iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9ypw6 ),
    .o(_al_u4909_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'h0a0c))
    _al_u491 (
    .a(uart0_txen_pad),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_rx_buf [0]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] ),
    .o(_al_u491_o));
  AL_MAP_LUT4 #(
    .EQN("(C*A*~(D*B))"),
    .INIT(16'h20a0))
    _al_u4910 (
    .a(_al_u4908_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A25iu6 ),
    .c(_al_u4909_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W8hbx6 ),
    .o(_al_u4910_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(~C*B))"),
    .INIT(8'h5d))
    _al_u4911 (
    .a(_al_u4910_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kq7iu6 ),
    .c(_al_u1865_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rhvhu6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u4912 (
    .a(_al_u4368_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J71iu6_lutinv ),
    .o(_al_u4912_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u4913 (
    .a(_al_u4912_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ay8iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/My0iu6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u4914 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E4yhu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qehbx6 ),
    .o(_al_u4914_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~((D*~C))*~(A)+B*(D*~C)*~(A)+~(B)*(D*~C)*A+B*(D*~C)*A)"),
    .INIT(16'h4e44))
    _al_u4915 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xg6iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/My0iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wqzhu6 ),
    .d(_al_u4914_o),
    .o(\u_cmsdk_mcu/HADDR [0]));
  AL_MAP_LUT4 #(
    .EQN("(A*~(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B))"),
    .INIT(16'h20a8))
    _al_u4916 (
    .a(_al_u4552_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xg6iu6 ),
    .c(_al_u4086_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bvfbx6 ),
    .o(_al_u4916_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u4917 (
    .a(_al_u4916_o),
    .b(_al_u4548_o),
    .c(_al_u4553_o),
    .o(_al_u4917_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u4918 (
    .a(_al_u4071_o),
    .b(_al_u4076_o),
    .c(_al_u4081_o),
    .o(_al_u4918_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u4919 (
    .a(_al_u4918_o),
    .b(_al_u4061_o),
    .c(_al_u4066_o),
    .o(_al_u4919_o));
  AL_MAP_LUT4 #(
    .EQN("(C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'ha0c0))
    _al_u492 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/apbsubsys_interrupt [1]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_buf_full ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] ),
    .o(_al_u492_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u4920 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jl3qw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ym3qw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yubbx6 ),
    .o(_al_u4920_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u4921 (
    .a(_al_u4920_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nwdbx6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufebx6 ),
    .o(_al_u4921_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u4922 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xg6iu6 ),
    .b(_al_u4919_o),
    .c(_al_u4921_o),
    .o(_al_u4922_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B))"),
    .INIT(16'h20a8))
    _al_u4923 (
    .a(_al_u4922_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xg6iu6 ),
    .c(_al_u4056_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dpwpw6 ),
    .o(_al_u4923_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u4924 (
    .a(_al_u4917_o),
    .b(_al_u4923_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/apbsys_hsel ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*~(B)*C*D)"),
    .INIT(16'h11f7))
    _al_u4925 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Am6iu6_lutinv ),
    .b(_al_u4438_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pg3qw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvabx6 ),
    .o(_al_u4925_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u4926 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dpwpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jl3qw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ym3qw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yubbx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mz6iu6 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C@B))"),
    .INIT(8'h82))
    _al_u4927 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mz6iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ad7ax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvabx6 ),
    .o(_al_u4927_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u4928 (
    .a(_al_u4927_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kl8ax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Su8ax6 ),
    .o(_al_u4928_o));
  AL_MAP_LUT4 #(
    .EQN("(C*A*~(D*~B))"),
    .INIT(16'h80a0))
    _al_u4929 (
    .a(_al_u4925_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Am6iu6_lutinv ),
    .c(_al_u4928_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pg3qw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X87iu6 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*~B))"),
    .INIT(8'ha8))
    _al_u493 (
    .a(_al_u473_o),
    .b(_al_u491_o),
    .c(_al_u492_o),
    .o(_al_u493_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*B*C*D)"),
    .INIT(16'h4b4d))
    _al_u4930 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Am6iu6_lutinv ),
    .b(_al_u4438_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bf3qw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pg3qw6 ),
    .o(_al_u4930_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*~A)"),
    .INIT(8'h04))
    _al_u4931 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kl8ax6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Su8ax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvabx6 ),
    .o(_al_u4931_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*~A)"),
    .INIT(16'h0040))
    _al_u4932 (
    .a(_al_u4930_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mz6iu6 ),
    .c(_al_u4931_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ad7ax6 ),
    .o(_al_u4932_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u4933 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ad7ax6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kl8ax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvabx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nw6iu6 ));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u4934 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Su8ax6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ym3qw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yubbx6 ),
    .o(_al_u4934_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u4935 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nw6iu6 ),
    .b(_al_u4934_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dpwpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jl3qw6 ),
    .o(_al_u4935_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u4936 (
    .a(_al_u4935_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pg3qw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J17iu6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(~D*~(~C*~A)))"),
    .INIT(16'h3301))
    _al_u4937 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X87iu6 ),
    .b(_al_u4932_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J17iu6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bf3qw6 ),
    .o(_al_u4937_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u4938 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nd3qw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vn9bx6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yf1qw6 ),
    .o(_al_u4938_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*~A)"),
    .INIT(16'h0004))
    _al_u4939 (
    .a(_al_u4937_o),
    .b(_al_u4938_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H4ypw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ke1qw6 ),
    .o(_al_u4939_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u494 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n7_lutinv ),
    .b(_al_u493_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [0]),
    .o(_al_u494_o));
  AL_MAP_LUT4 #(
    .EQN("(A*(B*~(C)*~(D)+~(B)*C*~(D)+B*~(C)*D))"),
    .INIT(16'h0828))
    _al_u4940 (
    .a(_al_u4927_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kl8ax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Su8ax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvabx6 ),
    .o(_al_u4940_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*~B)*~(~D*A))"),
    .INIT(16'hfc54))
    _al_u4941 (
    .a(_al_u4438_o),
    .b(_al_u4940_o),
    .c(_al_u4935_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bf3qw6 ),
    .o(_al_u4941_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(~C*~(D*B)))"),
    .INIT(16'ha8a0))
    _al_u4942 (
    .a(_al_u4941_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Am6iu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bf3qw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pg3qw6 ),
    .o(_al_u4942_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(D*C*~B))"),
    .INIT(16'h4555))
    _al_u4943 (
    .a(_al_u4942_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Am6iu6_lutinv ),
    .c(_al_u4438_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J17iu6_lutinv ),
    .o(_al_u4943_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*~A)"),
    .INIT(16'h4000))
    _al_u4944 (
    .a(_al_u4943_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nd3qw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vn9bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yf1qw6 ),
    .o(_al_u4944_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u4945 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nd3qw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pg3qw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vn9bx6 ),
    .o(_al_u4945_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(B*~A))"),
    .INIT(8'h0b))
    _al_u4946 (
    .a(_al_u4438_o),
    .b(_al_u4938_o),
    .c(_al_u4945_o),
    .o(_al_u4946_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(B@A))"),
    .INIT(8'h09))
    _al_u4947 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bf3qw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pg3qw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Su8ax6 ),
    .o(_al_u4947_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u4948 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nw6iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mz6iu6 ),
    .c(_al_u4947_o),
    .o(_al_u4948_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~A*~(~C*~B))"),
    .INIT(16'h5400))
    _al_u4949 (
    .a(_al_u4946_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Am6iu6_lutinv ),
    .c(_al_u4438_o),
    .d(_al_u4948_o),
    .o(_al_u4949_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*B))"),
    .INIT(8'hd5))
    _al_u495 (
    .a(_al_u494_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n27_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n28 [0]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/read_mux_byte0 [0]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u4950 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B79bx6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H4ypw6 ),
    .o(_al_u4950_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(D*~(~C*~B)))"),
    .INIT(16'h0155))
    _al_u4951 (
    .a(_al_u4939_o),
    .b(_al_u4944_o),
    .c(_al_u4949_o),
    .d(_al_u4950_o),
    .o(_al_u4951_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*A)"),
    .INIT(16'h0002))
    _al_u4952 (
    .a(_al_u4549_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bvfbx6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H7hbx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q4dbx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fs6iu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~(~B*A))"),
    .INIT(16'h000d))
    _al_u4953 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B79bx6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ke1qw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nwdbx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufebx6 ),
    .o(_al_u4953_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*~A)"),
    .INIT(16'h1000))
    _al_u4954 (
    .a(_al_u4951_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qc3pw6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fs6iu6 ),
    .d(_al_u4953_o),
    .o(_al_u4954_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*B))"),
    .INIT(8'ha2))
    _al_u4955 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nr4iu6_lutinv ),
    .b(_al_u4954_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Su8ax6 ),
    .o(_al_u4955_o));
  AL_MAP_LUT3 #(
    .EQN("~(~A*~(C*B))"),
    .INIT(8'hea))
    _al_u4956 (
    .a(_al_u4955_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hw8ax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y1xhu6 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*B))"),
    .INIT(8'ha2))
    _al_u4957 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nr4iu6_lutinv ),
    .b(_al_u4954_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yf1qw6 ),
    .o(_al_u4957_o));
  AL_MAP_LUT3 #(
    .EQN("~(~A*~(C*B))"),
    .INIT(8'hea))
    _al_u4958 (
    .a(_al_u4957_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Le2qw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F2xhu6 ));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*~(D@C)))"),
    .INIT(16'h2aa2))
    _al_u4959 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nr4iu6_lutinv ),
    .b(_al_u4954_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ad7ax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vn9bx6 ),
    .o(_al_u4959_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u496 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [9]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [10]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [11]),
    .o(_al_u496_o));
  AL_MAP_LUT3 #(
    .EQN("~(~A*~(C*B))"),
    .INIT(8'hea))
    _al_u4960 (
    .a(_al_u4959_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pe7ax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M2xhu6 ));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*(D@C)))"),
    .INIT(16'ha22a))
    _al_u4961 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nr4iu6_lutinv ),
    .b(_al_u4954_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Am6iu6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Su8ax6 ),
    .o(_al_u4961_o));
  AL_MAP_LUT3 #(
    .EQN("~(~A*~(C*B))"),
    .INIT(8'hea))
    _al_u4962 (
    .a(_al_u4961_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D43qw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T2xhu6 ));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*(D@C)))"),
    .INIT(16'ha22a))
    _al_u4963 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nr4iu6_lutinv ),
    .b(_al_u4954_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Am6iu6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pg3qw6 ),
    .o(_al_u4963_o));
  AL_MAP_LUT3 #(
    .EQN("~(~A*~(C*B))"),
    .INIT(8'hea))
    _al_u4964 (
    .a(_al_u4963_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Di3qw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A3xhu6 ));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*~(D@C)))"),
    .INIT(16'h2aa2))
    _al_u4965 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nr4iu6_lutinv ),
    .b(_al_u4954_o),
    .c(_al_u4438_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kl8ax6 ),
    .o(_al_u4965_o));
  AL_MAP_LUT3 #(
    .EQN("~(~A*~(C*B))"),
    .INIT(8'hea))
    _al_u4966 (
    .a(_al_u4965_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zm8ax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H3xhu6 ));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*~(D@C)))"),
    .INIT(16'h2aa2))
    _al_u4967 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nr4iu6_lutinv ),
    .b(_al_u4954_o),
    .c(_al_u4438_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bf3qw6 ),
    .o(_al_u4967_o));
  AL_MAP_LUT3 #(
    .EQN("~(~A*~(C*B))"),
    .INIT(8'hea))
    _al_u4968 (
    .a(_al_u4967_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sqwpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O3xhu6 ));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*B*A)"),
    .INIT(16'h0800))
    _al_u4969 (
    .a(_al_u4545_o),
    .b(_al_u4546_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/HADDR[27]_lutinv ),
    .d(_al_u4553_o),
    .o(_al_u4969_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u497 (
    .a(_al_u496_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [7]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [8]),
    .o(_al_u497_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*B*A)"),
    .INIT(16'h0800))
    _al_u4970 (
    .a(_al_u4923_o),
    .b(_al_u4969_o),
    .c(\u_cmsdk_mcu/HADDR [12]),
    .d(_al_u4544_o),
    .o(_al_u4970_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u4971 (
    .a(\u_cmsdk_mcu/HADDR [15]),
    .b(\u_cmsdk_mcu/HADDR [14]),
    .c(\u_cmsdk_mcu/HADDR [13]),
    .o(_al_u4971_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u4972 (
    .a(_al_u4916_o),
    .b(_al_u4970_o),
    .c(_al_u4971_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/sysrom_hsel ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u4973 (
    .a(\u_cmsdk_mcu/HADDR [13]),
    .b(\u_cmsdk_mcu/HADDR [12]),
    .o(_al_u4973_o));
  AL_MAP_LUT4 #(
    .EQN("(A*(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B))"),
    .INIT(16'h8a02))
    _al_u4974 (
    .a(_al_u4922_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xg6iu6 ),
    .c(_al_u4056_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dpwpw6 ),
    .o(_al_u4974_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u4975 (
    .a(_al_u4973_o),
    .b(_al_u4974_o),
    .c(\u_cmsdk_mcu/HADDR [15]),
    .d(\u_cmsdk_mcu/HADDR [14]),
    .o(_al_u4975_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u4976 (
    .a(_al_u4917_o),
    .b(_al_u4975_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/sysctrl_hsel ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u4977 (
    .a(_al_u4971_o),
    .b(_al_u4974_o),
    .o(_al_u4977_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u4978 (
    .a(_al_u4917_o),
    .b(_al_u4977_o),
    .c(\u_cmsdk_mcu/HADDR [12]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio1_hsel ));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u4979 (
    .a(_al_u4917_o),
    .b(_al_u4977_o),
    .c(\u_cmsdk_mcu/HADDR [12]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_hsel ));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u498 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [4]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [5]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [6]),
    .o(_al_u498_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(C*~A))"),
    .INIT(16'h8caf))
    _al_u4980 (
    .a(_al_u4539_o),
    .b(_al_u4912_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iiliu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ay8iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z18iu6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(D*~(~A*~(C*B)))"),
    .INIT(16'hea00))
    _al_u4981 (
    .a(_al_u3618_o),
    .b(_al_u1346_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Difiu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 ),
    .o(_al_u4981_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u4982 (
    .a(_al_u1266_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pthiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 ),
    .o(_al_u4982_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D*C*A))"),
    .INIT(16'h1333))
    _al_u4983 (
    .a(_al_u695_o),
    .b(_al_u4982_o),
    .c(_al_u1582_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Edapw6_lutinv ),
    .o(_al_u4983_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*~A)"),
    .INIT(16'h0004))
    _al_u4984 (
    .a(_al_u4981_o),
    .b(_al_u4983_o),
    .c(_al_u3187_o),
    .d(_al_u3995_o),
    .o(_al_u4984_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*~A))"),
    .INIT(8'h8c))
    _al_u4985 (
    .a(_al_u3103_o),
    .b(_al_u2868_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 ),
    .o(_al_u4985_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u4986 (
    .a(_al_u1266_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 ),
    .o(_al_u4986_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~A*~(~D*C))"),
    .INIT(16'h1101))
    _al_u4987 (
    .a(_al_u3118_o),
    .b(_al_u4986_o),
    .c(_al_u1271_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 ),
    .o(_al_u4987_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(D*C*~B))"),
    .INIT(16'h4555))
    _al_u4988 (
    .a(_al_u4985_o),
    .b(_al_u4987_o),
    .c(_al_u1269_o),
    .d(_al_u1342_o),
    .o(_al_u4988_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(~B*~(~D*~C)))"),
    .INIT(16'h888a))
    _al_u4989 (
    .a(_al_u4984_o),
    .b(_al_u4988_o),
    .c(_al_u3103_o),
    .d(_al_u1342_o),
    .o(_al_u4989_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u499 (
    .a(_al_u498_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_byte_strobe [0]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_write_enable ),
    .o(_al_u499_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(~D*~(B*~A)))"),
    .INIT(16'hf040))
    _al_u4990 (
    .a(_al_u4989_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V3xhu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vygax6 ),
    .o(_al_u4990_o));
  AL_MAP_LUT4 #(
    .EQN("~(~C*~(~D*~B*~A))"),
    .INIT(16'hf0f1))
    _al_u4991 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z18iu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n1465 ),
    .c(_al_u4990_o),
    .d(_al_u3797_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U8vhu6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u4992 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z18iu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S18iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E18iu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*B)*~(~D*A))"),
    .INIT(16'hf351))
    _al_u4993 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xg6iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W7cow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I7cow6 ),
    .d(_al_u4495_o),
    .o(_al_u4993_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*~A)"),
    .INIT(16'h0100))
    _al_u4994 (
    .a(_al_u3885_o),
    .b(_al_u3887_o),
    .c(_al_u3889_o),
    .d(_al_u4197_o),
    .o(_al_u4994_o));
  AL_MAP_LUT4 #(
    .EQN("~(B*~(~D*~C*A))"),
    .INIT(16'h333b))
    _al_u4995 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E18iu6 ),
    .b(_al_u4993_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W7cow6 ),
    .d(_al_u4994_o),
    .o(\u_cmsdk_mcu/HTRANS [1]));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u4996 (
    .a(\u_cmsdk_mcu/HADDR [0]),
    .b(\u_cmsdk_mcu/HADDR [1]),
    .o(\u_cmsdk_mcu/u_ahb_ram/n5 [0]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*~A))"),
    .INIT(8'hdc))
    _al_u4997 (
    .a(\u_cmsdk_mcu/HADDR [0]),
    .b(\u_cmsdk_mcu/HSIZE [1]),
    .c(\u_cmsdk_mcu/HADDR [1]),
    .o(\u_cmsdk_mcu/u_ahb_ram/n5 [16]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u4998 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio1_hsel ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_ahb_to_gpio/n0 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u4999 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_hsel ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_ahb_to_gpio/n0 ));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*B*A)"),
    .INIT(16'h0800))
    _al_u500 (
    .a(_al_u497_o),
    .b(_al_u499_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [2]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [3]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_lockupreset_write ));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(~D*C*B))"),
    .INIT(16'h5515))
    _al_u5000 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nr4iu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E18iu6 ),
    .c(_al_u4994_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n1465 ),
    .o(_al_u5000_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u5001 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wjyiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rzciu6_lutinv ),
    .o(_al_u5001_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~((D*C))*~(A)+B*(D*C)*~(A)+~(B)*(D*C)*A+B*(D*C)*A)"),
    .INIT(16'he444))
    _al_u5002 (
    .a(_al_u5000_o),
    .b(\u_cmsdk_mcu/HWRITE ),
    .c(_al_u5001_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C1wpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hyuhu6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u5003 (
    .a(\u_cmsdk_mcu/HTRANS [1]),
    .b(\u_cmsdk_mcu/HWRITE ),
    .o(_al_u5003_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u5004 (
    .a(\u_cmsdk_mcu/flash_hsel ),
    .b(_al_u5003_o),
    .o(\u_cmsdk_mcu/u_ahb_rom/n2 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0a5c))
    _al_u5005 (
    .a(_al_u4490_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iqzhu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sqfax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uofax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pkhpw6 [0]));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u5006 (
    .a(\u_cmsdk_mcu/HSIZE [0]),
    .b(\u_cmsdk_mcu/HADDR [0]),
    .o(_al_u5006_o));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(~C*~A))"),
    .INIT(8'hcd))
    _al_u5007 (
    .a(_al_u5006_o),
    .b(\u_cmsdk_mcu/HSIZE [1]),
    .c(\u_cmsdk_mcu/HADDR [1]),
    .o(\u_cmsdk_mcu/u_ahb_ram/n5 [10]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*~A))"),
    .INIT(8'hdc))
    _al_u5008 (
    .a(_al_u5006_o),
    .b(\u_cmsdk_mcu/HSIZE [1]),
    .c(\u_cmsdk_mcu/HADDR [1]),
    .o(\u_cmsdk_mcu/u_ahb_ram/n5 [24]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u5009 (
    .a(\u_cmsdk_mcu/HTRANS [1]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ),
    .o(_al_u5009_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    _al_u501 (
    .a(_al_u497_o),
    .b(_al_u499_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [2]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [3]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_remap_write ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u5010 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/sysrom_hsel ),
    .b(_al_u5009_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/trans_valid ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u5011 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/sysctrl_hsel ),
    .b(_al_u5009_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/ahb_access ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u5012 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/apbsys_hsel ),
    .b(_al_u5009_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/n1 ));
  AL_MAP_LUT3 #(
    .EQN("~(C*B*A)"),
    .INIT(8'h7f))
    _al_u5013 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V34iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iqzhu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gpqpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n382 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u5014 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/ahb_access ),
    .b(\u_cmsdk_mcu/HWRITE ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/ahb_read ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u5015 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/ahb_access ),
    .b(\u_cmsdk_mcu/HWRITE ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/ahb_write ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u5016 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/ahb_access ),
    .b(\u_cmsdk_mcu/u_ahb_ram/n5 [0]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/nxt_byte_strobe [0]));
  AL_MAP_LUT4 #(
    .EQN("(A*~(~D*~C*~B))"),
    .INIT(16'haaa8))
    _al_u5017 (
    .a(_al_u4917_o),
    .b(_al_u4975_o),
    .c(_al_u4977_o),
    .d(_al_u4923_o),
    .o(_al_u5017_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u5018 (
    .a(_al_u5017_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/sysrom_hsel ),
    .c(\u_cmsdk_mcu/flash_hsel ),
    .o(\u_cmsdk_mcu/sram_hsel ));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*~A)"),
    .INIT(8'h04))
    _al_u5019 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sf1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sq4iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J0gax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahwiu6_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+~(A)*B*~(C)+A*B*~(C)+A*B*C)"),
    .INIT(8'h8e))
    _al_u502 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cjqpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ehqpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T0ipw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yfxhu6 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*~B))"),
    .INIT(8'ha8))
    _al_u5020 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahwiu6_lutinv ),
    .b(_al_u4492_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nmfax6 ),
    .o(_al_u5020_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u5021 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vr1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ar1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dncax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F6dbx6 ),
    .o(_al_u5021_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u5022 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vowiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hw8ax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sqwpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zm8ax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iv1iu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u5023 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cs1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zt1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Krbax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z2aax6 ),
    .o(_al_u5023_o));
  AL_MAP_LUT4 #(
    .EQN("(C*A*~(D*B))"),
    .INIT(16'h20a0))
    _al_u5024 (
    .a(_al_u5021_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iv1iu6 ),
    .c(_al_u5023_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[29] ),
    .o(_al_u5024_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5025 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xs1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dw1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Peeax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Widax6 ),
    .o(_al_u5025_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u5026 (
    .a(_al_u5024_o),
    .b(_al_u5025_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kw1iu6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J59ax6 ),
    .o(_al_u5026_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u5027 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ur4iu6 ),
    .b(_al_u5001_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/St1iu6 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*~B))"),
    .INIT(8'h8a))
    _al_u5028 (
    .a(_al_u5026_o),
    .b(_al_u1286_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/St1iu6 ),
    .o(_al_u5028_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u5029 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U2fiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E1fiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qf4bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Unyax6 ),
    .o(_al_u5029_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u503 (
    .a(_al_u374_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Di3qw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Le2qw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vuciu6 ));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u5030 (
    .a(_al_u540_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ilwiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hw8ax6 ),
    .o(_al_u5030_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u5031 (
    .a(_al_u5030_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K5eiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xznow6 ),
    .o(_al_u5031_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u5032 (
    .a(_al_u5029_o),
    .b(_al_u5031_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q0fiu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E34bx6 ),
    .o(_al_u5032_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u5033 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K5eiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R9yax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W5ypw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F0eow6 ));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u5034 (
    .a(_al_u3779_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F0eow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rz0bx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fllow6_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u5035 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pjyiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R9yax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W5ypw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M0eow6 ));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u5036 (
    .a(_al_u5032_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fllow6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M0eow6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tcipw6 ),
    .o(_al_u5036_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u5037 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I3fiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G2fiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cwyax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M85bx6 ),
    .o(_al_u5037_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u5038 (
    .a(_al_u5037_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C0fiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aw4bx6 ),
    .o(_al_u5038_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5039 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tzdiu6 ),
    .b(_al_u546_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tl4bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uizax6 ),
    .o(_al_u5039_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*A)"),
    .INIT(16'h0200))
    _al_u504 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vuciu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hw8ax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sqwpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zm8ax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xs1iu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5040 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hqgiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S1fiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pczax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wgipw6 ),
    .o(_al_u5040_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u5041 (
    .a(_al_u5036_o),
    .b(_al_u5038_o),
    .c(_al_u5039_o),
    .d(_al_u5040_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bewiu6 ));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u5042 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D43qw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hw8ax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pe7ax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H2qiu6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u5043 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iv1iu6 ),
    .b(_al_u540_o),
    .c(_al_u1385_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H2qiu6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uvsiu6 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u5044 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uvsiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ymwiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K0xiu6 ),
    .o(_al_u5044_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u5045 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J3xiu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H2qiu6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mmqiu6 ));
  AL_MAP_LUT4 #(
    .EQN("(A*~(~D*~C*B))"),
    .INIT(16'haaa2))
    _al_u5046 (
    .a(_al_u5044_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mmqiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Di3qw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Le2qw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yw1iu6 ));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D*C*B))"),
    .INIT(16'h2aaa))
    _al_u5047 (
    .a(_al_u5020_o),
    .b(_al_u5028_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bewiu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yw1iu6 ),
    .o(_al_u5047_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u5048 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iqzhu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nmfax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nrqpw6 ),
    .o(_al_u5048_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*~(~D*B))"),
    .INIT(16'h5010))
    _al_u5049 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sf1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sq4iu6 ),
    .c(_al_u5048_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J0gax6 ),
    .o(_al_u5049_o));
  AL_MAP_LUT2 #(
    .EQN("~(B*A)"),
    .INIT(4'h7))
    _al_u505 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xs1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dg2qw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Td7iu6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u5050 (
    .a(_al_u5049_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gpqpw6 ),
    .o(_al_u5050_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~A*~(D*C))"),
    .INIT(16'h0111))
    _al_u5051 (
    .a(_al_u5047_o),
    .b(_al_u5050_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sf1iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X42qw6 ),
    .o(_al_u5051_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u5052 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahwiu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nmfax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nrqpw6 ),
    .o(_al_u5052_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u5053 (
    .a(_al_u5052_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gpqpw6 ),
    .o(_al_u5053_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*B))"),
    .INIT(8'hd5))
    _al_u5054 (
    .a(_al_u5051_o),
    .b(_al_u5053_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wc2qw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S6phu6 ));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u5055 (
    .a(_al_u5050_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sf1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rr3qw6 ),
    .o(_al_u5055_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u5056 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zt1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kw1iu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tchbx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wahbx6 ),
    .o(_al_u5056_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    _al_u5057 (
    .a(_al_u533_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hw8ax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sqwpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zm8ax6 ),
    .o(_al_u5057_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*A*~(D*B))"),
    .INIT(16'h020a))
    _al_u5058 (
    .a(_al_u5056_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ar1iu6 ),
    .c(_al_u5057_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sx3qw6 ),
    .o(_al_u5058_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u5059 (
    .a(_al_u3779_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F0eow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kojpw6 ),
    .o(_al_u5059_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u506 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sqwpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zm8ax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J3xiu6_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u5060 (
    .a(_al_u5059_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M0eow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bc3bx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U6wiu6 ));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u5061 (
    .a(_al_u5058_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U6wiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iv1iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[28] ),
    .o(_al_u5061_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*~C))"),
    .INIT(16'h8088))
    _al_u5062 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yw1iu6 ),
    .b(_al_u5061_o),
    .c(_al_u1862_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/St1iu6 ),
    .o(_al_u5062_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*B))"),
    .INIT(8'ha2))
    _al_u5063 (
    .a(_al_u5055_o),
    .b(_al_u5020_o),
    .c(_al_u5062_o),
    .o(_al_u5063_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*B))"),
    .INIT(8'hd5))
    _al_u5064 (
    .a(_al_u5063_o),
    .b(_al_u5053_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cq3qw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z6phu6 ));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u5065 (
    .a(_al_u3779_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F0eow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Usipw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pwfow6_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u5066 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pwfow6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M0eow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V73bx6 ),
    .o(_al_u5066_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u5067 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K5eiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dtjow6 ),
    .o(_al_u5067_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u5068 (
    .a(_al_u5066_o),
    .b(_al_u5067_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mnmpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I0wiu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u5069 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xs1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vr1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bngax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yogax6 ),
    .o(_al_u5069_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u507 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vuciu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J3xiu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hw8ax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vr1iu6 ));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u5070 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I0wiu6 ),
    .b(_al_u5069_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zt1iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Khgax6 ),
    .o(_al_u5070_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u5071 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cs1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kw1iu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hjgax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nfgax6 ),
    .o(_al_u5071_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u5072 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dw1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ar1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Elgax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ibqpw6 ),
    .o(_al_u5072_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*~(D*A))"),
    .INIT(16'h40c0))
    _al_u5073 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iv1iu6 ),
    .b(_al_u5071_o),
    .c(_al_u5072_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[27] ),
    .o(_al_u5073_o));
  AL_MAP_LUT4 #(
    .EQN("(C*A*~(~D*B))"),
    .INIT(16'ha020))
    _al_u5074 (
    .a(_al_u5070_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/St1iu6 ),
    .c(_al_u5073_o),
    .d(_al_u1859_o),
    .o(_al_u5074_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u5075 (
    .a(_al_u5020_o),
    .b(_al_u5074_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yw1iu6 ),
    .o(_al_u5075_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u5076 (
    .a(_al_u5075_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sf1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idqpw6 ),
    .o(_al_u5076_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*B))"),
    .INIT(8'hd5))
    _al_u5077 (
    .a(_al_u5076_o),
    .b(_al_u5053_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vqgax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G7phu6 ));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u5078 (
    .a(_al_u3779_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F0eow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qx0bx6 ),
    .o(_al_u5078_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u5079 (
    .a(_al_u5078_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M0eow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P33bx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wtviu6 ));
  AL_MAP_LUT2 #(
    .EQN("~(B*A)"),
    .INIT(4'h7))
    _al_u508 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vr1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dg2qw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Md7iu6 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*A))"),
    .INIT(8'hc4))
    _al_u5080 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/St1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wtviu6 ),
    .c(_al_u1856_o),
    .o(_al_u5080_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u5081 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cs1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kw1iu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cxcbx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Itcbx6 ),
    .o(_al_u5081_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u5082 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xs1iu6 ),
    .b(_al_u5081_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W0dbx6 ),
    .o(_al_u5082_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5083 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vr1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ar1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nybbx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T2dbx6 ),
    .o(_al_u5083_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5084 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dw1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zt1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fvcbx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zycbx6 ),
    .o(_al_u5084_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u5085 (
    .a(_al_u5082_o),
    .b(_al_u5083_o),
    .c(_al_u5084_o),
    .o(_al_u5085_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u5086 (
    .a(_al_u5080_o),
    .b(_al_u5085_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iv1iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[26] ),
    .o(_al_u5086_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u5087 (
    .a(_al_u5020_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yw1iu6 ),
    .c(_al_u5086_o),
    .o(_al_u5087_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u5088 (
    .a(_al_u5087_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sf1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N0cbx6 ),
    .o(_al_u5088_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*B))"),
    .INIT(8'hd5))
    _al_u5089 (
    .a(_al_u5088_o),
    .b(_al_u5053_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q4dbx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N7phu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    _al_u509 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D43qw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Di3qw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Le2qw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pe7ax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Avwiu6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u5090 (
    .a(_al_u5049_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gpqpw6 ),
    .o(_al_u5090_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u5091 (
    .a(_al_u5090_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sf1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cncbx6 ),
    .o(_al_u5091_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u5092 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M0eow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F0eow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jz2bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X5upw6 ),
    .o(_al_u5092_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u5093 (
    .a(_al_u5092_o),
    .b(_al_u5067_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zdtpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wmviu6 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*A))"),
    .INIT(8'hc4))
    _al_u5094 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/St1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wmviu6 ),
    .c(_al_u1854_o),
    .o(_al_u5094_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5095 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cs1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kw1iu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Facbx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zdcbx6 ),
    .o(_al_u5095_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u5096 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xs1iu6 ),
    .b(_al_u5095_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Thcbx6 ),
    .o(_al_u5096_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5097 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vr1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ar1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F8cbx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qjcbx6 ),
    .o(_al_u5097_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5098 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dw1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zt1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cccbx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wfcbx6 ),
    .o(_al_u5098_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u5099 (
    .a(_al_u5096_o),
    .b(_al_u5097_o),
    .c(_al_u5098_o),
    .o(_al_u5099_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u510 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J3xiu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Avwiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hw8ax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dw1iu6 ));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u5100 (
    .a(_al_u5094_o),
    .b(_al_u5099_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iv1iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[25] ),
    .o(_al_u5100_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*~(D*C)))"),
    .INIT(16'ha222))
    _al_u5101 (
    .a(_al_u5091_o),
    .b(_al_u5020_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yw1iu6 ),
    .d(_al_u5100_o),
    .o(_al_u5101_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*B))"),
    .INIT(8'hd5))
    _al_u5102 (
    .a(_al_u5101_o),
    .b(_al_u5053_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nlcbx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U7phu6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u5103 (
    .a(_al_u5052_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gpqpw6 ),
    .o(_al_u5103_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u5104 (
    .a(_al_u5103_o),
    .b(_al_u5052_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q2ibx6 ),
    .o(_al_u5104_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u5105 (
    .a(_al_u3779_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F0eow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pv0bx6 ),
    .o(_al_u5105_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u5106 (
    .a(_al_u5105_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M0eow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rm2bx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wfviu6 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*A))"),
    .INIT(8'hc4))
    _al_u5107 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/St1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wfviu6 ),
    .c(_al_u1852_o),
    .o(_al_u5107_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5108 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xs1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cs1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Htbax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tkdax6 ),
    .o(_al_u5108_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u5109 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vr1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dw1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Apcax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mgeax6 ),
    .o(_al_u5109_o));
  AL_MAP_LUT2 #(
    .EQN("~(B*A)"),
    .INIT(4'h7))
    _al_u511 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dw1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dg2qw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae7iu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u5110 (
    .a(_al_u927_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ar1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nj2qw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nwbbx6 ),
    .o(_al_u5110_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5111 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zt1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kw1iu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G79ax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4aax6 ),
    .o(_al_u5111_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u5112 (
    .a(_al_u5108_o),
    .b(_al_u5109_o),
    .c(_al_u5110_o),
    .d(_al_u5111_o),
    .o(_al_u5112_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u5113 (
    .a(_al_u5107_o),
    .b(_al_u5112_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iv1iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[24] ),
    .o(_al_u5113_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u5114 (
    .a(_al_u5020_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yw1iu6 ),
    .c(_al_u5113_o),
    .o(_al_u5114_o));
  AL_MAP_LUT4 #(
    .EQN("~(~B*A*~(D*C))"),
    .INIT(16'hfddd))
    _al_u5115 (
    .a(_al_u5104_o),
    .b(_al_u5114_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sf1iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fl2qw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B8phu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5116 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vr1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cs1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Evbax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xqcax6 ),
    .o(_al_u5116_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u5117 (
    .a(_al_u5116_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dw1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jieax6 ),
    .o(_al_u5117_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5118 (
    .a(_al_u927_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zt1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T6aax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uh2qw6 ),
    .o(_al_u5118_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u5119 (
    .a(_al_u5118_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eg7iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F4ibx6 ),
    .o(_al_u5119_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*A)"),
    .INIT(16'h0200))
    _al_u512 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Avwiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hw8ax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sqwpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zm8ax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cs1iu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5120 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xs1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kw1iu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D99ax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qmdax6 ),
    .o(_al_u5120_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u5121 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yc7iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ar1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sbfax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgkbx6 ),
    .o(_al_u5121_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u5122 (
    .a(_al_u5117_o),
    .b(_al_u5119_o),
    .c(_al_u5120_o),
    .d(_al_u5121_o),
    .o(_al_u5122_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u5123 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M0eow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F0eow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dv2bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oxkpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jgeow6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u5124 (
    .a(_al_u5031_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jgeow6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P8viu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5125 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ws4iu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iv1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[23] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vpkpw6 ),
    .o(_al_u5125_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*~(~D*A))"),
    .INIT(16'hc040))
    _al_u5126 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/St1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P8viu6 ),
    .c(_al_u5125_o),
    .d(_al_u1850_o),
    .o(_al_u5126_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D*C*B))"),
    .INIT(16'h2aaa))
    _al_u5127 (
    .a(_al_u5020_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yw1iu6 ),
    .c(_al_u5122_o),
    .d(_al_u5126_o),
    .o(_al_u5127_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u5128 (
    .a(_al_u5127_o),
    .b(_al_u5052_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/No3qw6 ),
    .o(_al_u5128_o));
  AL_MAP_LUT4 #(
    .EQN("~(~B*A*~(D*C))"),
    .INIT(16'hfddd))
    _al_u5129 (
    .a(_al_u5128_o),
    .b(_al_u5103_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sf1iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nrkpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I8phu6 ));
  AL_MAP_LUT2 #(
    .EQN("~(B*A)"),
    .INIT(4'h7))
    _al_u513 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cs1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dg2qw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/He7iu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u5130 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vr1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ar1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Etfbx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tlebx6 ),
    .o(_al_u5130_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u5131 (
    .a(_al_u5130_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xs1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hrfbx6 ),
    .o(_al_u5131_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(~C*A))"),
    .INIT(16'h31f5))
    _al_u5132 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/St1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iv1iu6 ),
    .c(_al_u1846_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[21] ),
    .o(_al_u5132_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u5133 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dw1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zt1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kpfbx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qlfbx6 ),
    .o(_al_u5133_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u5134 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cs1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kw1iu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nnfbx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tjfbx6 ),
    .o(_al_u5134_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u5135 (
    .a(_al_u5131_o),
    .b(_al_u5132_o),
    .c(_al_u5133_o),
    .d(_al_u5134_o),
    .o(_al_u5135_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5136 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M0eow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F0eow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B3gbx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y0gbx6 ),
    .o(_al_u5136_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5137 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I3fiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvgiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F9gbx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tngbx6 ),
    .o(_al_u5137_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u5138 (
    .a(_al_u5136_o),
    .b(_al_u5137_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S1fiu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nhgbx6 ),
    .o(_al_u5138_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u5139 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rk1bx6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rm2bx6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tcipw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U31bx6 ),
    .o(_al_u5139_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u514 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J3xiu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Avwiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hw8ax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zt1iu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u5140 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P12bx6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P33bx6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qo3bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rijbx6 ),
    .o(_al_u5140_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u5141 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xq2bx6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y0gbx6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yxrpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z71bx6 ),
    .o(_al_u5141_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u5142 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Us3bx6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V52bx6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V73bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xo1bx6 ),
    .o(_al_u5142_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u5143 (
    .a(_al_u5139_o),
    .b(_al_u5140_o),
    .c(_al_u5141_o),
    .d(_al_u5142_o),
    .o(_al_u5143_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u5144 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fc1bx6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fe2bx6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gihbx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hg3bx6 ),
    .o(_al_u5144_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u5145 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aa2bx6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bc3bx6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dt1bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dv2bx6 ),
    .o(_al_u5145_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u5146 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lr9bx6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mk3bx6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Muhbx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5bbx6 ),
    .o(_al_u5146_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u5147 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jx1bx6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jz2bx6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lg1bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Li2bx6 ),
    .o(_al_u5147_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u5148 (
    .a(_al_u5144_o),
    .b(_al_u5145_o),
    .c(_al_u5146_o),
    .d(_al_u5147_o),
    .o(_al_u5148_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u5149 (
    .a(_al_u5067_o),
    .b(_al_u5143_o),
    .c(_al_u5148_o),
    .o(_al_u5149_o));
  AL_MAP_LUT2 #(
    .EQN("~(B*A)"),
    .INIT(4'h7))
    _al_u515 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zt1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dg2qw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qf7iu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u5150 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6eiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E1fiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D7gbx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lfgbx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zpkow6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5151 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q0fiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C0fiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hbgbx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jdgbx6 ),
    .o(_al_u5151_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    _al_u5152 (
    .a(_al_u5149_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zpkow6 ),
    .c(_al_u5151_o),
    .o(_al_u5152_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5153 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hqgiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tzdiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C5gbx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vpgbx6 ),
    .o(_al_u5153_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5154 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U2fiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G2fiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pjgbx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rlgbx6 ),
    .o(_al_u5154_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u5155 (
    .a(_al_u5138_o),
    .b(_al_u5152_o),
    .c(_al_u5153_o),
    .d(_al_u5154_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ntuiu6 ));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D*C*B))"),
    .INIT(16'h2aaa))
    _al_u5156 (
    .a(_al_u5020_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yw1iu6 ),
    .c(_al_u5135_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ntuiu6 ),
    .o(_al_u5156_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~A*~(D*C))"),
    .INIT(16'h0111))
    _al_u5157 (
    .a(_al_u5156_o),
    .b(_al_u5090_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sf1iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qwfbx6 ),
    .o(_al_u5157_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*B))"),
    .INIT(8'hd5))
    _al_u5158 (
    .a(_al_u5157_o),
    .b(_al_u5053_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bvfbx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W8phu6 ));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u5159 (
    .a(_al_u5090_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sf1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jhebx6 ),
    .o(_al_u5159_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u516 (
    .a(_al_u374_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J3xiu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hw8ax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gkwiu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u5160 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M0eow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F0eow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Li2bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nr0bx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mdfow6 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u5161 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mdfow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvgiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tjkpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fdfow6 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u5162 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fdfow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6eiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rhkpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Umuiu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5163 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vr1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kw1iu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M4ebx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xdebx6 ),
    .o(_al_u5163_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u5164 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Umuiu6 ),
    .b(_al_u5163_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xs1iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Acebx6 ),
    .o(_al_u5164_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u5165 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zt1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ar1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J6ebx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M2ebx6 ),
    .o(_al_u5165_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u5166 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dw1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cs1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Daebx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G8ebx6 ),
    .o(_al_u5166_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*~(D*A))"),
    .INIT(16'h40c0))
    _al_u5167 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iv1iu6 ),
    .b(_al_u5165_o),
    .c(_al_u5166_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[20] ),
    .o(_al_u5167_o));
  AL_MAP_LUT4 #(
    .EQN("(C*A*~(~D*B))"),
    .INIT(16'ha020))
    _al_u5168 (
    .a(_al_u5164_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/St1iu6 ),
    .c(_al_u5167_o),
    .d(_al_u1844_o),
    .o(_al_u5168_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*~(D*C)))"),
    .INIT(16'ha222))
    _al_u5169 (
    .a(_al_u5159_o),
    .b(_al_u5020_o),
    .c(_al_u5168_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yw1iu6 ),
    .o(_al_u5169_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u517 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gkwiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Di3qw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Le2qw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eg7iu6 ));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*B))"),
    .INIT(8'hd5))
    _al_u5170 (
    .a(_al_u5169_o),
    .b(_al_u5053_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufebx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D9phu6 ));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u5171 (
    .a(_al_u5090_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sf1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cydbx6 ),
    .o(_al_u5171_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u5172 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M0eow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F0eow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fe2bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mp0bx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mrfow6 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u5173 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mrfow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6eiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X6jpw6 ),
    .o(_al_u5173_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u5174 (
    .a(_al_u5173_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvgiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z8jpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bguiu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u5175 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vr1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cs1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qudbx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zodbx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hcuiu6 ));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u5176 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bguiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hcuiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kw1iu6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fldbx6 ),
    .o(_al_u5176_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(~C*A))"),
    .INIT(16'h31f5))
    _al_u5177 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/St1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iv1iu6 ),
    .c(_al_u1841_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[19] ),
    .o(_al_u5177_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5178 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xs1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zt1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cndbx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tsdbx6 ),
    .o(_al_u5178_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5179 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dw1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ar1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fjdbx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wqdbx6 ),
    .o(_al_u5179_o));
  AL_MAP_LUT2 #(
    .EQN("~(B*A)"),
    .INIT(4'h7))
    _al_u518 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eg7iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dg2qw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xf7iu6 ));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u5180 (
    .a(_al_u5176_o),
    .b(_al_u5177_o),
    .c(_al_u5178_o),
    .d(_al_u5179_o),
    .o(_al_u5180_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*~(D*C)))"),
    .INIT(16'ha222))
    _al_u5181 (
    .a(_al_u5171_o),
    .b(_al_u5020_o),
    .c(_al_u5180_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yw1iu6 ),
    .o(_al_u5181_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*B))"),
    .INIT(8'hd5))
    _al_u5182 (
    .a(_al_u5181_o),
    .b(_al_u5053_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nwdbx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K9phu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5183 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M0eow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F0eow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ln0bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V52bx6 ),
    .o(_al_u5183_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u5184 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6eiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvgiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hhvpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nr7ax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E5jow6 ));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u5185 (
    .a(_al_u5031_o),
    .b(_al_u5183_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E5jow6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U8uiu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5186 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cs1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kw1iu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ab9ax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bxbax6 ),
    .o(_al_u5186_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u5187 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U8uiu6 ),
    .b(_al_u5186_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zt1iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q8aax6 ),
    .o(_al_u5187_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5188 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vr1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dw1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gkeax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uscax6 ),
    .o(_al_u5188_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u5189 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xs1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ar1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nodax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T6kbx6 ),
    .o(_al_u5189_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u519 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[2] ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[3] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M8row6_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*~B))"),
    .INIT(8'ha8))
    _al_u5190 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iv1iu6 ),
    .b(_al_u1385_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[18] ),
    .o(_al_u5190_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*A)"),
    .INIT(16'h0080))
    _al_u5191 (
    .a(_al_u5187_o),
    .b(_al_u5188_o),
    .c(_al_u5189_o),
    .d(_al_u5190_o),
    .o(_al_u5191_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*~B))"),
    .INIT(8'h8a))
    _al_u5192 (
    .a(_al_u5191_o),
    .b(_al_u1839_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/St1iu6 ),
    .o(_al_u5192_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(C*~(D*~B)))"),
    .INIT(16'h2a0a))
    _al_u5193 (
    .a(_al_u5020_o),
    .b(_al_u4284_o),
    .c(_al_u5192_o),
    .d(_al_u927_o),
    .o(_al_u5193_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~A*~(D*C))"),
    .INIT(16'h0111))
    _al_u5194 (
    .a(_al_u5193_o),
    .b(_al_u5050_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sf1iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gbvpw6 ),
    .o(_al_u5194_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*B))"),
    .INIT(8'hd5))
    _al_u5195 (
    .a(_al_u5194_o),
    .b(_al_u5053_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ym3qw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R9phu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u5196 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zt1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kw1iu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Naaax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xc9ax6 ),
    .o(_al_u5196_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u5197 (
    .a(_al_u5196_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cs1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yybax6 ),
    .o(_al_u5197_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*~B))"),
    .INIT(8'ha8))
    _al_u5198 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iv1iu6 ),
    .b(_al_u1385_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[17] ),
    .o(_al_u5198_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u5199 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vr1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ar1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rucax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Syjbx6 ),
    .o(_al_u5199_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*~B*A)"),
    .INIT(16'h0020))
    _al_u520 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M8row6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[4] ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[1] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[5] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B0biu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5200 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xs1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dw1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dmeax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kqdax6 ),
    .o(_al_u5200_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u5201 (
    .a(_al_u5197_o),
    .b(_al_u5198_o),
    .c(_al_u5199_o),
    .d(_al_u5200_o),
    .o(_al_u5201_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u5202 (
    .a(_al_u3779_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F0eow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kl0bx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hbpow6_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u5203 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hbpow6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M0eow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P12bx6 ),
    .o(_al_u5203_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u5204 (
    .a(_al_u5031_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvgiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N0xpw6 ),
    .o(_al_u5204_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u5205 (
    .a(_al_u5203_o),
    .b(_al_u5204_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6eiu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lywpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U1uiu6 ));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*~C))"),
    .INIT(16'h8088))
    _al_u5206 (
    .a(_al_u5201_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U1uiu6 ),
    .c(_al_u1836_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/St1iu6 ),
    .o(_al_u5206_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(C*~(D*~B)))"),
    .INIT(16'h2a0a))
    _al_u5207 (
    .a(_al_u5020_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qa5iu6 ),
    .c(_al_u5206_o),
    .d(_al_u927_o),
    .o(_al_u5207_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~A*~(D*C))"),
    .INIT(16'h0111))
    _al_u5208 (
    .a(_al_u5207_o),
    .b(_al_u5049_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sf1iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kswpw6 ),
    .o(_al_u5208_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*B))"),
    .INIT(8'hd5))
    _al_u5209 (
    .a(_al_u5208_o),
    .b(_al_u5053_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jl3qw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y9phu6 ));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    _al_u521 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R9yax6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W5ypw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztupw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dtjow6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5210 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M0eow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F0eow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D70bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lg1bx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fviow6 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u5211 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fviow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvgiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pt7ax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yuiow6 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u5212 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yuiow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6eiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ofmpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uosiu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u5213 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vr1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dw1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F59bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N19bx6 ),
    .o(_al_u5213_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u5214 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uosiu6 ),
    .b(_al_u5213_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zt1iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ux8bx6 ),
    .o(_al_u5214_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*~B))"),
    .INIT(8'ha8))
    _al_u5215 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iv1iu6 ),
    .b(_al_u1385_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[10] ),
    .o(_al_u5215_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5216 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xs1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ar1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C07bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J39bx6 ),
    .o(_al_u5216_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u5217 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cs1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kw1iu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rz8bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xv8bx6 ),
    .o(_al_u5217_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u5218 (
    .a(_al_u5214_o),
    .b(_al_u5215_o),
    .c(_al_u5216_o),
    .d(_al_u5217_o),
    .o(_al_u5218_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(C*~(D*~B)))"),
    .INIT(16'h2a0a))
    _al_u5219 (
    .a(_al_u5020_o),
    .b(_al_u4796_o),
    .c(_al_u5218_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/St1iu6 ),
    .o(_al_u5219_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u522 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pjyiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dtjow6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I3fiu6 ));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u5220 (
    .a(_al_u5219_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sf1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bu6bx6 ),
    .o(_al_u5220_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*B))"),
    .INIT(8'hd5))
    _al_u5221 (
    .a(_al_u5220_o),
    .b(_al_u5053_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B79bx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vbphu6 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*~B))"),
    .INIT(8'ha8))
    _al_u5222 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iv1iu6 ),
    .b(_al_u1385_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[9] ),
    .o(_al_u5222_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5223 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xs1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dw1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oveax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzdax6 ),
    .o(_al_u5223_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5224 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zt1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yc7iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hdfax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yjaax6 ),
    .o(_al_u5224_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    _al_u5225 (
    .a(_al_u5222_o),
    .b(_al_u5223_o),
    .c(_al_u5224_o),
    .o(_al_u5225_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5226 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M0eow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F0eow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C50bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fc1bx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L9mow6 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u5227 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L9mow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvgiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vrtpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E9mow6 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u5228 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E9mow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6eiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tptpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bisiu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u5229 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vr1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ar1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C4dax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gwxpw6 ),
    .o(_al_u5229_o));
  AL_MAP_LUT2 #(
    .EQN("~(B*A)"),
    .INIT(4'h7))
    _al_u523 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I3fiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C1wpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B3fiu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5230 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cs1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kw1iu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Im9ax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J8cax6 ),
    .o(_al_u5230_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u5231 (
    .a(_al_u5225_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bisiu6 ),
    .c(_al_u5229_o),
    .d(_al_u5230_o),
    .o(_al_u5231_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(C*~(D*~B)))"),
    .INIT(16'h2a0a))
    _al_u5232 (
    .a(_al_u5020_o),
    .b(_al_u4776_o),
    .c(_al_u5231_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/St1iu6 ),
    .o(_al_u5232_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u5233 (
    .a(_al_u5232_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sf1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gyxpw6 ),
    .o(_al_u5233_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*B))"),
    .INIT(8'hd5))
    _al_u5234 (
    .a(_al_u5233_o),
    .b(_al_u5053_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H4ypw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ccphu6 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*~B))"),
    .INIT(8'ha8))
    _al_u5235 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iv1iu6 ),
    .b(_al_u1385_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[8] ),
    .o(_al_u5235_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5236 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vr1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dw1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B9jbx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tcjbx6 ),
    .o(_al_u5236_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u5237 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zt1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ar1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J5jbx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kn1qw6 ),
    .o(_al_u5237_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    _al_u5238 (
    .a(_al_u5235_o),
    .b(_al_u5236_o),
    .c(_al_u5237_o),
    .o(_al_u5238_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5239 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xs1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kw1iu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N3jbx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xajbx6 ),
    .o(_al_u5239_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u524 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vynow6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dtjow6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E1fiu6 ));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u5240 (
    .a(_al_u5238_o),
    .b(_al_u5239_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cs1iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F7jbx6 ),
    .o(_al_u5240_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u5241 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M0eow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F0eow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rijbx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tkjbx6 ),
    .o(_al_u5241_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u5242 (
    .a(_al_u5241_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rzciu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dtjow6 ),
    .o(_al_u5242_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u5243 (
    .a(_al_u5031_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6eiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tmjbx6 ),
    .o(_al_u5243_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u5244 (
    .a(_al_u5242_o),
    .b(_al_u5243_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvgiu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uojbx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ibsiu6 ));
  AL_MAP_LUT4 #(
    .EQN("(C*B*~(D*~A))"),
    .INIT(16'h80c0))
    _al_u5245 (
    .a(_al_u4756_o),
    .b(_al_u5240_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ibsiu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/St1iu6 ),
    .o(_al_u5245_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(~C*A))"),
    .INIT(16'h31f5))
    _al_u5246 (
    .a(_al_u5020_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sf1iu6 ),
    .c(_al_u5245_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mh1qw6 ),
    .o(_al_u5246_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C*A))"),
    .INIT(8'hb3))
    _al_u5247 (
    .a(_al_u5053_o),
    .b(_al_u5246_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yf1qw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jcphu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5248 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M0eow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F0eow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C30bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Us3bx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dzdow6 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u5249 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dzdow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvgiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ss0qw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wydow6 ));
  AL_MAP_LUT2 #(
    .EQN("~(B*A)"),
    .INIT(4'h7))
    _al_u525 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E1fiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C1wpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X0fiu6 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u5250 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wydow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6eiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rq0qw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4siu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5251 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vr1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dw1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kxeax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y5dax6 ),
    .o(_al_u5251_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u5252 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4siu6 ),
    .b(_al_u5251_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zt1iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vlaax6 ),
    .o(_al_u5252_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*~B))"),
    .INIT(8'ha8))
    _al_u5253 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iv1iu6 ),
    .b(_al_u1385_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[7] ),
    .o(_al_u5253_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5254 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xs1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ar1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N61qw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R1eax6 ),
    .o(_al_u5254_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u5255 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cs1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kw1iu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Facax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fo9ax6 ),
    .o(_al_u5255_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u5256 (
    .a(_al_u5252_o),
    .b(_al_u5253_o),
    .c(_al_u5254_o),
    .d(_al_u5255_o),
    .o(_al_u5256_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(C*~(D*~B)))"),
    .INIT(16'h2a0a))
    _al_u5257 (
    .a(_al_u5020_o),
    .b(_al_u4836_o),
    .c(_al_u5256_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/St1iu6 ),
    .o(_al_u5257_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u5258 (
    .a(_al_u5257_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sf1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M81qw6 ),
    .o(_al_u5258_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*B))"),
    .INIT(8'hd5))
    _al_u5259 (
    .a(_al_u5258_o),
    .b(_al_u5053_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ke1qw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qcphu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(B*~(~D*~C)))"),
    .INIT(16'h1115))
    _al_u526 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n265 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iqzhu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gnqpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J0gax6 ),
    .o(_al_u526_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u5260 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vynow6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R9yax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W5ypw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztupw6 ),
    .o(_al_u5260_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u5261 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M0eow6 ),
    .b(_al_u5260_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qo3bx6 ),
    .o(_al_u5261_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5262 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q0fiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C0fiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sn4bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wu3bx6 ),
    .o(_al_u5262_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u5263 (
    .a(_al_u5261_o),
    .b(_al_u5262_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F0eow6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C10bx6 ),
    .o(_al_u5263_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5264 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6eiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I3fiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S3mpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Thxax6 ),
    .o(_al_u5264_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5265 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tzdiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E1fiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mfyax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yqzax6 ),
    .o(_al_u5265_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u5266 (
    .a(_al_u5263_o),
    .b(_al_u5264_o),
    .c(_al_u5265_o),
    .o(_al_u5266_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u5267 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G2fiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvgiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E05bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ujxax6 ),
    .o(_al_u5267_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u5268 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S1fiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U2fiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H4zax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I74bx6 ),
    .o(_al_u5268_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u5269 (
    .a(_al_u5266_o),
    .b(_al_u5267_o),
    .c(_al_u5268_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pxriu6 ));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*~(~D*~C)))"),
    .INIT(16'h222a))
    _al_u527 (
    .a(_al_u526_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iqzhu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nmfax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nrqpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V34iu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    _al_u5270 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hw8ax6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Le2qw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sqwpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zm8ax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wyqiu6 ));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u5271 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wyqiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D43qw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pe7ax6 ),
    .o(_al_u5271_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(C*A))"),
    .INIT(16'h5f13))
    _al_u5272 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iv1iu6 ),
    .b(_al_u5271_o),
    .c(_al_u1385_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Di3qw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wzpiu6 ));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u5273 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K0xiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ilwiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Le2qw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iqriu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(~A*~(C*B)))"),
    .INIT(16'h00ea))
    _al_u5274 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iqriu6 ),
    .b(_al_u374_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wyqiu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Di3qw6 ),
    .o(_al_u5274_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u5275 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Di3qw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Le2qw6 ),
    .o(_al_u5275_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(~A*~(D*B)))"),
    .INIT(16'he0a0))
    _al_u5276 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cvciu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K0xiu6 ),
    .c(_al_u5275_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pe7ax6 ),
    .o(_al_u5276_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u5277 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wzpiu6 ),
    .b(_al_u5274_o),
    .c(_al_u5276_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F0riu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5278 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vr1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ar1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Asupw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U7dax6 ),
    .o(_al_u5278_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u5279 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Di3qw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Le2qw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A2qiu6 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u528 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V34iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iqzhu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gpqpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M24iu6 ));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u5280 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K0xiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A2qiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D43qw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pe7ax6 ),
    .o(_al_u5280_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(~D*C*B))"),
    .INIT(16'h5515))
    _al_u5281 (
    .a(_al_u5280_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cvciu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A2qiu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D43qw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lariu6 ));
  AL_MAP_LUT4 #(
    .EQN("(C*A*~(D*B))"),
    .INIT(16'h20a0))
    _al_u5282 (
    .a(_al_u5278_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xs1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lariu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N3eax6 ),
    .o(_al_u5282_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5283 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dw1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kw1iu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bq9ax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gzeax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tsriu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u5284 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cs1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zt1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bccax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rnaax6 ),
    .o(_al_u5284_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*~(D*A))"),
    .INIT(16'h40c0))
    _al_u5285 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iv1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tsriu6 ),
    .c(_al_u5284_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[6] ),
    .o(_al_u5285_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u5286 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pxriu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F0riu6 ),
    .c(_al_u5282_o),
    .d(_al_u5285_o),
    .o(_al_u5286_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(C*~(D*~B)))"),
    .INIT(16'h2a0a))
    _al_u5287 (
    .a(_al_u5020_o),
    .b(_al_u4735_o),
    .c(_al_u5286_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/St1iu6 ),
    .o(_al_u5287_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u5288 (
    .a(_al_u5287_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sf1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nckbx6 ),
    .o(_al_u5288_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*B))"),
    .INIT(8'hd5))
    _al_u5289 (
    .a(_al_u5288_o),
    .b(_al_u5053_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nd3qw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xcphu6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u529 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bclpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sdlpw6 ),
    .o(_al_u529_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u5290 (
    .a(_al_u5275_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sqwpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zm8ax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ffqiu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*A)"),
    .INIT(16'h0080))
    _al_u5291 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ffqiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D43qw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hw8ax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pe7ax6 ),
    .o(_al_u5291_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u5292 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lariu6 ),
    .b(_al_u5291_o),
    .o(_al_u5292_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*~(~D*~C)))"),
    .INIT(16'h222a))
    _al_u5293 (
    .a(_al_u5292_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iv1iu6 ),
    .c(_al_u1385_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[5] ),
    .o(_al_u5293_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5294 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vr1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kw1iu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tc9bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zl9bx6 ),
    .o(_al_u5294_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u5295 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dw1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ar1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hi9bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ua9bx6 ),
    .o(_al_u5295_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*~(D*B))"),
    .INIT(16'h1050))
    _al_u5296 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ve7iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xs1iu6 ),
    .c(_al_u5295_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dk9bx6 ),
    .o(_al_u5296_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u5297 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cs1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zt1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lg9bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pe9bx6 ),
    .o(_al_u5297_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u5298 (
    .a(_al_u5293_o),
    .b(_al_u5294_o),
    .c(_al_u5296_o),
    .d(_al_u5297_o),
    .o(_al_u5298_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u5299 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6eiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E1fiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ox9bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T3abx6 ),
    .o(_al_u5299_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*(C@(D*A)))"),
    .INIT(16'h1230))
    _al_u530 (
    .a(_al_u529_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jflpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kalpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yklpw6 ),
    .o(_al_u530_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u5300 (
    .a(_al_u5299_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I3fiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bcabx6 ),
    .o(_al_u5300_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u5301 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M0eow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F0eow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lr9bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nt9bx6 ),
    .o(_al_u5301_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5302 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S1fiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q0fiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R1abx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V5abx6 ),
    .o(_al_u5302_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u5303 (
    .a(_al_u5301_o),
    .b(_al_u5302_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tzdiu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nv9bx6 ),
    .o(_al_u5303_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5304 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G2fiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvgiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rv7ax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X7abx6 ),
    .o(_al_u5304_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5305 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U2fiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C0fiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pz9bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z9abx6 ),
    .o(_al_u5305_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u5306 (
    .a(_al_u5300_o),
    .b(_al_u5303_o),
    .c(_al_u5304_o),
    .d(_al_u5305_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kkriu6 ));
  AL_MAP_LUT4 #(
    .EQN("(C*B*~(D*~A))"),
    .INIT(16'h80c0))
    _al_u5307 (
    .a(_al_u4712_o),
    .b(_al_u5298_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kkriu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/St1iu6 ),
    .o(_al_u5307_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*B)*~(D*A))"),
    .INIT(16'h51f3))
    _al_u5308 (
    .a(_al_u5052_o),
    .b(_al_u5020_o),
    .c(_al_u5307_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vn9bx6 ),
    .o(_al_u5308_o));
  AL_MAP_LUT4 #(
    .EQN("~(B*~A*~(D*C))"),
    .INIT(16'hfbbb))
    _al_u5309 (
    .a(_al_u5103_o),
    .b(_al_u5308_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sf1iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vefax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Edphu6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u531 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahlpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pmlpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U5yhu6 ));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u5310 (
    .a(_al_u5090_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sf1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ceabx6 ),
    .o(_al_u5310_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u5311 (
    .a(_al_u5292_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iv1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[4] ),
    .o(_al_u5311_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5312 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M0eow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F0eow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Czzax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mk3bx6 ),
    .o(_al_u5312_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5313 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6eiu6 ),
    .b(_al_u5067_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[5] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X5opw6 ),
    .o(_al_u5313_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u5314 (
    .a(_al_u5312_o),
    .b(_al_u5313_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvgiu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y7opw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eariu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u5315 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vr1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kw1iu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q9dax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xr9ax6 ),
    .o(_al_u5315_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u5316 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eariu6 ),
    .b(_al_u5315_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zt1iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Npaax6 ),
    .o(_al_u5316_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5317 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xs1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dw1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C1fax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J5eax6 ),
    .o(_al_u5317_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5318 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cs1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ar1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qc5bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xdcax6 ),
    .o(_al_u5318_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u5319 (
    .a(_al_u5311_o),
    .b(_al_u5316_o),
    .c(_al_u5317_o),
    .d(_al_u5318_o),
    .o(_al_u5319_o));
  AL_MAP_LUT2 #(
    .EQN("~(B*A)"),
    .INIT(4'h7))
    _al_u532 (
    .a(_al_u530_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U5yhu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U03iu6 ));
  AL_MAP_LUT4 #(
    .EQN("(C*B*~(D*~A))"),
    .INIT(16'h80c0))
    _al_u5320 (
    .a(_al_u4688_o),
    .b(_al_u5319_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F0riu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/St1iu6 ),
    .o(_al_u5320_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*B))"),
    .INIT(8'ha2))
    _al_u5321 (
    .a(_al_u5310_o),
    .b(_al_u5020_o),
    .c(_al_u5320_o),
    .o(_al_u5321_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*B))"),
    .INIT(8'hd5))
    _al_u5322 (
    .a(_al_u5321_o),
    .b(_al_u5053_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bf3qw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ldphu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u5323 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M0eow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F0eow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Muhbx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Owhbx6 ),
    .o(_al_u5323_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*A*~(D*C))"),
    .INIT(16'h0222))
    _al_u5324 (
    .a(_al_u5323_o),
    .b(_al_u5260_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rzciu6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dtjow6 ),
    .o(_al_u5324_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u5325 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6eiu6 ),
    .b(_al_u5067_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oyhbx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[3] ),
    .o(_al_u5325_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u5326 (
    .a(_al_u5324_o),
    .b(_al_u5325_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvgiu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0ibx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tmqiu6 ));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u5327 (
    .a(_al_u374_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fnwiu6 ),
    .c(_al_u5275_o),
    .o(_al_u5327_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u5328 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fgpiu6 ),
    .b(_al_u5327_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Thiax6 ),
    .o(_al_u5328_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u5329 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bt2qw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gr2qw6 ),
    .o(_al_u5329_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*A)"),
    .INIT(16'h0002))
    _al_u533 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D43qw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Di3qw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Le2qw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pe7ax6 ),
    .o(_al_u533_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5330 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vr1iu6 ),
    .b(_al_u927_o),
    .c(_al_u5329_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iddax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ogqiu6 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*~B))"),
    .INIT(8'ha8))
    _al_u5331 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iv1iu6 ),
    .b(_al_u1385_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[2] ),
    .o(_al_u5331_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*A)"),
    .INIT(16'h0080))
    _al_u5332 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tmqiu6 ),
    .b(_al_u5328_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ogqiu6 ),
    .d(_al_u5331_o),
    .o(_al_u5332_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u5333 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xs1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jf7iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B9eax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgbax6 ),
    .o(_al_u5333_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5334 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dw1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ar1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T5yax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U4fax6 ),
    .o(_al_u5334_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5335 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cs1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sg7iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P9bax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Phcax6 ),
    .o(_al_u5335_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u5336 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zt1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kw1iu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ftaax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pv9ax6 ),
    .o(_al_u5336_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u5337 (
    .a(_al_u5333_o),
    .b(_al_u5334_o),
    .c(_al_u5335_o),
    .d(_al_u5336_o),
    .o(_al_u5337_o));
  AL_MAP_LUT3 #(
    .EQN("(~(A)*~(B)*~(C)+A*B*~(C)+~(A)*~(B)*C+~(A)*B*C+A*B*C)"),
    .INIT(8'hd9))
    _al_u5338 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D43qw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hw8ax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pe7ax6 ),
    .o(_al_u5338_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u5339 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A2qiu6 ),
    .b(_al_u5338_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sqwpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zm8ax6 ),
    .o(_al_u5339_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u534 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hw8ax6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sqwpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zm8ax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cvciu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(~D*C*A))"),
    .INIT(16'h3313))
    _al_u5340 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ffqiu6 ),
    .b(_al_u5339_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ilwiu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hw8ax6 ),
    .o(_al_u5340_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u5341 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mmqiu6 ),
    .b(_al_u5275_o),
    .o(_al_u5341_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u5342 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J3xiu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ilwiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hw8ax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Le2qw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q3qiu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~B*A*~(D*C))"),
    .INIT(16'h0222))
    _al_u5343 (
    .a(_al_u5340_o),
    .b(_al_u5341_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q3qiu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Di3qw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vvpiu6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(D*(A*~(B)*~(C)+~(A)*B*~(C)+A*~(B)*C+~(A)*B*C+A*B*C))"),
    .INIT(16'he600))
    _al_u5344 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D43qw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hw8ax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pe7ax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zm8ax6 ),
    .o(_al_u5344_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*B*~(~D*~A))"),
    .INIT(16'h0c08))
    _al_u5345 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H2qiu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A2qiu6 ),
    .c(_al_u5344_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zm8ax6 ),
    .o(_al_u5345_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u5346 (
    .a(_al_u5345_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sqwpw6 ),
    .o(_al_u5346_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*A)"),
    .INIT(16'h0080))
    _al_u5347 (
    .a(_al_u5332_o),
    .b(_al_u5337_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vvpiu6_lutinv ),
    .d(_al_u5346_o),
    .o(_al_u5347_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*~(D*~C)))"),
    .INIT(16'h2a22))
    _al_u5348 (
    .a(_al_u5020_o),
    .b(_al_u5347_o),
    .c(_al_u4637_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/St1iu6 ),
    .o(_al_u5348_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u5349 (
    .a(_al_u5348_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sf1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xu2qw6 ),
    .o(_al_u5349_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u535 (
    .a(_al_u533_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cvciu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yc7iu6 ));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*B))"),
    .INIT(8'hd5))
    _al_u5350 (
    .a(_al_u5349_o),
    .b(_al_u5053_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P23qw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zdphu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u5351 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xs1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jf7iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahdax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dfbax6 ),
    .o(_al_u5351_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u5352 (
    .a(_al_u5351_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vr1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hlcax6 ),
    .o(_al_u5352_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*B)*~(D*A))"),
    .INIT(16'h51f3))
    _al_u5353 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dw1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q3qiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Di3qw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tceax6 ),
    .o(_al_u5353_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u5354 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zt1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kw1iu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bvaax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lx9ax6 ),
    .o(_al_u5354_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u5355 (
    .a(_al_u5352_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wzpiu6 ),
    .c(_al_u5353_o),
    .d(_al_u5354_o),
    .o(_al_u5355_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u5356 (
    .a(_al_u927_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gr2qw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K0qiu6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u5357 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K0qiu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eg7iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fm7ax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0bax6 ),
    .o(_al_u5357_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5358 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fgpiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cs1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Opbax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rkbax6 ),
    .o(_al_u5358_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u5359 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ws4iu6_lutinv ),
    .b(_al_u5345_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vz8ax6 ),
    .o(_al_u5359_o));
  AL_MAP_LUT2 #(
    .EQN("~(B*A)"),
    .INIT(4'h7))
    _al_u536 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yc7iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dg2qw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rc7iu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u5360 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sg7iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ar1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T7bax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xrxax6 ),
    .o(_al_u5360_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u5361 (
    .a(_al_u5358_o),
    .b(_al_u5359_o),
    .c(_al_u5360_o),
    .o(_al_u5361_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u5362 (
    .a(_al_u5357_o),
    .b(_al_u5361_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iv1iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[1] ),
    .o(_al_u5362_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u5363 (
    .a(_al_u5346_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ffqiu6 ),
    .c(_al_u5338_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qaqiu6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u5364 (
    .a(_al_u405_o),
    .b(_al_u5260_o),
    .o(_al_u5364_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5365 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M0eow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F0eow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L1bbx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5bbx6 ),
    .o(_al_u5365_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5366 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6eiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fpgiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I2zax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vlxax6 ),
    .o(_al_u5366_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5367 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvgiu6 ),
    .b(_al_u5067_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[2] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kzabx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dooow6 ));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u5368 (
    .a(_al_u5364_o),
    .b(_al_u5365_o),
    .c(_al_u5366_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dooow6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jaqiu6 ));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u5369 (
    .a(_al_u5355_o),
    .b(_al_u5362_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qaqiu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jaqiu6 ),
    .o(_al_u5369_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u537 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hw8ax6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sqwpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zm8ax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K0xiu6 ));
  AL_MAP_LUT4 #(
    .EQN("(A*~(C*~(D*~B)))"),
    .INIT(16'h2a0a))
    _al_u5370 (
    .a(_al_u5020_o),
    .b(_al_u4611_o),
    .c(_al_u5369_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/St1iu6 ),
    .o(_al_u5370_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u5371 (
    .a(_al_u5370_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sf1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hg7ax6 ),
    .o(_al_u5371_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*B))"),
    .INIT(8'hd5))
    _al_u5372 (
    .a(_al_u5371_o),
    .b(_al_u5053_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xn7ax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gephu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u5373 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vr1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cs1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bcgax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K6gax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mq1iu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u5374 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dw1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kw1iu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H8gax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q2gax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uu1iu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u5375 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zt1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ar1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N4gax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Usnpw6 ),
    .o(_al_u5375_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*~(D*A))"),
    .INIT(16'h40c0))
    _al_u5376 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iv1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uu1iu6 ),
    .c(_al_u5375_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[30] ),
    .o(_al_u5376_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u5377 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mq1iu6 ),
    .b(_al_u5376_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xs1iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eagax6 ),
    .o(_al_u5377_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*~B))"),
    .INIT(8'h8a))
    _al_u5378 (
    .a(_al_u5377_o),
    .b(_al_u1865_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/St1iu6 ),
    .o(_al_u5378_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u5379 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M0eow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F0eow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hg3bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S0kbx6 ),
    .o(_al_u5379_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u538 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Avwiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K0xiu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jf7iu6 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u5380 (
    .a(_al_u5379_o),
    .b(_al_u5067_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pdyax6 ),
    .o(_al_u5380_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5381 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tzdiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I3fiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eyyax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgzax6 ),
    .o(_al_u5381_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5382 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E1fiu6 ),
    .b(_al_u546_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uj4bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wpyax6 ),
    .o(_al_u5382_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u5383 (
    .a(_al_u5380_o),
    .b(_al_u5381_o),
    .c(_al_u5382_o),
    .o(_al_u5383_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5384 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hqgiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C0fiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cy4bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Elnpw6 ),
    .o(_al_u5384_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u5385 (
    .a(_al_u5384_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S1fiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rezax6 ),
    .o(_al_u5385_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u5386 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q0fiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G2fiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G54bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oa5bx6 ),
    .o(_al_u5386_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~B*~(D*A))"),
    .INIT(16'h0103))
    _al_u5387 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U2fiu6 ),
    .b(_al_u3779_o),
    .c(_al_u5260_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sh4bx6 ),
    .o(_al_u5387_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u5388 (
    .a(_al_u5383_o),
    .b(_al_u5385_o),
    .c(_al_u5386_o),
    .d(_al_u5387_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rw1iu6 ));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D*C*B))"),
    .INIT(16'h2aaa))
    _al_u5389 (
    .a(_al_u5020_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yw1iu6 ),
    .c(_al_u5378_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rw1iu6 ),
    .o(_al_u5389_o));
  AL_MAP_LUT2 #(
    .EQN("~(B*A)"),
    .INIT(4'h7))
    _al_u539 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jf7iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dg2qw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cf7iu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~B*~A*~(D*C))"),
    .INIT(16'h0111))
    _al_u5390 (
    .a(_al_u5389_o),
    .b(_al_u5050_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sf1iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uunpw6 ),
    .o(_al_u5390_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*B))"),
    .INIT(8'hd5))
    _al_u5391 (
    .a(_al_u5390_o),
    .b(_al_u5053_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydgax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H2yhu6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u5392 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E18iu6 ),
    .b(_al_u4368_o),
    .o(_al_u5392_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u5393 (
    .a(_al_u5392_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L18iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xipiu6 ));
  AL_MAP_LUT4 #(
    .EQN("(A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .INIT(16'ha280))
    _al_u5394 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xipiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fnpiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L2bax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tyaax6 ),
    .o(_al_u5394_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u5395 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gr2qw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0bax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sbfax6 ),
    .o(_al_u5395_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u5396 (
    .a(_al_u5395_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lbbax6 ),
    .o(_al_u5396_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u5397 (
    .a(_al_u5396_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P9bax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nvkbx6 [7]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u5398 (
    .a(_al_u5395_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T7bax6 ),
    .o(_al_u5398_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u5399 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L2bax6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tyaax6 ),
    .o(_al_u5399_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*~A)"),
    .INIT(16'h0100))
    _al_u540 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Di3qw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Le2qw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sqwpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zm8ax6 ),
    .o(_al_u540_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*A*~(~C*B))"),
    .INIT(16'h00a2))
    _al_u5400 (
    .a(_al_u5398_o),
    .b(_al_u5399_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[0] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X5bax6 ),
    .o(_al_u5400_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*~(~D*~A))"),
    .INIT(16'hc080))
    _al_u5401 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hz0iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nvkbx6 [7]),
    .c(_al_u5400_o),
    .d(_al_u5399_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Chkhu6 ));
  AL_MAP_LUT4 #(
    .EQN("(A@(D*~(~C*~B)))"),
    .INIT(16'h56aa))
    _al_u5402 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Chkhu6 ),
    .b(_al_u1888_o),
    .c(_al_u5399_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hz9ax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/eq1/xor_i0[1]_i1[1]_o_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u5403 (
    .a(_al_u5395_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P9bax6 ),
    .o(_al_u5403_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u5404 (
    .a(_al_u5403_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lbbax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T7bax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nvkbx6 [3]));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u5405 (
    .a(_al_u5395_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pkkbx6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X5bax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n6023_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*A)"),
    .INIT(16'h0080))
    _al_u5406 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/My0iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nvkbx6 [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n6023_lutinv ),
    .d(_al_u5399_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufkhu6 ));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u5407 (
    .a(_al_u5399_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lbbax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[3] ),
    .o(_al_u5407_o));
  AL_MAP_LUT4 #(
    .EQN("(D*B*~(~C*~A))"),
    .INIT(16'hc800))
    _al_u5408 (
    .a(_al_u5398_o),
    .b(_al_u5403_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n6023_lutinv ),
    .d(_al_u5407_o),
    .o(_al_u5408_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*A))"),
    .INIT(8'hc4))
    _al_u5409 (
    .a(_al_u4231_o),
    .b(_al_u5408_o),
    .c(_al_u5399_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Alkhu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*A)"),
    .INIT(16'h0080))
    _al_u541 (
    .a(_al_u540_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D43qw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hw8ax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pe7ax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sg7iu6 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u5410 (
    .a(_al_u5395_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T7bax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X5bax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n6021_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u5411 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n6021_lutinv ),
    .b(_al_u5395_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pkkbx6 ),
    .o(_al_u5411_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(~B*A))"),
    .INIT(8'h0d))
    _al_u5412 (
    .a(_al_u5399_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[5] ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lbbax6 ),
    .o(_al_u5412_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    _al_u5413 (
    .a(_al_u5411_o),
    .b(_al_u5403_o),
    .c(_al_u5412_o),
    .o(_al_u5413_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*A))"),
    .INIT(8'hc4))
    _al_u5414 (
    .a(_al_u4141_o),
    .b(_al_u5413_o),
    .c(_al_u5399_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qnkhu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*B)*~(D*~A))"),
    .INIT(16'ha2f3))
    _al_u5415 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Alkhu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qnkhu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tc9bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tt9ax6 ),
    .o(_al_u5415_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(~D*~C*A))"),
    .INIT(16'h3331))
    _al_u5416 (
    .a(_al_u5398_o),
    .b(_al_u5403_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pkkbx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X5bax6 ),
    .o(_al_u5416_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(~D*C))"),
    .INIT(16'h4404))
    _al_u5417 (
    .a(_al_u5416_o),
    .b(_al_u5396_o),
    .c(_al_u5399_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[7] ),
    .o(_al_u5417_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*A))"),
    .INIT(8'hc4))
    _al_u5418 (
    .a(_al_u4106_o),
    .b(_al_u5417_o),
    .c(_al_u5399_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gqkhu6 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C@B))"),
    .INIT(8'h82))
    _al_u5419 (
    .a(_al_u5415_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gqkhu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fo9ax6 ),
    .o(_al_u5419_o));
  AL_MAP_LUT2 #(
    .EQN("~(B*A)"),
    .INIT(4'h7))
    _al_u542 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sg7iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dg2qw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lg7iu6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u5420 (
    .a(_al_u5396_o),
    .b(_al_u5403_o),
    .o(_al_u5420_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u5421 (
    .a(_al_u5420_o),
    .b(_al_u5411_o),
    .o(_al_u5421_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*(~A*~(D)*~(C)+~A*D*~(C)+~(~A)*D*C+~A*D*C))"),
    .INIT(16'h3101))
    _al_u5422 (
    .a(_al_u3889_o),
    .b(_al_u5421_o),
    .c(_al_u5399_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[29] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uilhu6 ));
  AL_MAP_LUT4 #(
    .EQN("(B*(~A*~(D)*~(C)+~A*D*~(C)+~(~A)*D*C+~A*D*C))"),
    .INIT(16'hc404))
    _al_u5423 (
    .a(_al_u4121_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nvkbx6 [7]),
    .c(_al_u5399_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[6] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yokhu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*B)*~(~D*A))"),
    .INIT(16'hf351))
    _al_u5424 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uilhu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yokhu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bq9ax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J59ax6 ),
    .o(_al_u5424_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*B))"),
    .INIT(8'ha2))
    _al_u5425 (
    .a(_al_u5396_o),
    .b(_al_u5399_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[13] ),
    .o(_al_u5425_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u5426 (
    .a(_al_u5411_o),
    .b(_al_u5425_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P9bax6 ),
    .o(_al_u5426_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*A))"),
    .INIT(8'hc4))
    _al_u5427 (
    .a(_al_u4131_o),
    .b(_al_u5426_o),
    .c(_al_u5399_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cykhu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*~B)*~(D*~A))"),
    .INIT(16'h8acf))
    _al_u5428 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cykhu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yokhu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bq9ax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qkabx6 ),
    .o(_al_u5428_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u5429 (
    .a(_al_u5419_o),
    .b(_al_u5424_o),
    .c(_al_u5428_o),
    .o(_al_u5429_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u543 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wyiax6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuiax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ysiax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zqiax6 ),
    .o(_al_u543_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u5430 (
    .a(_al_u5398_o),
    .b(_al_u5403_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X5bax6 ),
    .o(_al_u5430_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u5431 (
    .a(_al_u5430_o),
    .b(_al_u5396_o),
    .o(_al_u5431_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*(~A*~(D)*~(C)+~A*D*~(C)+~(~A)*D*C+~A*D*C))"),
    .INIT(16'h3101))
    _al_u5432 (
    .a(_al_u4191_o),
    .b(_al_u5431_o),
    .c(_al_u5399_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[24] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lclhu6 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*A))"),
    .INIT(8'hc4))
    _al_u5433 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lclhu6 ),
    .b(_al_u5395_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G79ax6 ),
    .o(_al_u5433_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u5434 (
    .a(_al_u5403_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n6021_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n6006_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u5435 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n6006_lutinv ),
    .b(_al_u5396_o),
    .o(_al_u5435_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*(~A*~(D)*~(C)+~A*D*~(C)+~(~A)*D*C+~A*D*C))"),
    .INIT(16'h3101))
    _al_u5436 (
    .a(_al_u4081_o),
    .b(_al_u5435_o),
    .c(_al_u5399_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[20] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G7lhu6 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C@B))"),
    .INIT(8'h82))
    _al_u5437 (
    .a(_al_u5433_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G7lhu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M4ebx6 ),
    .o(_al_u5437_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*B))"),
    .INIT(8'ha2))
    _al_u5438 (
    .a(_al_u5396_o),
    .b(_al_u5399_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[12] ),
    .o(_al_u5438_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*~B))"),
    .INIT(8'ha8))
    _al_u5439 (
    .a(_al_u5438_o),
    .b(_al_u5403_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n6021_lutinv ),
    .o(_al_u5439_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u544 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E8iax6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W0jax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W2jax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wwiax6 ),
    .o(_al_u544_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*A))"),
    .INIT(8'hc4))
    _al_u5440 (
    .a(_al_u4126_o),
    .b(_al_u5439_o),
    .c(_al_u5399_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uwkhu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*~B)*~(D*~A))"),
    .INIT(16'h8acf))
    _al_u5441 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uwkhu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lclhu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G79ax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oi9ax6 ),
    .o(_al_u5441_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(~D*~C*B))"),
    .INIT(16'h5551))
    _al_u5442 (
    .a(_al_u5396_o),
    .b(_al_u5398_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P9bax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X5bax6 ),
    .o(_al_u5442_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*(~A*~(D)*~(C)+~A*D*~(C)+~(~A)*D*C+~A*D*C))"),
    .INIT(16'h3101))
    _al_u5443 (
    .a(_al_u4061_o),
    .b(_al_u5442_o),
    .c(_al_u5399_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[16] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A2lhu6 ));
  AL_MAP_LUT2 #(
    .EQN("~(B@A)"),
    .INIT(4'h9))
    _al_u5444 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A2lhu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qjbbx6 ),
    .o(_al_u5444_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u5445 (
    .a(_al_u5429_o),
    .b(_al_u5437_o),
    .c(_al_u5441_o),
    .d(_al_u5444_o),
    .o(_al_u5445_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u5446 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uilhu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J59ax6 ),
    .o(_al_u5446_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u5447 (
    .a(_al_u5398_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pkkbx6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X5bax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n6018_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u5448 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n6018_lutinv ),
    .b(_al_u5403_o),
    .o(_al_u5448_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u5449 (
    .a(_al_u5448_o),
    .b(_al_u5396_o),
    .o(_al_u5449_o));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B*A))"),
    .INIT(8'h8f))
    _al_u545 (
    .a(_al_u543_o),
    .b(_al_u544_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzjpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X5phu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~B*(~A*~(D)*~(C)+~A*D*~(C)+~(~A)*D*C+~A*D*C))"),
    .INIT(16'h3101))
    _al_u5450 (
    .a(_al_u4096_o),
    .b(_al_u5449_o),
    .c(_al_u5399_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[25] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sdlhu6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u5451 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sdlhu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Facbx6 ),
    .o(_al_u5451_o));
  AL_MAP_LUT3 #(
    .EQN("~(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'h2e))
    _al_u5452 (
    .a(_al_u3887_o),
    .b(_al_u5399_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[30] ),
    .o(_al_u5452_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~A*(D@C))"),
    .INIT(16'h0110))
    _al_u5453 (
    .a(_al_u5446_o),
    .b(_al_u5451_o),
    .c(_al_u5452_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q2gax6 ),
    .o(_al_u5453_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*B))"),
    .INIT(8'ha2))
    _al_u5454 (
    .a(_al_u5396_o),
    .b(_al_u5399_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[10] ),
    .o(_al_u5454_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*~B))"),
    .INIT(8'ha8))
    _al_u5455 (
    .a(_al_u5454_o),
    .b(_al_u5398_o),
    .c(_al_u5403_o),
    .o(_al_u5455_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*A))"),
    .INIT(8'hc4))
    _al_u5456 (
    .a(_al_u4116_o),
    .b(_al_u5455_o),
    .c(_al_u5399_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eukhu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*~B)*~(D@A))"),
    .INIT(16'h8a45))
    _al_u5457 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eukhu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sdlhu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Facbx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xv8bx6 ),
    .o(_al_u5457_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u5458 (
    .a(_al_u5396_o),
    .b(_al_u5398_o),
    .c(_al_u5403_o),
    .o(_al_u5458_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*(~A*~(D)*~(C)+~A*D*~(C)+~(~A)*D*C+~A*D*C))"),
    .INIT(16'h3101))
    _al_u5459 (
    .a(_al_u4101_o),
    .b(_al_u5458_o),
    .c(_al_u5399_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[26] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zelhu6 ));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*B*A)"),
    .INIT(16'h0800))
    _al_u546 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rzciu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R9yax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W5ypw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztupw6 ),
    .o(_al_u546_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u5460 (
    .a(_al_u5416_o),
    .b(_al_u5396_o),
    .o(_al_u5460_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*(~A*~(D)*~(C)+~A*D*~(C)+~(~A)*D*C+~A*D*C))"),
    .INIT(16'h3101))
    _al_u5461 (
    .a(_al_u4184_o),
    .b(_al_u5460_o),
    .c(_al_u5399_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[23] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eblhu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*B)*~(D*~A))"),
    .INIT(16'ha2f3))
    _al_u5462 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zelhu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eblhu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D99ax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Itcbx6 ),
    .o(_al_u5462_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*~A))"),
    .INIT(8'h23))
    _al_u5463 (
    .a(_al_u5411_o),
    .b(_al_u5396_o),
    .c(_al_u5403_o),
    .o(_al_u5463_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*(~A*~(D)*~(C)+~A*D*~(C)+~(~A)*D*C+~A*D*C))"),
    .INIT(16'h3101))
    _al_u5464 (
    .a(_al_u4086_o),
    .b(_al_u5463_o),
    .c(_al_u5399_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[21] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O8lhu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(C*~A))"),
    .INIT(16'haf23))
    _al_u5465 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eblhu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O8lhu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D99ax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tjfbx6 ),
    .o(_al_u5465_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u5466 (
    .a(_al_u5453_o),
    .b(_al_u5457_o),
    .c(_al_u5462_o),
    .d(_al_u5465_o),
    .o(_al_u5466_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u5467 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n6018_lutinv ),
    .b(_al_u5396_o),
    .o(_al_u5467_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u5468 (
    .a(_al_u5420_o),
    .b(_al_u5399_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[17] ),
    .o(_al_u5468_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~B*~(~D*A))"),
    .INIT(16'h3010))
    _al_u5469 (
    .a(_al_u4066_o),
    .b(_al_u5467_o),
    .c(_al_u5468_o),
    .d(_al_u5399_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I3lhu6 ));
  AL_MAP_LUT2 #(
    .EQN("~(B*A)"),
    .INIT(4'h7))
    _al_u547 (
    .a(_al_u546_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C1wpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mpgiu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(C*~A))"),
    .INIT(16'haf23))
    _al_u5470 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O8lhu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I3lhu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tjfbx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xc9ax6 ),
    .o(_al_u5470_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(~D*C))"),
    .INIT(16'h4404))
    _al_u5471 (
    .a(_al_u5448_o),
    .b(_al_u5396_o),
    .c(_al_u5399_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[9] ),
    .o(_al_u5471_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*A))"),
    .INIT(8'hc4))
    _al_u5472 (
    .a(_al_u4111_o),
    .b(_al_u5471_o),
    .c(_al_u5399_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wskhu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*B)*~(~D*A))"),
    .INIT(16'hf351))
    _al_u5473 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Alkhu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wskhu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Im9ax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tt9ax6 ),
    .o(_al_u5473_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u5474 (
    .a(_al_u5396_o),
    .b(_al_u5403_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T7bax6 ),
    .o(_al_u5474_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*(~A*~(D)*~(C)+~A*D*~(C)+~(~A)*D*C+~A*D*C))"),
    .INIT(16'h3101))
    _al_u5475 (
    .a(_al_u4071_o),
    .b(_al_u5474_o),
    .c(_al_u5399_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[18] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q4lhu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*B)*~(~D*A))"),
    .INIT(16'hf351))
    _al_u5476 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cykhu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q4lhu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ab9ax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qkabx6 ),
    .o(_al_u5476_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(C*~A))"),
    .INIT(16'h8caf))
    _al_u5477 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q4lhu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qnkhu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ab9ax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tc9bx6 ),
    .o(_al_u5477_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u5478 (
    .a(_al_u5470_o),
    .b(_al_u5473_o),
    .c(_al_u5476_o),
    .d(_al_u5477_o),
    .o(_al_u5478_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(C*~(~D*~B)))"),
    .INIT(16'h0515))
    _al_u5479 (
    .a(_al_u5396_o),
    .b(_al_u5398_o),
    .c(_al_u5403_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n6023_lutinv ),
    .o(_al_u5479_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*B*A)"),
    .INIT(16'h0800))
    _al_u548 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pjyiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R9yax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W5ypw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztupw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G2fiu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~B*(~A*~(D)*~(C)+~A*D*~(C)+~(~A)*D*C+~A*D*C))"),
    .INIT(16'h3101))
    _al_u5480 (
    .a(_al_u4076_o),
    .b(_al_u5479_o),
    .c(_al_u5399_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[19] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y5lhu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*~B)*~(D*~A))"),
    .INIT(16'h8acf))
    _al_u5481 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I3lhu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y5lhu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fldbx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xc9ax6 ),
    .o(_al_u5481_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(~D*C))"),
    .INIT(16'h4404))
    _al_u5482 (
    .a(_al_u5430_o),
    .b(_al_u5396_o),
    .c(_al_u5399_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[8] ),
    .o(_al_u5482_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*A))"),
    .INIT(8'hc4))
    _al_u5483 (
    .a(_al_u4237_o),
    .b(_al_u5482_o),
    .c(_al_u5399_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Orkhu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(~C*A))"),
    .INIT(16'hf531))
    _al_u5484 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zelhu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Orkhu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Itcbx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N3jbx6 ),
    .o(_al_u5484_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(C*~A))"),
    .INIT(16'h8caf))
    _al_u5485 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wskhu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Orkhu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Im9ax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N3jbx6 ),
    .o(_al_u5485_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(~C*A))"),
    .INIT(16'hf531))
    _al_u5486 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y5lhu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uwkhu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fldbx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oi9ax6 ),
    .o(_al_u5486_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u5487 (
    .a(_al_u5481_o),
    .b(_al_u5484_o),
    .c(_al_u5485_o),
    .d(_al_u5486_o),
    .o(_al_u5487_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u5488 (
    .a(_al_u5445_o),
    .b(_al_u5466_o),
    .c(_al_u5478_o),
    .d(_al_u5487_o),
    .o(_al_u5488_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*B))"),
    .INIT(8'ha2))
    _al_u5489 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nvkbx6 [7]),
    .b(_al_u5399_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[1] ),
    .o(_al_u5489_o));
  AL_MAP_LUT2 #(
    .EQN("~(B*A)"),
    .INIT(4'h7))
    _al_u549 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G2fiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C1wpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z1fiu6 ));
  AL_MAP_LUT4 #(
    .EQN("(C*B*~(~D*A))"),
    .INIT(16'hc040))
    _al_u5490 (
    .a(_al_u4423_o),
    .b(_al_u5489_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n6018_lutinv ),
    .d(_al_u5399_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kikhu6 ));
  AL_MAP_LUT4 #(
    .EQN("(B*(~A*~(D)*~(C)+~A*D*~(C)+~(~A)*D*C+~A*D*C))"),
    .INIT(16'hc404))
    _al_u5491 (
    .a(_al_u4136_o),
    .b(_al_u5396_o),
    .c(_al_u5399_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[14] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kzkhu6 ));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    _al_u5492 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kzkhu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rg9ax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/eq1/xor_i0[15]_i1[15]_o_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u5493 (
    .a(_al_u5396_o),
    .b(_al_u5403_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n6021_lutinv ),
    .o(_al_u5493_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*(~A*~(D)*~(C)+~A*D*~(C)+~(~A)*D*C+~A*D*C))"),
    .INIT(16'h3101))
    _al_u5494 (
    .a(_al_u3885_o),
    .b(_al_u5493_o),
    .c(_al_u5399_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[28] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nhlhu6 ));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u5495 (
    .a(_al_u5420_o),
    .b(_al_u5398_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n6023_lutinv ),
    .o(_al_u5495_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*(~A*~(D)*~(C)+~A*D*~(C)+~(~A)*D*C+~A*D*C))"),
    .INIT(16'h3101))
    _al_u5496 (
    .a(_al_u4197_o),
    .b(_al_u5495_o),
    .c(_al_u5399_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[27] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gglhu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C@B)*~(D@A))"),
    .INIT(16'h8241))
    _al_u5497 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nhlhu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gglhu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nfgax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wahbx6 ),
    .o(_al_u5497_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u5498 (
    .a(_al_u5474_o),
    .b(_al_u5399_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[15] ),
    .o(_al_u5498_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*~B))"),
    .INIT(8'ha8))
    _al_u5499 (
    .a(_al_u5498_o),
    .b(_al_u5396_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n6023_lutinv ),
    .o(_al_u5499_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*B*A)"),
    .INIT(16'h0800))
    _al_u550 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vynow6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R9yax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W5ypw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztupw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C0fiu6 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*A))"),
    .INIT(8'hc4))
    _al_u5500 (
    .a(_al_u4056_o),
    .b(_al_u5499_o),
    .c(_al_u5399_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S0lhu6 ));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(D@C))"),
    .INIT(16'h4004))
    _al_u5501 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/eq1/xor_i0[15]_i1[15]_o_lutinv ),
    .b(_al_u5497_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S0lhu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ue9ax6 ),
    .o(_al_u5501_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*(~A*~(D)*~(C)+~A*D*~(C)+~(~A)*D*C+~A*D*C))"),
    .INIT(16'h3101))
    _al_u5502 (
    .a(_al_u4091_o),
    .b(_al_u5420_o),
    .c(_al_u5399_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[22] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W9lhu6 ));
  AL_MAP_LUT4 #(
    .EQN("(B*(~A*~(D)*~(C)+~A*D*~(C)+~(~A)*D*C+~A*D*C))"),
    .INIT(16'hc404))
    _al_u5503 (
    .a(_al_u4225_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nvkbx6 [3]),
    .c(_al_u5399_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[2] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sjkhu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C@B)*~(D@A))"),
    .INIT(16'h8241))
    _al_u5504 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W9lhu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sjkhu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pv9ax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zvgbx6 ),
    .o(_al_u5504_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(~D*C))"),
    .INIT(16'h8808))
    _al_u5505 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n6006_lutinv ),
    .b(_al_u5396_o),
    .c(_al_u5399_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[4] ),
    .o(_al_u5505_o));
  AL_MAP_LUT4 #(
    .EQN("(D@(B*~(~C*A)))"),
    .INIT(16'h3bc4))
    _al_u5506 (
    .a(_al_u4219_o),
    .b(_al_u5505_o),
    .c(_al_u5399_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xr9ax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/eq1/xor_i0[5]_i1[5]_o_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u5507 (
    .a(_al_u5398_o),
    .b(_al_u5403_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n6023_lutinv ),
    .o(_al_u5507_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(~D*C))"),
    .INIT(16'h4404))
    _al_u5508 (
    .a(_al_u5507_o),
    .b(_al_u5396_o),
    .c(_al_u5399_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[11] ),
    .o(_al_u5508_o));
  AL_MAP_LUT4 #(
    .EQN("(D@(B*~(~C*A)))"),
    .INIT(16'h3bc4))
    _al_u5509 (
    .a(_al_u4035_o),
    .b(_al_u5508_o),
    .c(_al_u5399_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lk9ax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/eq1/xor_i0[12]_i1[12]_o_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("~(B*A)"),
    .INIT(4'h7))
    _al_u551 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C0fiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C1wpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzeiu6 ));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u5510 (
    .a(_al_u5504_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/eq1/xor_i0[5]_i1[5]_o_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/eq1/xor_i0[12]_i1[12]_o_lutinv ),
    .o(_al_u5510_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*~(D@A))"),
    .INIT(16'h8040))
    _al_u5511 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kikhu6 ),
    .b(_al_u5501_o),
    .c(_al_u5510_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lx9ax6 ),
    .o(_al_u5511_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u5512 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J71iu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N39ax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ttmhu6 ));
  AL_MAP_LUT4 #(
    .EQN("(C*B*~(D@A))"),
    .INIT(16'h8040))
    _al_u5513 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufkhu6 ),
    .b(_al_u5488_o),
    .c(_al_u5511_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ttmhu6 ),
    .o(_al_u5513_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*A)"),
    .INIT(16'h0080))
    _al_u5514 (
    .a(_al_u5399_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J0iax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6lax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 ),
    .o(_al_u5514_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~B*~(~D*~A))"),
    .INIT(16'h3020))
    _al_u5515 (
    .a(_al_u5394_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/eq1/xor_i0[1]_i1[1]_o_lutinv ),
    .c(_al_u5513_o),
    .d(_al_u5514_o),
    .o(_al_u5515_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u5516 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eg7iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dg2qw6 ),
    .o(_al_u5516_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B)*~(C)*~(D)+A*B*~(C)*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+A*B*C*D)"),
    .INIT(16'hbb8a))
    _al_u5517 (
    .a(_al_u5515_o),
    .b(_al_u5516_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F4ibx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uephu6 ));
  AL_MAP_LUT4 #(
    .EQN("(A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .INIT(16'ha280))
    _al_u5518 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xipiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fnpiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R19ax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zx8ax6 ),
    .o(_al_u5518_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u5519 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gr2qw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sbfax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vz8ax6 ),
    .o(_al_u5519_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u552 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_i [7]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_i [8]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_i [9]),
    .o(_al_u552_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u5520 (
    .a(_al_u5519_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vibax6 ),
    .o(_al_u5520_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u5521 (
    .a(_al_u5520_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgbax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ntkbx6 [7]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u5522 (
    .a(_al_u5519_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dfbax6 ),
    .o(_al_u5522_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u5523 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R19ax6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zx8ax6 ),
    .o(_al_u5523_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*A*~(~D*B))"),
    .INIT(16'h0a02))
    _al_u5524 (
    .a(_al_u5522_o),
    .b(_al_u5523_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hdbax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[0] ),
    .o(_al_u5524_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*~(~D*~A))"),
    .INIT(16'hc080))
    _al_u5525 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hz0iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ntkbx6 [7]),
    .c(_al_u5524_o),
    .d(_al_u5523_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oxhhu6 ));
  AL_MAP_LUT4 #(
    .EQN("(A@(D*~(~C*~B)))"),
    .INIT(16'h56aa))
    _al_u5526 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oxhhu6 ),
    .b(_al_u1888_o),
    .c(_al_u5523_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xwaax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/eq0/xor_i0[1]_i1[1]_o_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u5527 (
    .a(_al_u5522_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vibax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgbax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ntkbx6 [3]));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u5528 (
    .a(_al_u5519_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hdbax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tikbx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n5997_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*A)"),
    .INIT(16'h0080))
    _al_u5529 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/My0iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ntkbx6 [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n5997_lutinv ),
    .d(_al_u5523_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gwhhu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u553 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_i [3]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_i [4]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_i [5]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_i [6]),
    .o(_al_u553_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u5530 (
    .a(_al_u5519_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dfbax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hdbax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n5995_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u5531 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n5995_lutinv ),
    .b(_al_u5519_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tikbx6 ),
    .o(_al_u5531_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u5532 (
    .a(_al_u5519_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgbax6 ),
    .o(_al_u5532_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(~B*A))"),
    .INIT(8'h0d))
    _al_u5533 (
    .a(_al_u5523_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[5] ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vibax6 ),
    .o(_al_u5533_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    _al_u5534 (
    .a(_al_u5531_o),
    .b(_al_u5532_o),
    .c(_al_u5533_o),
    .o(_al_u5534_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*A))"),
    .INIT(8'hc4))
    _al_u5535 (
    .a(_al_u4141_o),
    .b(_al_u5534_o),
    .c(_al_u5523_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C4ihu6 ));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u5536 (
    .a(_al_u5523_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vibax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[3] ),
    .o(_al_u5536_o));
  AL_MAP_LUT4 #(
    .EQN("(C*A*~(D*~B))"),
    .INIT(16'h80a0))
    _al_u5537 (
    .a(_al_u5532_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n5997_lutinv ),
    .c(_al_u5536_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dfbax6 ),
    .o(_al_u5537_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*A))"),
    .INIT(8'hc4))
    _al_u5538 (
    .a(_al_u4231_o),
    .b(_al_u5537_o),
    .c(_al_u5523_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M1ihu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*B)*~(~D*A))"),
    .INIT(16'hf351))
    _al_u5539 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C4ihu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M1ihu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jraax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pe9bx6 ),
    .o(_al_u5539_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u554 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_i [13]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_i [14]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_i [15]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_i [2]),
    .o(_al_u554_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(~C*~(~D*B)))"),
    .INIT(16'ha0a8))
    _al_u5540 (
    .a(_al_u5520_o),
    .b(_al_u5522_o),
    .c(_al_u5532_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hdbax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ntkbx6 [9]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u5541 (
    .a(_al_u5519_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tikbx6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgbax6 ),
    .o(_al_u5541_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*B))"),
    .INIT(8'ha2))
    _al_u5542 (
    .a(_al_u5541_o),
    .b(_al_u5523_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[7] ),
    .o(_al_u5542_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*~(~D*A))"),
    .INIT(16'hc040))
    _al_u5543 (
    .a(_al_u4106_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ntkbx6 [9]),
    .c(_al_u5542_o),
    .d(_al_u5523_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S6ihu6 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C@B))"),
    .INIT(8'h82))
    _al_u5544 (
    .a(_al_u5539_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S6ihu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vlaax6 ),
    .o(_al_u5544_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*A*~(D*C))"),
    .INIT(16'h0222))
    _al_u5545 (
    .a(_al_u5519_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dfbax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hdbax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tikbx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n5992_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u5546 (
    .a(_al_u5523_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[17] ),
    .o(_al_u5546_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(~A*~(C*B)))"),
    .INIT(16'h00ea))
    _al_u5547 (
    .a(_al_u5520_o),
    .b(_al_u5532_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n5992_lutinv ),
    .d(_al_u5546_o),
    .o(_al_u5547_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*A))"),
    .INIT(8'hc4))
    _al_u5548 (
    .a(_al_u4066_o),
    .b(_al_u5547_o),
    .c(_al_u5523_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ujihu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*~B)*~(~D*A))"),
    .INIT(16'hcf45))
    _al_u5549 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ujihu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M1ihu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jraax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Naaax6 ),
    .o(_al_u5549_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u555 (
    .a(_al_u552_o),
    .b(_al_u553_o),
    .c(_al_u554_o),
    .o(_al_u555_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(~D*~C*B))"),
    .INIT(16'h5551))
    _al_u5550 (
    .a(_al_u5520_o),
    .b(_al_u5522_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hdbax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgbax6 ),
    .o(_al_u5550_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*(~A*~(D)*~(C)+~A*D*~(C)+~(~A)*D*C+~A*D*C))"),
    .INIT(16'h3101))
    _al_u5551 (
    .a(_al_u4061_o),
    .b(_al_u5550_o),
    .c(_al_u5523_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[16] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Miihu6 ));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D@C))"),
    .INIT(16'h8008))
    _al_u5552 (
    .a(_al_u5544_o),
    .b(_al_u5549_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Miihu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nlbbx6 ),
    .o(_al_u5552_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*B))"),
    .INIT(8'ha2))
    _al_u5553 (
    .a(_al_u5520_o),
    .b(_al_u5523_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[13] ),
    .o(_al_u5553_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u5554 (
    .a(_al_u5531_o),
    .b(_al_u5553_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgbax6 ),
    .o(_al_u5554_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*A))"),
    .INIT(8'hc4))
    _al_u5555 (
    .a(_al_u4131_o),
    .b(_al_u5554_o),
    .c(_al_u5523_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oeihu6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u5556 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oeihu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nmabx6 ),
    .o(_al_u5556_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(~A*~(D)*~(C)+~A*D*~(C)+~(~A)*D*C+~A*D*C))"),
    .INIT(16'hc404))
    _al_u5557 (
    .a(_al_u4121_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ntkbx6 [7]),
    .c(_al_u5523_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[6] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K5ihu6 ));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*~(D@B))"),
    .INIT(16'h4010))
    _al_u5558 (
    .a(_al_u5556_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K5ihu6 ),
    .c(_al_u5519_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rnaax6 ),
    .o(_al_u5558_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u5559 (
    .a(_al_u5520_o),
    .b(_al_u5522_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgbax6 ),
    .o(_al_u5559_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u556 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_i [1]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_i [10]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_i [11]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_i [12]),
    .o(_al_u556_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*(~A*~(D)*~(C)+~A*D*~(C)+~(~A)*D*C+~A*D*C))"),
    .INIT(16'h3101))
    _al_u5560 (
    .a(_al_u4071_o),
    .b(_al_u5559_o),
    .c(_al_u5523_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[18] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Clihu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(~C*A))"),
    .INIT(16'hf531))
    _al_u5561 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oeihu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Clihu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nmabx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q8aax6 ),
    .o(_al_u5561_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(B*~(D*~C)))"),
    .INIT(16'h1511))
    _al_u5562 (
    .a(_al_u5520_o),
    .b(_al_u5532_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n5997_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dfbax6 ),
    .o(_al_u5562_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*(~A*~(D)*~(C)+~A*D*~(C)+~(~A)*D*C+~A*D*C))"),
    .INIT(16'h3101))
    _al_u5563 (
    .a(_al_u4076_o),
    .b(_al_u5562_o),
    .c(_al_u5523_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[19] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kmihu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(C*~A))"),
    .INIT(16'h8caf))
    _al_u5564 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kmihu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Clihu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cndbx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q8aax6 ),
    .o(_al_u5564_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u5565 (
    .a(_al_u5552_o),
    .b(_al_u5558_o),
    .c(_al_u5561_o),
    .d(_al_u5564_o),
    .o(_al_u5565_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(~A*~(D)*~(C)+~A*D*~(C)+~(~A)*D*C+~A*D*C))"),
    .INIT(16'hc404))
    _al_u5566 (
    .a(_al_u4237_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ntkbx6 [9]),
    .c(_al_u5523_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[8] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A8ihu6 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*B))"),
    .INIT(8'ha2))
    _al_u5567 (
    .a(_al_u5520_o),
    .b(_al_u5523_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[12] ),
    .o(_al_u5567_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*~B))"),
    .INIT(8'ha8))
    _al_u5568 (
    .a(_al_u5567_o),
    .b(_al_u5532_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n5995_lutinv ),
    .o(_al_u5568_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*A))"),
    .INIT(8'hc4))
    _al_u5569 (
    .a(_al_u4126_o),
    .b(_al_u5568_o),
    .c(_al_u5523_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gdihu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*~B)*~(D*~A))"),
    .INIT(16'ha8fc))
    _al_u557 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n31 ),
    .b(uart0_txen_pad),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_ctrl [1]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_i [0]),
    .o(_al_u557_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*B)*~(D*~A))"),
    .INIT(16'ha2f3))
    _al_u5570 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A8ihu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gdihu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Egaax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J5jbx6 ),
    .o(_al_u5570_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u5571 (
    .a(_al_u5520_o),
    .b(_al_u5532_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n5992_lutinv ),
    .o(_al_u5571_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*(~A*~(D)*~(C)+~A*D*~(C)+~(~A)*D*C+~A*D*C))"),
    .INIT(16'h3101))
    _al_u5572 (
    .a(_al_u4096_o),
    .b(_al_u5571_o),
    .c(_al_u5523_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[25] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Guihu6 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C@B))"),
    .INIT(8'h82))
    _al_u5573 (
    .a(_al_u5570_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Guihu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cccbx6 ),
    .o(_al_u5573_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*B))"),
    .INIT(8'ha2))
    _al_u5574 (
    .a(_al_u5520_o),
    .b(_al_u5523_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[9] ),
    .o(_al_u5574_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*~B))"),
    .INIT(8'ha8))
    _al_u5575 (
    .a(_al_u5574_o),
    .b(_al_u5532_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n5992_lutinv ),
    .o(_al_u5575_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*A))"),
    .INIT(8'hc4))
    _al_u5576 (
    .a(_al_u4111_o),
    .b(_al_u5575_o),
    .c(_al_u5523_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I9ihu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*B)*~(D@A))"),
    .INIT(16'ha251))
    _al_u5577 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I9ihu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A8ihu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J5jbx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yjaax6 ),
    .o(_al_u5577_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*~A))"),
    .INIT(8'h23))
    _al_u5578 (
    .a(_al_u5531_o),
    .b(_al_u5520_o),
    .c(_al_u5532_o),
    .o(_al_u5578_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*(~A*~(D)*~(C)+~A*D*~(C)+~(~A)*D*C+~A*D*C))"),
    .INIT(16'h3101))
    _al_u5579 (
    .a(_al_u4086_o),
    .b(_al_u5578_o),
    .c(_al_u5523_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[21] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Apihu6 ));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u558 (
    .a(_al_u555_o),
    .b(_al_u556_o),
    .c(_al_u557_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reload_i ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(~C*A))"),
    .INIT(16'hc4f5))
    _al_u5580 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kmihu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Apihu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cndbx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qlfbx6 ),
    .o(_al_u5580_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(C*~A))"),
    .INIT(16'h8caf))
    _al_u5581 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ujihu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C4ihu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Naaax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pe9bx6 ),
    .o(_al_u5581_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u5582 (
    .a(_al_u5573_o),
    .b(_al_u5577_o),
    .c(_al_u5580_o),
    .d(_al_u5581_o),
    .o(_al_u5582_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u5583 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gdihu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Egaax6 ),
    .o(_al_u5583_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u5584 (
    .a(_al_u5520_o),
    .b(_al_u5532_o),
    .o(_al_u5584_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u5585 (
    .a(_al_u5531_o),
    .b(_al_u5584_o),
    .o(_al_u5585_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*(~A*~(D)*~(C)+~A*D*~(C)+~(~A)*D*C+~A*D*C))"),
    .INIT(16'h3101))
    _al_u5586 (
    .a(_al_u3889_o),
    .b(_al_u5585_o),
    .c(_al_u5523_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[29] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mzihu6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u5587 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mzihu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z2aax6 ),
    .o(_al_u5587_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~A*~(~D*B))"),
    .INIT(16'h0501))
    _al_u5588 (
    .a(_al_u5520_o),
    .b(_al_u5522_o),
    .c(_al_u5532_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hdbax6 ),
    .o(_al_u5588_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*(~A*~(D)*~(C)+~A*D*~(C)+~(~A)*D*C+~A*D*C))"),
    .INIT(16'h3101))
    _al_u5589 (
    .a(_al_u4191_o),
    .b(_al_u5588_o),
    .c(_al_u5523_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[24] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ysihu6 ));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    _al_u559 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_txd ),
    .b(uart0_txd_pad),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/update_reg_txd ));
  AL_MAP_LUT4 #(
    .EQN("(~B*~A*~(D@C))"),
    .INIT(16'h1001))
    _al_u5590 (
    .a(_al_u5583_o),
    .b(_al_u5587_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ysihu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4aax6 ),
    .o(_al_u5590_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u5591 (
    .a(_al_u5522_o),
    .b(_al_u5532_o),
    .o(_al_u5591_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(~D*C))"),
    .INIT(16'h4404))
    _al_u5592 (
    .a(_al_u5591_o),
    .b(_al_u5520_o),
    .c(_al_u5523_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[10] ),
    .o(_al_u5592_o));
  AL_MAP_LUT4 #(
    .EQN("~(D@(B*~(~C*A)))"),
    .INIT(16'hc43b))
    _al_u5593 (
    .a(_al_u4116_o),
    .b(_al_u5592_o),
    .c(_al_u5523_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ux8bx6 ),
    .o(_al_u5593_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u5594 (
    .a(_al_u5520_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n5997_lutinv ),
    .o(_al_u5594_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u5595 (
    .a(_al_u5591_o),
    .b(_al_u5594_o),
    .o(_al_u5595_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*(~A*~(D)*~(C)+~A*D*~(C)+~(~A)*D*C+~A*D*C))"),
    .INIT(16'h3101))
    _al_u5596 (
    .a(_al_u4197_o),
    .b(_al_u5595_o),
    .c(_al_u5523_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[27] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wwihu6 ));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D@C))"),
    .INIT(16'h8008))
    _al_u5597 (
    .a(_al_u5590_o),
    .b(_al_u5593_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wwihu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Khgax6 ),
    .o(_al_u5597_o));
  AL_MAP_LUT3 #(
    .EQN("~(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'h2e))
    _al_u5598 (
    .a(_al_u3887_o),
    .b(_al_u5523_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[30] ),
    .o(_al_u5598_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*~B)*~(~D*A))"),
    .INIT(16'hfc54))
    _al_u5599 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Apihu6 ),
    .b(_al_u5598_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N4gax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qlfbx6 ),
    .o(_al_u5599_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*B*~A)"),
    .INIT(16'h0400))
    _al_u560 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_state_inc ),
    .b(_al_u370_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_state [0]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_state [1]),
    .o(_al_u560_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u5600 (
    .a(_al_u5520_o),
    .b(_al_u5541_o),
    .o(_al_u5600_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~A*~(~D*C))"),
    .INIT(16'h1101))
    _al_u5601 (
    .a(_al_u5588_o),
    .b(_al_u5600_o),
    .c(_al_u5523_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[23] ),
    .o(_al_u5601_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*A))"),
    .INIT(8'hc4))
    _al_u5602 (
    .a(_al_u4184_o),
    .b(_al_u5601_o),
    .c(_al_u5523_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qrihu6 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C@B))"),
    .INIT(8'h82))
    _al_u5603 (
    .a(_al_u5599_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qrihu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T6aax6 ),
    .o(_al_u5603_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(~D*A))"),
    .INIT(16'h3f15))
    _al_u5604 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mzihu6 ),
    .b(_al_u5598_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N4gax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z2aax6 ),
    .o(_al_u5604_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u5605 (
    .a(_al_u5520_o),
    .b(_al_u5532_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n5995_lutinv ),
    .o(_al_u5605_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*(~A*~(D)*~(C)+~A*D*~(C)+~(~A)*D*C+~A*D*C))"),
    .INIT(16'h3101))
    _al_u5606 (
    .a(_al_u3885_o),
    .b(_al_u5605_o),
    .c(_al_u5523_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[28] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eyihu6 ));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D@C))"),
    .INIT(16'h8008))
    _al_u5607 (
    .a(_al_u5603_o),
    .b(_al_u5604_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eyihu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tchbx6 ),
    .o(_al_u5607_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u5608 (
    .a(_al_u5565_o),
    .b(_al_u5582_o),
    .c(_al_u5597_o),
    .d(_al_u5607_o),
    .o(_al_u5608_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*B))"),
    .INIT(8'ha2))
    _al_u5609 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ntkbx6 [7]),
    .b(_al_u5523_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[1] ),
    .o(_al_u5609_o));
  AL_MAP_LUT3 #(
    .EQN("~(~A*~(C*B))"),
    .INIT(8'hea))
    _al_u561 (
    .a(_al_u560_o),
    .b(_al_u364_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n102 [3]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_rx_state [3]));
  AL_MAP_LUT4 #(
    .EQN("(C*B*~(~D*A))"),
    .INIT(16'hc040))
    _al_u5610 (
    .a(_al_u4423_o),
    .b(_al_u5609_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n5992_lutinv ),
    .d(_al_u5523_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wyhhu6 ));
  AL_MAP_LUT4 #(
    .EQN("(B*(~A*~(D)*~(C)+~A*D*~(C)+~(~A)*D*C+~A*D*C))"),
    .INIT(16'hc404))
    _al_u5611 (
    .a(_al_u4225_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ntkbx6 [3]),
    .c(_al_u5523_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[2] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E0ihu6 ));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    _al_u5612 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E0ihu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ftaax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/eq0/xor_i0[3]_i1[3]_o_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(B*(~A*~(D)*~(C)+~A*D*~(C)+~(~A)*D*C+~A*D*C))"),
    .INIT(16'hc404))
    _al_u5613 (
    .a(_al_u4136_o),
    .b(_al_u5520_o),
    .c(_al_u5523_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[14] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wfihu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~B*~A*~(~D*C))"),
    .INIT(16'h1101))
    _al_u5614 (
    .a(_al_u5594_o),
    .b(_al_u5559_o),
    .c(_al_u5523_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[15] ),
    .o(_al_u5614_o));
  AL_MAP_LUT4 #(
    .EQN("(D@(B*~(~C*A)))"),
    .INIT(16'h3bc4))
    _al_u5615 (
    .a(_al_u4056_o),
    .b(_al_u5614_o),
    .c(_al_u5523_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kcaax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/eq0/xor_i0[16]_i1[16]_o_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C@A))"),
    .INIT(8'h21))
    _al_u5616 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wfihu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/eq0/xor_i0[16]_i1[16]_o_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Heaax6 ),
    .o(_al_u5616_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*(~A*~(D)*~(C)+~A*D*~(C)+~(~A)*D*C+~A*D*C))"),
    .INIT(16'h3101))
    _al_u5617 (
    .a(_al_u4091_o),
    .b(_al_u5584_o),
    .c(_al_u5523_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[22] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iqihu6 ));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(D@C))"),
    .INIT(16'h4004))
    _al_u5618 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/eq0/xor_i0[3]_i1[3]_o_lutinv ),
    .b(_al_u5616_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iqihu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wxgbx6 ),
    .o(_al_u5618_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*B))"),
    .INIT(8'ha2))
    _al_u5619 (
    .a(_al_u5520_o),
    .b(_al_u5523_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[4] ),
    .o(_al_u5619_o));
  AL_MAP_LUT3 #(
    .EQN("~(~A*~(C*B))"),
    .INIT(8'hea))
    _al_u562 (
    .a(_al_u560_o),
    .b(_al_u364_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n102 [1]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_rx_state [1]));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u5620 (
    .a(_al_u5619_o),
    .b(_al_u5532_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n5995_lutinv ),
    .o(_al_u5620_o));
  AL_MAP_LUT4 #(
    .EQN("(D@(B*~(~C*A)))"),
    .INIT(16'h3bc4))
    _al_u5621 (
    .a(_al_u4219_o),
    .b(_al_u5620_o),
    .c(_al_u5523_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Npaax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/eq0/xor_i0[5]_i1[5]_o_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*B))"),
    .INIT(8'ha2))
    _al_u5622 (
    .a(_al_u5520_o),
    .b(_al_u5523_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[11] ),
    .o(_al_u5622_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*A))"),
    .INIT(8'hc4))
    _al_u5623 (
    .a(_al_u5591_o),
    .b(_al_u5622_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n5997_lutinv ),
    .o(_al_u5623_o));
  AL_MAP_LUT4 #(
    .EQN("(D@(B*~(~C*A)))"),
    .INIT(16'h3bc4))
    _al_u5624 (
    .a(_al_u4035_o),
    .b(_al_u5623_o),
    .c(_al_u5523_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Biaax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/eq0/xor_i0[12]_i1[12]_o_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u5625 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/eq0/xor_i0[5]_i1[5]_o_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/eq0/xor_i0[12]_i1[12]_o_lutinv ),
    .o(_al_u5625_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u5626 (
    .a(_al_u5591_o),
    .b(_al_u5520_o),
    .o(_al_u5626_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*(~A*~(D)*~(C)+~A*D*~(C)+~(~A)*D*C+~A*D*C))"),
    .INIT(16'h3101))
    _al_u5627 (
    .a(_al_u4101_o),
    .b(_al_u5626_o),
    .c(_al_u5523_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[26] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ovihu6 ));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    _al_u5628 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ovihu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fvcbx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/eq0/xor_i0[27]_i1[27]_o_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u5629 (
    .a(_al_u5520_o),
    .b(_al_u5532_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n5995_lutinv ),
    .o(_al_u5629_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*A)"),
    .INIT(16'h0002))
    _al_u563 (
    .a(_al_u456_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/i_paddr [12]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/i_paddr [13]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/i_paddr [14]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_apb_slave_mux/n0 ));
  AL_MAP_LUT4 #(
    .EQN("(~B*(~A*~(D)*~(C)+~A*D*~(C)+~(~A)*D*C+~A*D*C))"),
    .INIT(16'h3101))
    _al_u5630 (
    .a(_al_u4081_o),
    .b(_al_u5629_o),
    .c(_al_u5523_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[20] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Snihu6 ));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    _al_u5631 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Snihu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J6ebx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/eq0/xor_i0[21]_i1[21]_o_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    _al_u5632 (
    .a(_al_u5618_o),
    .b(_al_u5625_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/eq0/xor_i0[27]_i1[27]_o_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/eq0/xor_i0[21]_i1[21]_o_lutinv ),
    .o(_al_u5632_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C@A))"),
    .INIT(8'h84))
    _al_u5633 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wyhhu6 ),
    .b(_al_u5632_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bvaax6 ),
    .o(_al_u5633_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u5634 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J71iu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D1aax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wbkhu6 ));
  AL_MAP_LUT4 #(
    .EQN("(C*B*~(D@A))"),
    .INIT(16'h8040))
    _al_u5635 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gwhhu6 ),
    .b(_al_u5608_o),
    .c(_al_u5633_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wbkhu6 ),
    .o(_al_u5635_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*A)"),
    .INIT(16'h0080))
    _al_u5636 (
    .a(_al_u5523_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J0iax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6lax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 ),
    .o(_al_u5636_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~B*~(~D*~A))"),
    .INIT(16'h3020))
    _al_u5637 (
    .a(_al_u5518_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/eq0/xor_i0[1]_i1[1]_o_lutinv ),
    .c(_al_u5635_o),
    .d(_al_u5636_o),
    .o(_al_u5637_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u5638 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ws4iu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dg2qw6 ),
    .o(_al_u5638_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B)*~(C)*~(D)+A*B*~(C)*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+A*B*C*D)"),
    .INIT(16'hbb8a))
    _al_u5639 (
    .a(_al_u5637_o),
    .b(_al_u5638_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vpkpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bfphu6 ));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u564 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/state_reg [0]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/state_reg [1]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/state_reg [2]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/apb_tran_end ));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+A*~(B)*C*D)"),
    .INIT(16'h2e3e))
    _al_u5640 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/n1 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/state_reg [0]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/state_reg [1]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/state_reg [2]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/next_state [1]));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*~A)"),
    .INIT(8'h04))
    _al_u5641 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/state_reg [0]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/state_reg [1]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/state_reg [2]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/next_state [0]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u5642 (
    .a(\u_cmsdk_mcu/sram_hsel ),
    .b(_al_u5003_o),
    .o(\u_cmsdk_mcu/u_ahb_ram/n2 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u5643 (
    .a(_al_u5515_o),
    .b(_al_u5637_o),
    .o(_al_u5643_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u5644 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Scbiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ud4iu6 ),
    .o(_al_u5644_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h7745))
    _al_u5645 (
    .a(_al_u5643_o),
    .b(_al_u5644_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rkbax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ifphu6 ));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~C*B*A)"),
    .INIT(16'hfff7))
    _al_u5646 (
    .a(_al_u5643_o),
    .b(_al_u4452_o),
    .c(_al_u1779_o),
    .d(_al_u1257_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dt4iu6 ));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u5647 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cvciu6 ),
    .b(_al_u5275_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D43qw6 ),
    .o(_al_u5647_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u5648 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gkwiu6 ),
    .b(_al_u5647_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A2qiu6 ),
    .o(_al_u5648_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*~B*~A)"),
    .INIT(16'h0010))
    _al_u5649 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K0qiu6_lutinv ),
    .b(_al_u5291_o),
    .c(_al_u5648_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q3qiu6 ),
    .o(_al_u5649_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u565 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_apb_slave_mux/n0 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/apb_tran_end ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PWRITE ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n68 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5650 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xs1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yc7iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eafax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xaeax6 ),
    .o(_al_u5650_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5651 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ve7iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vr1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Efdax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H4bax6 ),
    .o(_al_u5651_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5652 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dw1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zt1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D1aax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q6fax6 ),
    .o(_al_u5652_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5653 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cs1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ar1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I1lpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljcax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ktwiu6 ));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u5654 (
    .a(_al_u5650_o),
    .b(_al_u5651_o),
    .c(_al_u5652_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ktwiu6 ),
    .o(_al_u5654_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u5655 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fgpiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kw1iu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lmkbx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N39ax6 ),
    .o(_al_u5655_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5656 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jf7iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sg7iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pkkbx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tikbx6 ),
    .o(_al_u5656_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u5657 (
    .a(_al_u5649_o),
    .b(_al_u5654_o),
    .c(_al_u5655_o),
    .d(_al_u5656_o),
    .o(_al_u5657_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u5658 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F0eow6 ),
    .b(_al_u5260_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C3wpw6 ),
    .o(_al_u5658_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u5659 (
    .a(_al_u5658_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M0eow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U31bx6 ),
    .o(_al_u5659_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u566 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[4] ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[5] ),
    .o(_al_u566_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5660 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvgiu6 ),
    .b(_al_u5067_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[0] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N8rpw6 ),
    .o(_al_u5660_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u5661 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6eiu6 ),
    .b(_al_u405_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6rpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zszax6 ),
    .o(_al_u5661_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u5662 (
    .a(_al_u5659_o),
    .b(_al_u5660_o),
    .c(_al_u5661_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M1xiu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u5663 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eg7iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ws4iu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tyaax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zx8ax6 ),
    .o(_al_u5663_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*B*A)"),
    .INIT(16'h0800))
    _al_u5664 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qaqiu6 ),
    .b(_al_u5663_o),
    .c(_al_u5274_o),
    .d(_al_u5340_o),
    .o(_al_u5664_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u5665 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yw1iu6 ),
    .b(_al_u5657_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M1xiu6 ),
    .d(_al_u5664_o),
    .o(_al_u5665_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(C*~(D*~B)))"),
    .INIT(16'h2a0a))
    _al_u5666 (
    .a(_al_u5020_o),
    .b(_al_u4865_o),
    .c(_al_u5665_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/St1iu6 ),
    .o(_al_u5666_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~A*~(D*C))"),
    .INIT(16'h0111))
    _al_u5667 (
    .a(_al_u5666_o),
    .b(_al_u5049_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sf1iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H3lpw6 ),
    .o(_al_u5667_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u5668 (
    .a(_al_u5667_o),
    .b(_al_u5103_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ksgax6 ),
    .o(_al_u5668_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*B))"),
    .INIT(8'hd5))
    _al_u5669 (
    .a(_al_u5668_o),
    .b(_al_u5053_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qehbx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6phu6 ));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u567 (
    .a(_al_u566_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/mux4_b6_sel_is_13_o ));
  AL_MAP_LUT4 #(
    .EQN("(~C*~B*~(D*A))"),
    .INIT(16'h0103))
    _al_u5670 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xs1iu6 ),
    .b(_al_u5291_o),
    .c(_al_u5271_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F7eax6 ),
    .o(_al_u5670_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u5671 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fgpiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dw1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hmbax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y2fax6 ),
    .o(_al_u5671_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u5672 (
    .a(_al_u5670_o),
    .b(_al_u5671_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iv1iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[3] ),
    .o(_al_u5672_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u5673 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vr1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ar1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mbdax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wtxax6 ),
    .o(_al_u5673_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u5674 (
    .a(_al_u5673_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zt1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jraax6 ),
    .o(_al_u5674_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5675 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jf7iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kw1iu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tt9ax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vibax6 ),
    .o(_al_u5675_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5676 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cs1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sg7iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lbbax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tfcax6 ),
    .o(_al_u5676_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u5677 (
    .a(_al_u5672_o),
    .b(_al_u5674_o),
    .c(_al_u5675_o),
    .d(_al_u5676_o),
    .o(_al_u5677_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u5678 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M0eow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F0eow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gihbx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ikhbx6 ),
    .o(_al_u5678_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u5679 (
    .a(_al_u5678_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fpgiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kqhbx6 ),
    .o(_al_u5679_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'h0a0c))
    _al_u568 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_ctrl [6]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_rx_buf [6]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/mux3_b6/B1_0 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5680 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6eiu6 ),
    .b(_al_u5067_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[4] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Imhbx6 ),
    .o(_al_u5680_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u5681 (
    .a(_al_u5679_o),
    .b(_al_u5680_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvgiu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Johbx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yzqiu6 ));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u5682 (
    .a(_al_u5677_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F0riu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yzqiu6 ),
    .o(_al_u5682_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*~(D*~C)))"),
    .INIT(16'h2a22))
    _al_u5683 (
    .a(_al_u5020_o),
    .b(_al_u5682_o),
    .c(_al_u4663_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/St1iu6 ),
    .o(_al_u5683_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u5684 (
    .a(_al_u5683_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sf1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V53qw6 ),
    .o(_al_u5684_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u5685 (
    .a(_al_u5684_o),
    .b(_al_u5053_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pg3qw6 ),
    .o(_al_u5685_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*B))"),
    .INIT(8'hd5))
    _al_u5686 (
    .a(_al_u5685_o),
    .b(_al_u5103_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tb3qw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sdphu6 ));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u5687 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F0eow6 ),
    .b(_al_u5260_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cxzax6 ),
    .o(_al_u5687_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u5688 (
    .a(_al_u405_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvgiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Avzax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oarpw6 ),
    .o(_al_u5688_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u5689 (
    .a(_al_u5687_o),
    .b(_al_u5688_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M0eow6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aa2bx6 ),
    .o(_al_u5689_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u569 (
    .a(_al_u473_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n27_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/mux4_b6_sel_is_13_o ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/mux3_b6/B1_0 ),
    .o(_al_u569_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5690 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6eiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fpgiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G0zax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wnxax6 ),
    .o(_al_u5690_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u5691 (
    .a(_al_u5689_o),
    .b(_al_u5690_o),
    .c(_al_u5067_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[1] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ovpiu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5692 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ws4iu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iv1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[0] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R19ax6 ),
    .o(_al_u5692_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u5693 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ovpiu6 ),
    .b(_al_u5692_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eg7iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L2bax6 ),
    .o(_al_u5693_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u5694 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fgpiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zt1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xnbax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xwaax6 ),
    .o(_al_u5694_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u5695 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kw1iu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hz9ax6 ),
    .o(_al_u5695_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5696 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sg7iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ar1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nu5bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X5bax6 ),
    .o(_al_u5696_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~B*~(D*A))"),
    .INIT(16'h1030))
    _al_u5697 (
    .a(_al_u927_o),
    .b(_al_u5695_o),
    .c(_al_u5696_o),
    .d(_al_u1385_o),
    .o(_al_u5697_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u5698 (
    .a(_al_u5694_o),
    .b(_al_u5697_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jf7iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hdbax6 ),
    .o(_al_u5698_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u5699 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yw1iu6 ),
    .b(_al_u5693_o),
    .c(_al_u5698_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vvpiu6_lutinv ),
    .o(_al_u5699_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C*A))"),
    .INIT(8'hb3))
    _al_u570 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n7_lutinv ),
    .b(_al_u569_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [6]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/read_mux_byte0 [6]));
  AL_MAP_LUT4 #(
    .EQN("(A*~(C*~(D*~B)))"),
    .INIT(16'h2a0a))
    _al_u5700 (
    .a(_al_u5020_o),
    .b(_al_u4581_o),
    .c(_al_u5699_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/St1iu6 ),
    .o(_al_u5700_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~A*~(D*C))"),
    .INIT(16'h0111))
    _al_u5701 (
    .a(_al_u5700_o),
    .b(_al_u5050_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sf1iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L9bbx6 ),
    .o(_al_u5701_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u5702 (
    .a(_al_u5701_o),
    .b(_al_u5053_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vj3qw6 ),
    .o(_al_u5702_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*B))"),
    .INIT(8'hd5))
    _al_u5703 (
    .a(_al_u5702_o),
    .b(_al_u5103_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dugax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nephu6 ));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    _al_u5704 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gr2qw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H4bax6 ),
    .o(_al_u5704_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u5705 (
    .a(_al_u3885_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L18iu6 ),
    .c(_al_u5704_o),
    .o(_al_u5705_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*~A)"),
    .INIT(16'h4000))
    _al_u5706 (
    .a(_al_u5392_o),
    .b(_al_u5705_o),
    .c(_al_u3887_o),
    .d(_al_u3889_o),
    .o(_al_u5706_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u5707 (
    .a(_al_u4035_o),
    .b(_al_u4101_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F2dax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T2dbx6 ),
    .o(_al_u5707_o));
  AL_MAP_LUT3 #(
    .EQN("(A*(C@B))"),
    .INIT(8'h28))
    _al_u5708 (
    .a(_al_u5707_o),
    .b(_al_u4191_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Apcax6 ),
    .o(_al_u5708_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(~C*~A))"),
    .INIT(16'h32fa))
    _al_u5709 (
    .a(_al_u4061_o),
    .b(_al_u4225_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Btbbx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iddax6 ),
    .o(_al_u5709_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u571 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] ),
    .o(_al_u571_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*(D@C))"),
    .INIT(16'h0880))
    _al_u5710 (
    .a(_al_u5708_o),
    .b(_al_u5709_o),
    .c(_al_u4091_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K5hbx6 ),
    .o(_al_u5710_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*~B)*(D@A))"),
    .INIT(16'h54a8))
    _al_u5711 (
    .a(_al_u4066_o),
    .b(_al_u4126_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I0dax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rucax6 ),
    .o(_al_u5711_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*~B)*~(~D*~A))"),
    .INIT(16'hfca8))
    _al_u5712 (
    .a(_al_u4136_o),
    .b(_al_u4225_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iddax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lycax6 ),
    .o(_al_u5712_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(~D*~A))"),
    .INIT(16'h3f2a))
    _al_u5713 (
    .a(_al_u4071_o),
    .b(_al_u4126_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I0dax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uscax6 ),
    .o(_al_u5713_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u5714 (
    .a(_al_u5710_o),
    .b(_al_u5711_o),
    .c(_al_u5712_o),
    .d(_al_u5713_o),
    .o(_al_u5714_o));
  AL_MAP_LUT4 #(
    .EQN("((C@B)*(D@A))"),
    .INIT(16'h1428))
    _al_u5715 (
    .a(_al_u4081_o),
    .b(_al_u4131_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Buabx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xdebx6 ),
    .o(_al_u5715_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*~B)*~(~C*~A))"),
    .INIT(16'hfac8))
    _al_u5716 (
    .a(_al_u4035_o),
    .b(_al_u4237_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F2dax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tcjbx6 ),
    .o(_al_u5716_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*(D@C))"),
    .INIT(16'h0880))
    _al_u5717 (
    .a(_al_u5715_o),
    .b(_al_u5716_o),
    .c(_al_u4111_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C4dax6 ),
    .o(_al_u5717_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5718 (
    .a(_al_u4071_o),
    .b(_al_u4237_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tcjbx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uscax6 ),
    .o(_al_u5718_o));
  AL_MAP_LUT4 #(
    .EQN("((C@B)*(D@A))"),
    .INIT(16'h1428))
    _al_u5719 (
    .a(_al_u4197_o),
    .b(_al_u4231_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mbdax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yogax6 ),
    .o(_al_u5719_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*B*A)"),
    .INIT(16'h0800))
    _al_u572 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n27_lutinv ),
    .b(_al_u571_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[4] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[5] ),
    .o(_al_u572_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*(D@C))"),
    .INIT(16'h0880))
    _al_u5720 (
    .a(_al_u5718_o),
    .b(_al_u5719_o),
    .c(_al_u4056_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Owcax6 ),
    .o(_al_u5720_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u5721 (
    .a(_al_u5714_o),
    .b(_al_u5717_o),
    .c(_al_u5720_o),
    .o(_al_u5721_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(~D*~A))"),
    .INIT(16'h3f2a))
    _al_u5722 (
    .a(_al_u4101_o),
    .b(_al_u4136_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lycax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T2dbx6 ),
    .o(_al_u5722_o));
  AL_MAP_LUT4 #(
    .EQN("(D*A*~(C*B))"),
    .INIT(16'h2a00))
    _al_u5723 (
    .a(_al_u5722_o),
    .b(_al_u4061_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Btbbx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Efdax6 ),
    .o(_al_u5723_o));
  AL_MAP_LUT4 #(
    .EQN("((D@B)*(C@A))"),
    .INIT(16'h1248))
    _al_u5724 (
    .a(_al_u4086_o),
    .b(_al_u4219_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Etfbx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q9dax6 ),
    .o(_al_u5724_o));
  AL_MAP_LUT4 #(
    .EQN("((C@B)*(D@A))"),
    .INIT(16'h1428))
    _al_u5725 (
    .a(_al_u4076_o),
    .b(_al_u4096_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qjcbx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qudbx6 ),
    .o(_al_u5725_o));
  AL_MAP_LUT4 #(
    .EQN("((D@B)*(C@A))"),
    .INIT(16'h1248))
    _al_u5726 (
    .a(_al_u4116_o),
    .b(_al_u4184_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F59bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xqcax6 ),
    .o(_al_u5726_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u5727 (
    .a(_al_u5723_o),
    .b(_al_u5724_o),
    .c(_al_u5725_o),
    .d(_al_u5726_o),
    .o(_al_u5727_o));
  AL_MAP_LUT4 #(
    .EQN("((D@B)*(C@A))"),
    .INIT(16'h1248))
    _al_u5728 (
    .a(_al_u4106_o),
    .b(_al_u4141_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y5dax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zl9bx6 ),
    .o(_al_u5728_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*(D@C))"),
    .INIT(16'h0880))
    _al_u5729 (
    .a(_al_u5727_o),
    .b(_al_u5728_o),
    .c(_al_u4121_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U7dax6 ),
    .o(_al_u5729_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u573 (
    .a(_al_u470_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [1]),
    .o(_al_u573_o));
  AL_MAP_LUT4 #(
    .EQN("(C*A*(D@B))"),
    .INIT(16'h2080))
    _al_u5730 (
    .a(_al_u5721_o),
    .b(_al_u4423_o),
    .c(_al_u5729_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hlcax6 ),
    .o(_al_u5730_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u5731 (
    .a(_al_u4106_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Facax6 ),
    .o(_al_u5731_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u5732 (
    .a(_al_u4126_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P4cax6 ),
    .o(_al_u5732_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~A*(D@C))"),
    .INIT(16'h0110))
    _al_u5733 (
    .a(_al_u5731_o),
    .b(_al_u5732_o),
    .c(_al_u4191_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Htbax6 ),
    .o(_al_u5733_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*~B)*~(~C*~A))"),
    .INIT(16'hfac8))
    _al_u5734 (
    .a(_al_u4081_o),
    .b(_al_u4126_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G8ebx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P4cax6 ),
    .o(_al_u5734_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u5735 (
    .a(_al_u5733_o),
    .b(_al_u5734_o),
    .c(_al_u4035_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6cax6 ),
    .o(_al_u5735_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u5736 (
    .a(_al_u4096_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljcax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zdcbx6 ),
    .o(_al_u5736_o));
  AL_MAP_LUT3 #(
    .EQN("(A*(C@B))"),
    .INIT(8'h28))
    _al_u5737 (
    .a(_al_u5736_o),
    .b(_al_u4197_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hjgax6 ),
    .o(_al_u5737_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(~D*~A))"),
    .INIT(16'h3f2a))
    _al_u5738 (
    .a(_al_u4136_o),
    .b(_al_u4225_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Phcax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S2cax6 ),
    .o(_al_u5738_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*~B)*~(~D*~A))"),
    .INIT(16'hfca8))
    _al_u5739 (
    .a(_al_u4225_o),
    .b(_al_u4237_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F7jbx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Phcax6 ),
    .o(_al_u5739_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h3ff5))
    _al_u574 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_rx_buf [1]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/apbsubsys_interrupt [0]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] ),
    .o(_al_u574_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5740 (
    .a(_al_u4066_o),
    .b(_al_u4141_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lg9bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yybax6 ),
    .o(_al_u5740_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(~D*~A))"),
    .INIT(16'h3f2a))
    _al_u5741 (
    .a(_al_u4066_o),
    .b(_al_u4136_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S2cax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yybax6 ),
    .o(_al_u5741_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u5742 (
    .a(_al_u5738_o),
    .b(_al_u5739_o),
    .c(_al_u5740_o),
    .d(_al_u5741_o),
    .o(_al_u5742_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*~B)*~(~D*~A))"),
    .INIT(16'hfca8))
    _al_u5743 (
    .a(_al_u4096_o),
    .b(_al_u4111_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J8cax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zdcbx6 ),
    .o(_al_u5743_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*~B)*~(C*A))"),
    .INIT(16'h5f4c))
    _al_u5744 (
    .a(_al_u4111_o),
    .b(_al_u4141_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J8cax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lg9bx6 ),
    .o(_al_u5744_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u5745 (
    .a(_al_u5737_o),
    .b(_al_u5742_o),
    .c(_al_u5743_o),
    .d(_al_u5744_o),
    .o(_al_u5745_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5746 (
    .a(_al_u4081_o),
    .b(_al_u4101_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cxcbx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G8ebx6 ),
    .o(_al_u5746_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(~D*~A))"),
    .INIT(16'h3f2a))
    _al_u5747 (
    .a(_al_u4035_o),
    .b(_al_u4106_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Facax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6cax6 ),
    .o(_al_u5747_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(~D*~A))"),
    .INIT(16'h3f2a))
    _al_u5748 (
    .a(_al_u4091_o),
    .b(_al_u4237_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F7jbx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tzgbx6 ),
    .o(_al_u5748_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*~B)*~(D*A))"),
    .INIT(16'h54fc))
    _al_u5749 (
    .a(_al_u4091_o),
    .b(_al_u4101_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cxcbx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tzgbx6 ),
    .o(_al_u5749_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf53f))
    _al_u575 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_ctrl [1]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_buf_full ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] ),
    .o(_al_u575_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u5750 (
    .a(_al_u5746_o),
    .b(_al_u5747_o),
    .c(_al_u5748_o),
    .d(_al_u5749_o),
    .o(_al_u5750_o));
  AL_MAP_LUT4 #(
    .EQN("((C@B)*(D@A))"),
    .INIT(16'h1428))
    _al_u5751 (
    .a(_al_u4076_o),
    .b(_al_u4184_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Evbax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zodbx6 ),
    .o(_al_u5751_o));
  AL_MAP_LUT4 #(
    .EQN("((D@B)*(C@A))"),
    .INIT(16'h1248))
    _al_u5752 (
    .a(_al_u4071_o),
    .b(_al_u4231_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bxbax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tfcax6 ),
    .o(_al_u5752_o));
  AL_MAP_LUT4 #(
    .EQN("((C@B)*(D@A))"),
    .INIT(16'h1428))
    _al_u5753 (
    .a(_al_u4086_o),
    .b(_al_u4131_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Koabx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nnfbx6 ),
    .o(_al_u5753_o));
  AL_MAP_LUT4 #(
    .EQN("((D@B)*(C@A))"),
    .INIT(16'h1248))
    _al_u5754 (
    .a(_al_u4056_o),
    .b(_al_u4219_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V0cax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xdcax6 ),
    .o(_al_u5754_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u5755 (
    .a(_al_u5751_o),
    .b(_al_u5752_o),
    .c(_al_u5753_o),
    .d(_al_u5754_o),
    .o(_al_u5755_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u5756 (
    .a(_al_u5735_o),
    .b(_al_u5745_o),
    .c(_al_u5750_o),
    .d(_al_u5755_o),
    .o(_al_u5756_o));
  AL_MAP_LUT4 #(
    .EQN("((C@B)*(D@A))"),
    .INIT(16'h1428))
    _al_u5757 (
    .a(_al_u4116_o),
    .b(_al_u4121_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bccax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rz8bx6 ),
    .o(_al_u5757_o));
  AL_MAP_LUT3 #(
    .EQN("(A*(C@B))"),
    .INIT(8'h28))
    _al_u5758 (
    .a(_al_u5757_o),
    .b(_al_u4061_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Knbbx6 ),
    .o(_al_u5758_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u5759 (
    .a(_al_u4423_o),
    .b(_al_u5756_o),
    .c(_al_u5758_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Opbax6 ),
    .o(_al_u5759_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(B*A))"),
    .INIT(8'h07))
    _al_u576 (
    .a(_al_u574_o),
    .b(_al_u575_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[4] ),
    .o(_al_u576_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u5760 (
    .a(_al_u5730_o),
    .b(_al_u5759_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dncax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Krbax6 ),
    .o(_al_u5760_o));
  AL_MAP_LUT4 #(
    .EQN("((C@B)*(D@A))"),
    .INIT(16'h1428))
    _al_u5761 (
    .a(_al_u4096_o),
    .b(_al_u4219_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J5eax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Thcbx6 ),
    .o(_al_u5761_o));
  AL_MAP_LUT4 #(
    .EQN("((D@B)*(C@A))"),
    .INIT(16'h1248))
    _al_u5762 (
    .a(_al_u4061_o),
    .b(_al_u4091_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Erbbx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N3hbx6 ),
    .o(_al_u5762_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u5763 (
    .a(_al_u4423_o),
    .b(_al_u5761_o),
    .c(_al_u5762_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahdax6 ),
    .o(_al_u5763_o));
  AL_MAP_LUT4 #(
    .EQN("((C@B)*(D@A))"),
    .INIT(16'h1428))
    _al_u5764 (
    .a(_al_u4035_o),
    .b(_al_u4101_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W0dbx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yxdax6 ),
    .o(_al_u5764_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*~B)*~(C*A))"),
    .INIT(16'h5f4c))
    _al_u5765 (
    .a(_al_u4081_o),
    .b(_al_u4191_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Acebx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tkdax6 ),
    .o(_al_u5765_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*(D@C))"),
    .INIT(16'h0880))
    _al_u5766 (
    .a(_al_u5764_o),
    .b(_al_u5765_o),
    .c(_al_u4225_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B9eax6 ),
    .o(_al_u5766_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(~C*~A))"),
    .INIT(16'h32fa))
    _al_u5767 (
    .a(_al_u4081_o),
    .b(_al_u4191_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Acebx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tkdax6 ),
    .o(_al_u5767_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*(D@C))"),
    .INIT(16'h0880))
    _al_u5768 (
    .a(_al_u5766_o),
    .b(_al_u5767_o),
    .c(_al_u4106_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R1eax6 ),
    .o(_al_u5768_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*~B)*~(C*A))"),
    .INIT(16'h5f4c))
    _al_u5769 (
    .a(_al_u4197_o),
    .b(_al_u4231_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bngax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F7eax6 ),
    .o(_al_u5769_o));
  AL_MAP_LUT4 #(
    .EQN("~(~B*~((~D*~C))*~(A)+~B*(~D*~C)*~(A)+~(~B)*(~D*~C)*A+~B*(~D*~C)*A)"),
    .INIT(16'heee4))
    _al_u577 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n25_lutinv ),
    .b(_al_u572_o),
    .c(_al_u573_o),
    .d(_al_u576_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/read_mux_byte0 [1]));
  AL_MAP_LUT4 #(
    .EQN("((D@B)*(C@A))"),
    .INIT(16'h1248))
    _al_u5770 (
    .a(_al_u4066_o),
    .b(_al_u4121_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kqdax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N3eax6 ),
    .o(_al_u5770_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*(D@C))"),
    .INIT(16'h0880))
    _al_u5771 (
    .a(_al_u5769_o),
    .b(_al_u5770_o),
    .c(_al_u4136_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eudax6 ),
    .o(_al_u5771_o));
  AL_MAP_LUT4 #(
    .EQN("((D@B)*(C@A))"),
    .INIT(16'h1248))
    _al_u5772 (
    .a(_al_u4126_o),
    .b(_al_u4237_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bwdax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xajbx6 ),
    .o(_al_u5772_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5773 (
    .a(_al_u4184_o),
    .b(_al_u4231_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F7eax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qmdax6 ),
    .o(_al_u5773_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*~B)*~(~D*~A))"),
    .INIT(16'hfca8))
    _al_u5774 (
    .a(_al_u4184_o),
    .b(_al_u4197_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bngax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qmdax6 ),
    .o(_al_u5774_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u5775 (
    .a(_al_u5771_o),
    .b(_al_u5772_o),
    .c(_al_u5773_o),
    .d(_al_u5774_o),
    .o(_al_u5775_o));
  AL_MAP_LUT4 #(
    .EQN("((D@B)*(C@A))"),
    .INIT(16'h1248))
    _al_u5776 (
    .a(_al_u4071_o),
    .b(_al_u4111_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nodax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzdax6 ),
    .o(_al_u5776_o));
  AL_MAP_LUT4 #(
    .EQN("((C@B)*(D@A))"),
    .INIT(16'h1428))
    _al_u5777 (
    .a(_al_u4086_o),
    .b(_al_u4131_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Esabx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hrfbx6 ),
    .o(_al_u5777_o));
  AL_MAP_LUT4 #(
    .EQN("((D@B)*(C@A))"),
    .INIT(16'h1248))
    _al_u5778 (
    .a(_al_u4056_o),
    .b(_al_u4116_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hsdax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J39bx6 ),
    .o(_al_u5778_o));
  AL_MAP_LUT4 #(
    .EQN("((C@B)*(D@A))"),
    .INIT(16'h1428))
    _al_u5779 (
    .a(_al_u4076_o),
    .b(_al_u4141_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dk9bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tsdbx6 ),
    .o(_al_u5779_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u578 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vowiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J3xiu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hw8ax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ws4iu6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u5780 (
    .a(_al_u5776_o),
    .b(_al_u5777_o),
    .c(_al_u5778_o),
    .d(_al_u5779_o),
    .o(_al_u5780_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u5781 (
    .a(_al_u5763_o),
    .b(_al_u5768_o),
    .c(_al_u5775_o),
    .d(_al_u5780_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Drhhu6_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u5782 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Drhhu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Widax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xaeax6 ),
    .o(_al_u5782_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5783 (
    .a(_al_u4101_o),
    .b(_al_u4225_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U4fax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zycbx6 ),
    .o(_al_u5783_o));
  AL_MAP_LUT3 #(
    .EQN("(A*(C@B))"),
    .INIT(8'h28))
    _al_u5784 (
    .a(_al_u5783_o),
    .b(_al_u4056_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aoeax6 ),
    .o(_al_u5784_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*~B)*~(~C*~A))"),
    .INIT(16'hfac8))
    _al_u5785 (
    .a(_al_u4071_o),
    .b(_al_u4136_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gkeax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xpeax6 ),
    .o(_al_u5785_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*(D@C))"),
    .INIT(16'h0880))
    _al_u5786 (
    .a(_al_u5784_o),
    .b(_al_u5785_o),
    .c(_al_u4237_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B9jbx6 ),
    .o(_al_u5786_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u5787 (
    .a(_al_u4096_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wfcbx6 ),
    .o(_al_u5787_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~A*(C@B))"),
    .INIT(16'h1400))
    _al_u5788 (
    .a(_al_u5787_o),
    .b(_al_u4184_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jieax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q6fax6 ),
    .o(_al_u5788_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u5789 (
    .a(_al_u4071_o),
    .b(_al_u4096_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gkeax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wfcbx6 ),
    .o(_al_u5789_o));
  AL_MAP_LUT2 #(
    .EQN("~(B*A)"),
    .INIT(4'h7))
    _al_u579 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ws4iu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dg2qw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bs4iu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5790 (
    .a(_al_u4035_o),
    .b(_al_u4121_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gzeax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rteax6 ),
    .o(_al_u5790_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u5791 (
    .a(_al_u5786_o),
    .b(_al_u5788_o),
    .c(_al_u5789_o),
    .d(_al_u5790_o),
    .o(_al_u5791_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(~D*~A))"),
    .INIT(16'h3f2a))
    _al_u5792 (
    .a(_al_u4101_o),
    .b(_al_u4126_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ureax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zycbx6 ),
    .o(_al_u5792_o));
  AL_MAP_LUT3 #(
    .EQN("(A*(C@B))"),
    .INIT(8'h28))
    _al_u5793 (
    .a(_al_u5792_o),
    .b(_al_u4106_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kxeax6 ),
    .o(_al_u5793_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*~B)*(C@A))"),
    .INIT(16'h5a48))
    _al_u5794 (
    .a(_al_u4081_o),
    .b(_al_u4131_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Daebx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hqabx6 ),
    .o(_al_u5794_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*~B)*~(C*A))"),
    .INIT(16'h5f4c))
    _al_u5795 (
    .a(_al_u4061_o),
    .b(_al_u4225_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hpbbx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U4fax6 ),
    .o(_al_u5795_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u5796 (
    .a(_al_u4131_o),
    .b(_al_u4136_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hqabx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xpeax6 ),
    .o(_al_u5796_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u5797 (
    .a(_al_u5794_o),
    .b(_al_u5795_o),
    .c(_al_u5796_o),
    .o(_al_u5797_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*~B)*~(~C*~A))"),
    .INIT(16'hfac8))
    _al_u5798 (
    .a(_al_u4061_o),
    .b(_al_u4126_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hpbbx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ureax6 ),
    .o(_al_u5798_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*~B)*~(~D*~A))"),
    .INIT(16'hfca8))
    _al_u5799 (
    .a(_al_u4035_o),
    .b(_al_u4121_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gzeax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rteax6 ),
    .o(_al_u5799_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u580 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [7]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [8]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [9]),
    .o(_al_u580_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u5800 (
    .a(_al_u5793_o),
    .b(_al_u5797_o),
    .c(_al_u5798_o),
    .d(_al_u5799_o),
    .o(_al_u5800_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u5801 (
    .a(_al_u4423_o),
    .b(_al_u5791_o),
    .c(_al_u5800_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tceax6 ),
    .o(_al_u5801_o));
  AL_MAP_LUT4 #(
    .EQN("((C@B)*(D@A))"),
    .INIT(16'h1428))
    _al_u5802 (
    .a(_al_u4091_o),
    .b(_al_u4191_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mgeax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q1hbx6 ),
    .o(_al_u5802_o));
  AL_MAP_LUT4 #(
    .EQN("((D@B)*(C@A))"),
    .INIT(16'h1248))
    _al_u5803 (
    .a(_al_u4066_o),
    .b(_al_u4141_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dmeax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hi9bx6 ),
    .o(_al_u5803_o));
  AL_MAP_LUT4 #(
    .EQN("((C@B)*(D@A))"),
    .INIT(16'h1428))
    _al_u5804 (
    .a(_al_u4076_o),
    .b(_al_u4111_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oveax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wqdbx6 ),
    .o(_al_u5804_o));
  AL_MAP_LUT4 #(
    .EQN("((D@B)*(C@A))"),
    .INIT(16'h1248))
    _al_u5805 (
    .a(_al_u4219_o),
    .b(_al_u4231_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C1fax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y2fax6 ),
    .o(_al_u5805_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u5806 (
    .a(_al_u5802_o),
    .b(_al_u5803_o),
    .c(_al_u5804_o),
    .d(_al_u5805_o),
    .o(_al_u5806_o));
  AL_MAP_LUT4 #(
    .EQN("((C@B)*(D@A))"),
    .INIT(16'h1428))
    _al_u5807 (
    .a(_al_u4116_o),
    .b(_al_u4197_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Elgax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N19bx6 ),
    .o(_al_u5807_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*(D@C))"),
    .INIT(16'h0880))
    _al_u5808 (
    .a(_al_u5806_o),
    .b(_al_u5807_o),
    .c(_al_u4086_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kpfbx6 ),
    .o(_al_u5808_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u5809 (
    .a(_al_u5801_o),
    .b(_al_u5808_o),
    .o(_al_u5809_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u581 (
    .a(_al_u580_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [10]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [11]),
    .o(_al_u581_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*A*~(D*C))"),
    .INIT(16'h0222))
    _al_u5810 (
    .a(_al_u5760_o),
    .b(_al_u5782_o),
    .c(_al_u5809_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Peeax6 ),
    .o(_al_u5810_o));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*C)*~(~B*A))"),
    .INIT(16'hf222))
    _al_u5811 (
    .a(_al_u5706_o),
    .b(_al_u5810_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jvvpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dhvhu6 ));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u5812 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Drhhu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eagax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xaeax6 ),
    .o(_al_u5812_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u5813 (
    .a(_al_u5730_o),
    .b(_al_u5809_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bcgax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H8gax6 ),
    .o(_al_u5813_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(D*C))"),
    .INIT(16'h0444))
    _al_u5814 (
    .a(_al_u5812_o),
    .b(_al_u5813_o),
    .c(_al_u5759_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K6gax6 ),
    .o(_al_u5814_o));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*C)*~(~B*A))"),
    .INIT(16'hf222))
    _al_u5815 (
    .a(_al_u5706_o),
    .b(_al_u5814_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pexpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Khvhu6 ));
  AL_MAP_LUT4 #(
    .EQN("(D*~A*~(C*B))"),
    .INIT(16'h1500))
    _al_u5816 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lf1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iqzhu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nmfax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tb3qw6 ),
    .o(_al_u5816_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*A)"),
    .INIT(16'h0080))
    _al_u5817 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tszhu6 ),
    .b(_al_u5816_o),
    .c(_al_u4492_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J0gax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oa4iu6 ));
  AL_MAP_LUT4 #(
    .EQN("~((C*B)*~(D)*~(A)+(C*B)*D*~(A)+~((C*B))*D*A+(C*B)*D*A)"),
    .INIT(16'h15bf))
    _al_u5818 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oa4iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n382 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yf1qw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vrkbx6 [10]),
    .o(_al_u5818_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C*~A))"),
    .INIT(8'h73))
    _al_u5819 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n382 ),
    .b(_al_u5818_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ym4iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N6xhu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u582 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [5]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [6]),
    .o(_al_u582_o));
  AL_MAP_LUT4 #(
    .EQN("~((C*B)*~(D)*~(A)+(C*B)*D*~(A)+~((C*B))*D*A+(C*B)*D*A)"),
    .INIT(16'h15bf))
    _al_u5820 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oa4iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n382 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ke1qw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vrkbx6 [9]),
    .o(_al_u5820_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C*~A))"),
    .INIT(8'h73))
    _al_u5821 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n382 ),
    .b(_al_u5820_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pl4iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U6xhu6 ));
  AL_MAP_LUT4 #(
    .EQN("~((C*B)*~(D)*~(A)+(C*B)*D*~(A)+~((C*B))*D*A+(C*B)*D*A)"),
    .INIT(16'h15bf))
    _al_u5822 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oa4iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n382 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nd3qw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vrkbx6 [8]),
    .o(_al_u5822_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C*~A))"),
    .INIT(8'h73))
    _al_u5823 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n382 ),
    .b(_al_u5822_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gk4iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B7xhu6 ));
  AL_MAP_LUT4 #(
    .EQN("~((C*B)*~(D)*~(A)+(C*B)*D*~(A)+~((C*B))*D*A+(C*B)*D*A)"),
    .INIT(16'h15bf))
    _al_u5824 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oa4iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n382 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vn9bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vrkbx6 [7]),
    .o(_al_u5824_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C*~A))"),
    .INIT(8'h73))
    _al_u5825 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n382 ),
    .b(_al_u5824_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xi4iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I7xhu6 ));
  AL_MAP_LUT4 #(
    .EQN("~((C*B)*~(D)*~(A)+(C*B)*D*~(A)+~((C*B))*D*A+(C*B)*D*A)"),
    .INIT(16'h15bf))
    _al_u5826 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oa4iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n382 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bf3qw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vrkbx6 [6]),
    .o(_al_u5826_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C*~A))"),
    .INIT(8'h73))
    _al_u5827 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n382 ),
    .b(_al_u5826_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oh4iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P7xhu6 ));
  AL_MAP_LUT4 #(
    .EQN("~((C*B)*~(D)*~(A)+(C*B)*D*~(A)+~((C*B))*D*A+(C*B)*D*A)"),
    .INIT(16'h15bf))
    _al_u5828 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oa4iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n382 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pg3qw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vrkbx6 [5]),
    .o(_al_u5828_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C*~A))"),
    .INIT(8'h73))
    _al_u5829 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n382 ),
    .b(_al_u5828_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H34iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W7xhu6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u583 (
    .a(_al_u581_o),
    .b(_al_u582_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n24_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("~((C*B)*~(D)*~(A)+(C*B)*D*~(A)+~((C*B))*D*A+(C*B)*D*A)"),
    .INIT(16'h15bf))
    _al_u5830 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oa4iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n382 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P23qw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vrkbx6 [4]),
    .o(_al_u5830_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C*~A))"),
    .INIT(8'h73))
    _al_u5831 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n382 ),
    .b(_al_u5830_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Df4iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D8xhu6 ));
  AL_MAP_LUT4 #(
    .EQN("~((C*B)*~(D)*~(A)+(C*B)*D*~(A)+~((C*B))*D*A+(C*B)*D*A)"),
    .INIT(16'h15bf))
    _al_u5832 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oa4iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n382 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xn7ax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vrkbx6 [3]),
    .o(_al_u5832_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C*~A))"),
    .INIT(8'h73))
    _al_u5833 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n382 ),
    .b(_al_u5832_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ud4iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K8xhu6 ));
  AL_MAP_LUT4 #(
    .EQN("~((C*B)*~(D)*~(A)+(C*B)*D*~(A)+~((C*B))*D*A+(C*B)*D*A)"),
    .INIT(16'h15bf))
    _al_u5834 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oa4iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n382 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vj3qw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vrkbx6 [2]),
    .o(_al_u5834_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C*~A))"),
    .INIT(8'h73))
    _al_u5835 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n382 ),
    .b(_al_u5834_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O34iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R8xhu6 ));
  AL_MAP_LUT4 #(
    .EQN("~((C*~B)*~(D)*~(A)+(C*~B)*D*~(A)+~((C*~B))*D*A+(C*~B)*D*A)"),
    .INIT(16'h45ef))
    _al_u5836 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oa4iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n382 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T24iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vrkbx6 [1]),
    .o(_al_u5836_o));
  AL_MAP_LUT4 #(
    .EQN("~(A*~(D*C*~B))"),
    .INIT(16'h7555))
    _al_u5837 (
    .a(_al_u5836_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oa4iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n382 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qehbx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y8xhu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h5ff3))
    _al_u5838 (
    .a(_al_u696_o),
    .b(_al_u932_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ejaju6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C*~B*A))"),
    .INIT(16'hdf00))
    _al_u5839 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xiaju6 ),
    .b(_al_u4351_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ejaju6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vgjpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mt4ju6 ));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(~B*~(~C*~A)))"),
    .INIT(16'h00cd))
    _al_u584 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [0]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [1]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOSIZE [0]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOSIZE [1]),
    .o(_al_u584_o));
  AL_MAP_LUT4 #(
    .EQN("(A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hc8f8))
    _al_u5840 (
    .a(_al_u1344_o),
    .b(_al_u2403_o),
    .c(_al_u3826_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tt4ju6_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u5841 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mt4ju6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tt4ju6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wc5ju6_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u5842 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qyniu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nkaju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vgjpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ys4ju6 ));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~((C*A))*~(B)+~D*(C*A)*~(B)+~(~D)*(C*A)*B+~D*(C*A)*B)"),
    .INIT(16'h7f4c))
    _al_u5843 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D5epw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/To2ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wc5ju6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ys4ju6 ),
    .o(_al_u5843_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u5844 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mt4ju6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ys4ju6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cg5ju6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(A*~(~B*~(~D*C)))"),
    .INIT(16'h88a8))
    _al_u5845 (
    .a(_al_u5843_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D5epw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/To2ju6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cg5ju6_lutinv ),
    .o(_al_u5845_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*A)"),
    .INIT(16'h0080))
    _al_u5846 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vo3ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D31ju6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vgjpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T05ju6 ));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u5847 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T05ju6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rskax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ubypw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I55ju6 ));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u5848 (
    .a(_al_u606_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vgjpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ),
    .o(_al_u5848_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~B*~(D*A))"),
    .INIT(16'h0103))
    _al_u5849 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I55ju6 ),
    .b(_al_u5848_o),
    .c(n1[13]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_apsr_o[3] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N45ju6 ));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*~A)"),
    .INIT(16'h4000))
    _al_u585 (
    .a(_al_u584_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOTRANS ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOWRITE ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/IOSEL ),
    .o(_al_u585_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~A*~(~D*B))"),
    .INIT(16'h0501))
    _al_u5850 (
    .a(_al_u1296_o),
    .b(_al_u1329_o),
    .c(_al_u1662_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ),
    .o(_al_u5850_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(C*A))"),
    .INIT(16'h4c5f))
    _al_u5851 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Difiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 ),
    .o(_al_u5851_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(B*~(~C*~A)))"),
    .INIT(16'h3700))
    _al_u5852 (
    .a(_al_u5850_o),
    .b(_al_u5851_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vgjpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/By4ju6 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u5853 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N45ju6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/By4ju6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [32]),
    .o(_al_u5853_o));
  AL_MAP_LUT4 #(
    .EQN("(D*A*~(~C*~B))"),
    .INIT(16'ha800))
    _al_u5854 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yljiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Owoiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vgjpw6 ),
    .o(_al_u5854_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*~(D*~B))"),
    .INIT(16'h4050))
    _al_u5855 (
    .a(_al_u5845_o),
    .b(_al_u2281_o),
    .c(_al_u5853_o),
    .d(_al_u5854_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bbliu6 ));
  AL_MAP_LUT4 #(
    .EQN("(A*~(~D*~(C)*~(B)+~D*C*~(B)+~(~D)*C*B+~D*C*B))"),
    .INIT(16'h2a08))
    _al_u5856 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [30]),
    .b(_al_u1541_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wc5ju6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ys4ju6 ),
    .o(_al_u5856_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~B*~(D*A))"),
    .INIT(16'h0103))
    _al_u5857 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I55ju6 ),
    .b(_al_u5848_o),
    .c(n1[12]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_apsr_o[2] ),
    .o(_al_u5857_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u5858 (
    .a(_al_u5857_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/By4ju6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [31]),
    .o(_al_u5858_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*~A))"),
    .INIT(8'h8c))
    _al_u5859 (
    .a(_al_u2270_o),
    .b(_al_u5858_o),
    .c(_al_u5854_o),
    .o(_al_u5859_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~A*~(D*~C)))"),
    .INIT(16'h8c88))
    _al_u586 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n24_lutinv ),
    .b(_al_u585_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [10]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [11]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n39 ));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~D*C*~A))"),
    .INIT(16'hcc8c))
    _al_u5860 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [30]),
    .b(_al_u5859_o),
    .c(_al_u1541_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cg5ju6_lutinv ),
    .o(_al_u5860_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*~B*A)"),
    .INIT(16'h0020))
    _al_u5861 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bbliu6 ),
    .b(_al_u5856_o),
    .c(_al_u5860_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fpnpw6 ),
    .o(_al_u5861_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~C*~(D*A)))"),
    .INIT(16'hc8c0))
    _al_u5862 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [29]),
    .b(_al_u1533_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mt4ju6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tt4ju6_lutinv ),
    .o(_al_u5862_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~B*~(D*A))"),
    .INIT(16'h0103))
    _al_u5863 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I55ju6 ),
    .b(_al_u5848_o),
    .c(n1[11]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_apsr_o[1] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J77ju6 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u5864 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J77ju6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/By4ju6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [30]),
    .o(_al_u5864_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*~(D*~B))"),
    .INIT(16'h4050))
    _al_u5865 (
    .a(_al_u5862_o),
    .b(_al_u2429_o),
    .c(_al_u5864_o),
    .d(_al_u5854_o),
    .o(_al_u5865_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D*(C@B)))"),
    .INIT(16'h82aa))
    _al_u5866 (
    .a(_al_u5865_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [29]),
    .c(_al_u1533_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ys4ju6 ),
    .o(_al_u5866_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'h0213))
    _al_u5867 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [25]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mi8ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wc5ju6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cg5ju6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yh8ju6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(~C*~B*~(D*A))"),
    .INIT(16'h0103))
    _al_u5868 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/By4ju6 ),
    .b(_al_u5848_o),
    .c(n1[7]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [26]),
    .o(_al_u5868_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*~A))"),
    .INIT(8'h8c))
    _al_u5869 (
    .a(_al_u2261_o),
    .b(_al_u5868_o),
    .c(_al_u5854_o),
    .o(_al_u5869_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(~B*~(~C*A)))"),
    .INIT(16'h00ce))
    _al_u587 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [0]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [1]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOSIZE [0]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOSIZE [1]),
    .o(_al_u587_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(D*C*A))"),
    .INIT(16'h4ccc))
    _al_u5870 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [25]),
    .b(_al_u5869_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mi8ju6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ys4ju6 ),
    .o(_al_u5870_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u5871 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yh8ju6_lutinv ),
    .b(_al_u5870_o),
    .o(_al_u5871_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u5872 (
    .a(_al_u5861_o),
    .b(_al_u5866_o),
    .c(_al_u5871_o),
    .o(_al_u5872_o));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u5873 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [0]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Go0iu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ys4ju6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tt4ju6_lutinv ),
    .o(_al_u5873_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u5874 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T05ju6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rskax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ubypw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_primask_o ),
    .o(_al_u5874_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u5875 (
    .a(_al_u5874_o),
    .b(_al_u5848_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_0 ),
    .o(_al_u5875_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u5876 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T05ju6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sqkax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ubypw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pk4ju6 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u5877 (
    .a(_al_u5875_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pk4ju6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[0] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wy4ju6 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u5878 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wy4ju6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/By4ju6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [1]),
    .o(_al_u5878_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(D*~C))"),
    .INIT(16'h4044))
    _al_u5879 (
    .a(_al_u5873_o),
    .b(_al_u5878_o),
    .c(_al_u1882_o),
    .d(_al_u5854_o),
    .o(_al_u5879_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*~A)"),
    .INIT(16'h4000))
    _al_u588 (
    .a(_al_u587_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOTRANS ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOWRITE ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/IOSEL ),
    .o(_al_u588_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~C*~(D*~A)))"),
    .INIT(16'hc4c0))
    _al_u5880 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [0]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Go0iu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mt4ju6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ys4ju6 ),
    .o(_al_u5880_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u5881 (
    .a(_al_u5879_o),
    .b(_al_u5880_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ibliu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'h0213))
    _al_u5882 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q5phu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N18ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wc5ju6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cg5ju6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z08ju6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(~D*~B*~(C*A))"),
    .INIT(16'h0013))
    _al_u5883 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/By4ju6 ),
    .b(_al_u5848_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [10]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_9 ),
    .o(_al_u5883_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*~A))"),
    .INIT(8'h8c))
    _al_u5884 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I28ju6 ),
    .b(_al_u5883_o),
    .c(_al_u5854_o),
    .o(_al_u5884_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(D*C*A))"),
    .INIT(16'h4ccc))
    _al_u5885 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q5phu6 ),
    .b(_al_u5884_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N18ju6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ys4ju6 ),
    .o(_al_u5885_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u5886 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z08ju6_lutinv ),
    .b(_al_u5885_o),
    .o(_al_u5886_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u5887 (
    .a(_al_u5872_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ibliu6 ),
    .c(_al_u5886_o),
    .o(_al_u5887_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'h0213))
    _al_u5888 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E2epw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mk6ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wc5ju6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cg5ju6_lutinv ),
    .o(_al_u5888_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~B*~(C*A))"),
    .INIT(16'h0013))
    _al_u5889 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/By4ju6 ),
    .b(_al_u5848_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [7]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_6 ),
    .o(_al_u5889_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u589 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [10]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [11]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n26_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*~A))"),
    .INIT(8'h8c))
    _al_u5890 (
    .a(_al_u1952_o),
    .b(_al_u5889_o),
    .c(_al_u5854_o),
    .o(_al_u5890_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(D*C*A))"),
    .INIT(16'h4ccc))
    _al_u5891 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E2epw6 ),
    .b(_al_u5890_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mk6ju6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ys4ju6 ),
    .o(_al_u5891_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u5892 (
    .a(_al_u5888_o),
    .b(_al_u5891_o),
    .o(_al_u5892_o));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~((C*A))*~(B)+~D*(C*A)*~(B)+~(~D)*(C*A)*B+~D*(C*A)*B)"),
    .INIT(16'h7f4c))
    _al_u5893 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [24]),
    .b(_al_u1493_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wc5ju6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ys4ju6 ),
    .o(_al_u5893_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(~B*~(~D*C)))"),
    .INIT(16'h88a8))
    _al_u5894 (
    .a(_al_u5893_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [24]),
    .c(_al_u1493_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cg5ju6_lutinv ),
    .o(_al_u5894_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~B*~(D*A))"),
    .INIT(16'h0103))
    _al_u5895 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/By4ju6 ),
    .b(_al_u5848_o),
    .c(n1[6]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [25]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ww6ju6 ));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*~(D*~B))"),
    .INIT(16'h4050))
    _al_u5896 (
    .a(_al_u5894_o),
    .b(_al_u2439_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ww6ju6 ),
    .d(_al_u5854_o),
    .o(_al_u5896_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~C*~(D*A)))"),
    .INIT(16'hc8c0))
    _al_u5897 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [28]),
    .b(_al_u1525_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mt4ju6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tt4ju6_lutinv ),
    .o(_al_u5897_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~B*~(D*A))"),
    .INIT(16'h0103))
    _al_u5898 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I55ju6 ),
    .b(_al_u5848_o),
    .c(n1[10]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_apsr_o[0] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ok7ju6 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u5899 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ok7ju6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/By4ju6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [29]),
    .o(_al_u5899_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    _al_u590 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n24_lutinv ),
    .b(_al_u588_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n26_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n34 ));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*~(D*~B))"),
    .INIT(16'h4050))
    _al_u5900 (
    .a(_al_u5897_o),
    .b(_al_u2420_o),
    .c(_al_u5899_o),
    .d(_al_u5854_o),
    .o(_al_u5900_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D*(C@B)))"),
    .INIT(16'h82aa))
    _al_u5901 (
    .a(_al_u5900_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [28]),
    .c(_al_u1525_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ys4ju6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kgoiu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'h0213))
    _al_u5902 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [27]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F57ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wc5ju6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cg5ju6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R47ju6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(~C*~B*~(D*A))"),
    .INIT(16'h0103))
    _al_u5903 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/By4ju6 ),
    .b(_al_u5848_o),
    .c(n1[9]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [28]),
    .o(_al_u5903_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*~A))"),
    .INIT(8'h8c))
    _al_u5904 (
    .a(_al_u2447_o),
    .b(_al_u5903_o),
    .c(_al_u5854_o),
    .o(_al_u5904_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(D*C*A))"),
    .INIT(16'h4ccc))
    _al_u5905 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [27]),
    .b(_al_u5904_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F57ju6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ys4ju6 ),
    .o(_al_u5905_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u5906 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R47ju6_lutinv ),
    .b(_al_u5905_o),
    .o(_al_u5906_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'h0213))
    _al_u5907 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [26]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E17ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wc5ju6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cg5ju6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q07ju6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(~C*~B*~(D*A))"),
    .INIT(16'h0103))
    _al_u5908 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/By4ju6 ),
    .b(_al_u5848_o),
    .c(n1[8]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [27]),
    .o(_al_u5908_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*~A))"),
    .INIT(8'h8c))
    _al_u5909 (
    .a(_al_u2455_o),
    .b(_al_u5908_o),
    .c(_al_u5854_o),
    .o(_al_u5909_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*~A)"),
    .INIT(16'h4000))
    _al_u591 (
    .a(_al_u584_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOSEL ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOTRANS ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOWRITE ),
    .o(_al_u591_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(D*C*A))"),
    .INIT(16'h4ccc))
    _al_u5910 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [26]),
    .b(_al_u5909_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E17ju6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ys4ju6 ),
    .o(_al_u5910_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u5911 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q07ju6_lutinv ),
    .b(_al_u5910_o),
    .o(_al_u5911_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u5912 (
    .a(_al_u5896_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kgoiu6 ),
    .c(_al_u5906_o),
    .d(_al_u5911_o),
    .o(_al_u5912_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u5913 (
    .a(_al_u5887_o),
    .b(_al_u5892_o),
    .c(_al_u5912_o),
    .o(_al_u5913_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'h084c))
    _al_u5914 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4epw6 ),
    .b(_al_u1608_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wc5ju6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cg5ju6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cs7ju6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(~D*~B*~(C*A))"),
    .INIT(16'h0013))
    _al_u5915 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/By4ju6 ),
    .b(_al_u5848_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [9]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_8 ),
    .o(_al_u5915_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*~A))"),
    .INIT(8'h8c))
    _al_u5916 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cz7ju6 ),
    .b(_al_u5915_o),
    .c(_al_u5854_o),
    .o(_al_u5916_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D*~B*A))"),
    .INIT(16'hd0f0))
    _al_u5917 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4epw6 ),
    .b(_al_u1608_o),
    .c(_al_u5916_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ys4ju6 ),
    .o(_al_u5917_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u5918 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cs7ju6_lutinv ),
    .b(_al_u5917_o),
    .o(_al_u5918_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'h084c))
    _al_u5919 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z2epw6 ),
    .b(_al_u1429_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wc5ju6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cg5ju6_lutinv ),
    .o(_al_u5919_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~A*~(D*~C)))"),
    .INIT(16'h8c88))
    _al_u592 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n24_lutinv ),
    .b(_al_u591_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [10]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [11]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n39 ));
  AL_MAP_LUT4 #(
    .EQN("(~D*~B*~(C*A))"),
    .INIT(16'h0013))
    _al_u5920 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/By4ju6 ),
    .b(_al_u5848_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [17]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_16 ),
    .o(_al_u5920_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*~A))"),
    .INIT(8'h8c))
    _al_u5921 (
    .a(_al_u2289_o),
    .b(_al_u5920_o),
    .c(_al_u5854_o),
    .o(_al_u5921_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(D*~C*A))"),
    .INIT(16'hc4cc))
    _al_u5922 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z2epw6 ),
    .b(_al_u5921_o),
    .c(_al_u1429_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ys4ju6 ),
    .o(_al_u5922_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u5923 (
    .a(_al_u5919_o),
    .b(_al_u5922_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vdmiu6 ));
  AL_MAP_LUT4 #(
    .EQN("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'h084c))
    _al_u5924 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N3epw6 ),
    .b(_al_u1445_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wc5ju6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cg5ju6_lutinv ),
    .o(_al_u5924_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~B*~(D*A))"),
    .INIT(16'h0103))
    _al_u5925 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/By4ju6 ),
    .b(_al_u5848_o),
    .c(n1[0]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [19]),
    .o(_al_u5925_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*~A))"),
    .INIT(8'h8c))
    _al_u5926 (
    .a(_al_u2208_o),
    .b(_al_u5925_o),
    .c(_al_u5854_o),
    .o(_al_u5926_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(D*~C*A))"),
    .INIT(16'hc4cc))
    _al_u5927 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N3epw6 ),
    .b(_al_u5926_o),
    .c(_al_u1445_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ys4ju6 ),
    .o(_al_u5927_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u5928 (
    .a(_al_u5924_o),
    .b(_al_u5927_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X7miu6 ));
  AL_MAP_LUT4 #(
    .EQN("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'h084c))
    _al_u5929 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J1epw6 ),
    .b(_al_u1397_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wc5ju6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cg5ju6_lutinv ),
    .o(_al_u5929_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*~A)"),
    .INIT(16'h4000))
    _al_u593 (
    .a(_al_u587_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOSEL ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOTRANS ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOWRITE ),
    .o(_al_u593_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~B*~(C*A))"),
    .INIT(16'h0013))
    _al_u5930 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/By4ju6 ),
    .b(_al_u5848_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [13]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_12 ),
    .o(_al_u5930_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*~A))"),
    .INIT(8'h8c))
    _al_u5931 (
    .a(_al_u2084_o),
    .b(_al_u5930_o),
    .c(_al_u5854_o),
    .o(_al_u5931_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(D*~C*A))"),
    .INIT(16'hc4cc))
    _al_u5932 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J1epw6 ),
    .b(_al_u5931_o),
    .c(_al_u1397_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ys4ju6 ),
    .o(_al_u5932_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u5933 (
    .a(_al_u5929_o),
    .b(_al_u5932_o),
    .o(_al_u5933_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u5934 (
    .a(_al_u5918_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vdmiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X7miu6 ),
    .d(_al_u5933_o),
    .o(_al_u5934_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'h084c))
    _al_u5935 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U3epw6 ),
    .b(_al_u1453_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wc5ju6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cg5ju6_lutinv ),
    .o(_al_u5935_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~B*~(D*A))"),
    .INIT(16'h0103))
    _al_u5936 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/By4ju6 ),
    .b(_al_u5848_o),
    .c(n1[1]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [20]),
    .o(_al_u5936_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*~A))"),
    .INIT(8'h8c))
    _al_u5937 (
    .a(_al_u2217_o),
    .b(_al_u5936_o),
    .c(_al_u5854_o),
    .o(_al_u5937_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(D*~C*A))"),
    .INIT(16'hc4cc))
    _al_u5938 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U3epw6 ),
    .b(_al_u5937_o),
    .c(_al_u1453_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ys4ju6 ),
    .o(_al_u5938_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u5939 (
    .a(_al_u5935_o),
    .b(_al_u5938_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y4miu6 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    _al_u594 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n24_lutinv ),
    .b(_al_u593_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n26_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n34 ));
  AL_MAP_LUT4 #(
    .EQN("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'h084c))
    _al_u5940 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B4epw6 ),
    .b(_al_u1461_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wc5ju6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cg5ju6_lutinv ),
    .o(_al_u5940_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~B*~(D*A))"),
    .INIT(16'h0103))
    _al_u5941 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/By4ju6 ),
    .b(_al_u5848_o),
    .c(n1[2]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [21]),
    .o(_al_u5941_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*~A))"),
    .INIT(8'h8c))
    _al_u5942 (
    .a(_al_u2225_o),
    .b(_al_u5941_o),
    .c(_al_u5854_o),
    .o(_al_u5942_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(D*~C*A))"),
    .INIT(16'hc4cc))
    _al_u5943 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B4epw6 ),
    .b(_al_u5942_o),
    .c(_al_u1461_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ys4ju6 ),
    .o(_al_u5943_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u5944 (
    .a(_al_u5940_o),
    .b(_al_u5943_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z1miu6 ));
  AL_MAP_LUT4 #(
    .EQN("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'h084c))
    _al_u5945 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I4epw6 ),
    .b(_al_u1469_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wc5ju6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cg5ju6_lutinv ),
    .o(_al_u5945_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~B*~(D*A))"),
    .INIT(16'h0103))
    _al_u5946 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/By4ju6 ),
    .b(_al_u5848_o),
    .c(n1[3]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [22]),
    .o(_al_u5946_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*~A))"),
    .INIT(8'h8c))
    _al_u5947 (
    .a(_al_u2235_o),
    .b(_al_u5946_o),
    .c(_al_u5854_o),
    .o(_al_u5947_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(D*~C*A))"),
    .INIT(16'hc4cc))
    _al_u5948 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I4epw6 ),
    .b(_al_u5947_o),
    .c(_al_u1469_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ys4ju6 ),
    .o(_al_u5948_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u5949 (
    .a(_al_u5945_o),
    .b(_al_u5948_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Azliu6 ));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    _al_u595 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reload_i ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/BAUDTICK ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n48 ));
  AL_MAP_LUT4 #(
    .EQN("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'h084c))
    _al_u5950 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q1epw6 ),
    .b(_al_u1405_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wc5ju6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cg5ju6_lutinv ),
    .o(_al_u5950_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~B*~(C*A))"),
    .INIT(16'h0013))
    _al_u5951 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/By4ju6 ),
    .b(_al_u5848_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [14]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_13 ),
    .o(_al_u5951_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*~A))"),
    .INIT(8'h8c))
    _al_u5952 (
    .a(_al_u2106_o),
    .b(_al_u5951_o),
    .c(_al_u5854_o),
    .o(_al_u5952_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(D*~C*A))"),
    .INIT(16'hc4cc))
    _al_u5953 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q1epw6 ),
    .b(_al_u5952_o),
    .c(_al_u1405_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ys4ju6 ),
    .o(_al_u5953_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u5954 (
    .a(_al_u5950_o),
    .b(_al_u5953_o),
    .o(_al_u5954_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u5955 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y4miu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z1miu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Azliu6 ),
    .d(_al_u5954_o),
    .o(_al_u5955_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u5956 (
    .a(_al_u5913_o),
    .b(_al_u5934_o),
    .c(_al_u5955_o),
    .o(_al_u5956_o));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~((C*A))*~(B)+~D*(C*A)*~(B)+~(~D)*(C*A)*B+~D*(C*A)*B)"),
    .INIT(16'h7f4c))
    _al_u5957 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [3]),
    .b(_al_u1592_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wc5ju6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ys4ju6 ),
    .o(_al_u5957_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(~B*~(~D*C)))"),
    .INIT(16'h88a8))
    _al_u5958 (
    .a(_al_u5957_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [3]),
    .c(_al_u1592_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cg5ju6_lutinv ),
    .o(_al_u5958_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(B*A))"),
    .INIT(8'h07))
    _al_u5959 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hlliu6 ),
    .b(_al_u5848_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_3 ),
    .o(_al_u5959_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*A)"),
    .INIT(16'h0200))
    _al_u596 (
    .a(_al_u379_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_state [0]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_state [1]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_buf_full ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n61 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u5960 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pk4ju6 ),
    .b(_al_u5959_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[3] ),
    .o(_al_u5960_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u5961 (
    .a(_al_u5960_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/By4ju6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [4]),
    .o(_al_u5961_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*~(D*~B))"),
    .INIT(16'h4050))
    _al_u5962 (
    .a(_al_u5958_o),
    .b(_al_u1925_o),
    .c(_al_u5961_o),
    .d(_al_u5854_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dkkiu6 ));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~((C*A))*~(B)+~D*(C*A)*~(B)+~(~D)*(C*A)*B+~D*(C*A)*B)"),
    .INIT(16'h7f4c))
    _al_u5963 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [5]),
    .b(_al_u1600_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wc5ju6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ys4ju6 ),
    .o(_al_u5963_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(~B*~(~D*C)))"),
    .INIT(16'h88a8))
    _al_u5964 (
    .a(_al_u5963_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [5]),
    .c(_al_u1600_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cg5ju6_lutinv ),
    .o(_al_u5964_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~B*~(C*A))"),
    .INIT(16'h0013))
    _al_u5965 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pk4ju6 ),
    .b(_al_u5848_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[5] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_5 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I46ju6 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u5966 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I46ju6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/By4ju6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [6]),
    .o(_al_u5966_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*~(D*~B))"),
    .INIT(16'h4050))
    _al_u5967 (
    .a(_al_u5964_o),
    .b(_al_u1943_o),
    .c(_al_u5966_o),
    .d(_al_u5854_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lokiu6 ));
  AL_MAP_LUT4 #(
    .EQN("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'h084c))
    _al_u5968 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S2epw6 ),
    .b(_al_u1616_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wc5ju6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cg5ju6_lutinv ),
    .o(_al_u5968_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~B*~(C*A))"),
    .INIT(16'h0013))
    _al_u5969 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/By4ju6 ),
    .b(_al_u5848_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [8]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_7 ),
    .o(_al_u5969_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*C)*~(B*A))"),
    .INIT(16'h0777))
    _al_u597 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n61 ),
    .b(uart0_txen_pad),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_state [2]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_state [3]),
    .o(_al_u597_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*~A))"),
    .INIT(8'h8c))
    _al_u5970 (
    .a(_al_u1961_o),
    .b(_al_u5969_o),
    .c(_al_u5854_o),
    .o(_al_u5970_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(D*~C*A))"),
    .INIT(16'hc4cc))
    _al_u5971 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S2epw6 ),
    .b(_al_u5970_o),
    .c(_al_u1616_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ys4ju6 ),
    .o(_al_u5971_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u5972 (
    .a(_al_u5968_o),
    .b(_al_u5971_o),
    .o(_al_u5972_o));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~((C*A))*~(B)+~D*(C*A)*~(B)+~(~D)*(C*A)*B+~D*(C*A)*B)"),
    .INIT(16'h7f4c))
    _al_u5973 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [1]),
    .b(_al_u1354_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wc5ju6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ys4ju6 ),
    .o(_al_u5973_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(~B*~(~D*C)))"),
    .INIT(16'h88a8))
    _al_u5974 (
    .a(_al_u5973_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [1]),
    .c(_al_u1354_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cg5ju6_lutinv ),
    .o(_al_u5974_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u5975 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T05ju6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_control_o ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rskax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ubypw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rb7ju6 ));
  AL_MAP_LUT4 #(
    .EQN("(~D*~B*~(C*A))"),
    .INIT(16'h0013))
    _al_u5976 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pk4ju6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rb7ju6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[1] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_1 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pa7ju6 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u5977 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pa7ju6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/By4ju6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [2]),
    .o(_al_u5977_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*~(D*~B))"),
    .INIT(16'h4050))
    _al_u5978 (
    .a(_al_u5974_o),
    .b(_al_u1968_o),
    .c(_al_u5977_o),
    .d(_al_u5854_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bpliu6 ));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u5979 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dkkiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lokiu6 ),
    .c(_al_u5972_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bpliu6 ),
    .o(_al_u5979_o));
  AL_MAP_LUT2 #(
    .EQN("~(B*~A)"),
    .INIT(4'hb))
    _al_u598 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_state_inc ),
    .b(_al_u597_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_state_update ));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(B*~A))"),
    .INIT(8'h0b))
    _al_u5980 (
    .a(_al_u1581_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mt4ju6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ys4ju6 ),
    .o(_al_u5980_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hded4))
    _al_u5981 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [2]),
    .b(_al_u5980_o),
    .c(_al_u1581_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wc5ju6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Am5ju6_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u5982 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P8oiu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F26bx6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vgjpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rk5ju6 ));
  AL_MAP_LUT4 #(
    .EQN("(~D*~A*~(C*B))"),
    .INIT(16'h0015))
    _al_u5983 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rk5ju6 ),
    .b(_al_u5848_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_control_o ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_2 ),
    .o(_al_u5983_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u5984 (
    .a(_al_u5983_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pk4ju6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[2] ),
    .o(_al_u5984_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u5985 (
    .a(_al_u5984_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/By4ju6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [3]),
    .o(_al_u5985_o));
  AL_MAP_LUT4 #(
    .EQN("(C*A*~(D*~B))"),
    .INIT(16'h80a0))
    _al_u5986 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Am5ju6_lutinv ),
    .b(_al_u1916_o),
    .c(_al_u5985_o),
    .d(_al_u5854_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cgkiu6 ));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u5987 (
    .a(_al_u5956_o),
    .b(_al_u5979_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cgkiu6 ),
    .o(_al_u5987_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*~A))"),
    .INIT(16'h23af))
    _al_u5988 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N30iu6 ),
    .b(_al_u607_o),
    .c(_al_u932_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sqkax6 ),
    .o(_al_u5988_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*~A))"),
    .INIT(16'h23af))
    _al_u5989 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O00iu6 ),
    .b(_al_u607_o),
    .c(_al_u932_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R9mpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y1qow6 ));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*B)*~(C*A))"),
    .INIT(16'heca0))
    _al_u599 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n100 ),
    .b(_al_u364_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n88_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n102 [0]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_rx_state [0]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u5990 (
    .a(_al_u5988_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y1qow6 ),
    .o(_al_u5990_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*~A))"),
    .INIT(16'h23af))
    _al_u5991 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pxzhu6 ),
    .b(_al_u607_o),
    .c(_al_u932_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rskax6 ),
    .o(_al_u5991_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u5992 (
    .a(_al_u5990_o),
    .b(_al_u5991_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kupow6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*~A))"),
    .INIT(16'h23af))
    _al_u5993 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uwzhu6 ),
    .b(_al_u607_o),
    .c(_al_u932_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U1kpw6 ),
    .o(_al_u5993_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u5994 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kupow6_lutinv ),
    .b(_al_u5993_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J43ju6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*~A))"),
    .INIT(16'h23af))
    _al_u5995 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nwzhu6 ),
    .b(_al_u607_o),
    .c(_al_u932_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ubypw6 ),
    .o(_al_u5995_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u5996 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J43ju6_lutinv ),
    .b(_al_u5995_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N7pow6 ));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*~B))"),
    .INIT(8'h54))
    _al_u5997 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N7pow6 ),
    .b(_al_u604_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V2kow6_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(B@(C*~A))"),
    .INIT(8'h9c))
    _al_u5998 (
    .a(_al_u5990_o),
    .b(_al_u5991_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ),
    .o(_al_u5998_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A))"),
    .INIT(16'hb100))
    _al_u5999 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V2kow6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kupow6_lutinv ),
    .c(_al_u5998_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Queow6 ));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u600 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_apb_slave_mux/n4 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/state_reg [0]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PWRITE ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/write_enable ));
  AL_MAP_LUT4 #(
    .EQN("(A*~(C@(D*~B)))"),
    .INIT(16'h280a))
    _al_u6000 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V2kow6_lutinv ),
    .b(_al_u5988_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y1qow6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ),
    .o(_al_u6000_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u6001 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Queow6 ),
    .b(_al_u6000_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lolow6 ));
  AL_MAP_LUT3 #(
    .EQN("(~A*(C@B))"),
    .INIT(8'h14))
    _al_u6002 (
    .a(_al_u5988_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y1qow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ),
    .o(_al_u6002_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D*C*~B))"),
    .INIT(16'h8aaa))
    _al_u6003 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lolow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V2kow6_lutinv ),
    .c(_al_u5998_o),
    .d(_al_u6002_o),
    .o(_al_u6003_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'h3050))
    _al_u6004 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dc0iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y50iu6 ),
    .c(_al_u5988_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y1qow6 ),
    .o(_al_u6004_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u6005 (
    .a(_al_u6002_o),
    .b(_al_u6004_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R50iu6 ),
    .o(_al_u6005_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C@B))"),
    .INIT(8'h41))
    _al_u6006 (
    .a(_al_u5988_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y1qow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ),
    .o(_al_u6006_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*B))"),
    .INIT(8'ha2))
    _al_u6007 (
    .a(_al_u6005_o),
    .b(_al_u6006_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E90iu6 ),
    .o(_al_u6007_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'h3050))
    _al_u6008 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D50iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F60iu6 ),
    .c(_al_u5988_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y1qow6 ),
    .o(_al_u6008_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u6009 (
    .a(_al_u6002_o),
    .b(_al_u6008_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K50iu6 ),
    .o(_al_u6009_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u601 (
    .a(_al_u473_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/write_enable ),
    .c(_al_u467_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/write_enable00 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*B))"),
    .INIT(8'ha2))
    _al_u6010 (
    .a(_al_u6009_o),
    .b(_al_u6006_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W40iu6 ),
    .o(_al_u6010_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D))"),
    .INIT(16'h1105))
    _al_u6011 (
    .a(_al_u6003_o),
    .b(_al_u6007_o),
    .c(_al_u6010_o),
    .d(_al_u5998_o),
    .o(_al_u6011_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*B))"),
    .INIT(8'ha2))
    _al_u6012 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Queow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V2kow6_lutinv ),
    .c(_al_u5990_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V5oow6 ));
  AL_MAP_LUT4 #(
    .EQN("(C*~(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'h3050))
    _al_u6013 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E90iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R50iu6 ),
    .c(_al_u5988_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y1qow6 ),
    .o(_al_u6013_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u6014 (
    .a(_al_u6002_o),
    .b(_al_u6013_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dc0iu6 ),
    .o(_al_u6014_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*B))"),
    .INIT(8'ha2))
    _al_u6015 (
    .a(_al_u6014_o),
    .b(_al_u6006_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F60iu6 ),
    .o(_al_u6015_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'h5030))
    _al_u6016 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K50iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W40iu6 ),
    .c(_al_u5988_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y1qow6 ),
    .o(_al_u6016_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u6017 (
    .a(_al_u6002_o),
    .b(_al_u6016_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D50iu6 ),
    .o(_al_u6017_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*B))"),
    .INIT(8'ha2))
    _al_u6018 (
    .a(_al_u6017_o),
    .b(_al_u6006_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P40iu6 ),
    .o(_al_u6018_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'h53))
    _al_u6019 (
    .a(_al_u6015_o),
    .b(_al_u6018_o),
    .c(_al_u5998_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qb3ju6_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u602 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n7_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/write_enable ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/write_enable10 ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(C*A))"),
    .INIT(16'h4c5f))
    _al_u6020 (
    .a(_al_u1813_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xqpow6_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    _al_u6021 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R50iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xqpow6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fpnpw6 ),
    .o(_al_u6021_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u6022 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V5oow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qb3ju6_lutinv ),
    .c(_al_u6021_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mg3ju6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'h5030))
    _al_u6023 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dc0iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F60iu6 ),
    .c(_al_u5988_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y1qow6 ),
    .o(_al_u6023_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u6024 (
    .a(_al_u6006_o),
    .b(_al_u6023_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K50iu6 ),
    .o(_al_u6024_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*B))"),
    .INIT(8'ha2))
    _al_u6025 (
    .a(_al_u6024_o),
    .b(_al_u6002_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E90iu6 ),
    .o(_al_u6025_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h58fc))
    _al_u6026 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V2kow6_lutinv ),
    .b(_al_u6025_o),
    .c(_al_u5998_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 ),
    .o(_al_u6026_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~(B@A))"),
    .INIT(16'h0900))
    _al_u6027 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V2kow6_lutinv ),
    .b(_al_u5998_o),
    .c(_al_u6021_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 ),
    .o(_al_u6027_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'h5030))
    _al_u6028 (
    .a(_al_u823_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y50iu6 ),
    .c(_al_u5988_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y1qow6 ),
    .o(_al_u6028_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u6029 (
    .a(_al_u6006_o),
    .b(_al_u6028_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R50iu6 ),
    .o(_al_u6029_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u603 (
    .a(_al_u473_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/write_enable ),
    .c(_al_u571_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/write_enable08 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*B))"),
    .INIT(8'ha2))
    _al_u6030 (
    .a(_al_u6029_o),
    .b(_al_u6002_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M60iu6 ),
    .o(_al_u6030_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(A*~(D*~C)))"),
    .INIT(16'h1311))
    _al_u6031 (
    .a(_al_u6026_o),
    .b(_al_u6027_o),
    .c(_al_u6030_o),
    .d(_al_u5998_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xa4ju6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'h5030))
    _al_u6032 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V70iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H70iu6 ),
    .c(_al_u5988_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y1qow6 ),
    .o(_al_u6032_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u6033 (
    .a(_al_u6006_o),
    .b(_al_u6032_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A70iu6 ),
    .o(_al_u6033_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*B))"),
    .INIT(8'ha2))
    _al_u6034 (
    .a(_al_u6033_o),
    .b(_al_u6002_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O70iu6 ),
    .o(_al_u6034_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u6035 (
    .a(_al_u6030_o),
    .b(_al_u6034_o),
    .c(_al_u5998_o),
    .o(_al_u6035_o));
  AL_MAP_LUT4 #(
    .EQN("~(B*~(C)*~((D*A))+B*C*~((D*A))+~(B)*C*(D*A)+B*C*(D*A))"),
    .INIT(16'h1b33))
    _al_u6036 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V2kow6_lutinv ),
    .b(_al_u6035_o),
    .c(_al_u6021_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 ),
    .o(_al_u6036_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*B*~A)"),
    .INIT(16'h0400))
    _al_u6037 (
    .a(_al_u6011_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mg3ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xa4ju6_lutinv ),
    .d(_al_u6036_o),
    .o(_al_u6037_o));
  AL_MAP_LUT3 #(
    .EQN("(B@(C*~A))"),
    .INIT(8'h9c))
    _al_u6038 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J43ju6_lutinv ),
    .b(_al_u5995_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M93ju6_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(B@(C*~A))"),
    .INIT(8'h9c))
    _al_u6039 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kupow6_lutinv ),
    .b(_al_u5993_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ),
    .o(_al_u6039_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u604 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ),
    .o(_al_u604_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u6040 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M93ju6_lutinv ),
    .b(_al_u6039_o),
    .o(_al_u6040_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B*A))"),
    .INIT(8'h70))
    _al_u6041 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zvzhu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Svzhu6 ),
    .c(_al_u932_o),
    .o(_al_u6041_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u6042 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R9mpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rskax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sqkax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ubypw6 ),
    .o(_al_u6042_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    _al_u6043 (
    .a(_al_u607_o),
    .b(_al_u6042_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U1kpw6 ),
    .o(_al_u6043_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~A*~(D*~B))"),
    .INIT(16'h0405))
    _al_u6044 (
    .a(_al_u6041_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gwzhu6 ),
    .c(_al_u6043_o),
    .d(_al_u932_o),
    .o(_al_u6044_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u6045 (
    .a(_al_u6044_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 ),
    .o(_al_u6045_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u6046 (
    .a(_al_u6040_o),
    .b(_al_u6045_o),
    .o(_al_u6046_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*~B))"),
    .INIT(8'ha8))
    _al_u6047 (
    .a(_al_u6046_o),
    .b(_al_u604_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ),
    .o(_al_u6047_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u6048 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M93ju6_lutinv ),
    .b(_al_u6039_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R83ju6_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u6049 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R83ju6_lutinv ),
    .b(_al_u6045_o),
    .o(_al_u6049_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u605 (
    .a(_al_u604_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bi0iu6 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*~B))"),
    .INIT(8'ha8))
    _al_u6050 (
    .a(_al_u6049_o),
    .b(_al_u604_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ),
    .o(_al_u6050_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u6051 (
    .a(_al_u6047_o),
    .b(_al_u6050_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oh3ju6 ));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'h5030))
    _al_u6052 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S90iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X80iu6 ),
    .c(_al_u5988_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y1qow6 ),
    .o(_al_u6052_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u6053 (
    .a(_al_u6006_o),
    .b(_al_u6052_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q80iu6 ),
    .o(_al_u6053_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*B))"),
    .INIT(8'ha2))
    _al_u6054 (
    .a(_al_u6053_o),
    .b(_al_u6002_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L90iu6 ),
    .o(_al_u6054_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'h5030))
    _al_u6055 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z90iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L90iu6 ),
    .c(_al_u5988_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y1qow6 ),
    .o(_al_u6055_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u6056 (
    .a(_al_u6002_o),
    .b(_al_u6055_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S90iu6 ),
    .o(_al_u6056_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*B))"),
    .INIT(8'ha2))
    _al_u6057 (
    .a(_al_u6056_o),
    .b(_al_u6006_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X80iu6 ),
    .o(_al_u6057_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u6058 (
    .a(_al_u6054_o),
    .b(_al_u6057_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q34ju6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'h5030))
    _al_u6059 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ga0iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S90iu6 ),
    .c(_al_u5988_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y1qow6 ),
    .o(_al_u6059_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u606 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 ),
    .o(_al_u606_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u6060 (
    .a(_al_u6002_o),
    .b(_al_u6059_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z90iu6 ),
    .o(_al_u6060_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*B))"),
    .INIT(8'ha2))
    _al_u6061 (
    .a(_al_u6060_o),
    .b(_al_u6006_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L90iu6 ),
    .o(_al_u6061_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'h5030))
    _al_u6062 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Na0iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z90iu6 ),
    .c(_al_u5988_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y1qow6 ),
    .o(_al_u6062_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u6063 (
    .a(_al_u6002_o),
    .b(_al_u6062_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ga0iu6 ),
    .o(_al_u6063_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*B))"),
    .INIT(8'ha2))
    _al_u6064 (
    .a(_al_u6063_o),
    .b(_al_u6006_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S90iu6 ),
    .o(_al_u6064_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*A)"),
    .INIT(16'h0080))
    _al_u6065 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q34ju6_lutinv ),
    .b(_al_u6061_o),
    .c(_al_u6064_o),
    .d(_al_u5998_o),
    .o(_al_u6065_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'h3050))
    _al_u6066 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ib0iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wb0iu6 ),
    .c(_al_u5988_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y1qow6 ),
    .o(_al_u6066_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u6067 (
    .a(_al_u6002_o),
    .b(_al_u6066_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pb0iu6 ),
    .o(_al_u6067_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*B))"),
    .INIT(8'ha2))
    _al_u6068 (
    .a(_al_u6067_o),
    .b(_al_u6006_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bb0iu6 ),
    .o(_al_u6068_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'h5030))
    _al_u6069 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U30iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pb0iu6 ),
    .c(_al_u5988_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y1qow6 ),
    .o(_al_u6069_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u607 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 ),
    .o(_al_u607_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u6070 (
    .a(_al_u6006_o),
    .b(_al_u6069_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ib0iu6 ),
    .o(_al_u6070_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*B))"),
    .INIT(8'ha2))
    _al_u6071 (
    .a(_al_u6070_o),
    .b(_al_u6002_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wb0iu6 ),
    .o(_al_u6071_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u6072 (
    .a(_al_u6068_o),
    .b(_al_u6071_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ov3ju6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(C*~(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'h3050))
    _al_u6073 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bb0iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pb0iu6 ),
    .c(_al_u5988_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y1qow6 ),
    .o(_al_u6073_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u6074 (
    .a(_al_u6006_o),
    .b(_al_u6073_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ua0iu6 ),
    .o(_al_u6074_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*B))"),
    .INIT(8'ha2))
    _al_u6075 (
    .a(_al_u6074_o),
    .b(_al_u6002_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ib0iu6 ),
    .o(_al_u6075_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u6076 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ov3ju6_lutinv ),
    .b(_al_u6075_o),
    .o(_al_u6076_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'h5030))
    _al_u6077 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ib0iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ua0iu6 ),
    .c(_al_u5988_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y1qow6 ),
    .o(_al_u6077_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u6078 (
    .a(_al_u6002_o),
    .b(_al_u6077_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bb0iu6 ),
    .o(_al_u6078_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*B))"),
    .INIT(8'ha2))
    _al_u6079 (
    .a(_al_u6078_o),
    .b(_al_u6006_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Na0iu6 ),
    .o(_al_u6079_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u608 (
    .a(_al_u606_o),
    .b(_al_u607_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L0niu6 ));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'h5030))
    _al_u6080 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B40iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wb0iu6 ),
    .c(_al_u5988_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y1qow6 ),
    .o(_al_u6080_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u6081 (
    .a(_al_u6006_o),
    .b(_al_u6080_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pb0iu6 ),
    .o(_al_u6081_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*B))"),
    .INIT(8'ha2))
    _al_u6082 (
    .a(_al_u6081_o),
    .b(_al_u6002_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U30iu6 ),
    .o(_al_u6082_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u6083 (
    .a(_al_u6079_o),
    .b(_al_u6082_o),
    .c(_al_u5998_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gk3ju6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'h5030))
    _al_u6084 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L90iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q80iu6 ),
    .c(_al_u5988_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y1qow6 ),
    .o(_al_u6084_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u6085 (
    .a(_al_u6002_o),
    .b(_al_u6084_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X80iu6 ),
    .o(_al_u6085_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*B))"),
    .INIT(8'ha2))
    _al_u6086 (
    .a(_al_u6085_o),
    .b(_al_u6006_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J80iu6 ),
    .o(_al_u6086_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'h53))
    _al_u6087 (
    .a(_al_u6064_o),
    .b(_al_u6086_o),
    .c(_al_u5998_o),
    .o(_al_u6087_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'h5030))
    _al_u6088 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ua0iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ga0iu6 ),
    .c(_al_u5988_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y1qow6 ),
    .o(_al_u6088_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u6089 (
    .a(_al_u6002_o),
    .b(_al_u6088_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Na0iu6 ),
    .o(_al_u6089_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u609 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 ),
    .o(_al_u609_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*B))"),
    .INIT(8'ha2))
    _al_u6090 (
    .a(_al_u6089_o),
    .b(_al_u6006_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z90iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Id4ju6 ));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'h5030))
    _al_u6091 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bb0iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Na0iu6 ),
    .c(_al_u5988_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y1qow6 ),
    .o(_al_u6091_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u6092 (
    .a(_al_u6006_o),
    .b(_al_u6091_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ga0iu6 ),
    .o(_al_u6092_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*B))"),
    .INIT(8'ha2))
    _al_u6093 (
    .a(_al_u6092_o),
    .b(_al_u6002_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ua0iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uc4ju6 ));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*~A)"),
    .INIT(16'h1000))
    _al_u6094 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gk3ju6_lutinv ),
    .b(_al_u6087_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Id4ju6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uc4ju6 ),
    .o(_al_u6094_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u6095 (
    .a(_al_u6079_o),
    .b(_al_u5998_o),
    .o(_al_u6095_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(~A*~(D*B)))"),
    .INIT(16'he0a0))
    _al_u6096 (
    .a(_al_u6065_o),
    .b(_al_u6076_o),
    .c(_al_u6094_o),
    .d(_al_u6095_o),
    .o(_al_u6096_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u6097 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M93ju6_lutinv ),
    .b(_al_u6045_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jfmow6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u6098 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N7pow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3how6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(A*~(~D*C)))"),
    .INIT(16'h1131))
    _al_u6099 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oh3ju6 ),
    .b(_al_u6096_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jfmow6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3how6_lutinv ),
    .o(_al_u6099_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~(~B*~A))"),
    .INIT(16'h0e00))
    _al_u610 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bi0iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L0niu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ),
    .d(_al_u609_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jzmiu6 ));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u6100 (
    .a(_al_u6040_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3how6_lutinv ),
    .c(_al_u6045_o),
    .o(_al_u6100_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'h5030))
    _al_u6101 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X80iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J80iu6 ),
    .c(_al_u5988_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y1qow6 ),
    .o(_al_u6101_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u6102 (
    .a(_al_u6006_o),
    .b(_al_u6101_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C80iu6 ),
    .o(_al_u6102_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*B))"),
    .INIT(8'ha2))
    _al_u6103 (
    .a(_al_u6102_o),
    .b(_al_u6002_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q80iu6 ),
    .o(_al_u6103_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'h53))
    _al_u6104 (
    .a(_al_u6061_o),
    .b(_al_u6103_o),
    .c(_al_u5998_o),
    .o(_al_u6104_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'h5030))
    _al_u6105 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A70iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M60iu6 ),
    .c(_al_u5988_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y1qow6 ),
    .o(_al_u6105_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u6106 (
    .a(_al_u6006_o),
    .b(_al_u6105_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y50iu6 ),
    .o(_al_u6106_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*B))"),
    .INIT(8'ha2))
    _al_u6107 (
    .a(_al_u6106_o),
    .b(_al_u6002_o),
    .c(_al_u823_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Csnow6 ));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'h5030))
    _al_u6108 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C80iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O70iu6 ),
    .c(_al_u5988_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y1qow6 ),
    .o(_al_u6108_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u6109 (
    .a(_al_u6002_o),
    .b(_al_u6108_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V70iu6 ),
    .o(_al_u6109_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u611 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D43qw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pe7ax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ilwiu6 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*B))"),
    .INIT(8'ha2))
    _al_u6110 (
    .a(_al_u6109_o),
    .b(_al_u6006_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H70iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C34ju6 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    _al_u6111 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Csnow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C34ju6 ),
    .c(_al_u5998_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ha3ju6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'h5030))
    _al_u6112 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J80iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V70iu6 ),
    .c(_al_u5988_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y1qow6 ),
    .o(_al_u6112_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u6113 (
    .a(_al_u6006_o),
    .b(_al_u6112_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O70iu6 ),
    .o(_al_u6113_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*B))"),
    .INIT(8'ha2))
    _al_u6114 (
    .a(_al_u6113_o),
    .b(_al_u6002_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C80iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R04ju6 ));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'h5030))
    _al_u6115 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q80iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C80iu6 ),
    .c(_al_u5988_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y1qow6 ),
    .o(_al_u6115_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u6116 (
    .a(_al_u6006_o),
    .b(_al_u6115_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V70iu6 ),
    .o(_al_u6116_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*B))"),
    .INIT(8'ha2))
    _al_u6117 (
    .a(_al_u6116_o),
    .b(_al_u6002_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J80iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F14ju6 ));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*~A)"),
    .INIT(16'h4000))
    _al_u6118 (
    .a(_al_u6104_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ha3ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R04ju6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F14ju6 ),
    .o(_al_u6118_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u6119 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q34ju6_lutinv ),
    .b(_al_u6086_o),
    .c(_al_u6103_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M14ju6 ));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u612 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ilwiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Di3qw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Le2qw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ymwiu6 ));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'h5030))
    _al_u6120 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H70iu6 ),
    .b(_al_u823_o),
    .c(_al_u5988_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y1qow6 ),
    .o(_al_u6120_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u6121 (
    .a(_al_u6002_o),
    .b(_al_u6120_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A70iu6 ),
    .o(_al_u6121_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*B))"),
    .INIT(8'ha2))
    _al_u6122 (
    .a(_al_u6121_o),
    .b(_al_u6006_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M60iu6 ),
    .o(_al_u6122_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'h5030))
    _al_u6123 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O70iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A70iu6 ),
    .c(_al_u5988_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y1qow6 ),
    .o(_al_u6123_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u6124 (
    .a(_al_u6006_o),
    .b(_al_u6123_o),
    .c(_al_u823_o),
    .o(_al_u6124_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*B))"),
    .INIT(8'ha2))
    _al_u6125 (
    .a(_al_u6124_o),
    .b(_al_u6002_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H70iu6 ),
    .o(_al_u6125_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u6126 (
    .a(_al_u6122_o),
    .b(_al_u6125_o),
    .c(_al_u6034_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C34ju6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T14ju6 ));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D))"),
    .INIT(16'h88a0))
    _al_u6127 (
    .a(_al_u6118_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M14ju6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T14ju6 ),
    .d(_al_u5998_o),
    .o(_al_u6127_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(~B*~A))"),
    .INIT(8'h0e))
    _al_u6128 (
    .a(_al_u6047_o),
    .b(_al_u6100_o),
    .c(_al_u6127_o),
    .o(_al_u6128_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u6129 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M93ju6_lutinv ),
    .b(_al_u6039_o),
    .c(_al_u6045_o),
    .o(_al_u6129_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    _al_u613 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hw8ax6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sqwpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zm8ax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fnwiu6 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*~B))"),
    .INIT(8'ha8))
    _al_u6130 (
    .a(_al_u6129_o),
    .b(_al_u604_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ),
    .o(_al_u6130_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u6131 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M93ju6_lutinv ),
    .b(_al_u6039_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rupow6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(~D*C*~B))"),
    .INIT(16'h5545))
    _al_u6132 (
    .a(_al_u6130_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3how6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rupow6_lutinv ),
    .d(_al_u6045_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gy3ju6 ));
  AL_MAP_LUT4 #(
    .EQN("(C*~(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'h3050))
    _al_u6133 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P40iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D50iu6 ),
    .c(_al_u5988_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y1qow6 ),
    .o(_al_u6133_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u6134 (
    .a(_al_u6006_o),
    .b(_al_u6133_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I40iu6 ),
    .o(_al_u6134_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*B))"),
    .INIT(8'ha2))
    _al_u6135 (
    .a(_al_u6134_o),
    .b(_al_u6002_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W40iu6 ),
    .o(_al_u6135_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'h53))
    _al_u6136 (
    .a(_al_u6025_o),
    .b(_al_u6135_o),
    .c(_al_u5998_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lj3ju6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(C*~(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'h3050))
    _al_u6137 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U30iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I40iu6 ),
    .c(_al_u5988_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y1qow6 ),
    .o(_al_u6137_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u6138 (
    .a(_al_u6006_o),
    .b(_al_u6137_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wb0iu6 ),
    .o(_al_u6138_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*B))"),
    .INIT(8'ha2))
    _al_u6139 (
    .a(_al_u6138_o),
    .b(_al_u6002_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B40iu6 ),
    .o(_al_u6139_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u614 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ymwiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fnwiu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fgpiu6 ));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u6140 (
    .a(_al_u6075_o),
    .b(_al_u6139_o),
    .c(_al_u5998_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jb3ju6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'h5030))
    _al_u6141 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P40iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B40iu6 ),
    .c(_al_u5988_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y1qow6 ),
    .o(_al_u6141_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u6142 (
    .a(_al_u6006_o),
    .b(_al_u6141_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U30iu6 ),
    .o(_al_u6142_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*B))"),
    .INIT(8'ha2))
    _al_u6143 (
    .a(_al_u6142_o),
    .b(_al_u6002_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I40iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yt3ju6 ));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'h5030))
    _al_u6144 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W40iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I40iu6 ),
    .c(_al_u5988_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y1qow6 ),
    .o(_al_u6144_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u6145 (
    .a(_al_u6002_o),
    .b(_al_u6144_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P40iu6 ),
    .o(_al_u6145_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*B))"),
    .INIT(8'ha2))
    _al_u6146 (
    .a(_al_u6145_o),
    .b(_al_u6006_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B40iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mu3ju6 ));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*~A)"),
    .INIT(16'h1000))
    _al_u6147 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lj3ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jb3ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yt3ju6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mu3ju6 ),
    .o(_al_u6147_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u6148 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ov3ju6_lutinv ),
    .b(_al_u6082_o),
    .c(_al_u6139_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Av3ju6 ));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'h5030))
    _al_u6149 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E90iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K50iu6 ),
    .c(_al_u5988_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y1qow6 ),
    .o(_al_u6149_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u615 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fgpiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dg2qw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Scbiu6 ));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u6150 (
    .a(_al_u6002_o),
    .b(_al_u6149_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F60iu6 ),
    .o(_al_u6150_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*B))"),
    .INIT(8'ha2))
    _al_u6151 (
    .a(_al_u6150_o),
    .b(_al_u6006_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D50iu6 ),
    .o(_al_u6151_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u6152 (
    .a(_al_u6151_o),
    .b(_al_u6018_o),
    .c(_al_u6010_o),
    .d(_al_u6135_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tu3ju6 ));
  AL_MAP_LUT4 #(
    .EQN("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'ha088))
    _al_u6153 (
    .a(_al_u6147_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Av3ju6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tu3ju6 ),
    .d(_al_u5998_o),
    .o(_al_u6153_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(~D*~(C*A)))"),
    .INIT(16'h3320))
    _al_u6154 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oh3ju6 ),
    .b(_al_u6128_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gy3ju6 ),
    .d(_al_u6153_o),
    .o(_al_u6154_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*B*~A)"),
    .INIT(16'h0400))
    _al_u6155 (
    .a(_al_u6099_o),
    .b(_al_u6154_o),
    .c(_al_u6021_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fpnpw6 ),
    .o(_al_u6155_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u6156 (
    .a(_al_u5988_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y1qow6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gweow6_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u6157 (
    .a(_al_u6002_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gweow6_lutinv ),
    .o(_al_u6157_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*~A)"),
    .INIT(8'h04))
    _al_u6158 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V2kow6_lutinv ),
    .b(_al_u5998_o),
    .c(_al_u6157_o),
    .o(_al_u6158_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*A*~(~D*C))"),
    .INIT(16'h2202))
    _al_u6159 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Queow6 ),
    .b(_al_u6158_o),
    .c(_al_u6000_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gweow6_lutinv ),
    .o(_al_u6159_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B*A))"),
    .INIT(8'h70))
    _al_u616 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Scbiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H34iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hmbax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n853 ));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'h5030))
    _al_u6160 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M60iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R50iu6 ),
    .c(_al_u5988_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y1qow6 ),
    .o(_al_u6160_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u6161 (
    .a(_al_u6002_o),
    .b(_al_u6160_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y50iu6 ),
    .o(_al_u6161_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*B))"),
    .INIT(8'ha2))
    _al_u6162 (
    .a(_al_u6161_o),
    .b(_al_u6006_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dc0iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nweow6 ));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D))"),
    .INIT(16'h1105))
    _al_u6163 (
    .a(_al_u6159_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nweow6 ),
    .c(_al_u6151_o),
    .d(_al_u5998_o),
    .o(_al_u6163_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u6164 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V2kow6_lutinv ),
    .b(_al_u5998_o),
    .c(_al_u5990_o),
    .o(_al_u6164_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(~A*~(~C*~B)))"),
    .INIT(16'hab00))
    _al_u6165 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V2kow6_lutinv ),
    .b(_al_u5998_o),
    .c(_al_u5990_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jbjow6 ));
  AL_MAP_LUT4 #(
    .EQN("(B*(~A*~(C)*~(D)+~A*C*~(D)+~(~A)*C*D+~A*C*D))"),
    .INIT(16'hc044))
    _al_u6166 (
    .a(_al_u6164_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jbjow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V2kow6_lutinv ),
    .d(_al_u6002_o),
    .o(_al_u6166_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D))"),
    .INIT(16'h1105))
    _al_u6167 (
    .a(_al_u6166_o),
    .b(_al_u6122_o),
    .c(_al_u6007_o),
    .d(_al_u5998_o),
    .o(_al_u6167_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u6168 (
    .a(_al_u6164_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jbjow6 ),
    .o(_al_u6168_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D))"),
    .INIT(16'h1105))
    _al_u6169 (
    .a(_al_u6168_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Csnow6 ),
    .c(_al_u6015_o),
    .d(_al_u5998_o),
    .o(_al_u6169_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u617 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n3685 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X5phu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Daiax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ajohu6 ));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))"),
    .INIT(16'h44c0))
    _al_u6170 (
    .a(_al_u6164_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jbjow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V2kow6_lutinv ),
    .d(_al_u6157_o),
    .o(_al_u6170_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'h0511))
    _al_u6171 (
    .a(_al_u6170_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nweow6 ),
    .c(_al_u6125_o),
    .d(_al_u5998_o),
    .o(_al_u6171_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u6172 (
    .a(_al_u6163_o),
    .b(_al_u6167_o),
    .c(_al_u6169_o),
    .d(_al_u6171_o),
    .o(_al_u6172_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~D*~(C*A)))"),
    .INIT(16'hcc80))
    _al_u6173 (
    .a(_al_u6037_o),
    .b(_al_u6155_o),
    .c(_al_u6172_o),
    .d(_al_u6045_o),
    .o(_al_u6173_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'h084c))
    _al_u6174 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L2epw6 ),
    .b(_al_u1421_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wc5ju6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cg5ju6_lutinv ),
    .o(_al_u6174_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~B*~(C*A))"),
    .INIT(16'h0013))
    _al_u6175 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/By4ju6 ),
    .b(_al_u5848_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [16]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_15 ),
    .o(_al_u6175_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*~A))"),
    .INIT(8'h8c))
    _al_u6176 (
    .a(_al_u2150_o),
    .b(_al_u6175_o),
    .c(_al_u5854_o),
    .o(_al_u6176_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(D*~C*A))"),
    .INIT(16'hc4cc))
    _al_u6177 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L2epw6 ),
    .b(_al_u6176_o),
    .c(_al_u1421_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ys4ju6 ),
    .o(_al_u6177_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u6178 (
    .a(_al_u6174_o),
    .b(_al_u6177_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ngmiu6 ));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .INIT(16'h082a))
    _al_u6179 (
    .a(_al_u1624_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [10]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wc5ju6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cg5ju6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I98ju6_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    _al_u618 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reload_i ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/baud_updated ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n44 ));
  AL_MAP_LUT4 #(
    .EQN("(~D*~B*~(C*A))"),
    .INIT(16'h0013))
    _al_u6180 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/By4ju6 ),
    .b(_al_u5848_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [11]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_10 ),
    .o(_al_u6180_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*~A))"),
    .INIT(8'h8c))
    _al_u6181 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ka8ju6 ),
    .b(_al_u6180_o),
    .c(_al_u5854_o),
    .o(_al_u6181_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D*B*~A))"),
    .INIT(16'hb0f0))
    _al_u6182 (
    .a(_al_u1624_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [10]),
    .c(_al_u6181_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ys4ju6 ),
    .o(_al_u6182_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u6183 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I98ju6_lutinv ),
    .b(_al_u6182_o),
    .o(_al_u6183_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .INIT(16'h082a))
    _al_u6184 (
    .a(_al_u1632_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C1epw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wc5ju6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cg5ju6_lutinv ),
    .o(_al_u6184_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~B*~(C*A))"),
    .INIT(16'h0013))
    _al_u6185 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/By4ju6 ),
    .b(_al_u5848_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [12]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_11 ),
    .o(_al_u6185_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*~A))"),
    .INIT(8'h8c))
    _al_u6186 (
    .a(_al_u2062_o),
    .b(_al_u6185_o),
    .c(_al_u5854_o),
    .o(_al_u6186_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D*B*~A))"),
    .INIT(16'hb0f0))
    _al_u6187 (
    .a(_al_u1632_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C1epw6 ),
    .c(_al_u6186_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ys4ju6 ),
    .o(_al_u6187_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u6188 (
    .a(_al_u6184_o),
    .b(_al_u6187_o),
    .o(_al_u6188_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .INIT(16'h082a))
    _al_u6189 (
    .a(_al_u1413_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X1epw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wc5ju6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cg5ju6_lutinv ),
    .o(_al_u6189_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u619 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n44 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [13]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n37 [9]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_baud_cntr_i [9]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~B*~(C*A))"),
    .INIT(16'h0013))
    _al_u6190 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/By4ju6 ),
    .b(_al_u5848_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [15]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_14 ),
    .o(_al_u6190_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*~A))"),
    .INIT(8'h8c))
    _al_u6191 (
    .a(_al_u2128_o),
    .b(_al_u6190_o),
    .c(_al_u5854_o),
    .o(_al_u6191_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D*B*~A))"),
    .INIT(16'hb0f0))
    _al_u6192 (
    .a(_al_u1413_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X1epw6 ),
    .c(_al_u6191_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ys4ju6 ),
    .o(_al_u6192_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u6193 (
    .a(_al_u6189_o),
    .b(_al_u6192_o),
    .o(_al_u6193_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u6194 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ngmiu6 ),
    .b(_al_u6183_o),
    .c(_al_u6188_o),
    .d(_al_u6193_o),
    .o(_al_u6194_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'h084c))
    _al_u6195 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [23]),
    .b(_al_u1485_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wc5ju6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cg5ju6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Of5ju6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(~C*~B*~(D*A))"),
    .INIT(16'h0103))
    _al_u6196 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/By4ju6 ),
    .b(_al_u5848_o),
    .c(n1[5]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [24]),
    .o(_al_u6196_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*~A))"),
    .INIT(8'h8c))
    _al_u6197 (
    .a(_al_u2252_o),
    .b(_al_u6196_o),
    .c(_al_u5854_o),
    .o(_al_u6197_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(D*~C*A))"),
    .INIT(16'hc4cc))
    _al_u6198 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [23]),
    .b(_al_u6197_o),
    .c(_al_u1485_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ys4ju6 ),
    .o(_al_u6198_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u6199 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Of5ju6_lutinv ),
    .b(_al_u6198_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Evkiu6 ));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u620 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n44 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [12]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n37 [8]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_baud_cntr_i [8]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'h084c))
    _al_u6200 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G3epw6 ),
    .b(_al_u1437_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wc5ju6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cg5ju6_lutinv ),
    .o(_al_u6200_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~B*~(C*A))"),
    .INIT(16'h0013))
    _al_u6201 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/By4ju6 ),
    .b(_al_u5848_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [18]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_17 ),
    .o(_al_u6201_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*~A))"),
    .INIT(8'h8c))
    _al_u6202 (
    .a(_al_u2171_o),
    .b(_al_u6201_o),
    .c(_al_u5854_o),
    .o(_al_u6202_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(D*~C*A))"),
    .INIT(16'hc4cc))
    _al_u6203 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G3epw6 ),
    .b(_al_u6202_o),
    .c(_al_u1437_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ys4ju6 ),
    .o(_al_u6203_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u6204 (
    .a(_al_u6200_o),
    .b(_al_u6203_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wamiu6 ));
  AL_MAP_LUT4 #(
    .EQN("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'h084c))
    _al_u6205 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P4epw6 ),
    .b(_al_u1477_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wc5ju6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cg5ju6_lutinv ),
    .o(_al_u6205_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~B*~(D*A))"),
    .INIT(16'h0103))
    _al_u6206 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/By4ju6 ),
    .b(_al_u5848_o),
    .c(n1[4]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [23]),
    .o(_al_u6206_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*~A))"),
    .INIT(8'h8c))
    _al_u6207 (
    .a(_al_u2244_o),
    .b(_al_u6206_o),
    .c(_al_u5854_o),
    .o(_al_u6207_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(D*~C*A))"),
    .INIT(16'hc4cc))
    _al_u6208 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P4epw6 ),
    .b(_al_u6207_o),
    .c(_al_u1477_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ys4ju6 ),
    .o(_al_u6208_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u6209 (
    .a(_al_u6205_o),
    .b(_al_u6208_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uvliu6 ));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u621 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n44 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [11]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n37 [7]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_baud_cntr_i [7]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u6210 (
    .a(_al_u6194_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Evkiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wamiu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uvliu6 ),
    .o(_al_u6210_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(B*A))"),
    .INIT(8'h07))
    _al_u6211 (
    .a(_al_u1573_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mt4ju6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ys4ju6 ),
    .o(_al_u6211_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hed4d))
    _al_u6212 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [4]),
    .b(_al_u6211_o),
    .c(_al_u1573_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wc5ju6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kl4ju6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(~D*~B*~(C*A))"),
    .INIT(16'h0013))
    _al_u6213 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pk4ju6 ),
    .b(_al_u5848_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[4] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_4 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uj4ju6 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u6214 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uj4ju6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/By4ju6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [5]),
    .o(_al_u6214_o));
  AL_MAP_LUT4 #(
    .EQN("(C*A*~(D*~B))"),
    .INIT(16'h80a0))
    _al_u6215 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kl4ju6_lutinv ),
    .b(_al_u1934_o),
    .c(_al_u6214_o),
    .d(_al_u5854_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kkkiu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D*C*A))"),
    .INIT(16'h1333))
    _al_u6216 (
    .a(_al_u5987_o),
    .b(_al_u6173_o),
    .c(_al_u6210_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kkkiu6 ),
    .o(_al_u6216_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    _al_u6217 (
    .a(_al_u6216_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fhoiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_apsr_o[2] ),
    .o(_al_u6217_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*(~(A)*~(C)*~(D)+A*C*~(D)+A*C*D))"),
    .INIT(16'h2021))
    _al_u6218 (
    .a(_al_u6217_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rwjax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6 ),
    .o(_al_u6218_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u6219 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jfmow6 ),
    .b(_al_u6039_o),
    .o(_al_u6219_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u622 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n44 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [10]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n37 [6]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_baud_cntr_i [6]));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*A)"),
    .INIT(16'h0200))
    _al_u6220 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oh3ju6 ),
    .b(_al_u6130_o),
    .c(_al_u6219_o),
    .d(_al_u6021_o),
    .o(_al_u6220_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(~D*A))"),
    .INIT(16'h3f15))
    _al_u6221 (
    .a(_al_u6047_o),
    .b(_al_u6050_o),
    .c(_al_u6087_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ha3ju6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nd3ju6 ));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(D*C))"),
    .INIT(16'h0444))
    _al_u6222 (
    .a(_al_u6220_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nd3ju6 ),
    .c(_al_u6130_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jb3ju6_lutinv ),
    .o(_al_u6222_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*~B))"),
    .INIT(8'h8a))
    _al_u6223 (
    .a(_al_u6222_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mg3ju6_lutinv ),
    .c(_al_u6219_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ru2ju6 ));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u6224 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N7pow6 ),
    .b(_al_u6044_o),
    .c(_al_u6041_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P73ju6 ));
  AL_MAP_LUT4 #(
    .EQN("(D*~B*~(~C*A))"),
    .INIT(16'h3100))
    _al_u6225 (
    .a(_al_u6040_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P73ju6 ),
    .c(_al_u6035_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ),
    .o(_al_u6225_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hfadd))
    _al_u6226 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M93ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gk3ju6_lutinv ),
    .c(_al_u6104_o),
    .d(_al_u6039_o),
    .o(_al_u6226_o));
  AL_MAP_LUT4 #(
    .EQN("(C*A*~(~D*B))"),
    .INIT(16'ha020))
    _al_u6227 (
    .a(_al_u6225_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rupow6_lutinv ),
    .c(_al_u6226_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lj3ju6_lutinv ),
    .o(_al_u6227_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u6228 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N7pow6 ),
    .b(_al_u6044_o),
    .o(_al_u6228_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~B*~(C*~A))"),
    .INIT(16'h0023))
    _al_u6229 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ru2ju6 ),
    .b(_al_u6227_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P73ju6 ),
    .d(_al_u6228_o),
    .o(_al_u6229_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u623 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n44 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [9]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n37 [5]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_baud_cntr_i [5]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h770c))
    _al_u6230 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qb3ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M93ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jb3ju6_lutinv ),
    .d(_al_u6039_o),
    .o(_al_u6230_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u6231 (
    .a(_al_u6230_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M93ju6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ha3ju6_lutinv ),
    .o(_al_u6231_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u6232 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P73ju6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 ),
    .o(_al_u6232_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~A*~(D*C)))"),
    .INIT(16'hc888))
    _al_u6233 (
    .a(_al_u6231_o),
    .b(_al_u6232_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R83ju6_lutinv ),
    .d(_al_u6087_o),
    .o(_al_u6233_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u6234 (
    .a(_al_u6229_o),
    .b(_al_u6233_o),
    .o(_al_u6234_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u6235 (
    .a(_al_u6228_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_apsr_o[1] ),
    .o(_al_u6235_o));
  AL_MAP_LUT4 #(
    .EQN("~(D*~((~B*~A))*~(C)+D*(~B*~A)*~(C)+~(D)*(~B*~A)*C+D*(~B*~A)*C)"),
    .INIT(16'he0ef))
    _al_u6236 (
    .a(_al_u6234_o),
    .b(_al_u6235_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fpnpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [33]),
    .o(_al_u6236_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*(B@A))"),
    .INIT(8'h06))
    _al_u6237 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rwjax6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6 ),
    .o(_al_u6237_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(~A*~(D)*~(B)+~A*D*~(B)+~(~A)*D*B+~A*D*B))"),
    .INIT(16'h20e0))
    _al_u6238 (
    .a(_al_u6236_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ng8iu6 ),
    .c(_al_u6237_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_apsr_o[1] ),
    .o(_al_u6238_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u6239 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ru2ju6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bbliu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fpnpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vioiu6_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u624 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n44 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [8]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n37 [4]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_baud_cntr_i [4]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    _al_u6240 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rwjax6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6 ),
    .o(_al_u6240_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(~A*~(D)*~(B)+~A*D*~(B)+~(~A)*D*B+~A*D*B))"),
    .INIT(16'h020e))
    _al_u6241 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vioiu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fhoiu6 ),
    .c(_al_u6240_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_apsr_o[3] ),
    .o(_al_u6241_o));
  AL_MAP_LUT3 #(
    .EQN("(~(A)*~(B)*~(C)+A*~(B)*~(C)+~(A)*B*~(C)+A*~(B)*C+~(A)*B*C+A*B*C)"),
    .INIT(8'he7))
    _al_u6242 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [31]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D5epw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [32]),
    .o(_al_u6242_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u6243 (
    .a(_al_u1662_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 ),
    .o(_al_u6243_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u6244 (
    .a(_al_u6243_o),
    .b(_al_u932_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 ),
    .o(_al_u6244_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*A*~(D*C))"),
    .INIT(16'h0222))
    _al_u6245 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Im2ju6 ),
    .b(_al_u6244_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ldoiu6_lutinv ),
    .d(_al_u1660_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P9niu6 ));
  AL_MAP_LUT3 #(
    .EQN("(A*B*~(C)+A*~(B)*C+~(A)*B*C+A*B*C)"),
    .INIT(8'he8))
    _al_u6246 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rwjax6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6 ),
    .o(_al_u6246_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(~A*~(D)*~(B)+~A*D*~(B)+~(~A)*D*B+~A*D*B))"),
    .INIT(16'h20e0))
    _al_u6247 (
    .a(_al_u6242_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P9niu6 ),
    .c(_al_u6246_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_apsr_o[0] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qj2ju6 ));
  AL_MAP_LUT4 #(
    .EQN("(~B*~A*~(D@C))"),
    .INIT(16'h1001))
    _al_u6248 (
    .a(_al_u6218_o),
    .b(_al_u6238_o),
    .c(_al_u6241_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qj2ju6 ),
    .o(_al_u6248_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*A))"),
    .INIT(8'hc4))
    _al_u6249 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yo1ju6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rwjax6 ),
    .o(_al_u6249_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u625 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n44 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [7]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n37 [3]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_baud_cntr_i [3]));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(B*A)))"),
    .INIT(16'h080f))
    _al_u6250 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cwiiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rwjax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ai2ju6_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u6251 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Htyiu6 ),
    .b(_al_u2771_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ai2ju6_lutinv ),
    .o(_al_u6251_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~B*~(~C*A))"),
    .INIT(16'h0031))
    _al_u6252 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yo1ju6 ),
    .b(_al_u6251_o),
    .c(_al_u2380_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 ),
    .o(_al_u6252_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*A)"),
    .INIT(16'h0002))
    _al_u6253 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mldpw6 ),
    .b(_al_u1812_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F6ziu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vygax6 ),
    .o(_al_u6253_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'he4fc))
    _al_u6254 (
    .a(_al_u6248_o),
    .b(_al_u6249_o),
    .c(_al_u6252_o),
    .d(_al_u6253_o),
    .o(_al_u6254_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u6255 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U98iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N98iu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ),
    .o(_al_u6255_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~A*~(~D*C))"),
    .INIT(16'h1101))
    _al_u6256 (
    .a(_al_u3208_o),
    .b(_al_u6255_o),
    .c(_al_u1782_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ),
    .o(_al_u6256_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D*C*~B))"),
    .INIT(16'h8aaa))
    _al_u6257 (
    .a(_al_u6256_o),
    .b(_al_u1643_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U98iu6 ),
    .d(_al_u1907_o),
    .o(_al_u6257_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(~D*~C*B))"),
    .INIT(16'haaa2))
    _al_u6258 (
    .a(_al_u3233_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jckax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N4kax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4jax6 ),
    .o(_al_u6258_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+A*~(B)*C*D)"),
    .INIT(16'h23e3))
    _al_u6259 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nsaiu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 ),
    .o(_al_u6259_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u626 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n44 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [6]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n37 [2]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_baud_cntr_i [2]));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D*~C*~B))"),
    .INIT(16'ha8aa))
    _al_u6260 (
    .a(_al_u3191_o),
    .b(_al_u6259_o),
    .c(_al_u606_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ),
    .o(_al_u6260_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~B*~(~D*A))"),
    .INIT(16'h0301))
    _al_u6261 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yo1ju6 ),
    .b(_al_u6258_o),
    .c(_al_u6260_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6 ),
    .o(_al_u6261_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(~D*A))"),
    .INIT(16'h3f15))
    _al_u6262 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I82ju6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ls1ju6 ),
    .c(_al_u609_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ),
    .o(_al_u6262_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*~C))"),
    .INIT(16'h8088))
    _al_u6263 (
    .a(_al_u6257_o),
    .b(_al_u6261_o),
    .c(_al_u6262_o),
    .d(_al_u3109_o),
    .o(_al_u6263_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(D*~C*A))"),
    .INIT(16'hc4cc))
    _al_u6264 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eoyiu6_lutinv ),
    .b(_al_u682_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ),
    .o(_al_u6264_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u6265 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xc2ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vygax6 ),
    .o(_al_u6265_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h5507))
    _al_u6266 (
    .a(_al_u3109_o),
    .b(_al_u6265_o),
    .c(_al_u2829_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ),
    .o(_al_u6266_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*B*~(~D*~A))"),
    .INIT(16'h0c08))
    _al_u6267 (
    .a(_al_u1385_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/SLEEPHOLDACKn ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z9opw6 ),
    .o(_al_u6267_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~(~B*~A))"),
    .INIT(16'h000e))
    _al_u6268 (
    .a(_al_u6264_o),
    .b(_al_u6266_o),
    .c(_al_u6267_o),
    .d(_al_u1907_o),
    .o(_al_u6268_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*~C))"),
    .INIT(16'h8088))
    _al_u6269 (
    .a(_al_u6254_o),
    .b(_al_u6263_o),
    .c(_al_u6268_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qe8iu6_lutinv ),
    .o(_al_u6269_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u627 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n44 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [19]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n37 [15]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_baud_cntr_i [15]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hfd05))
    _al_u6270 (
    .a(_al_u6269_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yv1ju6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Buohu6 ));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*~A)"),
    .INIT(16'h0100))
    _al_u6271 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dt4iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tu4iu6 ),
    .c(_al_u933_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/DBGRESTARTED ),
    .o(_al_u6271_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u6272 (
    .a(_al_u6271_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kt4iu6 ));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u6273 (
    .a(\u_cmsdk_mcu/HADDR [10]),
    .b(\u_cmsdk_mcu/HADDR [8]),
    .c(\u_cmsdk_mcu/HADDR [7]),
    .o(_al_u6273_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*B))"),
    .INIT(8'ha2))
    _al_u6274 (
    .a(_al_u6273_o),
    .b(\u_cmsdk_mcu/HADDR [3]),
    .c(\u_cmsdk_mcu/HADDR [2]),
    .o(_al_u6274_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(~B*~(~D*~C)))"),
    .INIT(16'h4445))
    _al_u6275 (
    .a(\u_cmsdk_mcu/HADDR [9]),
    .b(\u_cmsdk_mcu/HADDR [7]),
    .c(\u_cmsdk_mcu/HADDR [4]),
    .d(\u_cmsdk_mcu/HADDR [3]),
    .o(_al_u6275_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(~D*~(~C*B)))"),
    .INIT(16'h5504))
    _al_u6276 (
    .a(_al_u6274_o),
    .b(_al_u6275_o),
    .c(\u_cmsdk_mcu/HADDR [8]),
    .d(\u_cmsdk_mcu/HADDR [11]),
    .o(_al_u6276_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u6277 (
    .a(\u_cmsdk_mcu/HADDR [9]),
    .b(\u_cmsdk_mcu/HADDR [8]),
    .c(\u_cmsdk_mcu/HADDR [11]),
    .o(_al_u6277_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u6278 (
    .a(\u_cmsdk_mcu/HADDR [10]),
    .b(\u_cmsdk_mcu/HADDR [4]),
    .c(\u_cmsdk_mcu/HADDR [3]),
    .d(\u_cmsdk_mcu/HADDR [2]),
    .o(_al_u6278_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~(B*A))"),
    .INIT(16'h0007))
    _al_u6279 (
    .a(\u_cmsdk_mcu/HADDR [9]),
    .b(\u_cmsdk_mcu/HADDR [8]),
    .c(\u_cmsdk_mcu/HADDR [6]),
    .d(\u_cmsdk_mcu/HADDR [5]),
    .o(_al_u6279_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u628 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n44 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [18]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n37 [14]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_baud_cntr_i [14]));
  AL_MAP_LUT4 #(
    .EQN("(D*~A*~(~C*~B))"),
    .INIT(16'h5400))
    _al_u6280 (
    .a(_al_u6276_o),
    .b(_al_u6277_o),
    .c(_al_u6278_o),
    .d(_al_u6279_o),
    .o(_al_u6280_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*A))"),
    .INIT(8'hc4))
    _al_u6281 (
    .a(\u_cmsdk_mcu/HADDR [4]),
    .b(\u_cmsdk_mcu/HADDR [3]),
    .c(\u_cmsdk_mcu/HADDR [2]),
    .o(_al_u6281_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*~B))"),
    .INIT(8'ha8))
    _al_u6282 (
    .a(\u_cmsdk_mcu/HADDR [5]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xg6iu6 ),
    .c(_al_u4423_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bg9iu6 ));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(D*~C))"),
    .INIT(16'h4044))
    _al_u6283 (
    .a(_al_u6281_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bg9iu6 ),
    .c(\u_cmsdk_mcu/HADDR [6]),
    .d(\u_cmsdk_mcu/HADDR [4]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uf9iu6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u6284 (
    .a(\u_cmsdk_mcu/HADDR [8]),
    .b(\u_cmsdk_mcu/HADDR [5]),
    .o(_al_u6284_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D*C*B))"),
    .INIT(16'h2aaa))
    _al_u6285 (
    .a(\u_cmsdk_mcu/HADDR [7]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xg6iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B79bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pg3qw6 ),
    .o(_al_u6285_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*A)"),
    .INIT(16'h0200))
    _al_u6286 (
    .a(_al_u6277_o),
    .b(_al_u6284_o),
    .c(_al_u6285_o),
    .d(\u_cmsdk_mcu/HADDR [10]),
    .o(_al_u6286_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(A*~(~D*~C)))"),
    .INIT(16'h444c))
    _al_u6287 (
    .a(\u_cmsdk_mcu/HADDR [7]),
    .b(\u_cmsdk_mcu/HADDR [6]),
    .c(\u_cmsdk_mcu/HADDR [3]),
    .d(\u_cmsdk_mcu/HADDR [2]),
    .o(_al_u6287_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*B*~(D*~A))"),
    .INIT(16'h080c))
    _al_u6288 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uf9iu6 ),
    .b(_al_u6286_o),
    .c(_al_u6287_o),
    .d(\u_cmsdk_mcu/HADDR [11]),
    .o(_al_u6288_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u6289 (
    .a(_al_u4921_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dpwpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kl8ax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvabx6 ),
    .o(_al_u6289_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u629 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n44 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [17]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n37 [13]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_baud_cntr_i [13]));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*A)"),
    .INIT(16'h0080))
    _al_u6290 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xg6iu6 ),
    .b(_al_u6289_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fs6iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Su8ax6 ),
    .o(_al_u6290_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    _al_u6291 (
    .a(_al_u4091_o),
    .b(_al_u4101_o),
    .c(_al_u4126_o),
    .d(_al_u4131_o),
    .o(_al_u6291_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u6292 (
    .a(_al_u4551_o),
    .b(_al_u6291_o),
    .c(_al_u4035_o),
    .d(_al_u4086_o),
    .o(_al_u6292_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*~A)"),
    .INIT(16'h4000))
    _al_u6293 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xg6iu6 ),
    .b(_al_u4919_o),
    .c(_al_u6292_o),
    .d(_al_u4056_o),
    .o(_al_u6293_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(~D*~C))"),
    .INIT(16'h8880))
    _al_u6294 (
    .a(\u_cmsdk_mcu/HADDR [15]),
    .b(\u_cmsdk_mcu/HSIZE [1]),
    .c(_al_u6290_o),
    .d(_al_u6293_o),
    .o(_al_u6294_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(~B*~A)))"),
    .INIT(16'h010f))
    _al_u6295 (
    .a(_al_u6280_o),
    .b(_al_u6288_o),
    .c(_al_u5000_o),
    .d(_al_u6294_o),
    .o(_al_u6295_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*(C@B))"),
    .INIT(8'h14))
    _al_u6296 (
    .a(_al_u5000_o),
    .b(\u_cmsdk_mcu/HADDR [10]),
    .c(\u_cmsdk_mcu/HADDR [3]),
    .o(_al_u6296_o));
  AL_MAP_LUT4 #(
    .EQN("~(~B*~A*~(D*C))"),
    .INIT(16'hfeee))
    _al_u6297 (
    .a(_al_u6295_o),
    .b(_al_u6296_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W5ypw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yavhu6 ));
  AL_MAP_LUT3 #(
    .EQN("(~A*(C@B))"),
    .INIT(8'h14))
    _al_u6298 (
    .a(_al_u5000_o),
    .b(\u_cmsdk_mcu/HADDR [7]),
    .c(\u_cmsdk_mcu/HADDR [2]),
    .o(_al_u6298_o));
  AL_MAP_LUT4 #(
    .EQN("~(~B*~A*~(D*C))"),
    .INIT(16'hfeee))
    _al_u6299 (
    .a(_al_u6295_o),
    .b(_al_u6298_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztupw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fbvhu6 ));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u630 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n44 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [16]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n37 [12]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_baud_cntr_i [12]));
  AL_MAP_LUT3 #(
    .EQN("(~A*(C@B))"),
    .INIT(8'h14))
    _al_u6300 (
    .a(_al_u5000_o),
    .b(\u_cmsdk_mcu/HADDR [5]),
    .c(\u_cmsdk_mcu/HADDR [3]),
    .o(_al_u6300_o));
  AL_MAP_LUT4 #(
    .EQN("~(~B*~A*~(D*C))"),
    .INIT(16'hfeee))
    _al_u6301 (
    .a(_al_u6295_o),
    .b(_al_u6300_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R9yax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mbvhu6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u6302 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I5xax6 ),
    .o(_al_u6302_o));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~A*~(~C*~B))"),
    .INIT(16'hffab))
    _al_u6303 (
    .a(_al_u6295_o),
    .b(_al_u5000_o),
    .c(\u_cmsdk_mcu/HADDR [4]),
    .d(_al_u6302_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hcvhu6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u6304 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yzspw6 ),
    .o(_al_u6304_o));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~A*~(~C*~B))"),
    .INIT(16'hffab))
    _al_u6305 (
    .a(_al_u6295_o),
    .b(_al_u5000_o),
    .c(\u_cmsdk_mcu/HADDR [8]),
    .d(_al_u6304_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tivhu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~D*~B*(C@A))"),
    .INIT(16'h0012))
    _al_u6306 (
    .a(_al_u6248_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F6ziu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P14qw6 ),
    .o(_al_u6306_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*B*A)"),
    .INIT(16'h0800))
    _al_u6307 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wh0ju6 ),
    .b(_al_u4376_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jckax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 ),
    .o(_al_u6307_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B*~A))"),
    .INIT(8'hb0))
    _al_u6308 (
    .a(_al_u6307_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rwjax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6 ),
    .o(_al_u6308_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~D*~C*~A))"),
    .INIT(16'hccc8))
    _al_u6309 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P14qw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rwjax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T6ziu6 ));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u631 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n44 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [15]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n37 [11]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_baud_cntr_i [11]));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(B*~A))"),
    .INIT(8'h0b))
    _al_u6310 (
    .a(_al_u6308_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T6ziu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 ),
    .o(_al_u6310_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(~B*~A))"),
    .INIT(8'he0))
    _al_u6311 (
    .a(_al_u6306_o),
    .b(_al_u6310_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W0piu6_lutinv ),
    .o(_al_u6311_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~(B@A))"),
    .INIT(16'h0009))
    _al_u6312 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dcziu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rwjax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Skjax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6 ),
    .o(_al_u6312_o));
  AL_MAP_LUT4 #(
    .EQN("(A*(B*~(C)*~(D)+~(B)*C*~(D)+B*~(C)*D+~(B)*C*D+B*C*D))"),
    .INIT(16'ha828))
    _al_u6313 (
    .a(_al_u6312_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N4kax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4jax6 ),
    .o(_al_u6313_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~B*~(C*~A))"),
    .INIT(16'h0023))
    _al_u6314 (
    .a(_al_u6313_o),
    .b(_al_u3419_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P14qw6 ),
    .o(_al_u6314_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(~A*~(~C*B)))"),
    .INIT(16'hae00))
    _al_u6315 (
    .a(_al_u6311_o),
    .b(_al_u3183_o),
    .c(_al_u6314_o),
    .d(_al_u2868_o),
    .o(_al_u6315_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*A)"),
    .INIT(16'h0080))
    _al_u6316 (
    .a(_al_u3223_o),
    .b(_al_u1367_o),
    .c(_al_u3124_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 ),
    .o(_al_u6316_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*~B*~A)"),
    .INIT(16'h0010))
    _al_u6317 (
    .a(_al_u1784_o),
    .b(_al_u1801_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oeziu6 ),
    .d(_al_u6316_o),
    .o(_al_u6317_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(~D*C))"),
    .INIT(16'h8808))
    _al_u6318 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Veziu6 ),
    .b(_al_u6317_o),
    .c(_al_u3202_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 ),
    .o(_al_u6318_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*~A))"),
    .INIT(8'h8c))
    _al_u6319 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z37ow6_lutinv ),
    .b(_al_u4161_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ),
    .o(_al_u6319_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u632 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n44 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [14]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n37 [10]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_baud_cntr_i [10]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u6320 (
    .a(_al_u903_o),
    .b(_al_u3094_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 ),
    .o(_al_u6320_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(D*C*B))"),
    .INIT(16'h1555))
    _al_u6321 (
    .a(_al_u6320_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D6kiu6_lutinv ),
    .d(_al_u1266_o),
    .o(_al_u6321_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    _al_u6322 (
    .a(_al_u3664_o),
    .b(_al_u6319_o),
    .c(_al_u6321_o),
    .o(_al_u6322_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*~B))"),
    .INIT(8'h8a))
    _al_u6323 (
    .a(_al_u6322_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wxyiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gebow6_lutinv ),
    .o(_al_u6323_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u6324 (
    .a(_al_u2364_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 ),
    .o(_al_u6324_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(~D*B*A))"),
    .INIT(16'h0f07))
    _al_u6325 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuyiu6_lutinv ),
    .b(_al_u4393_o),
    .c(_al_u6324_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6 ),
    .o(_al_u6325_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(~D*C))"),
    .INIT(16'h8808))
    _al_u6326 (
    .a(_al_u6318_o),
    .b(_al_u6323_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Htyiu6 ),
    .d(_al_u6325_o),
    .o(_al_u6326_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~A*~(D*B))"),
    .INIT(16'h0105))
    _al_u6327 (
    .a(_al_u3101_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N3ziu6 ),
    .c(_al_u3236_o),
    .d(_al_u1271_o),
    .o(_al_u6327_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*A*~(D*B))"),
    .INIT(16'h020a))
    _al_u6328 (
    .a(_al_u6327_o),
    .b(_al_u2361_o),
    .c(_al_u3078_o),
    .d(_al_u3401_o),
    .o(_al_u6328_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(~D*~C))"),
    .INIT(16'h8880))
    _al_u6329 (
    .a(_al_u6326_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rcziu6 ),
    .c(_al_u6328_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vygax6 ),
    .o(_al_u6329_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u633 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n44 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [5]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n37 [1]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_baud_cntr_i [1]));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*C)*~(B*~A))"),
    .INIT(16'hbb0b))
    _al_u6330 (
    .a(_al_u6315_o),
    .b(_al_u6329_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vgjpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oxohu6 ));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*~(~D*B))"),
    .INIT(16'h5010))
    _al_u6331 (
    .a(_al_u5329_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gz6ax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mnmpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uj4bx6 ),
    .o(_al_u6331_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(C*~A))"),
    .INIT(16'haf23))
    _al_u6332 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gz6ax6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tl4bx6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uj4bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vpgbx6 ),
    .o(_al_u6332_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(~B*A))"),
    .INIT(8'hd0))
    _al_u6333 (
    .a(_al_u6331_o),
    .b(_al_u6332_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F17ax6 ),
    .o(_al_u6333_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u6334 (
    .a(_al_u6333_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gz6ax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uj4bx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rerow6_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u6335 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F17ax6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mnmpw6 ),
    .o(_al_u6335_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u6336 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rerow6_lutinv ),
    .b(_al_u6335_o),
    .o(_al_u6336_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u6337 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C10bx6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qo3bx6 ),
    .o(_al_u6337_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u6338 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lr9bx6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nt9bx6 ),
    .o(_al_u6338_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(C)*~((D*~B))+~(A)*C*~((D*~B))+A*C*~((D*~B))+~(A)*C*(D*~B))"),
    .INIT(16'hd4f5))
    _al_u6339 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Auyax6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cwyax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eyyax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tngbx6 ),
    .o(_al_u6339_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u634 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n44 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [4]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n37 [0]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_baud_cntr_i [0]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*A))"),
    .INIT(8'hc4))
    _al_u6340 (
    .a(_al_u6337_o),
    .b(_al_u6338_o),
    .c(_al_u6339_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hkgow6 ));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    _al_u6341 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hkgow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Auyax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eyyax6 ),
    .o(_al_u6341_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u6342 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Czzax6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mk3bx6 ),
    .o(_al_u6342_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u6343 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gihbx6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ikhbx6 ),
    .o(_al_u6343_o));
  AL_MAP_LUT4 #(
    .EQN("(~(B)*~((~C*A))*~(D)+~(B)*~((~C*A))*D+B*~((~C*A))*D+~(B)*(~C*A)*D)"),
    .INIT(16'hf731))
    _al_u6344 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bcabx6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S3mpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vbspw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yryax6 ),
    .o(_al_u6344_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*A))"),
    .INIT(8'hc4))
    _al_u6345 (
    .a(_al_u6342_o),
    .b(_al_u6343_o),
    .c(_al_u6344_o),
    .o(_al_u6345_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u6346 (
    .a(_al_u6345_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S3mpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yryax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oltow6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(B*~(~C*A)))"),
    .INIT(16'h003b))
    _al_u6347 (
    .a(_al_u6342_o),
    .b(_al_u6343_o),
    .c(_al_u6344_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vbspw6 ),
    .o(_al_u6347_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*B*~(~C*A))"),
    .INIT(16'h00c4))
    _al_u6348 (
    .a(_al_u6342_o),
    .b(_al_u6343_o),
    .c(_al_u6344_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bcabx6 ),
    .o(_al_u6348_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(B*~(~C*A)))"),
    .INIT(16'h003b))
    _al_u6349 (
    .a(_al_u6337_o),
    .b(_al_u6338_o),
    .c(_al_u6339_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cwyax6 ),
    .o(_al_u6349_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u635 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_state [0]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_state [1]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/lt2/o_1_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(~D*B*~(~C*A))"),
    .INIT(16'h00c4))
    _al_u6350 (
    .a(_al_u6337_o),
    .b(_al_u6338_o),
    .c(_al_u6339_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tngbx6 ),
    .o(_al_u6350_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~A*~(~D*~C))"),
    .INIT(16'h1110))
    _al_u6351 (
    .a(_al_u6347_o),
    .b(_al_u6348_o),
    .c(_al_u6349_o),
    .d(_al_u6350_o),
    .o(_al_u6351_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u6352 (
    .a(_al_u6337_o),
    .b(_al_u6338_o),
    .o(_al_u6352_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(A*B*~(C)+A*~(B)*C+~(A)*B*C+A*B*C))"),
    .INIT(16'h00e8))
    _al_u6353 (
    .a(_al_u6341_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oltow6_lutinv ),
    .c(_al_u6351_o),
    .d(_al_u6352_o),
    .o(_al_u6353_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u6354 (
    .a(_al_u6342_o),
    .b(_al_u6343_o),
    .o(_al_u6354_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C)*~((~D*~A))+~B*C*~((~D*~A))+~(~B)*C*(~D*~A)+~B*C*(~D*~A))"),
    .INIT(16'h3372))
    _al_u6355 (
    .a(_al_u6353_o),
    .b(_al_u6341_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oltow6_lutinv ),
    .d(_al_u6354_o),
    .o(_al_u6355_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(~C*A))"),
    .INIT(16'hc4f5))
    _al_u6356 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C5gbx6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgzax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uizax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vkzax6 ),
    .o(_al_u6356_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(~D*C))"),
    .INIT(16'h8808))
    _al_u6357 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Muhbx6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Owhbx6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgzax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vkzax6 ),
    .o(_al_u6357_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u6358 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L1bbx6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5bbx6 ),
    .o(_al_u6358_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B*~A))"),
    .INIT(8'hb0))
    _al_u6359 (
    .a(_al_u6356_o),
    .b(_al_u6357_o),
    .c(_al_u6358_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mjgow6 ));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u636 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/lt2/o_1_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_state [2]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_state [3]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_buf_full ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n63 ));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u6360 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mjgow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Muhbx6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Owhbx6 ),
    .o(_al_u6360_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u6361 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mjgow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgzax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vkzax6 ),
    .o(_al_u6361_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u6362 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C3wpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U31bx6 ),
    .o(_al_u6362_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(~C*A))"),
    .INIT(16'hc4f5))
    _al_u6363 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nv9bx6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wmzax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xozax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yqzax6 ),
    .o(_al_u6363_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(~D*C))"),
    .INIT(16'h8808))
    _al_u6364 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aa2bx6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cxzax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wmzax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yqzax6 ),
    .o(_al_u6364_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*~B))"),
    .INIT(8'h8a))
    _al_u6365 (
    .a(_al_u6362_o),
    .b(_al_u6363_o),
    .c(_al_u6364_o),
    .o(_al_u6365_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u6366 (
    .a(_al_u6365_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wmzax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yqzax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xttow6_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(~B*A))"),
    .INIT(8'h0d))
    _al_u6367 (
    .a(_al_u6362_o),
    .b(_al_u6364_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xozax6 ),
    .o(_al_u6367_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*A*~(C*~B))"),
    .INIT(16'h008a))
    _al_u6368 (
    .a(_al_u6362_o),
    .b(_al_u6363_o),
    .c(_al_u6364_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nv9bx6 ),
    .o(_al_u6368_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(B*~A))"),
    .INIT(8'h0b))
    _al_u6369 (
    .a(_al_u6357_o),
    .b(_al_u6358_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uizax6 ),
    .o(_al_u6369_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u637 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_state_inc ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n61 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n63 ),
    .o(_al_u637_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*~(B*~A))"),
    .INIT(16'h00b0))
    _al_u6370 (
    .a(_al_u6356_o),
    .b(_al_u6357_o),
    .c(_al_u6358_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C5gbx6 ),
    .o(_al_u6370_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~A*~(~D*~C))"),
    .INIT(16'h1110))
    _al_u6371 (
    .a(_al_u6367_o),
    .b(_al_u6368_o),
    .c(_al_u6369_o),
    .d(_al_u6370_o),
    .o(_al_u6371_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*(B*C*~(D)+B*~(C)*D+~(B)*C*D+B*C*D))"),
    .INIT(16'h5440))
    _al_u6372 (
    .a(_al_u6360_o),
    .b(_al_u6361_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xttow6_lutinv ),
    .d(_al_u6371_o),
    .o(_al_u6372_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u6373 (
    .a(_al_u6362_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aa2bx6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cxzax6 ),
    .o(_al_u6373_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C)*~((~D*~A))+~B*C*~((~D*~A))+~(~B)*C*(~D*~A)+~B*C*(~D*~A))"),
    .INIT(16'h3372))
    _al_u6374 (
    .a(_al_u6372_o),
    .b(_al_u6361_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xttow6_lutinv ),
    .d(_al_u6373_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oetow6_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u6375 (
    .a(_al_u6347_o),
    .b(_al_u6348_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rjtow6_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u6376 (
    .a(_al_u6349_o),
    .b(_al_u6350_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yjtow6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B)*~((~D*~A))+C*B*~((~D*~A))+~(C)*B*(~D*~A)+C*B*(~D*~A))"),
    .INIT(16'hf0e4))
    _al_u6377 (
    .a(_al_u6353_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rjtow6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yjtow6_lutinv ),
    .d(_al_u6354_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q8tow6_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u6378 (
    .a(_al_u6367_o),
    .b(_al_u6368_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iwtow6_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u6379 (
    .a(_al_u6369_o),
    .b(_al_u6370_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tktow6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("~(A*~(B*~(~D*C)))"),
    .INIT(16'hdd5d))
    _al_u638 (
    .a(_al_u637_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_state_inc ),
    .c(_al_u379_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/lt2/o_1_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n74 ));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B)*~((~D*~A))+C*B*~((~D*~A))+~(C)*B*(~D*~A)+C*B*(~D*~A))"),
    .INIT(16'hf0e4))
    _al_u6380 (
    .a(_al_u6372_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iwtow6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tktow6_lutinv ),
    .d(_al_u6373_o),
    .o(_al_u6380_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~C)*~(B*~A))"),
    .INIT(16'hb0bb))
    _al_u6381 (
    .a(_al_u6355_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oetow6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q8tow6_lutinv ),
    .d(_al_u6380_o),
    .o(_al_u6381_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u6382 (
    .a(_al_u6352_o),
    .b(_al_u6354_o),
    .o(_al_u6382_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(~B*A))"),
    .INIT(8'h0d))
    _al_u6383 (
    .a(_al_u6355_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oetow6_lutinv ),
    .c(_al_u6382_o),
    .o(_al_u6383_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u6384 (
    .a(_al_u6360_o),
    .b(_al_u6373_o),
    .o(_al_u6384_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(B*~A))"),
    .INIT(8'h0b))
    _al_u6385 (
    .a(_al_u6381_o),
    .b(_al_u6383_o),
    .c(_al_u6384_o),
    .o(_al_u6385_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u6386 (
    .a(_al_u6385_o),
    .b(_al_u6355_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oetow6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Irrow6_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u6387 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D70bx6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lg1bx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F5uow6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u6388 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C50bx6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fc1bx6 ),
    .o(_al_u6388_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~((C*~B))*~(D)+~(A)*~((C*~B))*D+A*~((C*~B))*D+~(A)*(C*~B)*D)"),
    .INIT(16'hdf45))
    _al_u6389 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Od4bx6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qf4bx6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rlgbx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sh4bx6 ),
    .o(_al_u6389_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    _al_u639 (
    .a(_al_u637_o),
    .b(uart0_txen_pad),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_ctrl [2]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/intr_stat_set [0]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*A))"),
    .INIT(8'hc4))
    _al_u6390 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F5uow6 ),
    .b(_al_u6388_o),
    .c(_al_u6389_o),
    .o(_al_u6390_o));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    _al_u6391 (
    .a(_al_u6390_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Od4bx6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sh4bx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Phuow6_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u6392 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rijbx6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tkjbx6 ),
    .o(_al_u6392_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u6393 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C30bx6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Us3bx6 ),
    .o(_al_u6393_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(C)*~((D*~B))+~(A)*C*~((D*~B))+A*C*~((D*~B))+~(A)*C*(D*~B))"),
    .INIT(16'hd4f5))
    _al_u6394 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I74bx6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K94bx6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mb4bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z9abx6 ),
    .o(_al_u6394_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*A))"),
    .INIT(8'hc4))
    _al_u6395 (
    .a(_al_u6392_o),
    .b(_al_u6393_o),
    .c(_al_u6394_o),
    .o(_al_u6395_o));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    _al_u6396 (
    .a(_al_u6395_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I74bx6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mb4bx6 ),
    .o(_al_u6396_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(B*~(~C*A)))"),
    .INIT(16'h003b))
    _al_u6397 (
    .a(_al_u6392_o),
    .b(_al_u6393_o),
    .c(_al_u6394_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K94bx6 ),
    .o(_al_u6397_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*B*~(~C*A))"),
    .INIT(16'h00c4))
    _al_u6398 (
    .a(_al_u6392_o),
    .b(_al_u6393_o),
    .c(_al_u6394_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z9abx6 ),
    .o(_al_u6398_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(B*~(~C*A)))"),
    .INIT(16'h003b))
    _al_u6399 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F5uow6 ),
    .b(_al_u6388_o),
    .c(_al_u6389_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qf4bx6 ),
    .o(_al_u6399_o));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    _al_u640 (
    .a(_al_u637_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_tx_buf [7]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_tx_shift_buf [7]));
  AL_MAP_LUT4 #(
    .EQN("(~D*B*~(~C*A))"),
    .INIT(16'h00c4))
    _al_u6400 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F5uow6 ),
    .b(_al_u6388_o),
    .c(_al_u6389_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rlgbx6 ),
    .o(_al_u6400_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~A*~(~D*~C))"),
    .INIT(16'h1110))
    _al_u6401 (
    .a(_al_u6397_o),
    .b(_al_u6398_o),
    .c(_al_u6399_o),
    .d(_al_u6400_o),
    .o(_al_u6401_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u6402 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F5uow6 ),
    .b(_al_u6388_o),
    .o(_al_u6402_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(A*~(B)*~(C)+~(A)*~(B)*C+A*~(B)*C+A*B*C))"),
    .INIT(16'h00b2))
    _al_u6403 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Phuow6_lutinv ),
    .b(_al_u6396_o),
    .c(_al_u6401_o),
    .d(_al_u6402_o),
    .o(_al_u6403_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u6404 (
    .a(_al_u6392_o),
    .b(_al_u6393_o),
    .o(_al_u6404_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(C)*~((~D*~A))+B*C*~((~D*~A))+~(B)*C*(~D*~A)+B*C*(~D*~A))"),
    .INIT(16'hccd8))
    _al_u6405 (
    .a(_al_u6403_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Phuow6_lutinv ),
    .c(_al_u6396_o),
    .d(_al_u6404_o),
    .o(_al_u6405_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u6406 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fb0bx6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rk1bx6 ),
    .o(_al_u6406_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u6407 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E90bx6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z71bx6 ),
    .o(_al_u6407_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(C)*~((D*~B))+~(A)*C*~((D*~B))+A*C*~((D*~B))+~(A)*C*(D*~B))"),
    .INIT(16'hd4f5))
    _al_u6408 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E05bx6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G25bx6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I45bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X7abx6 ),
    .o(_al_u6408_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*A))"),
    .INIT(8'hc4))
    _al_u6409 (
    .a(_al_u6406_o),
    .b(_al_u6407_o),
    .c(_al_u6408_o),
    .o(_al_u6409_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u641 (
    .a(_al_u637_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_tx_buf [6]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_shift_buf [7]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_tx_shift_buf [6]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u6410 (
    .a(_al_u6409_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E05bx6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I45bx6 ),
    .o(_al_u6410_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u6411 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hf0bx6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yxrpw6 ),
    .o(_al_u6411_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u6412 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gd0bx6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xo1bx6 ),
    .o(_al_u6412_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(C)*~((D*~B))+~(A)*C*~((D*~B))+A*C*~((D*~B))+~(A)*C*(D*~B))"),
    .INIT(16'hd4f5))
    _al_u6413 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K65bx6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M85bx6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oa5bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pjgbx6 ),
    .o(_al_u6413_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*A))"),
    .INIT(8'hc4))
    _al_u6414 (
    .a(_al_u6411_o),
    .b(_al_u6412_o),
    .c(_al_u6413_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Whgow6 ));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    _al_u6415 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Whgow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K65bx6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oa5bx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G9uow6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(B*~(~C*A)))"),
    .INIT(16'h003b))
    _al_u6416 (
    .a(_al_u6406_o),
    .b(_al_u6407_o),
    .c(_al_u6408_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G25bx6 ),
    .o(_al_u6416_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*B*~(~C*A))"),
    .INIT(16'h00c4))
    _al_u6417 (
    .a(_al_u6406_o),
    .b(_al_u6407_o),
    .c(_al_u6408_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X7abx6 ),
    .o(_al_u6417_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(B*~(~C*A)))"),
    .INIT(16'h003b))
    _al_u6418 (
    .a(_al_u6411_o),
    .b(_al_u6412_o),
    .c(_al_u6413_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M85bx6 ),
    .o(_al_u6418_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*B*~(~C*A))"),
    .INIT(16'h00c4))
    _al_u6419 (
    .a(_al_u6411_o),
    .b(_al_u6412_o),
    .c(_al_u6413_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pjgbx6 ),
    .o(_al_u6419_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u642 (
    .a(_al_u637_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_tx_buf [5]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_shift_buf [6]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_tx_shift_buf [5]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~A*~(~D*~C))"),
    .INIT(16'h1110))
    _al_u6420 (
    .a(_al_u6416_o),
    .b(_al_u6417_o),
    .c(_al_u6418_o),
    .d(_al_u6419_o),
    .o(_al_u6420_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u6421 (
    .a(_al_u6411_o),
    .b(_al_u6412_o),
    .o(_al_u6421_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(A*B*~(C)+A*~(B)*C+~(A)*B*C+A*B*C))"),
    .INIT(16'h00e8))
    _al_u6422 (
    .a(_al_u6410_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G9uow6_lutinv ),
    .c(_al_u6420_o),
    .d(_al_u6421_o),
    .o(_al_u6422_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u6423 (
    .a(_al_u6406_o),
    .b(_al_u6407_o),
    .o(_al_u6423_o));
  AL_MAP_LUT4 #(
    .EQN("~(~C*~(B)*~((~D*~A))+~C*B*~((~D*~A))+~(~C)*B*(~D*~A)+~C*B*(~D*~A))"),
    .INIT(16'hf0b1))
    _al_u6424 (
    .a(_al_u6422_o),
    .b(_al_u6410_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G9uow6_lutinv ),
    .d(_al_u6423_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tdtow6_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u6425 (
    .a(_al_u6397_o),
    .b(_al_u6398_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Akuow6_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u6426 (
    .a(_al_u6399_o),
    .b(_al_u6400_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L8uow6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B)*~((~D*~A))+C*B*~((~D*~A))+~(C)*B*(~D*~A)+C*B*(~D*~A))"),
    .INIT(16'hf0e4))
    _al_u6427 (
    .a(_al_u6403_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Akuow6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L8uow6_lutinv ),
    .d(_al_u6404_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yctow6_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u6428 (
    .a(_al_u6416_o),
    .b(_al_u6417_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q7uow6_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u6429 (
    .a(_al_u6418_o),
    .b(_al_u6419_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E8uow6_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u643 (
    .a(_al_u637_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_tx_buf [4]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_shift_buf [5]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_tx_shift_buf [4]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B)*~((~D*~A))+C*B*~((~D*~A))+~(C)*B*(~D*~A)+C*B*(~D*~A))"),
    .INIT(16'hf0e4))
    _al_u6430 (
    .a(_al_u6422_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q7uow6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E8uow6_lutinv ),
    .d(_al_u6423_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P3uow6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*C)*~(B*~A))"),
    .INIT(16'hbb0b))
    _al_u6431 (
    .a(_al_u6405_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tdtow6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yctow6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P3uow6_lutinv ),
    .o(_al_u6431_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u6432 (
    .a(_al_u6421_o),
    .b(_al_u6423_o),
    .o(_al_u6432_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(~B*A))"),
    .INIT(8'h0d))
    _al_u6433 (
    .a(_al_u6405_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tdtow6_lutinv ),
    .c(_al_u6432_o),
    .o(_al_u6433_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u6434 (
    .a(_al_u6404_o),
    .b(_al_u6402_o),
    .o(_al_u6434_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(B*~A))"),
    .INIT(8'h0b))
    _al_u6435 (
    .a(_al_u6431_o),
    .b(_al_u6433_o),
    .c(_al_u6434_o),
    .o(_al_u6435_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u6436 (
    .a(_al_u6435_o),
    .b(_al_u6405_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tdtow6_lutinv ),
    .o(_al_u6436_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(~D*~(B*~A)))"),
    .INIT(16'hf040))
    _al_u6437 (
    .a(_al_u6381_o),
    .b(_al_u6383_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q8tow6_lutinv ),
    .d(_al_u6384_o),
    .o(_al_u6437_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*~(B*~A))"),
    .INIT(16'h00b0))
    _al_u6438 (
    .a(_al_u6381_o),
    .b(_al_u6383_o),
    .c(_al_u6380_o),
    .d(_al_u6384_o),
    .o(_al_u6438_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*~A))"),
    .INIT(8'h32))
    _al_u6439 (
    .a(_al_u6433_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P3uow6_lutinv ),
    .c(_al_u6434_o),
    .o(_al_u6439_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u644 (
    .a(_al_u637_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_tx_buf [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_shift_buf [4]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_tx_shift_buf [3]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~(B*~A))"),
    .INIT(16'h000b))
    _al_u6440 (
    .a(_al_u6431_o),
    .b(_al_u6433_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yctow6_lutinv ),
    .d(_al_u6434_o),
    .o(_al_u6440_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*~C)*~(~B*~A))"),
    .INIT(16'heee0))
    _al_u6441 (
    .a(_al_u6437_o),
    .b(_al_u6438_o),
    .c(_al_u6439_o),
    .d(_al_u6440_o),
    .o(_al_u6441_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u6442 (
    .a(_al_u6435_o),
    .b(_al_u6432_o),
    .o(_al_u6442_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(A*B*~(C)+A*~(B)*C+~(A)*B*C+A*B*C))"),
    .INIT(16'h00e8))
    _al_u6443 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Irrow6_lutinv ),
    .b(_al_u6436_o),
    .c(_al_u6441_o),
    .d(_al_u6442_o),
    .o(_al_u6443_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u6444 (
    .a(_al_u6384_o),
    .b(_al_u6382_o),
    .o(_al_u6444_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u6445 (
    .a(_al_u6443_o),
    .b(_al_u6444_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B4fow6 ));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    _al_u6446 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B4fow6 ),
    .b(_al_u6435_o),
    .c(_al_u6432_o),
    .o(_al_u6446_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(~C*A))"),
    .INIT(16'hf531))
    _al_u6447 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pz9bx6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sn4bx6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Up4bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wr4bx6 ),
    .o(_al_u6447_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*~C))"),
    .INIT(16'h8088))
    _al_u6448 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bc3bx6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kojpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sn4bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wr4bx6 ),
    .o(_al_u6448_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u6449 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Usipw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V73bx6 ),
    .o(_al_u6449_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u645 (
    .a(_al_u637_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_tx_buf [2]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_shift_buf [3]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_tx_shift_buf [2]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B*~A))"),
    .INIT(8'hb0))
    _al_u6450 (
    .a(_al_u6447_o),
    .b(_al_u6448_o),
    .c(_al_u6449_o),
    .o(_al_u6450_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u6451 (
    .a(_al_u6450_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sn4bx6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wr4bx6 ),
    .o(_al_u6451_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(C*~A))"),
    .INIT(16'h8caf))
    _al_u6452 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aw4bx6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cy4bx6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hbgbx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yt4bx6 ),
    .o(_al_u6452_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*~(~D*A))"),
    .INIT(16'hc040))
    _al_u6453 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cy4bx6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hg3bx6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S0kbx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yt4bx6 ),
    .o(_al_u6453_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u6454 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rz0bx6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tcipw6 ),
    .o(_al_u6454_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B*~A))"),
    .INIT(8'hb0))
    _al_u6455 (
    .a(_al_u6452_o),
    .b(_al_u6453_o),
    .c(_al_u6454_o),
    .o(_al_u6455_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u6456 (
    .a(_al_u6455_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cy4bx6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yt4bx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gpsow6_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(B*~A))"),
    .INIT(8'h0b))
    _al_u6457 (
    .a(_al_u6448_o),
    .b(_al_u6449_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Up4bx6 ),
    .o(_al_u6457_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*~(B*~A))"),
    .INIT(16'h00b0))
    _al_u6458 (
    .a(_al_u6447_o),
    .b(_al_u6448_o),
    .c(_al_u6449_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pz9bx6 ),
    .o(_al_u6458_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(B*~A))"),
    .INIT(8'h0b))
    _al_u6459 (
    .a(_al_u6453_o),
    .b(_al_u6454_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aw4bx6 ),
    .o(_al_u6459_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u646 (
    .a(_al_u637_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_tx_buf [1]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_shift_buf [2]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_tx_shift_buf [1]));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*~(B*~A))"),
    .INIT(16'h00b0))
    _al_u6460 (
    .a(_al_u6452_o),
    .b(_al_u6453_o),
    .c(_al_u6454_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hbgbx6 ),
    .o(_al_u6460_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~A*~(~D*~C))"),
    .INIT(16'h1110))
    _al_u6461 (
    .a(_al_u6457_o),
    .b(_al_u6458_o),
    .c(_al_u6459_o),
    .d(_al_u6460_o),
    .o(_al_u6461_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u6462 (
    .a(_al_u6455_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hg3bx6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S0kbx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tmrow6 ));
  AL_MAP_LUT4 #(
    .EQN("(~D*(A*B*~(C)+A*~(B)*C+~(A)*B*C+A*B*C))"),
    .INIT(16'h00e8))
    _al_u6463 (
    .a(_al_u6451_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gpsow6_lutinv ),
    .c(_al_u6461_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tmrow6 ),
    .o(_al_u6463_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u6464 (
    .a(_al_u6450_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bc3bx6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kojpw6 ),
    .o(_al_u6464_o));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~(B)*~((~C*~A))+~D*B*~((~C*~A))+~(~D)*B*(~C*~A)+~D*B*(~C*~A))"),
    .INIT(16'hfb01))
    _al_u6465 (
    .a(_al_u6463_o),
    .b(_al_u6451_o),
    .c(_al_u6464_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gpsow6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxrow6_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u6466 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P33bx6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qx0bx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Amsow6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u6467 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jz2bx6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X5upw6 ),
    .o(_al_u6467_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(C)*~((D*~B))+~(A)*C*~((D*~B))+A*C*~((D*~B))+~(A)*C*(D*~B))"),
    .INIT(16'hd4f5))
    _al_u6468 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C14bx6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E34bx6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G54bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jdgbx6 ),
    .o(_al_u6468_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*A))"),
    .INIT(8'hc4))
    _al_u6469 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Amsow6 ),
    .b(_al_u6467_o),
    .c(_al_u6468_o),
    .o(_al_u6469_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u647 (
    .a(_al_u637_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_tx_buf [0]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_shift_buf [1]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_tx_shift_buf [0]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    _al_u6470 (
    .a(_al_u6469_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C14bx6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G54bx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Upsow6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(C*~A))"),
    .INIT(16'haf23))
    _al_u6471 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Az3bx6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R1abx6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wu3bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yw3bx6 ),
    .o(_al_u6471_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*~(~D*A))"),
    .INIT(16'hc040))
    _al_u6472 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Az3bx6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pv0bx6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rm2bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wu3bx6 ),
    .o(_al_u6472_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u6473 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dv2bx6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oxkpw6 ),
    .o(_al_u6473_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B*~A))"),
    .INIT(8'hb0))
    _al_u6474 (
    .a(_al_u6471_o),
    .b(_al_u6472_o),
    .c(_al_u6473_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Odgow6 ));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u6475 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Odgow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Az3bx6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wu3bx6 ),
    .o(_al_u6475_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(B*~A))"),
    .INIT(8'h0b))
    _al_u6476 (
    .a(_al_u6472_o),
    .b(_al_u6473_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yw3bx6 ),
    .o(_al_u6476_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*~(B*~A))"),
    .INIT(16'h00b0))
    _al_u6477 (
    .a(_al_u6471_o),
    .b(_al_u6472_o),
    .c(_al_u6473_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R1abx6 ),
    .o(_al_u6477_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(B*~(~C*A)))"),
    .INIT(16'h003b))
    _al_u6478 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Amsow6 ),
    .b(_al_u6467_o),
    .c(_al_u6468_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E34bx6 ),
    .o(_al_u6478_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*B*~(~C*A))"),
    .INIT(16'h00c4))
    _al_u6479 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Amsow6 ),
    .b(_al_u6467_o),
    .c(_al_u6468_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jdgbx6 ),
    .o(_al_u6479_o));
  AL_MAP_LUT2 #(
    .EQN("~(B*~A)"),
    .INIT(4'hb))
    _al_u648 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/write_enable00 ),
    .b(_al_u637_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n50 ));
  AL_MAP_LUT4 #(
    .EQN("(~B*~A*~(~D*~C))"),
    .INIT(16'h1110))
    _al_u6480 (
    .a(_al_u6476_o),
    .b(_al_u6477_o),
    .c(_al_u6478_o),
    .d(_al_u6479_o),
    .o(_al_u6480_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u6481 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Amsow6 ),
    .b(_al_u6467_o),
    .o(_al_u6481_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(A*~(B)*~(C)+~(A)*~(B)*C+A*~(B)*C+A*B*C))"),
    .INIT(16'h00b2))
    _al_u6482 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Upsow6_lutinv ),
    .b(_al_u6475_o),
    .c(_al_u6480_o),
    .d(_al_u6481_o),
    .o(_al_u6482_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u6483 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Odgow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pv0bx6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rm2bx6 ),
    .o(_al_u6483_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((~B*~A))+C*D*~((~B*~A))+~(C)*D*(~B*~A)+C*D*(~B*~A))"),
    .INIT(16'hf1e0))
    _al_u6484 (
    .a(_al_u6482_o),
    .b(_al_u6483_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Upsow6_lutinv ),
    .d(_al_u6475_o),
    .o(_al_u6484_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u6485 (
    .a(_al_u6476_o),
    .b(_al_u6477_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iqsow6_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u6486 (
    .a(_al_u6478_o),
    .b(_al_u6479_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pqsow6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C)*~((~B*~A))+D*C*~((~B*~A))+~(D)*C*(~B*~A)+D*C*(~B*~A))"),
    .INIT(16'hfe10))
    _al_u6487 (
    .a(_al_u6482_o),
    .b(_al_u6483_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iqsow6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pqsow6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yksow6_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u6488 (
    .a(_al_u6457_o),
    .b(_al_u6458_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tzsow6_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u6489 (
    .a(_al_u6459_o),
    .b(_al_u6460_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fzsow6_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    _al_u649 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/write_enable10 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/baud_updated ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n46 ));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C)*~((~B*~A))+D*C*~((~B*~A))+~(D)*C*(~B*~A)+D*C*(~B*~A))"),
    .INIT(16'hfe10))
    _al_u6490 (
    .a(_al_u6463_o),
    .b(_al_u6464_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tzsow6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fzsow6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rksow6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*C)*~(~B*A))"),
    .INIT(16'hdd0d))
    _al_u6491 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxrow6_lutinv ),
    .b(_al_u6484_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yksow6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rksow6_lutinv ),
    .o(_al_u6491_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u6492 (
    .a(_al_u6464_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tmrow6 ),
    .o(_al_u6492_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(B*~A))"),
    .INIT(8'h0b))
    _al_u6493 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxrow6_lutinv ),
    .b(_al_u6484_o),
    .c(_al_u6492_o),
    .o(_al_u6493_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u6494 (
    .a(_al_u6483_o),
    .b(_al_u6481_o),
    .o(_al_u6494_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(B*~A))"),
    .INIT(8'h0b))
    _al_u6495 (
    .a(_al_u6491_o),
    .b(_al_u6493_o),
    .c(_al_u6494_o),
    .o(_al_u6495_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u6496 (
    .a(_al_u6495_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxrow6_lutinv ),
    .c(_al_u6484_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gqrow6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*B)*~(~D*A))"),
    .INIT(16'hf351))
    _al_u6497 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nazax6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nhgbx6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pczax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rezax6 ),
    .o(_al_u6497_o));
  AL_MAP_LUT4 #(
    .EQN("(D*A*~(C*~B))"),
    .INIT(16'h8a00))
    _al_u6498 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ln0bx6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nazax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rezax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V52bx6 ),
    .o(_al_u6498_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u6499 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kl0bx6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P12bx6 ),
    .o(_al_u6499_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*A)"),
    .INIT(16'h0080))
    _al_u650 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/read_enable ),
    .b(_al_u473_o),
    .c(_al_u467_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/state_reg [0]),
    .o(_al_u650_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B*~A))"),
    .INIT(8'hb0))
    _al_u6500 (
    .a(_al_u6497_o),
    .b(_al_u6498_o),
    .c(_al_u6499_o),
    .o(_al_u6500_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u6501 (
    .a(_al_u6500_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nazax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rezax6 ),
    .o(_al_u6501_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(~C*A))"),
    .INIT(16'hc4f5))
    _al_u6502 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H4zax6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J6zax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L8zax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V5abx6 ),
    .o(_al_u6502_o));
  AL_MAP_LUT4 #(
    .EQN("(C*A*~(D*~B))"),
    .INIT(16'h80a0))
    _al_u6503 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dt1bx6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H4zax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jj0bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L8zax6 ),
    .o(_al_u6503_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u6504 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ih0bx6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jx1bx6 ),
    .o(_al_u6504_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B*~A))"),
    .INIT(8'hb0))
    _al_u6505 (
    .a(_al_u6502_o),
    .b(_al_u6503_o),
    .c(_al_u6504_o),
    .o(_al_u6505_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u6506 (
    .a(_al_u6505_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H4zax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L8zax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J2sow6_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(B*~A))"),
    .INIT(8'h0b))
    _al_u6507 (
    .a(_al_u6498_o),
    .b(_al_u6499_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pczax6 ),
    .o(_al_u6507_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*~(B*~A))"),
    .INIT(16'h00b0))
    _al_u6508 (
    .a(_al_u6497_o),
    .b(_al_u6498_o),
    .c(_al_u6499_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nhgbx6 ),
    .o(_al_u6508_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(B*~A))"),
    .INIT(8'h0b))
    _al_u6509 (
    .a(_al_u6503_o),
    .b(_al_u6504_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J6zax6 ),
    .o(_al_u6509_o));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    _al_u651 (
    .a(_al_u650_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rxbuf_sample ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n106 ));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*~(B*~A))"),
    .INIT(16'h00b0))
    _al_u6510 (
    .a(_al_u6502_o),
    .b(_al_u6503_o),
    .c(_al_u6504_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V5abx6 ),
    .o(_al_u6510_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~(~B*~A))"),
    .INIT(16'h000e))
    _al_u6511 (
    .a(_al_u6507_o),
    .b(_al_u6508_o),
    .c(_al_u6509_o),
    .d(_al_u6510_o),
    .o(_al_u6511_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u6512 (
    .a(_al_u6500_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ln0bx6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V52bx6 ),
    .o(_al_u6512_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(~(A)*B*~(C)+~(A)*~(B)*C+~(A)*B*C+A*B*C))"),
    .INIT(16'h00d4))
    _al_u6513 (
    .a(_al_u6501_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J2sow6_lutinv ),
    .c(_al_u6511_o),
    .d(_al_u6512_o),
    .o(_al_u6513_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u6514 (
    .a(_al_u6507_o),
    .b(_al_u6508_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E3sow6_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u6515 (
    .a(_al_u6505_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dt1bx6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jj0bx6 ),
    .o(_al_u6515_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u6516 (
    .a(_al_u6509_o),
    .b(_al_u6510_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L3sow6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(B*~(D)*~((~C*~A))+B*D*~((~C*~A))+~(B)*D*(~C*~A)+B*D*(~C*~A))"),
    .INIT(16'hcdc8))
    _al_u6517 (
    .a(_al_u6513_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E3sow6_lutinv ),
    .c(_al_u6515_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L3sow6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ewrow6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(~C*A))"),
    .INIT(16'hf531))
    _al_u6518 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lfgbx6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Slyax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Unyax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wpyax6 ),
    .o(_al_u6518_o));
  AL_MAP_LUT4 #(
    .EQN("(D*A*~(C*~B))"),
    .INIT(16'h8a00))
    _al_u6519 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ot0bx6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Slyax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wpyax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xq2bx6 ),
    .o(_al_u6519_o));
  AL_MAP_LUT4 #(
    .EQN("~(~(C*B)*~(D*A))"),
    .INIT(16'heac0))
    _al_u652 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/read_enable ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_apb_slave_mux/n0 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gpio0_prdata [7]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/read_mux_byte0_reg [7]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_apb_slave_mux/n118 [7]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u6520 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B3gbx6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y0gbx6 ),
    .o(_al_u6520_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B*~A))"),
    .INIT(8'hb0))
    _al_u6521 (
    .a(_al_u6518_o),
    .b(_al_u6519_o),
    .c(_al_u6520_o),
    .o(_al_u6521_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u6522 (
    .a(_al_u6521_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ot0bx6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xq2bx6 ),
    .o(_al_u6522_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u6523 (
    .a(_al_u6521_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Slyax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wpyax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V1sow6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(~C*A))"),
    .INIT(16'hc4f5))
    _al_u6524 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mfyax6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ohyax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qjyax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T3abx6 ),
    .o(_al_u6524_o));
  AL_MAP_LUT4 #(
    .EQN("(C*A*~(D*~B))"),
    .INIT(16'h80a0))
    _al_u6525 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Li2bx6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mfyax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nr0bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qjyax6 ),
    .o(_al_u6525_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u6526 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fe2bx6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mp0bx6 ),
    .o(_al_u6526_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B*~A))"),
    .INIT(8'hb0))
    _al_u6527 (
    .a(_al_u6524_o),
    .b(_al_u6525_o),
    .c(_al_u6526_o),
    .o(_al_u6527_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u6528 (
    .a(_al_u6527_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mfyax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qjyax6 ),
    .o(_al_u6528_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(B*~A))"),
    .INIT(8'h0b))
    _al_u6529 (
    .a(_al_u6519_o),
    .b(_al_u6520_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Unyax6 ),
    .o(_al_u6529_o));
  AL_MAP_LUT4 #(
    .EQN("~(~(C*B)*~(D*A))"),
    .INIT(16'heac0))
    _al_u653 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/read_enable ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_apb_slave_mux/n0 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gpio0_prdata [6]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/read_mux_byte0_reg [6]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_apb_slave_mux/n118 [6]));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*~(B*~A))"),
    .INIT(16'h00b0))
    _al_u6530 (
    .a(_al_u6518_o),
    .b(_al_u6519_o),
    .c(_al_u6520_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lfgbx6 ),
    .o(_al_u6530_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(B*~A))"),
    .INIT(8'h0b))
    _al_u6531 (
    .a(_al_u6525_o),
    .b(_al_u6526_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ohyax6 ),
    .o(_al_u6531_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*~(B*~A))"),
    .INIT(16'h00b0))
    _al_u6532 (
    .a(_al_u6524_o),
    .b(_al_u6525_o),
    .c(_al_u6526_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T3abx6 ),
    .o(_al_u6532_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~(~B*~A))"),
    .INIT(16'h000e))
    _al_u6533 (
    .a(_al_u6529_o),
    .b(_al_u6530_o),
    .c(_al_u6531_o),
    .d(_al_u6532_o),
    .o(_al_u6533_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*(~(B)*C*~(D)+~(B)*~(C)*D+~(B)*C*D+B*C*D))"),
    .INIT(16'h5110))
    _al_u6534 (
    .a(_al_u6522_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V1sow6_lutinv ),
    .c(_al_u6528_o),
    .d(_al_u6533_o),
    .o(_al_u6534_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u6535 (
    .a(_al_u6527_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Li2bx6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nr0bx6 ),
    .o(_al_u6535_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u6536 (
    .a(_al_u6529_o),
    .b(_al_u6530_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D6sow6_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u6537 (
    .a(_al_u6531_o),
    .b(_al_u6532_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z3sow6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((~B*~A))+C*D*~((~B*~A))+~(C)*D*(~B*~A)+C*D*(~B*~A))"),
    .INIT(16'hf1e0))
    _al_u6538 (
    .a(_al_u6534_o),
    .b(_al_u6535_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D6sow6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z3sow6_lutinv ),
    .o(_al_u6538_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((~B*~A))+C*D*~((~B*~A))+~(C)*D*(~B*~A)+C*D*(~B*~A))"),
    .INIT(16'hf1e0))
    _al_u6539 (
    .a(_al_u6513_o),
    .b(_al_u6515_o),
    .c(_al_u6501_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J2sow6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gxrow6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("~(~(C*B)*~(D*A))"),
    .INIT(16'heac0))
    _al_u654 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/read_enable ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_apb_slave_mux/n0 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gpio0_prdata [5]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/read_mux_byte0_reg [5]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_apb_slave_mux/n118 [5]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((~B*~A))+C*D*~((~B*~A))+~(C)*D*(~B*~A)+C*D*(~B*~A))"),
    .INIT(16'hf1e0))
    _al_u6540 (
    .a(_al_u6534_o),
    .b(_al_u6535_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V1sow6_lutinv ),
    .d(_al_u6528_o),
    .o(_al_u6540_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*C)*~(~B*A))"),
    .INIT(16'hdd0d))
    _al_u6541 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ewrow6_lutinv ),
    .b(_al_u6538_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gxrow6_lutinv ),
    .d(_al_u6540_o),
    .o(_al_u6541_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u6542 (
    .a(_al_u6522_o),
    .b(_al_u6535_o),
    .o(_al_u6542_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(B*~A))"),
    .INIT(8'h0b))
    _al_u6543 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gxrow6_lutinv ),
    .b(_al_u6540_o),
    .c(_al_u6542_o),
    .o(_al_u6543_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u6544 (
    .a(_al_u6515_o),
    .b(_al_u6512_o),
    .o(_al_u6544_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(B*~A))"),
    .INIT(8'h0b))
    _al_u6545 (
    .a(_al_u6541_o),
    .b(_al_u6543_o),
    .c(_al_u6544_o),
    .o(_al_u6545_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u6546 (
    .a(_al_u6545_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gxrow6_lutinv ),
    .c(_al_u6540_o),
    .o(_al_u6546_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*~(B*~A))"),
    .INIT(16'h00b0))
    _al_u6547 (
    .a(_al_u6541_o),
    .b(_al_u6543_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ewrow6_lutinv ),
    .d(_al_u6544_o),
    .o(_al_u6547_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(~D*~(B*~A)))"),
    .INIT(16'hf040))
    _al_u6548 (
    .a(_al_u6541_o),
    .b(_al_u6543_o),
    .c(_al_u6538_o),
    .d(_al_u6544_o),
    .o(_al_u6548_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*~A))"),
    .INIT(8'h32))
    _al_u6549 (
    .a(_al_u6493_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rksow6_lutinv ),
    .c(_al_u6494_o),
    .o(_al_u6549_o));
  AL_MAP_LUT4 #(
    .EQN("~(~(C*B)*~(D*A))"),
    .INIT(16'heac0))
    _al_u655 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/read_enable ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_apb_slave_mux/n0 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gpio0_prdata [4]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/read_mux_byte0_reg [4]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_apb_slave_mux/n118 [4]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~(B*~A))"),
    .INIT(16'h000b))
    _al_u6550 (
    .a(_al_u6491_o),
    .b(_al_u6493_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yksow6_lutinv ),
    .d(_al_u6494_o),
    .o(_al_u6550_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*~C)*~(~B*~A))"),
    .INIT(16'heee0))
    _al_u6551 (
    .a(_al_u6547_o),
    .b(_al_u6548_o),
    .c(_al_u6549_o),
    .d(_al_u6550_o),
    .o(_al_u6551_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u6552 (
    .a(_al_u6495_o),
    .b(_al_u6492_o),
    .o(_al_u6552_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(A*B*~(C)+A*~(B)*C+~(A)*B*C+A*B*C))"),
    .INIT(16'h00e8))
    _al_u6553 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gqrow6_lutinv ),
    .b(_al_u6546_o),
    .c(_al_u6551_o),
    .d(_al_u6552_o),
    .o(_al_u6553_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u6554 (
    .a(_al_u6545_o),
    .b(_al_u6542_o),
    .o(_al_u6554_o));
  AL_MAP_LUT4 #(
    .EQN("~(~B*~(D)*~((~C*~A))+~B*D*~((~C*~A))+~(~B)*D*(~C*~A)+~B*D*(~C*~A))"),
    .INIT(16'hc8cd))
    _al_u6555 (
    .a(_al_u6553_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gqrow6_lutinv ),
    .c(_al_u6554_o),
    .d(_al_u6546_o),
    .o(_al_u6555_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(B)*~((~D*~A))+~C*B*~((~D*~A))+~(~C)*B*(~D*~A)+~C*B*(~D*~A))"),
    .INIT(16'h0f4e))
    _al_u6556 (
    .a(_al_u6443_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Irrow6_lutinv ),
    .c(_al_u6436_o),
    .d(_al_u6444_o),
    .o(_al_u6556_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u6557 (
    .a(_al_u6555_o),
    .b(_al_u6556_o),
    .o(_al_u6557_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u6558 (
    .a(_al_u6553_o),
    .b(_al_u6554_o),
    .o(_al_u6558_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u6559 (
    .a(_al_u6549_o),
    .b(_al_u6550_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mtrow6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("~(~(C*B)*~(D*A))"),
    .INIT(16'heac0))
    _al_u656 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/read_enable ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_apb_slave_mux/n0 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gpio0_prdata [3]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/read_mux_byte0_reg [3]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_apb_slave_mux/n118 [3]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0a1f))
    _al_u6560 (
    .a(_al_u6553_o),
    .b(_al_u6554_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mtrow6_lutinv ),
    .d(_al_u6547_o),
    .o(_al_u6560_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u6561 (
    .a(_al_u6437_o),
    .b(_al_u6438_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kctow6_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u6562 (
    .a(_al_u6439_o),
    .b(_al_u6440_o),
    .o(_al_u6562_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(B)*~((~D*~A))+~C*B*~((~D*~A))+~(~C)*B*(~D*~A)+~C*B*(~D*~A))"),
    .INIT(16'h0f4e))
    _al_u6563 (
    .a(_al_u6443_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kctow6_lutinv ),
    .c(_al_u6562_o),
    .d(_al_u6444_o),
    .o(_al_u6563_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*B*~(D*A))"),
    .INIT(16'h040c))
    _al_u6564 (
    .a(_al_u6558_o),
    .b(_al_u6560_o),
    .c(_al_u6563_o),
    .d(_al_u6548_o),
    .o(_al_u6564_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*~B)*~(D*~A))"),
    .INIT(16'ha8fc))
    _al_u6565 (
    .a(_al_u6558_o),
    .b(_al_u6555_o),
    .c(_al_u6556_o),
    .d(_al_u6552_o),
    .o(_al_u6565_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(D*~(~C*~B)))"),
    .INIT(16'h0155))
    _al_u6566 (
    .a(_al_u6446_o),
    .b(_al_u6557_o),
    .c(_al_u6564_o),
    .d(_al_u6565_o),
    .o(_al_u6566_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u6567 (
    .a(_al_u6566_o),
    .b(_al_u6555_o),
    .c(_al_u6556_o),
    .o(_al_u6567_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u6568 (
    .a(_al_u6558_o),
    .b(_al_u6560_o),
    .c(_al_u6548_o),
    .o(_al_u6568_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A))"),
    .INIT(16'he400))
    _al_u6569 (
    .a(_al_u6566_o),
    .b(_al_u6568_o),
    .c(_al_u6563_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wgipw6 ),
    .o(_al_u6569_o));
  AL_MAP_LUT4 #(
    .EQN("~(~(C*B)*~(D*A))"),
    .INIT(16'heac0))
    _al_u657 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/read_enable ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_apb_slave_mux/n0 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gpio0_prdata [2]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/read_mux_byte0_reg [2]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_apb_slave_mux/n118 [2]));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u6570 (
    .a(_al_u6446_o),
    .b(_al_u6558_o),
    .c(_al_u6552_o),
    .o(_al_u6570_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*(~(A)*B*~(D)+~(A)*~(B)*D+~(A)*B*D+A*B*D))"),
    .INIT(16'h0d04))
    _al_u6571 (
    .a(_al_u6567_o),
    .b(_al_u6569_o),
    .c(_al_u6570_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Elnpw6 ),
    .o(_al_u6571_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u6572 (
    .a(_al_u5329_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zdtpw6 ),
    .o(_al_u6572_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u6573 (
    .a(_al_u6571_o),
    .b(_al_u6572_o),
    .o(_al_u6573_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(D)*~((C*~A))+B*D*~((C*~A))+~(B)*D*(C*~A)+B*D*(C*~A))"),
    .INIT(16'hdc8c))
    _al_u6574 (
    .a(_al_u6571_o),
    .b(_al_u6567_o),
    .c(_al_u6572_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Elnpw6 ),
    .o(_al_u6574_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u6575 (
    .a(_al_u6570_o),
    .b(_al_u5329_o),
    .o(_al_u6575_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(~C*~A))"),
    .INIT(16'hfa32))
    _al_u6576 (
    .a(_al_u6573_o),
    .b(_al_u6574_o),
    .c(_al_u6575_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rerow6_lutinv ),
    .o(_al_u6576_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u6577 (
    .a(_al_u6576_o),
    .b(_al_u6574_o),
    .o(_al_u6577_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    _al_u6578 (
    .a(_al_u6336_o),
    .b(_al_u6577_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sbrow6 ),
    .o(_al_u6578_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u6579 (
    .a(_al_u6566_o),
    .b(_al_u6568_o),
    .c(_al_u6563_o),
    .o(_al_u6579_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u658 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n7_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/read_enable ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/mux9_b10_sel_is_3_o ));
  AL_MAP_LUT4 #(
    .EQN("(B*~(D)*~((C*~A))+B*D*~((C*~A))+~(B)*D*(C*~A)+B*D*(C*~A))"),
    .INIT(16'hdc8c))
    _al_u6580 (
    .a(_al_u6571_o),
    .b(_al_u6579_o),
    .c(_al_u6572_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wgipw6 ),
    .o(_al_u6580_o));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    _al_u6581 (
    .a(_al_u6333_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tl4bx6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vpgbx6 ),
    .o(_al_u6581_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*~B)*~(C*~A))"),
    .INIT(16'haf8c))
    _al_u6582 (
    .a(_al_u6574_o),
    .b(_al_u6580_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rerow6_lutinv ),
    .d(_al_u6581_o),
    .o(_al_u6582_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~(B*~A))"),
    .INIT(16'h000b))
    _al_u6583 (
    .a(_al_u6582_o),
    .b(_al_u6576_o),
    .c(_al_u6333_o),
    .d(_al_u6335_o),
    .o(_al_u6583_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(~D*~(B*~A)))"),
    .INIT(16'hf040))
    _al_u6584 (
    .a(_al_u6582_o),
    .b(_al_u6576_o),
    .c(_al_u6580_o),
    .d(_al_u6335_o),
    .o(_al_u6584_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u6585 (
    .a(_al_u6333_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tl4bx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ffrow6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(B*~A)))"),
    .INIT(16'h040f))
    _al_u6586 (
    .a(_al_u6582_o),
    .b(_al_u6576_o),
    .c(_al_u3722_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ffrow6_lutinv ),
    .o(_al_u6586_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~B*~(D*A))"),
    .INIT(16'h1030))
    _al_u6587 (
    .a(_al_u6583_o),
    .b(_al_u6584_o),
    .c(_al_u6586_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vpgbx6 ),
    .o(_al_u6587_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(~C*~(~B*~A)))"),
    .INIT(16'h00f1))
    _al_u6588 (
    .a(_al_u6336_o),
    .b(_al_u6577_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sbrow6 ),
    .d(_al_u3749_o),
    .o(_al_u6588_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*~A))"),
    .INIT(8'h23))
    _al_u6589 (
    .a(_al_u5329_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F17ax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mnmpw6 ),
    .o(_al_u6589_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u659 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/mux9_b10_sel_is_3_o ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [9]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_apb_slave_mux/n117 [9]));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    _al_u6590 (
    .a(_al_u6573_o),
    .b(_al_u6575_o),
    .c(_al_u6589_o),
    .o(_al_u6590_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u6591 (
    .a(_al_u6590_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B0biu6 ),
    .o(_al_u6591_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C*~(B*~A)))"),
    .INIT(16'h4f00))
    _al_u6592 (
    .a(_al_u6578_o),
    .b(_al_u6587_o),
    .c(_al_u6588_o),
    .d(_al_u6591_o),
    .o(_al_u6592_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(~C*~(D*~A)))"),
    .INIT(16'h3130))
    _al_u6593 (
    .a(_al_u1774_o),
    .b(_al_u1791_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pdyax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T8kbx6 ),
    .o(_al_u6593_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~B*~A)*~(D)*~(C)+~(~B*~A)*D*~(C)+~(~(~B*~A))*D*C+~(~B*~A)*D*C)"),
    .INIT(16'hfe0e))
    _al_u6594 (
    .a(_al_u6592_o),
    .b(_al_u6593_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fnnpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Puohu6 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u6595 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cz8iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oy8iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_primask_o ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K7row6_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(~B*A))"),
    .INIT(8'h0d))
    _al_u6596 (
    .a(_al_u6592_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K7row6_lutinv ),
    .c(_al_u6593_o),
    .o(_al_u6596_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*~A))"),
    .INIT(8'h23))
    _al_u6597 (
    .a(_al_u2855_o),
    .b(_al_u1385_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fnnpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J3row6 ));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u6598 (
    .a(_al_u6596_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Usaiu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J3row6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V2row6 ));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(~D*~(B*~A)))"),
    .INIT(16'h0f04))
    _al_u6599 (
    .a(_al_u6582_o),
    .b(_al_u6576_o),
    .c(_al_u6573_o),
    .d(_al_u6335_o),
    .o(_al_u6599_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u660 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/mux9_b10_sel_is_3_o ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [8]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_apb_slave_mux/n117 [8]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u6600 (
    .a(_al_u6599_o),
    .b(_al_u6566_o),
    .o(_al_u6600_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*~B))"),
    .INIT(8'ha8))
    _al_u6601 (
    .a(_al_u6385_o),
    .b(_al_u6372_o),
    .c(_al_u6373_o),
    .o(_al_u6601_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0a1f))
    _al_u6602 (
    .a(_al_u6353_o),
    .b(_al_u6354_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hkgow6 ),
    .d(_al_u6345_o),
    .o(_al_u6602_o));
  AL_MAP_LUT4 #(
    .EQN("~(~B*~((D*~C))*~(A)+~B*(D*~C)*~(A)+~(~B)*(D*~C)*A+~B*(D*~C)*A)"),
    .INIT(16'he4ee))
    _al_u6603 (
    .a(_al_u6385_o),
    .b(_al_u6602_o),
    .c(_al_u6372_o),
    .d(_al_u6365_o),
    .o(_al_u6603_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u6604 (
    .a(_al_u6601_o),
    .b(_al_u6603_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mjgow6 ),
    .o(_al_u6604_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u6605 (
    .a(_al_u6422_o),
    .b(_al_u6423_o),
    .o(_al_u6605_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u6606 (
    .a(_al_u6605_o),
    .b(_al_u6409_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Whgow6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zfgow6_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u6607 (
    .a(_al_u6403_o),
    .b(_al_u6404_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4fow6 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u6608 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4fow6 ),
    .b(_al_u6390_o),
    .c(_al_u6395_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gggow6_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u6609 (
    .a(_al_u6435_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zfgow6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gggow6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lfgow6_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u661 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/mux9_b10_sel_is_3_o ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [19]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_apb_slave_mux/n117 [19]));
  AL_MAP_LUT4 #(
    .EQN("(A*~(~D*~(C)*~(B)+~D*C*~(B)+~(~D)*C*B+~D*C*B))"),
    .INIT(16'h2a08))
    _al_u6610 (
    .a(_al_u6600_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B4fow6 ),
    .c(_al_u6604_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lfgow6_lutinv ),
    .o(_al_u6610_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u6611 (
    .a(_al_u6599_o),
    .b(_al_u6566_o),
    .o(_al_u6611_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u6612 (
    .a(_al_u6583_o),
    .b(_al_u6590_o),
    .o(_al_u6612_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*~B))"),
    .INIT(8'ha8))
    _al_u6613 (
    .a(_al_u6495_o),
    .b(_al_u6482_o),
    .c(_al_u6483_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J8fow6_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u6614 (
    .a(_al_u6463_o),
    .b(_al_u6464_o),
    .o(_al_u6614_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u6615 (
    .a(_al_u6482_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Odgow6 ),
    .o(_al_u6615_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(C)*~(A)+~(~D*B)*C*~(A)+~(~(~D*B))*C*A+~(~D*B)*C*A)"),
    .INIT(16'hf5b1))
    _al_u6616 (
    .a(_al_u6495_o),
    .b(_al_u6614_o),
    .c(_al_u6615_o),
    .d(_al_u6450_o),
    .o(_al_u6616_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u6617 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J8fow6_lutinv ),
    .b(_al_u6616_o),
    .c(_al_u6469_o),
    .o(_al_u6617_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u6618 (
    .a(_al_u6495_o),
    .b(_al_u6614_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C8fow6 ));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u6619 (
    .a(_al_u6617_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C8fow6 ),
    .c(_al_u6455_o),
    .o(_al_u6619_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u662 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/mux9_b10_sel_is_3_o ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [18]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_apb_slave_mux/n117 [18]));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u6620 (
    .a(_al_u6513_o),
    .b(_al_u6515_o),
    .o(_al_u6620_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u6621 (
    .a(_al_u6620_o),
    .b(_al_u6500_o),
    .c(_al_u6505_o),
    .o(_al_u6621_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0a1f))
    _al_u6622 (
    .a(_al_u6534_o),
    .b(_al_u6535_o),
    .c(_al_u6521_o),
    .d(_al_u6527_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pagow6_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(B)*~(A)+~C*B*~(A)+~(~C)*B*A+~C*B*A)"),
    .INIT(8'h72))
    _al_u6623 (
    .a(_al_u6545_o),
    .b(_al_u6621_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pagow6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bagow6_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'h4e))
    _al_u6624 (
    .a(_al_u6558_o),
    .b(_al_u6619_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bagow6_lutinv ),
    .o(_al_u6624_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*~(D*B))"),
    .INIT(16'h1050))
    _al_u6625 (
    .a(_al_u6610_o),
    .b(_al_u6611_o),
    .c(_al_u6612_o),
    .d(_al_u6624_o),
    .o(_al_u6625_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*~A))"),
    .INIT(8'h32))
    _al_u6626 (
    .a(_al_u6625_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pdyax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T8kbx6 ),
    .o(_al_u6626_o));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    _al_u6627 (
    .a(_al_u6626_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xdspw6 ),
    .o(_al_u6627_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u6628 (
    .a(_al_u6596_o),
    .b(_al_u1299_o),
    .o(_al_u6628_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u6629 (
    .a(_al_u6600_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B4fow6 ),
    .o(_al_u6629_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u663 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/mux9_b10_sel_is_3_o ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [17]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_apb_slave_mux/n117 [17]));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u6630 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pdyax6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T8kbx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A0fow6_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u6631 (
    .a(_al_u6590_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A0fow6_lutinv ),
    .o(_al_u6631_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u6632 (
    .a(_al_u6611_o),
    .b(_al_u6631_o),
    .c(_al_u6558_o),
    .o(_al_u6632_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u6633 (
    .a(_al_u6629_o),
    .b(_al_u6632_o),
    .o(_al_u6633_o));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u6634 (
    .a(_al_u6600_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B4fow6 ),
    .c(_al_u6435_o),
    .d(_al_u6385_o),
    .o(_al_u6634_o));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u6635 (
    .a(_al_u6611_o),
    .b(_al_u6558_o),
    .c(_al_u6495_o),
    .d(_al_u6545_o),
    .o(_al_u6635_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D*~(C*~B)))"),
    .INIT(16'h20aa))
    _al_u6636 (
    .a(_al_u6631_o),
    .b(_al_u6582_o),
    .c(_al_u6576_o),
    .d(_al_u6333_o),
    .o(_al_u6636_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    _al_u6637 (
    .a(_al_u6634_o),
    .b(_al_u6635_o),
    .c(_al_u6636_o),
    .o(_al_u6637_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C@B)*~(D@A))"),
    .INIT(16'h8241))
    _al_u6638 (
    .a(_al_u6633_o),
    .b(_al_u6637_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jpmpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xiipw6 ),
    .o(_al_u6638_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u6639 (
    .a(_al_u6558_o),
    .b(_al_u6545_o),
    .o(_al_u6639_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u664 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/mux9_b10_sel_is_3_o ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [16]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_apb_slave_mux/n117 [16]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u6640 (
    .a(_al_u6545_o),
    .b(_al_u6620_o),
    .o(_al_u6640_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*~B)*~(D)*~(A)+~(~C*~B)*D*~(A)+~(~(~C*~B))*D*A+~(~C*~B)*D*A)"),
    .INIT(16'hfe54))
    _al_u6641 (
    .a(_al_u6558_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C8fow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J8fow6_lutinv ),
    .d(_al_u6640_o),
    .o(_al_u6641_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(A*~(~D*~C)))"),
    .INIT(16'h1113))
    _al_u6642 (
    .a(_al_u6639_o),
    .b(_al_u6641_o),
    .c(_al_u6534_o),
    .d(_al_u6535_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q1fow6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u6643 (
    .a(_al_u6611_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q1fow6 ),
    .o(_al_u6643_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u6644 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B4fow6 ),
    .b(_al_u6385_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z2fow6 ));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    _al_u6645 (
    .a(_al_u6435_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4fow6 ),
    .c(_al_u6605_o),
    .o(_al_u6645_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u6646 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B4fow6 ),
    .b(_al_u6601_o),
    .c(_al_u6645_o),
    .o(_al_u6646_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u6647 (
    .a(_al_u6353_o),
    .b(_al_u6354_o),
    .o(_al_u6647_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*A*~(~D*B))"),
    .INIT(16'h0a02))
    _al_u6648 (
    .a(_al_u6600_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z2fow6 ),
    .c(_al_u6646_o),
    .d(_al_u6647_o),
    .o(_al_u6648_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(~C*~B*~A))"),
    .INIT(16'hfe00))
    _al_u6649 (
    .a(_al_u6643_o),
    .b(_al_u6648_o),
    .c(_al_u6590_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A0fow6_lutinv ),
    .o(_al_u6649_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u665 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/mux9_b10_sel_is_3_o ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [15]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_apb_slave_mux/n117 [15]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u6650 (
    .a(_al_u6600_o),
    .b(_al_u6631_o),
    .o(_al_u6650_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(~B*A))"),
    .INIT(8'hd0))
    _al_u6651 (
    .a(_al_u6650_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G2iax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzjpw6 ),
    .o(_al_u6651_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u6652 (
    .a(_al_u6611_o),
    .b(_al_u6631_o),
    .o(_al_u6652_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C@B)*~(D*~A))"),
    .INIT(16'h82c3))
    _al_u6653 (
    .a(_al_u6650_o),
    .b(_al_u6652_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F4iax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G2iax6 ),
    .o(_al_u6653_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u6654 (
    .a(_al_u6649_o),
    .b(_al_u6651_o),
    .c(_al_u6653_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T5mpw6 ),
    .o(_al_u6654_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(D*C*~A))"),
    .INIT(16'h8ccc))
    _al_u6655 (
    .a(_al_u6627_o),
    .b(_al_u6628_o),
    .c(_al_u6638_o),
    .d(_al_u6654_o),
    .o(_al_u6655_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u6656 (
    .a(_al_u6596_o),
    .b(_al_u1777_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ),
    .o(_al_u6656_o));
  AL_MAP_LUT4 #(
    .EQN("~(~A*~(D*C*~B))"),
    .INIT(16'hbaaa))
    _al_u6657 (
    .a(_al_u6655_o),
    .b(_al_u6656_o),
    .c(_al_u1299_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzjpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fivhu6 ));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u6658 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F0eow6 ),
    .b(_al_u5260_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jj0bx6 ),
    .o(_al_u6658_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u6659 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6eiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvgiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Amupw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yjupw6 ),
    .o(_al_u6659_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u666 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/mux9_b10_sel_is_3_o ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [14]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_apb_slave_mux/n117 [14]));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u6660 (
    .a(_al_u6658_o),
    .b(_al_u6659_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M0eow6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dt1bx6 ),
    .o(_al_u6660_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u6661 (
    .a(_al_u6652_o),
    .b(_al_u6660_o),
    .c(_al_u5067_o),
    .o(_al_u6661_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u6662 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xs1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dw1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Erbbx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hpbbx6 ),
    .o(_al_u6662_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u6663 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zt1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ar1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nlbbx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pbbbx6 ),
    .o(_al_u6663_o));
  AL_MAP_LUT4 #(
    .EQN("(C*A*~(D*B))"),
    .INIT(16'h20a0))
    _al_u6664 (
    .a(_al_u6662_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iv1iu6 ),
    .c(_al_u6663_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[16] ),
    .o(_al_u6664_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u6665 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vr1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kw1iu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Btbbx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qjbbx6 ),
    .o(_al_u6665_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u6666 (
    .a(_al_u6664_o),
    .b(_al_u6665_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cs1iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Knbbx6 ),
    .o(_al_u6666_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(~C*~(~B*A)))"),
    .INIT(16'hf200))
    _al_u6667 (
    .a(_al_u927_o),
    .b(_al_u1299_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iv1iu6 ),
    .d(_al_u1385_o),
    .o(_al_u6667_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*A*~(C*~B))"),
    .INIT(16'h008a))
    _al_u6668 (
    .a(_al_u6666_o),
    .b(_al_u1833_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/St1iu6 ),
    .d(_al_u6667_o),
    .o(_al_u6668_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u6669 (
    .a(_al_u5020_o),
    .b(_al_u6661_o),
    .c(_al_u6668_o),
    .o(_al_u6669_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u667 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/mux9_b10_sel_is_3_o ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [13]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_apb_slave_mux/n117 [13]));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u6670 (
    .a(_al_u5049_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sf1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pdbbx6 ),
    .o(_al_u6670_o));
  AL_MAP_LUT4 #(
    .EQN("~(C*~B*~(D*A))"),
    .INIT(16'hefcf))
    _al_u6671 (
    .a(_al_u5053_o),
    .b(_al_u6669_o),
    .c(_al_u6670_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yubbx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Faphu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u6672 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M0eow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F0eow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ih0bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jx1bx6 ),
    .o(_al_u6672_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u6673 (
    .a(_al_u6672_o),
    .b(_al_u3779_o),
    .c(_al_u5260_o),
    .o(_al_u6673_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u6674 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6eiu6 ),
    .b(_al_u405_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T2kbx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ujspw6 ),
    .o(_al_u6674_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u6675 (
    .a(_al_u6673_o),
    .b(_al_u6674_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvgiu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wlspw6 ),
    .o(_al_u6675_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u6676 (
    .a(_al_u6650_o),
    .b(_al_u6675_o),
    .c(_al_u5067_o),
    .o(_al_u6676_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u6677 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xs1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kw1iu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hsdax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ue9ax6 ),
    .o(_al_u6677_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u6678 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vr1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cs1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Owcax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V0cax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mjtiu6 ));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u6679 (
    .a(_al_u6677_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mjtiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iv1iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[15] ),
    .o(_al_u6679_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u668 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/mux9_b10_sel_is_3_o ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [12]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_apb_slave_mux/n117 [12]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u6680 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zt1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ar1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Chwpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kcaax6 ),
    .o(_al_u6680_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u6681 (
    .a(_al_u6679_o),
    .b(_al_u6680_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dw1iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aoeax6 ),
    .o(_al_u6681_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*A*~(C*~B))"),
    .INIT(16'h008a))
    _al_u6682 (
    .a(_al_u6681_o),
    .b(_al_u1868_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/St1iu6 ),
    .d(_al_u6667_o),
    .o(_al_u6682_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u6683 (
    .a(_al_u5020_o),
    .b(_al_u6676_o),
    .c(_al_u6682_o),
    .o(_al_u6683_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u6684 (
    .a(_al_u5049_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sf1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cjwpw6 ),
    .o(_al_u6684_o));
  AL_MAP_LUT4 #(
    .EQN("~(C*~B*~(D*A))"),
    .INIT(16'hefcf))
    _al_u6685 (
    .a(_al_u5053_o),
    .b(_al_u6683_o),
    .c(_al_u6684_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dpwpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Maphu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u6686 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M0eow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F0eow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hf0bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yxrpw6 ),
    .o(_al_u6686_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u6687 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U2fiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E1fiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mb4bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qjyax6 ),
    .o(_al_u6687_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u6688 (
    .a(_al_u6686_o),
    .b(_al_u6687_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvgiu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nbxax6 ),
    .o(_al_u6688_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u6689 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S1fiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G2fiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I45bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L8zax6 ),
    .o(_al_u6689_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u669 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/mux9_b10_sel_is_3_o ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [11]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_apb_slave_mux/n117 [11]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u6690 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I3fiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C0fiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wr4bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yryax6 ),
    .o(_al_u6690_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u6691 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tzdiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q0fiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Az3bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wmzax6 ),
    .o(_al_u6691_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u6692 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6eiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xrgiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F17ax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L9xax6 ),
    .o(_al_u6692_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u6693 (
    .a(_al_u6689_o),
    .b(_al_u6690_o),
    .c(_al_u6691_o),
    .d(_al_u6692_o),
    .o(_al_u6693_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*A)"),
    .INIT(16'h0080))
    _al_u6694 (
    .a(_al_u6688_o),
    .b(_al_u6693_o),
    .c(_al_u5031_o),
    .d(_al_u5260_o),
    .o(_al_u6694_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D*B*~A))"),
    .INIT(16'hb0f0))
    _al_u6695 (
    .a(_al_u6629_o),
    .b(_al_u6632_o),
    .c(_al_u6694_o),
    .d(_al_u5067_o),
    .o(_al_u6695_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u6696 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xs1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vr1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eudax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lycax6 ),
    .o(_al_u6696_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u6697 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dw1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ar1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xpeax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z47ax6 ),
    .o(_al_u6697_o));
  AL_MAP_LUT4 #(
    .EQN("(C*A*~(D*B))"),
    .INIT(16'h20a0))
    _al_u6698 (
    .a(_al_u6696_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iv1iu6 ),
    .c(_al_u6697_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[14] ),
    .o(_al_u6698_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u6699 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cs1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kw1iu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rg9ax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S2cax6 ),
    .o(_al_u6699_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u670 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/mux9_b10_sel_is_3_o ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [10]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_apb_slave_mux/n117 [10]));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u6700 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uvsiu6 ),
    .b(_al_u6699_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zt1iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Heaax6 ),
    .o(_al_u6700_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*~(D*~A))"),
    .INIT(16'h80c0))
    _al_u6701 (
    .a(_al_u4906_o),
    .b(_al_u6698_o),
    .c(_al_u6700_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/St1iu6 ),
    .o(_al_u6701_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u6702 (
    .a(_al_u5020_o),
    .b(_al_u6695_o),
    .c(_al_u6701_o),
    .o(_al_u6702_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u6703 (
    .a(_al_u5050_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sf1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z67ax6 ),
    .o(_al_u6703_o));
  AL_MAP_LUT4 #(
    .EQN("~(C*~B*~(D*A))"),
    .INIT(16'hefcf))
    _al_u6704 (
    .a(_al_u5053_o),
    .b(_al_u6702_o),
    .c(_al_u6703_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ad7ax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Taphu6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u6705 (
    .a(_al_u1781_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Difiu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qaciu6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(B*~(~C*~A)))"),
    .INIT(16'h0037))
    _al_u6706 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uzaiu6 ),
    .b(_al_u1299_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qaciu6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ),
    .o(_al_u6706_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(~D*~(~C*~A)))"),
    .INIT(16'h3301))
    _al_u6707 (
    .a(_al_u6596_o),
    .b(_al_u6706_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bciax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P2vhu6 ));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u6708 (
    .a(_al_u5050_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sf1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sd8ax6 ),
    .o(_al_u6708_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u6709 (
    .a(_al_u5053_o),
    .b(_al_u6708_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvabx6 ),
    .o(_al_u6709_o));
  AL_MAP_LUT4 #(
    .EQN("~(~(C*B)*~(D*A))"),
    .INIT(16'heac0))
    _al_u671 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/read_enable ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_apb_slave_mux/n0 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gpio0_prdata [1]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/read_mux_byte0_reg [1]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_apb_slave_mux/n118 [1]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u6710 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I3fiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvgiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rfxax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vbspw6 ),
    .o(_al_u6710_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u6711 (
    .a(_al_u6710_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q0fiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yw3bx6 ),
    .o(_al_u6711_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u6712 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6eiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U2fiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K94bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pdxax6 ),
    .o(_al_u6712_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u6713 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G2fiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C0fiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G25bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Up4bx6 ),
    .o(_al_u6713_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u6714 (
    .a(_al_u6711_o),
    .b(_al_u6712_o),
    .c(_al_u6713_o),
    .o(_al_u6714_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u6715 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M0eow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F0eow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gd0bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xo1bx6 ),
    .o(_al_u6715_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u6716 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tzdiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E1fiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ohyax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xozax6 ),
    .o(_al_u6716_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u6717 (
    .a(_al_u6715_o),
    .b(_al_u6716_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S1fiu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J6zax6 ),
    .o(_al_u6717_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*A)"),
    .INIT(16'h0080))
    _al_u6718 (
    .a(_al_u6714_o),
    .b(_al_u6717_o),
    .c(_al_u5031_o),
    .d(_al_u5260_o),
    .o(_al_u6718_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u6719 (
    .a(_al_u6637_o),
    .b(_al_u6718_o),
    .c(_al_u5067_o),
    .o(_al_u6719_o));
  AL_MAP_LUT4 #(
    .EQN("~(~(C*B)*~(D*A))"),
    .INIT(16'heac0))
    _al_u672 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/read_enable ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_apb_slave_mux/n0 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gpio0_prdata [0]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/read_mux_byte0_reg [0]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_apb_slave_mux/n118 [0]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u6720 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xs1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cs1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Esabx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Koabx6 ),
    .o(_al_u6720_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u6721 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dw1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zt1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hqabx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nmabx6 ),
    .o(_al_u6721_o));
  AL_MAP_LUT4 #(
    .EQN("(C*A*~(D*B))"),
    .INIT(16'h20a0))
    _al_u6722 (
    .a(_al_u6720_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iv1iu6 ),
    .c(_al_u6721_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[13] ),
    .o(_al_u6722_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u6723 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vr1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kw1iu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Buabx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qkabx6 ),
    .o(_al_u6723_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u6724 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uvsiu6 ),
    .b(_al_u6723_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ar1iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sb8ax6 ),
    .o(_al_u6724_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*~(D*~A))"),
    .INIT(16'h80c0))
    _al_u6725 (
    .a(_al_u4529_o),
    .b(_al_u6722_o),
    .c(_al_u6724_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/St1iu6 ),
    .o(_al_u6725_o));
  AL_MAP_LUT4 #(
    .EQN("~(A*~(C*~(D*B)))"),
    .INIT(16'h75f5))
    _al_u6726 (
    .a(_al_u6709_o),
    .b(_al_u6719_o),
    .c(_al_u5020_o),
    .d(_al_u6725_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Abphu6 ));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u6727 (
    .a(_al_u5050_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sf1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ggabx6 ),
    .o(_al_u6727_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u6728 (
    .a(_al_u5053_o),
    .b(_al_u6727_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kl8ax6 ),
    .o(_al_u6728_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u6729 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M0eow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F0eow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fb0bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rk1bx6 ),
    .o(_al_u6729_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u673 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J3xiu6_lutinv ),
    .b(_al_u533_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hw8ax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kw1iu6_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u6730 (
    .a(_al_u6729_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6eiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R7kpw6 ),
    .o(_al_u6730_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u6731 (
    .a(_al_u6730_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvgiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T9kpw6 ),
    .o(_al_u6731_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*~A))"),
    .INIT(8'h8c))
    _al_u6732 (
    .a(_al_u6649_o),
    .b(_al_u6731_o),
    .c(_al_u5067_o),
    .o(_al_u6732_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u6733 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xs1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vr1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bwdax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I0dax6 ),
    .o(_al_u6733_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u6734 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cs1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ar1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P4cax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xpxax6 ),
    .o(_al_u6734_o));
  AL_MAP_LUT4 #(
    .EQN("(C*A*~(D*B))"),
    .INIT(16'h20a0))
    _al_u6735 (
    .a(_al_u6733_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iv1iu6 ),
    .c(_al_u6734_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[12] ),
    .o(_al_u6735_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u6736 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dw1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kw1iu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oi9ax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ureax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S1tiu6 ));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u6737 (
    .a(_al_u6735_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S1tiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zt1iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Egaax6 ),
    .o(_al_u6737_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*~(D*~A))"),
    .INIT(16'h80c0))
    _al_u6738 (
    .a(_al_u4886_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yw1iu6 ),
    .c(_al_u6737_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/St1iu6 ),
    .o(_al_u6738_o));
  AL_MAP_LUT4 #(
    .EQN("~(A*~(C*~(D*B)))"),
    .INIT(16'h75f5))
    _al_u6739 (
    .a(_al_u6728_o),
    .b(_al_u6732_o),
    .c(_al_u5020_o),
    .d(_al_u6738_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hbphu6 ));
  AL_MAP_LUT2 #(
    .EQN("~(B*A)"),
    .INIT(4'h7))
    _al_u674 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kw1iu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dg2qw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zg7iu6 ));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u6740 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J0iax6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6lax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 ),
    .o(_al_u6740_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    _al_u6741 (
    .a(_al_u4169_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qqhiu6 ),
    .c(_al_u6740_o),
    .o(_al_u6741_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u6742 (
    .a(_al_u6741_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzjpw6 ),
    .o(_al_u6742_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u6743 (
    .a(_al_u6628_o),
    .b(_al_u6742_o),
    .o(_al_u6743_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u6744 (
    .a(_al_u6743_o),
    .b(_al_u4533_o),
    .o(_al_u6744_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u6745 (
    .a(_al_u6628_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzjpw6 ),
    .o(_al_u6745_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u6746 (
    .a(_al_u6745_o),
    .b(_al_u6741_o),
    .o(_al_u6746_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u6747 (
    .a(_al_u6744_o),
    .b(_al_u6746_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L4lax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wfphu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*B)*~(~D*A))"),
    .INIT(16'hf351))
    _al_u6748 (
    .a(_al_u6746_o),
    .b(_al_u6743_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sn7iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W8hbx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yhvhu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*B*A))"),
    .INIT(16'h070f))
    _al_u6749 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R05iu6 ),
    .b(_al_u4170_o),
    .c(_al_u6741_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X7ypw6 ),
    .o(_al_u6749_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u675 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bciax6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/SLEEPHOLDACKn ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u6750 (
    .a(_al_u6745_o),
    .b(_al_u6749_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L0vhu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u6751 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vr1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ar1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dm6bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F2dax6 ),
    .o(_al_u6751_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u6752 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cs1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zt1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Biaax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6cax6 ),
    .o(_al_u6752_o));
  AL_MAP_LUT4 #(
    .EQN("(C*A*~(D*B))"),
    .INIT(16'h20a0))
    _al_u6753 (
    .a(_al_u6751_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iv1iu6 ),
    .c(_al_u6752_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[11] ),
    .o(_al_u6753_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u6754 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dw1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kw1iu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lk9ax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rteax6 ),
    .o(_al_u6754_o));
  AL_MAP_LUT4 #(
    .EQN("(C*A*~(D*B))"),
    .INIT(16'h20a0))
    _al_u6755 (
    .a(_al_u6753_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xs1iu6 ),
    .c(_al_u6754_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yxdax6 ),
    .o(_al_u6755_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*~(D*~A))"),
    .INIT(16'h80c0))
    _al_u6756 (
    .a(_al_u4816_o),
    .b(_al_u6755_o),
    .c(_al_u5044_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/St1iu6 ),
    .o(_al_u6756_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u6757 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F0eow6 ),
    .b(_al_u5260_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E90bx6 ),
    .o(_al_u6757_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u6758 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6eiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvgiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tyipw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V0jpw6 ),
    .o(_al_u6758_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u6759 (
    .a(_al_u6757_o),
    .b(_al_u6758_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M0eow6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z71bx6 ),
    .o(_al_u6759_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u676 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I6row6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(C*B*~(D*A))"),
    .INIT(16'h40c0))
    _al_u6760 (
    .a(_al_u6626_o),
    .b(_al_u6756_o),
    .c(_al_u6759_o),
    .d(_al_u5067_o),
    .o(_al_u6760_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u6761 (
    .a(_al_u5050_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sf1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ro8ax6 ),
    .o(_al_u6761_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u6762 (
    .a(_al_u5053_o),
    .b(_al_u6761_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Su8ax6 ),
    .o(_al_u6762_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C*~A))"),
    .INIT(8'h73))
    _al_u6763 (
    .a(_al_u6760_o),
    .b(_al_u6762_o),
    .c(_al_u5020_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Obphu6 ));
  AL_MAP_LUT4 #(
    .EQN("~(~(~C*B)*~(D*A))"),
    .INIT(16'hae0c))
    _al_u6764 (
    .a(_al_u6746_o),
    .b(_al_u6743_o),
    .c(_al_u4530_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E6iax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H5vhu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~C)*~(B)*~(A)+~(D*~C)*B*~(A)+~(~(D*~C))*B*A+~(D*~C)*B*A)"),
    .INIT(16'hd8dd))
    _al_u6765 (
    .a(_al_u6628_o),
    .b(_al_u6649_o),
    .c(_al_u6742_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T5mpw6 ),
    .o(_al_u6765_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(~C*A))"),
    .INIT(8'h3b))
    _al_u6766 (
    .a(_al_u6744_o),
    .b(_al_u6765_o),
    .c(_al_u4581_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z0vhu6 ));
  AL_MAP_LUT4 #(
    .EQN("~((D*~C)*~(B)*~(A)+(D*~C)*B*~(A)+~((D*~C))*B*A+(D*~C)*B*A)"),
    .INIT(16'h7277))
    _al_u6767 (
    .a(_al_u6628_o),
    .b(_al_u6637_o),
    .c(_al_u6742_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jpmpw6 ),
    .o(_al_u6767_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(~C*A))"),
    .INIT(8'h3b))
    _al_u6768 (
    .a(_al_u6744_o),
    .b(_al_u6767_o),
    .c(_al_u4611_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N1vhu6 ));
  AL_MAP_LUT4 #(
    .EQN("~((D*~C)*~(B)*~(A)+(D*~C)*B*~(A)+~((D*~C))*B*A+(D*~C)*B*A)"),
    .INIT(16'h7277))
    _al_u6769 (
    .a(_al_u6628_o),
    .b(_al_u6633_o),
    .c(_al_u6742_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xiipw6 ),
    .o(_al_u6769_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u677 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I6row6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vygax6 ),
    .o(_al_u677_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(~C*A))"),
    .INIT(8'h3b))
    _al_u6770 (
    .a(_al_u6744_o),
    .b(_al_u6769_o),
    .c(_al_u4637_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U1vhu6 ));
  AL_MAP_LUT4 #(
    .EQN("~((D*~C)*~(B)*~(A)+(D*~C)*B*~(A)+~((D*~C))*B*A+(D*~C)*B*A)"),
    .INIT(16'h7277))
    _al_u6771 (
    .a(_al_u6628_o),
    .b(_al_u6650_o),
    .c(_al_u6742_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G2iax6 ),
    .o(_al_u6771_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(~C*A))"),
    .INIT(8'h3b))
    _al_u6772 (
    .a(_al_u6744_o),
    .b(_al_u6771_o),
    .c(_al_u4663_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B2vhu6 ));
  AL_MAP_LUT4 #(
    .EQN("~((D*~C)*~(B)*~(A)+(D*~C)*B*~(A)+~((D*~C))*B*A+(D*~C)*B*A)"),
    .INIT(16'h7277))
    _al_u6773 (
    .a(_al_u6628_o),
    .b(_al_u6652_o),
    .c(_al_u6742_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F4iax6 ),
    .o(_al_u6773_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(~C*A))"),
    .INIT(8'h3b))
    _al_u6774 (
    .a(_al_u6744_o),
    .b(_al_u6773_o),
    .c(_al_u4688_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I2vhu6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u6775 (
    .a(_al_u6655_o),
    .b(_al_u6745_o),
    .o(_al_u6775_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(~C*A))"),
    .INIT(16'h31f5))
    _al_u6776 (
    .a(_al_u6744_o),
    .b(_al_u6746_o),
    .c(_al_u4712_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E8iax6 ),
    .o(_al_u6776_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C*A))"),
    .INIT(8'hb3))
    _al_u6777 (
    .a(_al_u6775_o),
    .b(_al_u6776_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xlfpw6 [1]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D3vhu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(~C*A))"),
    .INIT(16'h31f5))
    _al_u6778 (
    .a(_al_u6744_o),
    .b(_al_u6746_o),
    .c(_al_u4735_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zqiax6 ),
    .o(_al_u6778_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C*A))"),
    .INIT(8'hb3))
    _al_u6779 (
    .a(_al_u6775_o),
    .b(_al_u6778_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xlfpw6 [2]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K3vhu6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u678 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 ),
    .o(_al_u678_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(~C*A))"),
    .INIT(16'h31f5))
    _al_u6780 (
    .a(_al_u6744_o),
    .b(_al_u6746_o),
    .c(_al_u4836_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ysiax6 ),
    .o(_al_u6780_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C*A))"),
    .INIT(8'hb3))
    _al_u6781 (
    .a(_al_u6775_o),
    .b(_al_u6780_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xlfpw6 [3]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vhu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(~C*A))"),
    .INIT(16'h31f5))
    _al_u6782 (
    .a(_al_u6744_o),
    .b(_al_u6746_o),
    .c(_al_u4756_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuiax6 ),
    .o(_al_u6782_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C*A))"),
    .INIT(8'hb3))
    _al_u6783 (
    .a(_al_u6775_o),
    .b(_al_u6782_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xlfpw6 [4]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y3vhu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(~C*A))"),
    .INIT(16'h31f5))
    _al_u6784 (
    .a(_al_u6744_o),
    .b(_al_u6746_o),
    .c(_al_u4776_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wwiax6 ),
    .o(_al_u6784_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C*A))"),
    .INIT(8'hb3))
    _al_u6785 (
    .a(_al_u6775_o),
    .b(_al_u6784_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xlfpw6 [5]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F4vhu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(~C*A))"),
    .INIT(16'h31f5))
    _al_u6786 (
    .a(_al_u6744_o),
    .b(_al_u6746_o),
    .c(_al_u4796_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wyiax6 ),
    .o(_al_u6786_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C*A))"),
    .INIT(8'hb3))
    _al_u6787 (
    .a(_al_u6775_o),
    .b(_al_u6786_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xlfpw6 [6]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M4vhu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(~C*A))"),
    .INIT(16'h31f5))
    _al_u6788 (
    .a(_al_u6744_o),
    .b(_al_u6746_o),
    .c(_al_u4816_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W0jax6 ),
    .o(_al_u6788_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C*A))"),
    .INIT(8'hb3))
    _al_u6789 (
    .a(_al_u6775_o),
    .b(_al_u6788_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xlfpw6 [7]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T4vhu6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u679 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ),
    .o(_al_u679_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(~C*A))"),
    .INIT(16'h31f5))
    _al_u6790 (
    .a(_al_u6744_o),
    .b(_al_u6746_o),
    .c(_al_u4886_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W2jax6 ),
    .o(_al_u6790_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C*A))"),
    .INIT(8'hb3))
    _al_u6791 (
    .a(_al_u6775_o),
    .b(_al_u6790_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xlfpw6 [8]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A5vhu6 ));
  AL_MAP_LUT4 #(
    .EQN("~((D*~C)*~(B)*~(A)+(D*~C)*B*~(A)+~((D*~C))*B*A+(D*~C)*B*A)"),
    .INIT(16'h7277))
    _al_u6792 (
    .a(_al_u6628_o),
    .b(_al_u6626_o),
    .c(_al_u6742_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xdspw6 ),
    .o(_al_u6792_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(~C*A))"),
    .INIT(8'h3b))
    _al_u6793 (
    .a(_al_u6744_o),
    .b(_al_u6792_o),
    .c(_al_u4865_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O5vhu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u6794 (
    .a(_al_u5053_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sf1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F8dbx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H7hbx6 ),
    .o(_al_u6794_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(~C*~(~B*A)))"),
    .INIT(16'hf200))
    _al_u6795 (
    .a(_al_u6592_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K7row6_lutinv ),
    .c(_al_u6593_o),
    .d(_al_u5067_o),
    .o(_al_u6795_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(~C*A))"),
    .INIT(16'h31f5))
    _al_u6796 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/St1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iv1iu6 ),
    .c(_al_u1848_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[22] ),
    .o(_al_u6796_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u6797 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dw1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zt1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q1hbx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wxgbx6 ),
    .o(_al_u6797_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u6798 (
    .a(_al_u6797_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ar1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztgbx6 ),
    .o(_al_u6798_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u6799 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xs1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vr1iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K5hbx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N3hbx6 ),
    .o(_al_u6799_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u680 (
    .a(_al_u677_o),
    .b(_al_u678_o),
    .c(_al_u679_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 ),
    .o(_al_u680_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u6800 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cs1iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kw1iu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tzgbx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zvgbx6 ),
    .o(_al_u6800_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u6801 (
    .a(_al_u6796_o),
    .b(_al_u6798_o),
    .c(_al_u6799_o),
    .d(_al_u6800_o),
    .o(_al_u6801_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u6802 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yw1iu6 ),
    .b(_al_u6801_o),
    .o(_al_u6802_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u6803 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M0eow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F0eow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ot0bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xq2bx6 ),
    .o(_al_u6803_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u6804 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U2fiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G2fiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K65bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Od4bx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Smnow6 ));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u6805 (
    .a(_al_u6803_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Smnow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C0fiu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yt4bx6 ),
    .o(_al_u6805_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u6806 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hqgiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q0fiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C14bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gz6ax6 ),
    .o(_al_u6806_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u6807 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tzdiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvgiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Coupw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vkzax6 ),
    .o(_al_u6807_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u6808 (
    .a(_al_u6805_o),
    .b(_al_u6806_o),
    .c(_al_u6807_o),
    .o(_al_u6808_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u6809 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6eiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I3fiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Auyax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J7xax6 ),
    .o(_al_u6809_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u681 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 ),
    .o(_al_u681_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u6810 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S1fiu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E1fiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nazax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Slyax6 ),
    .o(_al_u6810_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u6811 (
    .a(_al_u6808_o),
    .b(_al_u6809_o),
    .c(_al_u6810_o),
    .o(_al_u6811_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D*C*~B))"),
    .INIT(16'h8aaa))
    _al_u6812 (
    .a(_al_u5020_o),
    .b(_al_u6795_o),
    .c(_al_u6802_o),
    .d(_al_u6811_o),
    .o(_al_u6812_o));
  AL_MAP_LUT2 #(
    .EQN("~(~B*A)"),
    .INIT(4'hd))
    _al_u6813 (
    .a(_al_u6794_o),
    .b(_al_u6812_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P8phu6 ));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(B*A))"),
    .INIT(8'h07))
    _al_u6814 (
    .a(_al_u1658_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ldiow6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 ),
    .o(_al_u6814_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C*~B*~A))"),
    .INIT(16'hef00))
    _al_u6815 (
    .a(_al_u677_o),
    .b(_al_u3115_o),
    .c(_al_u6814_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fpnpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hemow6_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u6816 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hemow6_lutinv ),
    .b(_al_u5001_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q2eow6 ));
  AL_MAP_LUT4 #(
    .EQN("(C*~(~B*~(D*~A)))"),
    .INIT(16'hd0c0))
    _al_u6817 (
    .a(_al_u3103_o),
    .b(_al_u1329_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fpnpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 ),
    .o(_al_u6817_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(C*~A))"),
    .INIT(16'haf23))
    _al_u6818 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ha3ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q2eow6 ),
    .c(_al_u6817_o),
    .d(_al_u1848_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mjnow6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u6819 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hemow6_lutinv ),
    .b(_al_u5001_o),
    .o(_al_u6819_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u682 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 ),
    .o(_al_u682_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(D*~(C*~A)))"),
    .INIT(16'h40cc))
    _al_u6820 (
    .a(_al_u6795_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mjnow6 ),
    .c(_al_u6811_o),
    .d(_al_u6819_o),
    .o(_al_u6820_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*C)*~(B*~A))"),
    .INIT(16'hbb0b))
    _al_u6821 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rw1iu6 ),
    .b(_al_u6819_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q2eow6 ),
    .d(_al_u1865_o),
    .o(_al_u6821_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*~A))"),
    .INIT(8'h8c))
    _al_u6822 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mg3ju6_lutinv ),
    .b(_al_u6821_o),
    .c(_al_u6817_o),
    .o(_al_u6822_o));
  AL_MAP_LUT4 #(
    .EQN("~((C*~B)*~(A)*~(D)+(C*~B)*A*~(D)+~((C*~B))*A*D+(C*~B)*A*D)"),
    .INIT(16'h55cf))
    _al_u6823 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ldiow6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S4kbx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 ),
    .o(_al_u6823_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u6824 (
    .a(_al_u6822_o),
    .b(_al_u6823_o),
    .o(_al_u6824_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u6825 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qyniu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S4kbx6 ),
    .o(_al_u6825_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(~B*~(C*~A)))"),
    .INIT(16'hdc00))
    _al_u6826 (
    .a(_al_u6820_o),
    .b(_al_u6824_o),
    .c(_al_u6825_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ms5bx6 ),
    .o(_al_u6826_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u6827 (
    .a(_al_u6695_o),
    .b(_al_u6819_o),
    .o(_al_u6827_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*~B)*~(D*~A))"),
    .INIT(16'h8acf))
    _al_u6828 (
    .a(_al_u4735_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pxriu6 ),
    .c(_al_u6819_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q2eow6 ),
    .o(_al_u6828_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u6829 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jb3ju6_lutinv ),
    .b(_al_u6828_o),
    .c(_al_u6817_o),
    .o(_al_u6829_o));
  AL_MAP_LUT4 #(
    .EQN("~(~A*~(D*C*B))"),
    .INIT(16'heaaa))
    _al_u683 (
    .a(_al_u680_o),
    .b(_al_u681_o),
    .c(_al_u682_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mihow6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u6830 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hemow6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V3xhu6 ),
    .o(_al_u6830_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u6831 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ms5bx6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S4kbx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qdhow6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0cdd))
    _al_u6832 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qdhow6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 ),
    .o(_al_u6832_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~B*~(~D*~A))"),
    .INIT(16'h0302))
    _al_u6833 (
    .a(_al_u6829_o),
    .b(_al_u6021_o),
    .c(_al_u6830_o),
    .d(_al_u6832_o),
    .o(_al_u6833_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*~B)*~(D*A))"),
    .INIT(16'h45cf))
    _al_u6834 (
    .a(_al_u6087_o),
    .b(_al_u4906_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q2eow6 ),
    .d(_al_u6817_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iimow6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(~C*~A))"),
    .INIT(16'h32fa))
    _al_u6835 (
    .a(_al_u6823_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S2ziu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ms5bx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bimow6 ));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~D*~(C*~A)))"),
    .INIT(16'hcc40))
    _al_u6836 (
    .a(_al_u6827_o),
    .b(_al_u6833_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iimow6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bimow6 ),
    .o(_al_u6836_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(~B*~A)))"),
    .INIT(16'h010f))
    _al_u6837 (
    .a(_al_u1269_o),
    .b(_al_u2868_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tucow6_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u6838 (
    .a(_al_u1887_o),
    .b(_al_u698_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D31ju6 ),
    .o(_al_u6838_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(A)*~(C)+~(D*~B)*A*~(C)+~(~(D*~B))*A*C+~(D*~B)*A*C)"),
    .INIT(16'hacaf))
    _al_u6839 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oh3ju6 ),
    .b(_al_u6830_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tucow6_lutinv ),
    .d(_al_u6838_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wxlow6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u684 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_f [0]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_f [1]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_f [2]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_f [3]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n40_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u6840 (
    .a(_al_u6219_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tucow6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hvcow6_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u6841 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hvcow6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3how6_lutinv ),
    .o(_al_u6841_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u6842 (
    .a(_al_u6129_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tucow6_lutinv ),
    .o(_al_u6842_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u6843 (
    .a(_al_u6841_o),
    .b(_al_u6842_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pxlow6 ));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~(B*~A))"),
    .INIT(16'hb000))
    _al_u6844 (
    .a(_al_u6826_o),
    .b(_al_u6836_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wxlow6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pxlow6 ),
    .o(_al_u6844_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*B)*~(D*A))"),
    .INIT(16'h51f3))
    _al_u6845 (
    .a(_al_u6104_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q2eow6 ),
    .c(_al_u1868_o),
    .d(_al_u6817_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J9eow6 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*~A))"),
    .INIT(8'h8c))
    _al_u6846 (
    .a(_al_u6676_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J9eow6 ),
    .c(_al_u6819_o),
    .o(_al_u6846_o));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'h47))
    _al_u6847 (
    .a(_al_u6047_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tucow6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vo3ju6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vacow6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u6848 (
    .a(_al_u6049_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tucow6_lutinv ),
    .o(_al_u6848_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*~B))"),
    .INIT(8'ha8))
    _al_u6849 (
    .a(_al_u6848_o),
    .b(_al_u604_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xbcow6_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(B*A))"),
    .INIT(8'h07))
    _al_u685 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reload_i ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n40_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/baud_updated ),
    .o(_al_u685_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*~B)*~(D*~A))"),
    .INIT(16'h8acf))
    _al_u6850 (
    .a(_al_u4836_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4siu6 ),
    .c(_al_u6819_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q2eow6 ),
    .o(_al_u6850_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u6851 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gk3ju6_lutinv ),
    .b(_al_u6850_o),
    .c(_al_u6817_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rcliu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*~B)*~(D*~A))"),
    .INIT(16'h8acf))
    _al_u6852 (
    .a(_al_u4865_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M1xiu6 ),
    .c(_al_u6819_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q2eow6 ),
    .o(_al_u6852_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u6853 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lj3ju6_lutinv ),
    .b(_al_u6852_o),
    .c(_al_u6817_o),
    .o(_al_u6853_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(~C*~A))"),
    .INIT(16'hfa32))
    _al_u6854 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vacow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xbcow6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rcliu6 ),
    .d(_al_u6853_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ogdow6 ));
  AL_MAP_LUT4 #(
    .EQN("(B*~(A*~(D)*~(C)+A*D*~(C)+~(A)*D*C+A*D*C))"),
    .INIT(16'h04c4))
    _al_u6855 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P8viu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hemow6_lutinv ),
    .c(_al_u5001_o),
    .d(_al_u1850_o),
    .o(_al_u6855_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*~A))"),
    .INIT(8'h23))
    _al_u6856 (
    .a(_al_u6036_o),
    .b(_al_u6855_o),
    .c(_al_u6817_o),
    .o(_al_u6856_o));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'h47))
    _al_u6857 (
    .a(_al_u6129_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tucow6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vxniu6_lutinv ),
    .o(_al_u6857_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*~B))"),
    .INIT(8'ha8))
    _al_u6858 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ogdow6 ),
    .b(_al_u6856_o),
    .c(_al_u6857_o),
    .o(_al_u6858_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(D*C*~B))"),
    .INIT(16'h4555))
    _al_u6859 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tucow6_lutinv ),
    .b(_al_u2647_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 ),
    .o(_al_u6859_o));
  AL_MAP_LUT2 #(
    .EQN("~(~B*A)"),
    .INIT(4'hd))
    _al_u686 (
    .a(_al_u685_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n43 [3]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_baud_cntr_f [3]));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u6860 (
    .a(_al_u6841_o),
    .b(_al_u6859_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eccow6 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    _al_u6861 (
    .a(_al_u6846_o),
    .b(_al_u6858_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eccow6 ),
    .o(_al_u6861_o));
  AL_MAP_LUT3 #(
    .EQN("~(C*B*~A)"),
    .INIT(8'hbf))
    _al_u6862 (
    .a(_al_u6844_o),
    .b(_al_u6861_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vdmiu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Admiu6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u6863 (
    .a(_al_u5998_o),
    .b(_al_u6817_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qtfow6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*C)*~(B*~A))"),
    .INIT(16'hbb0b))
    _al_u6864 (
    .a(_al_u6057_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qtfow6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q2eow6 ),
    .d(_al_u1833_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z4kow6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u6865 (
    .a(_al_u5998_o),
    .b(_al_u6817_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dyeow6_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*~B))"),
    .INIT(8'h8a))
    _al_u6866 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z4kow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F14ju6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dyeow6_lutinv ),
    .o(_al_u6866_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*~A))"),
    .INIT(8'h8c))
    _al_u6867 (
    .a(_al_u6661_o),
    .b(_al_u6866_o),
    .c(_al_u6819_o),
    .o(_al_u6867_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(~A*~(C*B)))"),
    .INIT(16'hea00))
    _al_u6868 (
    .a(_al_u6171_o),
    .b(_al_u6170_o),
    .c(_al_u6021_o),
    .d(_al_u6817_o),
    .o(_al_u6868_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(A*~(D)*~(C)+A*D*~(C)+~(A)*D*C+A*D*C))"),
    .INIT(16'h04c4))
    _al_u6869 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wfviu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hemow6_lutinv ),
    .c(_al_u5001_o),
    .d(_al_u1852_o),
    .o(_al_u6869_o));
  AL_MAP_LUT2 #(
    .EQN("~(~B*A)"),
    .INIT(4'hd))
    _al_u687 (
    .a(_al_u685_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n43 [2]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_baud_cntr_f [2]));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u6870 (
    .a(_al_u6868_o),
    .b(_al_u6869_o),
    .o(_al_u6870_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*~B)*~(D*~A))"),
    .INIT(16'h8acf))
    _al_u6871 (
    .a(_al_u4756_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ibsiu6 ),
    .c(_al_u6819_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q2eow6 ),
    .o(_al_u6871_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*~B))"),
    .INIT(8'h8a))
    _al_u6872 (
    .a(_al_u6871_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uc4ju6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dyeow6_lutinv ),
    .o(_al_u6872_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*~B))"),
    .INIT(8'h8a))
    _al_u6873 (
    .a(_al_u6872_o),
    .b(_al_u6071_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qtfow6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xv6ow6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*~B)*~(D*~A))"),
    .INIT(16'h8acf))
    _al_u6874 (
    .a(_al_u4581_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ovpiu6 ),
    .c(_al_u6819_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q2eow6 ),
    .o(_al_u6874_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*~B))"),
    .INIT(8'h8a))
    _al_u6875 (
    .a(_al_u6874_o),
    .b(_al_u6151_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qtfow6_lutinv ),
    .o(_al_u6875_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*~B))"),
    .INIT(8'h8a))
    _al_u6876 (
    .a(_al_u6875_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mu3ju6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dyeow6_lutinv ),
    .o(_al_u6876_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(~C*~A))"),
    .INIT(16'hfa32))
    _al_u6877 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vacow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xbcow6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xv6ow6 ),
    .d(_al_u6876_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bddow6 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    _al_u6878 (
    .a(_al_u6870_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bddow6 ),
    .c(_al_u6857_o),
    .o(_al_u6878_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    _al_u6879 (
    .a(_al_u6867_o),
    .b(_al_u6878_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eccow6 ),
    .o(_al_u6879_o));
  AL_MAP_LUT2 #(
    .EQN("~(~B*A)"),
    .INIT(4'hd))
    _al_u688 (
    .a(_al_u685_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n43 [1]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_baud_cntr_f [1]));
  AL_MAP_LUT3 #(
    .EQN("~(C*B*~A)"),
    .INIT(8'hbf))
    _al_u6880 (
    .a(_al_u6844_o),
    .b(_al_u6879_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wamiu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bamiu6 ));
  AL_MAP_LUT4 #(
    .EQN("(D*~(~A*~(C*B)))"),
    .INIT(16'hea00))
    _al_u6881 (
    .a(_al_u6167_o),
    .b(_al_u6166_o),
    .c(_al_u6021_o),
    .d(_al_u6817_o),
    .o(_al_u6881_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(A*~(D)*~(C)+A*D*~(C)+~(A)*D*C+A*D*C))"),
    .INIT(16'h04c4))
    _al_u6882 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wmviu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hemow6_lutinv ),
    .c(_al_u5001_o),
    .d(_al_u1854_o),
    .o(_al_u6882_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u6883 (
    .a(_al_u6881_o),
    .b(_al_u6882_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ukcow6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*~B)*~(D*~A))"),
    .INIT(16'h8acf))
    _al_u6884 (
    .a(_al_u4776_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bisiu6 ),
    .c(_al_u6819_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q2eow6 ),
    .o(_al_u6884_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*~B))"),
    .INIT(8'h8a))
    _al_u6885 (
    .a(_al_u6884_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Id4ju6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dyeow6_lutinv ),
    .o(_al_u6885_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*~B))"),
    .INIT(8'h8a))
    _al_u6886 (
    .a(_al_u6885_o),
    .b(_al_u6068_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qtfow6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Plcow6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(C*~A))"),
    .INIT(16'haf23))
    _al_u6887 (
    .a(_al_u4611_o),
    .b(_al_u6819_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q2eow6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jaqiu6 ),
    .o(_al_u6887_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*~B))"),
    .INIT(8'h8a))
    _al_u6888 (
    .a(_al_u6887_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yt3ju6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dyeow6_lutinv ),
    .o(_al_u6888_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*~B))"),
    .INIT(8'h8a))
    _al_u6889 (
    .a(_al_u6888_o),
    .b(_al_u6010_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qtfow6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gkcow6 ));
  AL_MAP_LUT2 #(
    .EQN("~(~B*A)"),
    .INIT(4'hd))
    _al_u689 (
    .a(_al_u685_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n43 [0]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_baud_cntr_f [0]));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(~C*~A))"),
    .INIT(16'hfa32))
    _al_u6890 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vacow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xbcow6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Plcow6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gkcow6 ),
    .o(_al_u6890_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*C)*~(B*~A))"),
    .INIT(16'hbb0b))
    _al_u6891 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U1uiu6 ),
    .b(_al_u6819_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q2eow6 ),
    .d(_al_u1836_o),
    .o(_al_u6891_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B*~A))"),
    .INIT(8'hb0))
    _al_u6892 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R04ju6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dyeow6_lutinv ),
    .c(_al_u6891_o),
    .o(_al_u6892_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*~B))"),
    .INIT(8'h8a))
    _al_u6893 (
    .a(_al_u6892_o),
    .b(_al_u6054_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qtfow6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wlcow6 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    _al_u6894 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eccow6 ),
    .b(_al_u6890_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wlcow6 ),
    .o(_al_u6894_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    _al_u6895 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ukcow6 ),
    .b(_al_u6894_o),
    .c(_al_u6857_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q7miu6 ));
  AL_MAP_LUT3 #(
    .EQN("~(C*B*~A)"),
    .INIT(8'hbf))
    _al_u6896 (
    .a(_al_u6844_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q7miu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X7miu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C7miu6 ));
  AL_MAP_LUT4 #(
    .EQN("(D*~(~A*~(C*B)))"),
    .INIT(16'hea00))
    _al_u6897 (
    .a(_al_u6169_o),
    .b(_al_u6168_o),
    .c(_al_u6021_o),
    .d(_al_u6817_o),
    .o(_al_u6897_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(A*~(D)*~(C)+A*D*~(C)+~(A)*D*C+A*D*C))"),
    .INIT(16'h04c4))
    _al_u6898 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wtviu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hemow6_lutinv ),
    .c(_al_u5001_o),
    .d(_al_u1856_o),
    .o(_al_u6898_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u6899 (
    .a(_al_u6897_o),
    .b(_al_u6898_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yfcow6 ));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u690 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_apb_slave_mux/n0 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/apb_tran_end ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PWRITE ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*~B)*~(D*~A))"),
    .INIT(16'h8acf))
    _al_u6900 (
    .a(_al_u4796_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uosiu6 ),
    .c(_al_u6819_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q2eow6 ),
    .o(_al_u6900_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*~B))"),
    .INIT(8'h8a))
    _al_u6901 (
    .a(_al_u6900_o),
    .b(_al_u6064_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dyeow6_lutinv ),
    .o(_al_u6901_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*~B))"),
    .INIT(8'h8a))
    _al_u6902 (
    .a(_al_u6901_o),
    .b(_al_u6075_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qtfow6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgcow6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*~B)*~(D*~A))"),
    .INIT(16'h8acf))
    _al_u6903 (
    .a(_al_u4637_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tmqiu6 ),
    .c(_al_u6819_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q2eow6 ),
    .o(_al_u6903_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B*~A))"),
    .INIT(8'hb0))
    _al_u6904 (
    .a(_al_u6139_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dyeow6_lutinv ),
    .c(_al_u6903_o),
    .o(_al_u6904_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*~B))"),
    .INIT(8'h8a))
    _al_u6905 (
    .a(_al_u6904_o),
    .b(_al_u6018_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qtfow6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kfcow6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(~C*~A))"),
    .INIT(16'hfa32))
    _al_u6906 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vacow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xbcow6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgcow6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kfcow6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B6dow6 ));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'h5030))
    _al_u6907 (
    .a(_al_u1839_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U8uiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hemow6_lutinv ),
    .d(_al_u5001_o),
    .o(_al_u6907_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(B*~A))"),
    .INIT(8'h0b))
    _al_u6908 (
    .a(_al_u6086_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qtfow6_lutinv ),
    .c(_al_u6907_o),
    .o(_al_u6908_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*~B))"),
    .INIT(8'h8a))
    _al_u6909 (
    .a(_al_u6908_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C34ju6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dyeow6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahcow6 ));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u691 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n6 ),
    .b(_al_u467_o),
    .c(_al_u472_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n40 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    _al_u6910 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eccow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B6dow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahcow6 ),
    .o(_al_u6910_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    _al_u6911 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yfcow6 ),
    .b(_al_u6910_o),
    .c(_al_u6857_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R4miu6 ));
  AL_MAP_LUT3 #(
    .EQN("~(C*B*~A)"),
    .INIT(8'hbf))
    _al_u6912 (
    .a(_al_u6844_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R4miu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y4miu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D4miu6 ));
  AL_MAP_LUT4 #(
    .EQN("(B*~(C*~(D*A)))"),
    .INIT(16'h8c0c))
    _al_u6913 (
    .a(_al_u6626_o),
    .b(_al_u6819_o),
    .c(_al_u6759_o),
    .d(_al_u5067_o),
    .o(_al_u6913_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*C)*~(B*~A))"),
    .INIT(16'hbb0b))
    _al_u6914 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bguiu6 ),
    .b(_al_u6819_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q2eow6 ),
    .d(_al_u1841_o),
    .o(_al_u6914_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B*~A))"),
    .INIT(8'hb0))
    _al_u6915 (
    .a(_al_u6034_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dyeow6_lutinv ),
    .c(_al_u6914_o),
    .o(_al_u6915_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*~B))"),
    .INIT(8'h8a))
    _al_u6916 (
    .a(_al_u6915_o),
    .b(_al_u6103_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qtfow6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K1cow6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*~B)*~(D*~A))"),
    .INIT(16'h8acf))
    _al_u6917 (
    .a(_al_u4663_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yzqiu6 ),
    .c(_al_u6819_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q2eow6 ),
    .o(_al_u6917_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B*~A))"),
    .INIT(8'hb0))
    _al_u6918 (
    .a(_al_u6135_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qtfow6_lutinv ),
    .c(_al_u6917_o),
    .o(_al_u6918_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*~B))"),
    .INIT(8'h8a))
    _al_u6919 (
    .a(_al_u6918_o),
    .b(_al_u6082_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dyeow6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B0cow6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u692 (
    .a(_al_u566_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[6] ),
    .o(_al_u692_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(~C*~A))"),
    .INIT(16'hfa32))
    _al_u6920 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eccow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xbcow6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K1cow6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B0cow6 ),
    .o(_al_u6920_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*C)*~(B*~A))"),
    .INIT(16'hbb0b))
    _al_u6921 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I0wiu6 ),
    .b(_al_u6819_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q2eow6 ),
    .d(_al_u1859_o),
    .o(_al_u6921_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u6922 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xa4ju6_lutinv ),
    .b(_al_u6921_o),
    .c(_al_u6817_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0cow6 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*~B))"),
    .INIT(8'ha8))
    _al_u6923 (
    .a(_al_u6920_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0cow6 ),
    .c(_al_u6857_o),
    .o(_al_u6923_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h3500))
    _al_u6924 (
    .a(_al_u6061_o),
    .b(_al_u6079_o),
    .c(_al_u5998_o),
    .d(_al_u6817_o),
    .o(_al_u6924_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u6925 (
    .a(_al_u6924_o),
    .b(_al_u4816_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q2eow6 ),
    .o(_al_u6925_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~C*~(D*~A)))"),
    .INIT(16'hc4c0))
    _al_u6926 (
    .a(_al_u6913_o),
    .b(_al_u6923_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vacow6 ),
    .d(_al_u6925_o),
    .o(_al_u6926_o));
  AL_MAP_LUT3 #(
    .EQN("~(C*B*~A)"),
    .INIT(8'hbf))
    _al_u6927 (
    .a(_al_u6844_o),
    .b(_al_u6926_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z1miu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E1miu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~C)*~(B*~A))"),
    .INIT(16'hb0bb))
    _al_u6928 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uc4ju6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qtfow6_lutinv ),
    .c(_al_u4886_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q2eow6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bxeow6 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*~B))"),
    .INIT(8'h8a))
    _al_u6929 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bxeow6 ),
    .b(_al_u6057_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dyeow6_lutinv ),
    .o(_al_u6929_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u693 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n6 ),
    .b(_al_u692_o),
    .c(_al_u467_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n49 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*~A))"),
    .INIT(8'h8c))
    _al_u6930 (
    .a(_al_u6732_o),
    .b(_al_u6929_o),
    .c(_al_u6819_o),
    .o(_al_u6930_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(~A*~(C*B)))"),
    .INIT(16'hea00))
    _al_u6931 (
    .a(_al_u6163_o),
    .b(_al_u6159_o),
    .c(_al_u6021_o),
    .d(_al_u6817_o),
    .o(_al_u6931_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'h5030))
    _al_u6932 (
    .a(_al_u1862_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U6wiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hemow6_lutinv ),
    .d(_al_u5001_o),
    .o(_al_u6932_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u6933 (
    .a(_al_u6931_o),
    .b(_al_u6932_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rjziu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(C*~A))"),
    .INIT(16'haf23))
    _al_u6934 (
    .a(_al_u4688_o),
    .b(_al_u6819_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q2eow6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eariu6 ),
    .o(_al_u6934_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*~B))"),
    .INIT(8'h8a))
    _al_u6935 (
    .a(_al_u6934_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mu3ju6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qtfow6_lutinv ),
    .o(_al_u6935_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*~B))"),
    .INIT(8'h8a))
    _al_u6936 (
    .a(_al_u6935_o),
    .b(_al_u6071_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dyeow6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Piziu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*C)*~(B*~A))"),
    .INIT(16'hbb0b))
    _al_u6937 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Umuiu6 ),
    .b(_al_u6819_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q2eow6 ),
    .d(_al_u1844_o),
    .o(_al_u6937_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B*~A))"),
    .INIT(8'hb0))
    _al_u6938 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F14ju6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qtfow6_lutinv ),
    .c(_al_u6937_o),
    .o(_al_u6938_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*~B))"),
    .INIT(8'h8a))
    _al_u6939 (
    .a(_al_u6938_o),
    .b(_al_u6125_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dyeow6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Alziu6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u694 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sq3ju6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*B)*~(~D*~A))"),
    .INIT(16'hf3a2))
    _al_u6940 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eccow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xbcow6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Piziu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Alziu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nycow6 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    _al_u6941 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rjziu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nycow6 ),
    .c(_al_u6857_o),
    .o(_al_u6941_o));
  AL_MAP_LUT4 #(
    .EQN("(D*B*~(~C*~A))"),
    .INIT(16'hc800))
    _al_u6942 (
    .a(_al_u6930_o),
    .b(_al_u6941_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vacow6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Azliu6 ),
    .o(_al_u6942_o));
  AL_MAP_LUT2 #(
    .EQN("~(B*~A)"),
    .INIT(4'hb))
    _al_u6943 (
    .a(_al_u6844_o),
    .b(_al_u6942_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fyliu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~C)*~(B*~A))"),
    .INIT(16'hb0bb))
    _al_u6944 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Id4ju6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qtfow6_lutinv ),
    .c(_al_u4529_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q2eow6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V1low6 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*~B))"),
    .INIT(8'h8a))
    _al_u6945 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V1low6 ),
    .b(_al_u6054_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dyeow6_lutinv ),
    .o(_al_u6945_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*~A))"),
    .INIT(8'h8c))
    _al_u6946 (
    .a(_al_u6719_o),
    .b(_al_u6945_o),
    .c(_al_u6819_o),
    .o(_al_u6946_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(~A*~(C*B)))"),
    .INIT(16'hea00))
    _al_u6947 (
    .a(_al_u6011_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lolow6 ),
    .c(_al_u6021_o),
    .d(_al_u6817_o),
    .o(_al_u6947_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*C)*~(B*~A))"),
    .INIT(16'hbb0b))
    _al_u6948 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bewiu6 ),
    .b(_al_u6819_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q2eow6 ),
    .d(_al_u1286_o),
    .o(_al_u6948_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u6949 (
    .a(_al_u6947_o),
    .b(_al_u6948_o),
    .o(_al_u6949_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u695 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sq3ju6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ),
    .o(_al_u695_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*~B)*~(D*~A))"),
    .INIT(16'h8acf))
    _al_u6950 (
    .a(_al_u4712_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kkriu6 ),
    .c(_al_u6819_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q2eow6 ),
    .o(_al_u6950_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*~B))"),
    .INIT(8'h8a))
    _al_u6951 (
    .a(_al_u6950_o),
    .b(_al_u6068_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dyeow6_lutinv ),
    .o(_al_u6951_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*~B))"),
    .INIT(8'h8a))
    _al_u6952 (
    .a(_al_u6951_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yt3ju6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qtfow6_lutinv ),
    .o(_al_u6952_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*C)*~(B*~A))"),
    .INIT(16'hbb0b))
    _al_u6953 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ntuiu6 ),
    .b(_al_u6819_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q2eow6 ),
    .d(_al_u1846_o),
    .o(_al_u6953_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B*~A))"),
    .INIT(8'hb0))
    _al_u6954 (
    .a(_al_u6122_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dyeow6_lutinv ),
    .c(_al_u6953_o),
    .o(_al_u6954_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*~B))"),
    .INIT(8'h8a))
    _al_u6955 (
    .a(_al_u6954_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R04ju6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qtfow6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G6cow6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*B)*~(~D*~A))"),
    .INIT(16'hf3a2))
    _al_u6956 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eccow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xbcow6_lutinv ),
    .c(_al_u6952_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G6cow6 ),
    .o(_al_u6956_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    _al_u6957 (
    .a(_al_u6949_o),
    .b(_al_u6956_o),
    .c(_al_u6857_o),
    .o(_al_u6957_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    _al_u6958 (
    .a(_al_u6946_o),
    .b(_al_u6957_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vacow6 ),
    .o(_al_u6958_o));
  AL_MAP_LUT3 #(
    .EQN("~(C*B*~A)"),
    .INIT(8'hbf))
    _al_u6959 (
    .a(_al_u6844_o),
    .b(_al_u6958_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uvliu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zuliu6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u696 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 ),
    .o(_al_u696_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(~C*~A))"),
    .INIT(16'hfa32))
    _al_u6960 (
    .a(_al_u6822_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xbcow6_lutinv ),
    .c(_al_u6857_o),
    .d(_al_u6829_o),
    .o(_al_u6960_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~C*~(D*~A)))"),
    .INIT(16'hc4c0))
    _al_u6961 (
    .a(_al_u6827_o),
    .b(_al_u6960_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vacow6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iimow6 ),
    .o(_al_u6961_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*~B))"),
    .INIT(8'ha8))
    _al_u6962 (
    .a(_al_u6961_o),
    .b(_al_u6820_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eccow6 ),
    .o(_al_u6962_o));
  AL_MAP_LUT3 #(
    .EQN("~(C*B*~A)"),
    .INIT(8'hbf))
    _al_u6963 (
    .a(_al_u6844_o),
    .b(_al_u6962_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Evkiu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vx9iu6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u6964 (
    .a(_al_u6842_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3how6_lutinv ),
    .o(_al_u6964_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u6965 (
    .a(_al_u6047_o),
    .b(_al_u6964_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tucow6_lutinv ),
    .o(_al_u6965_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~A*~(D*C))"),
    .INIT(16'h0111))
    _al_u6966 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tucow6_lutinv ),
    .b(_al_u6243_o),
    .c(_al_u609_o),
    .d(_al_u698_o),
    .o(_al_u6966_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*~A)"),
    .INIT(16'h0004))
    _al_u6967 (
    .a(_al_u6841_o),
    .b(_al_u6965_o),
    .c(_al_u6848_o),
    .d(_al_u6966_o),
    .o(_al_u6967_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u6968 (
    .a(_al_u6967_o),
    .b(_al_u6830_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tucow6_lutinv ),
    .o(_al_u6968_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(B*~A))"),
    .INIT(8'h0b))
    _al_u6969 (
    .a(_al_u6826_o),
    .b(_al_u6836_o),
    .c(_al_u6968_o),
    .o(_al_u6969_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u697 (
    .a(_al_u695_o),
    .b(_al_u696_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 ),
    .o(_al_u697_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u6970 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T23ju6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 ),
    .o(_al_u6970_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u6971 (
    .a(_al_u6970_o),
    .b(_al_u1582_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B4mow6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*~(C)*D))"),
    .INIT(16'h0144))
    _al_u6972 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ms5bx6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 ),
    .o(_al_u6972_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(~B*~(~D*C)))"),
    .INIT(16'h88a8))
    _al_u6973 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eccow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tucow6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B4mow6_lutinv ),
    .d(_al_u6972_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pkdow6 ));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u6974 (
    .a(_al_u6964_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tucow6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vo3ju6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kldow6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*~B)*~(~C*~A))"),
    .INIT(16'hfac8))
    _al_u6975 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pkdow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kldow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Plcow6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wlcow6 ),
    .o(_al_u6975_o));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'h47))
    _al_u6976 (
    .a(_al_u6047_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tucow6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vxniu6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hlziu6 ));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D*C*~B))"),
    .INIT(16'h8aaa))
    _al_u6977 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hlziu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tucow6_lutinv ),
    .c(_al_u1658_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pthiu6 ),
    .o(_al_u6977_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*~B))"),
    .INIT(8'ha8))
    _al_u6978 (
    .a(_al_u6975_o),
    .b(_al_u6977_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gkcow6 ),
    .o(_al_u6978_o));
  AL_MAP_LUT4 #(
    .EQN("(~(B)*~((~C*A))*~(D)+~(B)*(~C*A)*~(D)+~(B)*~((~C*A))*D+B*~((~C*A))*D+B*(~C*A)*D)"),
    .INIT(16'hfd33))
    _al_u6979 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 ),
    .o(_al_u6979_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u698 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 ),
    .o(_al_u698_o));
  AL_MAP_LUT4 #(
    .EQN("~((D*~C)*~(A)*~(B)+(D*~C)*A*~(B)+~((D*~C))*A*B+(D*~C)*A*B)"),
    .INIT(16'h7477))
    _al_u6980 (
    .a(_al_u6049_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tucow6_lutinv ),
    .c(_al_u6979_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ms5bx6 ),
    .o(_al_u6980_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*~B))"),
    .INIT(8'ha8))
    _al_u6981 (
    .a(_al_u6978_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ukcow6 ),
    .c(_al_u6980_o),
    .o(_al_u6981_o));
  AL_MAP_LUT3 #(
    .EQN("~(C*B*~A)"),
    .INIT(8'hbf))
    _al_u6982 (
    .a(_al_u6969_o),
    .b(_al_u6981_o),
    .c(_al_u6183_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hymiu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*~B)*~(~C*~A))"),
    .INIT(16'hfac8))
    _al_u6983 (
    .a(_al_u6822_o),
    .b(_al_u6977_o),
    .c(_al_u6980_o),
    .d(_al_u6829_o),
    .o(_al_u6983_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(~B*~(D*~A)))"),
    .INIT(16'hd0c0))
    _al_u6984 (
    .a(_al_u6827_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pkdow6 ),
    .c(_al_u6983_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iimow6 ),
    .o(_al_u6984_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*~B))"),
    .INIT(8'ha8))
    _al_u6985 (
    .a(_al_u6984_o),
    .b(_al_u6820_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kldow6 ),
    .o(_al_u6985_o));
  AL_MAP_LUT3 #(
    .EQN("~(C*B*~A)"),
    .INIT(8'hbf))
    _al_u6986 (
    .a(_al_u6969_o),
    .b(_al_u6985_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ngmiu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zfmiu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*~B)*~(~C*~A))"),
    .INIT(16'hfac8))
    _al_u6987 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pkdow6 ),
    .b(_al_u6977_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xv6ow6 ),
    .d(_al_u6876_o),
    .o(_al_u6987_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*~B))"),
    .INIT(8'ha8))
    _al_u6988 (
    .a(_al_u6987_o),
    .b(_al_u6870_o),
    .c(_al_u6980_o),
    .o(_al_u6988_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    _al_u6989 (
    .a(_al_u6867_o),
    .b(_al_u6988_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kldow6 ),
    .o(_al_u6989_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u699 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Np7ow6_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("~(C*B*~A)"),
    .INIT(8'hbf))
    _al_u6990 (
    .a(_al_u6969_o),
    .b(_al_u6989_o),
    .c(_al_u5886_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K3niu6 ));
  AL_MAP_LUT4 #(
    .EQN("~((B*~A)*~(C)*~(D)+(B*~A)*C*~(D)+~((B*~A))*C*D+(B*~A)*C*D)"),
    .INIT(16'h0fbb))
    _al_u6991 (
    .a(_al_u6969_o),
    .b(_al_u6989_o),
    .c(_al_u1581_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uzaiu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Czmiu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*~B)*~(~D*~A))"),
    .INIT(16'hfca8))
    _al_u6992 (
    .a(_al_u6977_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kldow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahcow6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kfcow6 ),
    .o(_al_u6992_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    _al_u6993 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pkdow6 ),
    .b(_al_u6992_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgcow6 ),
    .o(_al_u6993_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*~B))"),
    .INIT(8'ha8))
    _al_u6994 (
    .a(_al_u6993_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yfcow6 ),
    .c(_al_u6980_o),
    .o(_al_u6994_o));
  AL_MAP_LUT3 #(
    .EQN("~(C*B*~A)"),
    .INIT(8'hbf))
    _al_u6995 (
    .a(_al_u6969_o),
    .b(_al_u6994_o),
    .c(_al_u6188_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vrmiu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*~B)*~(~C*~A))"),
    .INIT(16'hfac8))
    _al_u6996 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pkdow6 ),
    .b(_al_u6977_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rcliu6 ),
    .d(_al_u6853_o),
    .o(_al_u6996_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*~B))"),
    .INIT(8'ha8))
    _al_u6997 (
    .a(_al_u6996_o),
    .b(_al_u6856_o),
    .c(_al_u6980_o),
    .o(_al_u6997_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    _al_u6998 (
    .a(_al_u6846_o),
    .b(_al_u6997_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kldow6 ),
    .o(_al_u6998_o));
  AL_MAP_LUT3 #(
    .EQN("~(C*B*~A)"),
    .INIT(8'hbf))
    _al_u6999 (
    .a(_al_u6969_o),
    .b(_al_u6998_o),
    .c(_al_u5918_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X6niu6 ));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u700 (
    .a(_al_u698_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Np7ow6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 ),
    .o(_al_u700_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*~B)*~(~D*~A))"),
    .INIT(16'hfca8))
    _al_u7000 (
    .a(_al_u6977_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kldow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K1cow6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B0cow6 ),
    .o(_al_u7000_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*~B))"),
    .INIT(8'ha8))
    _al_u7001 (
    .a(_al_u7000_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0cow6 ),
    .c(_al_u6980_o),
    .o(_al_u7001_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~C*~(D*~A)))"),
    .INIT(16'hc4c0))
    _al_u7002 (
    .a(_al_u6913_o),
    .b(_al_u7001_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pkdow6 ),
    .d(_al_u6925_o),
    .o(_al_u7002_o));
  AL_MAP_LUT3 #(
    .EQN("~(C*B*~A)"),
    .INIT(8'hbf))
    _al_u7003 (
    .a(_al_u6969_o),
    .b(_al_u7002_o),
    .c(_al_u5933_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bomiu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*~B)*~(~C*~A))"),
    .INIT(16'hfac8))
    _al_u7004 (
    .a(_al_u6977_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kldow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Piziu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Alziu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qodow6 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    _al_u7005 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rjziu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qodow6 ),
    .c(_al_u6980_o),
    .o(_al_u7005_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    _al_u7006 (
    .a(_al_u6930_o),
    .b(_al_u7005_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pkdow6 ),
    .o(_al_u7006_o));
  AL_MAP_LUT3 #(
    .EQN("~(C*B*~A)"),
    .INIT(8'hbf))
    _al_u7007 (
    .a(_al_u6969_o),
    .b(_al_u7006_o),
    .c(_al_u5954_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jlmiu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*~B)*~(~C*~A))"),
    .INIT(16'hfac8))
    _al_u7008 (
    .a(_al_u6977_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kldow6 ),
    .c(_al_u6952_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G6cow6 ),
    .o(_al_u7008_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    _al_u7009 (
    .a(_al_u6949_o),
    .b(_al_u7008_o),
    .c(_al_u6980_o),
    .o(_al_u7009_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u701 (
    .a(_al_u697_o),
    .b(_al_u700_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    _al_u7010 (
    .a(_al_u6946_o),
    .b(_al_u7009_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pkdow6 ),
    .o(_al_u7010_o));
  AL_MAP_LUT3 #(
    .EQN("~(C*B*~A)"),
    .INIT(8'hbf))
    _al_u7011 (
    .a(_al_u6969_o),
    .b(_al_u7010_o),
    .c(_al_u6193_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rimiu6 ));
  AL_MAP_LUT4 #(
    .EQN("~(C*~((~B*~A))*~(D)+C*(~B*~A)*~(D)+~(C)*(~B*~A)*D+C*(~B*~A)*D)"),
    .INIT(16'hee0f))
    _al_u7012 (
    .a(_al_u6046_o),
    .b(_al_u6100_o),
    .c(_al_u6830_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tucow6_lutinv ),
    .o(_al_u7012_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(B*~A))"),
    .INIT(8'h0b))
    _al_u7013 (
    .a(_al_u6826_o),
    .b(_al_u6836_o),
    .c(_al_u7012_o),
    .o(_al_u7013_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*~(D*B))"),
    .INIT(16'h1050))
    _al_u7014 (
    .a(_al_u6970_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ),
    .o(_al_u7014_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*~A))"),
    .INIT(8'h8c))
    _al_u7015 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ldiow6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qdhow6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 ),
    .o(_al_u7015_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(~B*~(~D*C)))"),
    .INIT(16'h88a8))
    _al_u7016 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eccow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tucow6_lutinv ),
    .c(_al_u7014_o),
    .d(_al_u7015_o),
    .o(_al_u7016_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    _al_u7017 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tucow6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mbhow6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S4kbx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G8how6 ));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(~B*~(D*C)))"),
    .INIT(16'h5444))
    _al_u7018 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tucow6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vxniu6_lutinv ),
    .c(_al_u1658_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pthiu6 ),
    .o(_al_u7018_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~A*~(~D*B))"),
    .INIT(16'h0501))
    _al_u7019 (
    .a(_al_u6964_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G8how6 ),
    .c(_al_u7018_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ms5bx6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ycliu6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u702 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Shopw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wxjpw6 ),
    .o(_al_u702_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*~B)*~(~D*~A))"),
    .INIT(16'hfca8))
    _al_u7020 (
    .a(_al_u7016_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ycliu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rcliu6 ),
    .d(_al_u6853_o),
    .o(_al_u7020_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u7021 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G8how6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ms5bx6 ),
    .o(_al_u7021_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    .INIT(16'h1013))
    _al_u7022 (
    .a(_al_u6046_o),
    .b(_al_u7021_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tucow6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vo3ju6_lutinv ),
    .o(_al_u7022_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*~B))"),
    .INIT(8'ha8))
    _al_u7023 (
    .a(_al_u7020_o),
    .b(_al_u6856_o),
    .c(_al_u7022_o),
    .o(_al_u7023_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(C*A))"),
    .INIT(16'h5f13))
    _al_u7024 (
    .a(_al_u1658_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mbhow6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ldiow6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S4kbx6 ),
    .o(_al_u7024_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    _al_u7025 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tucow6_lutinv ),
    .b(_al_u7024_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ms5bx6 ),
    .o(_al_u7025_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(~B*A))"),
    .INIT(8'h0d))
    _al_u7026 (
    .a(_al_u6848_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3how6_lutinv ),
    .c(_al_u7025_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cfliu6 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    _al_u7027 (
    .a(_al_u6846_o),
    .b(_al_u7023_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cfliu6 ),
    .o(_al_u7027_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u7028 (
    .a(_al_u7013_o),
    .b(_al_u7027_o),
    .o(_al_u7028_o));
  AL_MAP_LUT2 #(
    .EQN("~(B*A)"),
    .INIT(4'h7))
    _al_u7029 (
    .a(_al_u7028_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ibliu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tx8iu6 ));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u703 (
    .a(_al_u702_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dzvpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6kax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X7now6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*~B)*~(~D*~A))"),
    .INIT(16'hfca8))
    _al_u7030 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cfliu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ycliu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Plcow6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wlcow6 ),
    .o(_al_u7030_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    _al_u7031 (
    .a(_al_u7016_o),
    .b(_al_u7030_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gkcow6 ),
    .o(_al_u7031_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(~D*~C))"),
    .INIT(16'h4440))
    _al_u7032 (
    .a(_al_u7013_o),
    .b(_al_u7031_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ukcow6 ),
    .d(_al_u7022_o),
    .o(_al_u7032_o));
  AL_MAP_LUT2 #(
    .EQN("~(B*A)"),
    .INIT(4'h7))
    _al_u7033 (
    .a(_al_u7032_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cgkiu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qcaiu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*~B)*~(~D*~A))"),
    .INIT(16'hfca8))
    _al_u7034 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cfliu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ycliu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgcow6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahcow6 ),
    .o(_al_u7034_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    _al_u7035 (
    .a(_al_u7016_o),
    .b(_al_u7034_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kfcow6 ),
    .o(_al_u7035_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(~D*~C))"),
    .INIT(16'h4440))
    _al_u7036 (
    .a(_al_u7013_o),
    .b(_al_u7035_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yfcow6 ),
    .d(_al_u7022_o),
    .o(_al_u7036_o));
  AL_MAP_LUT2 #(
    .EQN("~(B*A)"),
    .INIT(4'h7))
    _al_u7037 (
    .a(_al_u7036_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dkkiu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jgkiu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*~B)*~(~D*~A))"),
    .INIT(16'hfca8))
    _al_u7038 (
    .a(_al_u7016_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cfliu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K1cow6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B0cow6 ),
    .o(_al_u7038_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*~B))"),
    .INIT(8'ha8))
    _al_u7039 (
    .a(_al_u7038_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0cow6 ),
    .c(_al_u7022_o),
    .o(_al_u7039_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u704 (
    .a(_al_u702_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dzvpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6kax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N9now6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~C*~(D*~A)))"),
    .INIT(16'hc4c0))
    _al_u7040 (
    .a(_al_u6913_o),
    .b(_al_u7039_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ycliu6 ),
    .d(_al_u6925_o),
    .o(_al_u7040_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u7041 (
    .a(_al_u7013_o),
    .b(_al_u7040_o),
    .o(_al_u7041_o));
  AL_MAP_LUT2 #(
    .EQN("~(B*A)"),
    .INIT(4'h7))
    _al_u7042 (
    .a(_al_u7041_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kkkiu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ef8iu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*~B)*~(~C*~A))"),
    .INIT(16'hfac8))
    _al_u7043 (
    .a(_al_u7016_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cfliu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Piziu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Alziu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gpeow6 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*~B))"),
    .INIT(8'ha8))
    _al_u7044 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gpeow6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rjziu6 ),
    .c(_al_u7022_o),
    .o(_al_u7044_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*~(~D*~B))"),
    .INIT(16'h5040))
    _al_u7045 (
    .a(_al_u7013_o),
    .b(_al_u6930_o),
    .c(_al_u7044_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ycliu6 ),
    .o(_al_u7045_o));
  AL_MAP_LUT2 #(
    .EQN("~(B*A)"),
    .INIT(4'h7))
    _al_u7046 (
    .a(_al_u7045_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lokiu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rkkiu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*~B)*~(~C*~A))"),
    .INIT(16'hfac8))
    _al_u7047 (
    .a(_al_u7016_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cfliu6 ),
    .c(_al_u6952_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G6cow6 ),
    .o(_al_u7047_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    _al_u7048 (
    .a(_al_u6949_o),
    .b(_al_u7047_o),
    .c(_al_u7022_o),
    .o(_al_u7048_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*~(~D*~B))"),
    .INIT(16'h5040))
    _al_u7049 (
    .a(_al_u7013_o),
    .b(_al_u6946_o),
    .c(_al_u7048_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ycliu6 ),
    .o(_al_u7049_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u705 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X7now6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N9now6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[0] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[0] ),
    .o(_al_u705_o));
  AL_MAP_LUT2 #(
    .EQN("~(B*A)"),
    .INIT(4'h7))
    _al_u7050 (
    .a(_al_u7049_o),
    .b(_al_u5892_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sokiu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*~B)*~(~D*~A))"),
    .INIT(16'hfca8))
    _al_u7051 (
    .a(_al_u7016_o),
    .b(_al_u6822_o),
    .c(_al_u7022_o),
    .d(_al_u6829_o),
    .o(_al_u7051_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~C*~(D*~A)))"),
    .INIT(16'hc4c0))
    _al_u7052 (
    .a(_al_u6827_o),
    .b(_al_u7051_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ycliu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iimow6 ),
    .o(_al_u7052_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(~D*~C))"),
    .INIT(16'h4440))
    _al_u7053 (
    .a(_al_u7013_o),
    .b(_al_u7052_o),
    .c(_al_u6820_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cfliu6 ),
    .o(_al_u7053_o));
  AL_MAP_LUT2 #(
    .EQN("~(B*A)"),
    .INIT(4'h7))
    _al_u7054 (
    .a(_al_u7053_o),
    .b(_al_u5972_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Drkiu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*~B)*~(~D*~A))"),
    .INIT(16'hfca8))
    _al_u7055 (
    .a(_al_u7016_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ycliu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xv6ow6 ),
    .d(_al_u6876_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mt6ow6 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*~B))"),
    .INIT(8'ha8))
    _al_u7056 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mt6ow6 ),
    .b(_al_u6870_o),
    .c(_al_u7022_o),
    .o(_al_u7056_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*~(~D*~B))"),
    .INIT(16'h5040))
    _al_u7057 (
    .a(_al_u7013_o),
    .b(_al_u6867_o),
    .c(_al_u7056_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cfliu6 ),
    .o(_al_u7057_o));
  AL_MAP_LUT2 #(
    .EQN("~(B*A)"),
    .INIT(4'h7))
    _al_u7058 (
    .a(_al_u7057_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bpliu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uoliu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7059 (
    .a(_al_u1774_o),
    .b(_al_u1791_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Halax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qakbx6 ),
    .o(_al_u7059_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*~A)"),
    .INIT(16'h0100))
    _al_u706 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dzvpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6kax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Shopw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wxjpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V6now6_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u7060 (
    .a(_al_u4284_o),
    .b(_al_u4289_o),
    .c(_al_u7059_o),
    .o(_al_u7060_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u7061 (
    .a(_al_u4289_o),
    .b(_al_u4172_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgziu6_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u7062 (
    .a(_al_u6844_o),
    .b(_al_u7060_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgziu6_lutinv ),
    .o(_al_u7062_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u7063 (
    .a(_al_u4289_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Et8iu6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Egziu6 ));
  AL_MAP_LUT4 #(
    .EQN("~(C*~((D*B))*~(A)+C*(D*B)*~(A)+~(C)*(D*B)*A+C*(D*B)*A)"),
    .INIT(16'h27af))
    _al_u7064 (
    .a(_al_u4289_o),
    .b(_al_u4290_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[21] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [21]),
    .o(_al_u7064_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u7065 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Egziu6 ),
    .b(_al_u7064_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [23]),
    .o(_al_u7065_o));
  AL_MAP_LUT4 #(
    .EQN("~(C*A*~(D*~B))"),
    .INIT(16'h7f5f))
    _al_u7066 (
    .a(_al_u7062_o),
    .b(_al_u6958_o),
    .c(_al_u7065_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgziu6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ocohu6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u7067 (
    .a(_al_u4289_o),
    .b(_al_u4290_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cmziu6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("~(C*~((D*B))*~(A)+C*(D*B)*~(A)+~(C)*(D*B)*A+C*(D*B)*A)"),
    .INIT(16'h27af))
    _al_u7068 (
    .a(_al_u4289_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Et8iu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[15] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [17]),
    .o(_al_u7068_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u7069 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cmziu6_lutinv ),
    .b(_al_u7068_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [15]),
    .o(_al_u7069_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*A)"),
    .INIT(16'h0200))
    _al_u707 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dzvpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6kax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Shopw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wxjpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C7now6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("~(C*A*~(D*~B))"),
    .INIT(16'h7f5f))
    _al_u7070 (
    .a(_al_u7062_o),
    .b(_al_u6861_o),
    .c(_al_u7069_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgziu6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zlohu6 ));
  AL_MAP_LUT4 #(
    .EQN("~(C*~((D*B))*~(A)+C*(D*B)*~(A)+~(C)*(D*B)*A+C*(D*B)*A)"),
    .INIT(16'h27af))
    _al_u7071 (
    .a(_al_u4289_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Et8iu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[16] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [18]),
    .o(_al_u7071_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u7072 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cmziu6_lutinv ),
    .b(_al_u7071_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [16]),
    .o(_al_u7072_o));
  AL_MAP_LUT4 #(
    .EQN("~(C*A*~(D*~B))"),
    .INIT(16'h7f5f))
    _al_u7073 (
    .a(_al_u7062_o),
    .b(_al_u6879_o),
    .c(_al_u7072_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgziu6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gmohu6 ));
  AL_MAP_LUT4 #(
    .EQN("~(C*~((D*B))*~(A)+C*(D*B)*~(A)+~(C)*(D*B)*A+C*(D*B)*A)"),
    .INIT(16'h27af))
    _al_u7074 (
    .a(_al_u4289_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Et8iu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[17] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [19]),
    .o(_al_u7074_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u7075 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cmziu6_lutinv ),
    .b(_al_u7074_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [17]),
    .o(_al_u7075_o));
  AL_MAP_LUT4 #(
    .EQN("~(C*A*~(D*~B))"),
    .INIT(16'h7f5f))
    _al_u7076 (
    .a(_al_u7062_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q7miu6 ),
    .c(_al_u7075_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgziu6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nmohu6 ));
  AL_MAP_LUT4 #(
    .EQN("~(C*~((D*B))*~(A)+C*(D*B)*~(A)+~(C)*(D*B)*A+C*(D*B)*A)"),
    .INIT(16'h27af))
    _al_u7077 (
    .a(_al_u4289_o),
    .b(_al_u4290_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[18] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [18]),
    .o(_al_u7077_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u7078 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Egziu6 ),
    .b(_al_u7077_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [20]),
    .o(_al_u7078_o));
  AL_MAP_LUT4 #(
    .EQN("~(C*A*~(D*~B))"),
    .INIT(16'h7f5f))
    _al_u7079 (
    .a(_al_u7062_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R4miu6 ),
    .c(_al_u7078_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgziu6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Umohu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u708 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V6now6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C7now6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[0] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[0] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yv9pw6 ));
  AL_MAP_LUT4 #(
    .EQN("~(C*~((D*B))*~(A)+C*(D*B)*~(A)+~(C)*(D*B)*A+C*(D*B)*A)"),
    .INIT(16'h27af))
    _al_u7080 (
    .a(_al_u4289_o),
    .b(_al_u4290_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[19] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [19]),
    .o(_al_u7080_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u7081 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Egziu6 ),
    .b(_al_u7080_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [21]),
    .o(_al_u7081_o));
  AL_MAP_LUT4 #(
    .EQN("~(C*A*~(D*~B))"),
    .INIT(16'h7f5f))
    _al_u7082 (
    .a(_al_u7062_o),
    .b(_al_u6926_o),
    .c(_al_u7081_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgziu6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bnohu6 ));
  AL_MAP_LUT4 #(
    .EQN("(D*~(B*~(~C*~A)))"),
    .INIT(16'h3700))
    _al_u7083 (
    .a(_al_u6930_o),
    .b(_al_u6941_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vacow6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgziu6_lutinv ),
    .o(_al_u7083_o));
  AL_MAP_LUT4 #(
    .EQN("~(C*~((D*B))*~(A)+C*(D*B)*~(A)+~(C)*(D*B)*A+C*(D*B)*A)"),
    .INIT(16'h27af))
    _al_u7084 (
    .a(_al_u4289_o),
    .b(_al_u4290_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[20] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [20]),
    .o(_al_u7084_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u7085 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Egziu6 ),
    .b(_al_u7084_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [22]),
    .o(_al_u7085_o));
  AL_MAP_LUT3 #(
    .EQN("~(C*~B*A)"),
    .INIT(8'hdf))
    _al_u7086 (
    .a(_al_u7062_o),
    .b(_al_u7083_o),
    .c(_al_u7085_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Inohu6 ));
  AL_MAP_LUT4 #(
    .EQN("~(C*~((D*B))*~(A)+C*(D*B)*~(A)+~(C)*(D*B)*A+C*(D*B)*A)"),
    .INIT(16'h27af))
    _al_u7087 (
    .a(_al_u4289_o),
    .b(_al_u4290_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[22] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [22]),
    .o(_al_u7087_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u7088 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Egziu6 ),
    .b(_al_u7087_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [24]),
    .o(_al_u7088_o));
  AL_MAP_LUT4 #(
    .EQN("~(C*A*~(D*~B))"),
    .INIT(16'h7f5f))
    _al_u7089 (
    .a(_al_u7062_o),
    .b(_al_u6962_o),
    .c(_al_u7088_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgziu6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Roohu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u709 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dzvpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6kax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Shopw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wxjpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9now6_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*~B))"),
    .INIT(8'ha8))
    _al_u7090 (
    .a(_al_u6842_o),
    .b(_al_u604_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ),
    .o(_al_u7090_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u7091 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hvcow6_lutinv ),
    .b(_al_u7090_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fucow6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~(B*~A))"),
    .INIT(16'hb000))
    _al_u7092 (
    .a(_al_u6826_o),
    .b(_al_u6836_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wxlow6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fucow6_lutinv ),
    .o(_al_u7092_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u7093 (
    .a(_al_u7090_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tucow6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vo3ju6_lutinv ),
    .o(_al_u7093_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*~B)*~(~D*~A))"),
    .INIT(16'hfca8))
    _al_u7094 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hlziu6 ),
    .b(_al_u7093_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Piziu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Alziu6 ),
    .o(_al_u7094_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u7095 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hvcow6_lutinv ),
    .b(_al_u6859_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kjziu6_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    _al_u7096 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rjziu6 ),
    .b(_al_u7094_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kjziu6_lutinv ),
    .o(_al_u7096_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*~A))"),
    .INIT(8'h8c))
    _al_u7097 (
    .a(_al_u6930_o),
    .b(_al_u7096_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xbcow6_lutinv ),
    .o(_al_u7097_o));
  AL_MAP_LUT3 #(
    .EQN("~(C*B*~A)"),
    .INIT(8'hbf))
    _al_u7098 (
    .a(_al_u7092_o),
    .b(_al_u7097_o),
    .c(_al_u5866_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P4liu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*~B)*~(~C*A))"),
    .INIT(16'hf5c4))
    _al_u7099 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xbcow6_lutinv ),
    .b(_al_u7093_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rcliu6 ),
    .d(_al_u6853_o),
    .o(_al_u7099_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*~A)"),
    .INIT(16'h1000))
    _al_u710 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dzvpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6kax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Shopw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wxjpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Panow6_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*~B))"),
    .INIT(8'ha8))
    _al_u7100 (
    .a(_al_u7099_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kjziu6_lutinv ),
    .c(_al_u6856_o),
    .o(_al_u7100_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*~(~D*~B))"),
    .INIT(16'h5040))
    _al_u7101 (
    .a(_al_u7092_o),
    .b(_al_u6846_o),
    .c(_al_u7100_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hlziu6 ),
    .o(_al_u7101_o));
  AL_MAP_LUT2 #(
    .EQN("~(B*A)"),
    .INIT(4'h7))
    _al_u7102 (
    .a(_al_u7101_o),
    .b(_al_u5896_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zvkiu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*~B)*~(~C*A))"),
    .INIT(16'hf5c4))
    _al_u7103 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xbcow6_lutinv ),
    .b(_al_u7093_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xv6ow6 ),
    .d(_al_u6876_o),
    .o(_al_u7103_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    _al_u7104 (
    .a(_al_u6870_o),
    .b(_al_u7103_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kjziu6_lutinv ),
    .o(_al_u7104_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*~(~D*~B))"),
    .INIT(16'h5040))
    _al_u7105 (
    .a(_al_u7092_o),
    .b(_al_u6867_o),
    .c(_al_u7104_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hlziu6 ),
    .o(_al_u7105_o));
  AL_MAP_LUT2 #(
    .EQN("~(B*A)"),
    .INIT(4'h7))
    _al_u7106 (
    .a(_al_u7105_o),
    .b(_al_u5871_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hsliu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*~B)*~(~C*A))"),
    .INIT(16'hf5c4))
    _al_u7107 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xbcow6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hlziu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Plcow6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wlcow6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ejcow6 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*~B))"),
    .INIT(8'ha8))
    _al_u7108 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ejcow6 ),
    .b(_al_u7093_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gkcow6 ),
    .o(_al_u7108_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    _al_u7109 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ukcow6 ),
    .b(_al_u7108_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kjziu6_lutinv ),
    .o(_al_u7109_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u711 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9now6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Panow6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[0] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[0] ),
    .o(_al_u711_o));
  AL_MAP_LUT3 #(
    .EQN("~(C*B*~A)"),
    .INIT(8'hbf))
    _al_u7110 (
    .a(_al_u7092_o),
    .b(_al_u7109_o),
    .c(_al_u5911_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fzkiu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*~B)*~(~C*A))"),
    .INIT(16'hf5c4))
    _al_u7111 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xbcow6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hlziu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgcow6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahcow6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iecow6 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*~B))"),
    .INIT(8'ha8))
    _al_u7112 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iecow6 ),
    .b(_al_u7093_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kfcow6 ),
    .o(_al_u7112_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    _al_u7113 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yfcow6 ),
    .b(_al_u7112_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kjziu6_lutinv ),
    .o(_al_u7113_o));
  AL_MAP_LUT3 #(
    .EQN("~(C*B*~A)"),
    .INIT(8'hbf))
    _al_u7114 (
    .a(_al_u7092_o),
    .b(_al_u7113_o),
    .c(_al_u5906_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X1liu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*~B)*~(~D*~A))"),
    .INIT(16'hfca8))
    _al_u7115 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hlziu6 ),
    .b(_al_u7093_o),
    .c(_al_u6952_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G6cow6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V3cow6 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    _al_u7116 (
    .a(_al_u6949_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V3cow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kjziu6_lutinv ),
    .o(_al_u7116_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*~A))"),
    .INIT(8'h8c))
    _al_u7117 (
    .a(_al_u6946_o),
    .b(_al_u7116_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xbcow6_lutinv ),
    .o(_al_u7117_o));
  AL_MAP_LUT4 #(
    .EQN("~(D*~C*B*~A)"),
    .INIT(16'hfbff))
    _al_u7118 (
    .a(_al_u7092_o),
    .b(_al_u7117_o),
    .c(_al_u5856_o),
    .d(_al_u5860_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K39iu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*~B)*~(~C*~A))"),
    .INIT(16'hfac8))
    _al_u7119 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hlziu6 ),
    .b(_al_u7093_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K1cow6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B0cow6 ),
    .o(_al_u7119_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u712 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dzvpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6kax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Shopw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wxjpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wanow6_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*~B))"),
    .INIT(8'ha8))
    _al_u7120 (
    .a(_al_u7119_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0cow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kjziu6_lutinv ),
    .o(_al_u7120_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(C*~(D*~A)))"),
    .INIT(16'h4c0c))
    _al_u7121 (
    .a(_al_u6913_o),
    .b(_al_u7120_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xbcow6_lutinv ),
    .d(_al_u6925_o),
    .o(_al_u7121_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u7122 (
    .a(_al_u7092_o),
    .b(_al_u7121_o),
    .o(_al_u7122_o));
  AL_MAP_LUT2 #(
    .EQN("~(B*A)"),
    .INIT(4'h7))
    _al_u7123 (
    .a(_al_u7122_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kgoiu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gfniu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*~C)*~(~B*~A))"),
    .INIT(16'heee0))
    _al_u7124 (
    .a(_al_u6822_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kjziu6_lutinv ),
    .c(_al_u7093_o),
    .d(_al_u6829_o),
    .o(_al_u7124_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(C*~(D*~A)))"),
    .INIT(16'h4c0c))
    _al_u7125 (
    .a(_al_u6827_o),
    .b(_al_u7124_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xbcow6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iimow6 ),
    .o(_al_u7125_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*~B))"),
    .INIT(8'ha8))
    _al_u7126 (
    .a(_al_u7125_o),
    .b(_al_u6820_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hlziu6 ),
    .o(_al_u7126_o));
  AL_MAP_LUT3 #(
    .EQN("~(C*B*~A)"),
    .INIT(8'hbf))
    _al_u7127 (
    .a(_al_u7092_o),
    .b(_al_u7126_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bbliu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D39iu6 ));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(B*~A))"),
    .INIT(8'h0b))
    _al_u7128 (
    .a(_al_u3874_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uzaiu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ),
    .o(_al_u7128_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*A)"),
    .INIT(16'h0200))
    _al_u7129 (
    .a(_al_u7128_o),
    .b(_al_u3874_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qaciu6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzjpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xibiu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*A)"),
    .INIT(16'h0002))
    _al_u713 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dzvpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6kax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Shopw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wxjpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E8now6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*~B)*~(D*A))"),
    .INIT(16'h45cf))
    _al_u7130 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xibiu6 ),
    .b(_al_u7128_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[0] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xdspw6 ),
    .o(_al_u7130_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u7131 (
    .a(_al_u3874_o),
    .b(_al_u4295_o),
    .o(_al_u7131_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C*~A))"),
    .INIT(8'h73))
    _al_u7132 (
    .a(_al_u7028_o),
    .b(_al_u7130_o),
    .c(_al_u7131_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W2vhu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*~B)*~(D*A))"),
    .INIT(16'h45cf))
    _al_u7133 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xibiu6 ),
    .b(_al_u7128_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[2] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jpmpw6 ),
    .o(_al_u7133_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C*~A))"),
    .INIT(8'h73))
    _al_u7134 (
    .a(_al_u7032_o),
    .b(_al_u7133_o),
    .c(_al_u7131_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G1vhu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*~B)*~(D*A))"),
    .INIT(16'h45cf))
    _al_u7135 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xibiu6 ),
    .b(_al_u7128_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[3] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xiipw6 ),
    .o(_al_u7135_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C*~A))"),
    .INIT(8'h73))
    _al_u7136 (
    .a(_al_u7036_o),
    .b(_al_u7135_o),
    .c(_al_u7131_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mrthu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(C*A))"),
    .INIT(16'h4c5f))
    _al_u7137 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xibiu6 ),
    .b(_al_u7128_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G2iax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[4] ),
    .o(_al_u7137_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C*~A))"),
    .INIT(8'h73))
    _al_u7138 (
    .a(_al_u7041_o),
    .b(_al_u7137_o),
    .c(_al_u7131_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ctthu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(C*A))"),
    .INIT(16'h4c5f))
    _al_u7139 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xibiu6 ),
    .b(_al_u7128_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F4iax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[5] ),
    .o(_al_u7139_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u714 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wanow6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E8now6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[0] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[0] ),
    .o(_al_u714_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C*~A))"),
    .INIT(8'h73))
    _al_u7140 (
    .a(_al_u7045_o),
    .b(_al_u7139_o),
    .c(_al_u7131_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C6vhu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*~B)*~(D*A))"),
    .INIT(16'h45cf))
    _al_u7141 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xibiu6 ),
    .b(_al_u7128_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[1] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T5mpw6 ),
    .o(_al_u7141_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C*~A))"),
    .INIT(8'h73))
    _al_u7142 (
    .a(_al_u7057_o),
    .b(_al_u7141_o),
    .c(_al_u7131_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S0vhu6 ));
  AL_MAP_LUT4 #(
    .EQN("~(C*~((D*B))*~(A)+C*(D*B)*~(A)+~(C)*(D*B)*A+C*(D*B)*A)"),
    .INIT(16'h27af))
    _al_u7143 (
    .a(_al_u4289_o),
    .b(_al_u4290_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[14] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [14]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idkow6 ));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*~(D*B))"),
    .INIT(16'h1050))
    _al_u7144 (
    .a(_al_u7060_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Egziu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idkow6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [16]),
    .o(_al_u7144_o));
  AL_MAP_LUT4 #(
    .EQN("~(C*~(D*~(B*~A)))"),
    .INIT(16'hbf0f))
    _al_u7145 (
    .a(_al_u6969_o),
    .b(_al_u6985_o),
    .c(_al_u7144_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgziu6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vcohu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*~A)*~(B)*~(C)+~(~D*~A)*B*~(C)+~(~(~D*~A))*B*C+~(~D*~A)*B*C)"),
    .INIT(16'hcfca))
    _al_u7146 (
    .a(_al_u6216_o),
    .b(_al_u2270_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ph8iu6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yi8iu6_lutinv ),
    .o(_al_u7146_o));
  AL_MAP_LUT4 #(
    .EQN("~(C*~(D*~(B*~A)))"),
    .INIT(16'hbf0f))
    _al_u7147 (
    .a(_al_u7092_o),
    .b(_al_u7117_o),
    .c(_al_u7146_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yi8iu6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R5liu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*~A)*~(C)*~(B)+~(~D*~A)*C*~(B)+~(~(~D*~A))*C*B+~(~D*~A)*C*B)"),
    .INIT(16'hf3e2))
    _al_u7148 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vioiu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ph8iu6_lutinv ),
    .c(_al_u2281_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yi8iu6_lutinv ),
    .o(_al_u7148_o));
  AL_MAP_LUT4 #(
    .EQN("~(C*~(D*~(B*~A)))"),
    .INIT(16'hbf0f))
    _al_u7149 (
    .a(_al_u7092_o),
    .b(_al_u7126_o),
    .c(_al_u7148_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yi8iu6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rgoiu6 ));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u715 (
    .a(_al_u705_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yv9pw6 ),
    .c(_al_u711_o),
    .d(_al_u714_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dc0iu6 ));
  AL_MAP_LUT4 #(
    .EQN("~(C*~((D*B))*~(A)+C*(D*B)*~(A)+~(C)*(D*B)*A+C*(D*B)*A)"),
    .INIT(16'h27af))
    _al_u7150 (
    .a(_al_u4289_o),
    .b(_al_u4290_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[1] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [1]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L0how6 ));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*~(D*B))"),
    .INIT(16'h1050))
    _al_u7151 (
    .a(_al_u7060_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Egziu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L0how6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [3]),
    .o(_al_u7151_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C*~A))"),
    .INIT(8'h73))
    _al_u7152 (
    .a(_al_u7032_o),
    .b(_al_u7151_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgziu6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ojohu6 ));
  AL_MAP_LUT4 #(
    .EQN("~(C*~((D*B))*~(A)+C*(D*B)*~(A)+~(C)*(D*B)*A+C*(D*B)*A)"),
    .INIT(16'h27af))
    _al_u7153 (
    .a(_al_u4289_o),
    .b(_al_u4290_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[2] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [2]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rwgow6 ));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*~(D*B))"),
    .INIT(16'h1050))
    _al_u7154 (
    .a(_al_u7060_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Egziu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rwgow6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [4]),
    .o(_al_u7154_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C*~A))"),
    .INIT(8'h73))
    _al_u7155 (
    .a(_al_u7036_o),
    .b(_al_u7154_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgziu6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vjohu6 ));
  AL_MAP_LUT4 #(
    .EQN("~(C*~((D*B))*~(A)+C*(D*B)*~(A)+~(C)*(D*B)*A+C*(D*B)*A)"),
    .INIT(16'h27af))
    _al_u7156 (
    .a(_al_u4289_o),
    .b(_al_u4290_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[3] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [3]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tkfow6 ));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*~(D*B))"),
    .INIT(16'h1050))
    _al_u7157 (
    .a(_al_u7060_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Egziu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tkfow6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [5]),
    .o(_al_u7157_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C*~A))"),
    .INIT(8'h73))
    _al_u7158 (
    .a(_al_u7041_o),
    .b(_al_u7157_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgziu6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ckohu6 ));
  AL_MAP_LUT4 #(
    .EQN("~(C*~((D*B))*~(A)+C*(D*B)*~(A)+~(C)*(D*B)*A+C*(D*B)*A)"),
    .INIT(16'h27af))
    _al_u7159 (
    .a(_al_u4289_o),
    .b(_al_u4290_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[4] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [4]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xneow6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u716 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dc0iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mifpw6 [0]));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*~(D*B))"),
    .INIT(16'h1050))
    _al_u7160 (
    .a(_al_u7060_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Egziu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xneow6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [6]),
    .o(_al_u7160_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C*~A))"),
    .INIT(8'h73))
    _al_u7161 (
    .a(_al_u7045_o),
    .b(_al_u7160_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgziu6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jkohu6 ));
  AL_MAP_LUT4 #(
    .EQN("~(C*~((D*B))*~(A)+C*(D*B)*~(A)+~(C)*(D*B)*A+C*(D*B)*A)"),
    .INIT(16'h27af))
    _al_u7162 (
    .a(_al_u4289_o),
    .b(_al_u4290_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[0] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [0]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wr6ow6 ));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*~(D*B))"),
    .INIT(16'h1050))
    _al_u7163 (
    .a(_al_u7060_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Egziu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wr6ow6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [2]),
    .o(_al_u7163_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C*~A))"),
    .INIT(8'h73))
    _al_u7164 (
    .a(_al_u7057_o),
    .b(_al_u7163_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgziu6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gtohu6 ));
  AL_MAP_LUT4 #(
    .EQN("~(C*~((D*B))*~(A)+C*(D*B)*~(A)+~(C)*(D*B)*A+C*(D*B)*A)"),
    .INIT(16'h27af))
    _al_u7165 (
    .a(_al_u4289_o),
    .b(_al_u4290_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[29] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [29]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M2cow6 ));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*~(D*B))"),
    .INIT(16'h1050))
    _al_u7166 (
    .a(_al_u7060_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Egziu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M2cow6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [31]),
    .o(_al_u7166_o));
  AL_MAP_LUT4 #(
    .EQN("~(C*~(D*~(B*~A)))"),
    .INIT(16'hbf0f))
    _al_u7167 (
    .a(_al_u7092_o),
    .b(_al_u7117_o),
    .c(_al_u7166_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgziu6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fpohu6 ));
  AL_MAP_LUT4 #(
    .EQN("~(C*~((D*B))*~(A)+C*(D*B)*~(A)+~(C)*(D*B)*A+C*(D*B)*A)"),
    .INIT(16'h27af))
    _al_u7168 (
    .a(_al_u4289_o),
    .b(_al_u4290_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[27] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [27]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qxbow6 ));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*~(D*B))"),
    .INIT(16'h1050))
    _al_u7169 (
    .a(_al_u7060_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Egziu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qxbow6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [29]),
    .o(_al_u7169_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u717 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N9now6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C7now6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[12] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[12] ),
    .o(_al_u717_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C*~A))"),
    .INIT(8'h73))
    _al_u7170 (
    .a(_al_u7122_o),
    .b(_al_u7169_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgziu6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mpohu6 ));
  AL_MAP_LUT4 #(
    .EQN("~(C*~((D*B))*~(A)+C*(D*B)*~(A)+~(C)*(D*B)*A+C*(D*B)*A)"),
    .INIT(16'h27af))
    _al_u7171 (
    .a(_al_u4289_o),
    .b(_al_u4290_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[30] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [30]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S98ow6 ));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*~(D*B))"),
    .INIT(16'h1050))
    _al_u7172 (
    .a(_al_u7060_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Egziu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S98ow6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [32]),
    .o(_al_u7172_o));
  AL_MAP_LUT4 #(
    .EQN("~(C*~(D*~(B*~A)))"),
    .INIT(16'hbf0f))
    _al_u7173 (
    .a(_al_u7092_o),
    .b(_al_u7126_o),
    .c(_al_u7172_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgziu6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xrohu6 ));
  AL_MAP_LUT4 #(
    .EQN("~(C*~((D*B))*~(A)+C*(D*B)*~(A)+~(C)*(D*B)*A+C*(D*B)*A)"),
    .INIT(16'h27af))
    _al_u7174 (
    .a(_al_u4289_o),
    .b(_al_u4290_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[9] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [9]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A0mow6 ));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*~(D*B))"),
    .INIT(16'h1050))
    _al_u7175 (
    .a(_al_u7060_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Egziu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A0mow6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [11]),
    .o(_al_u7175_o));
  AL_MAP_LUT4 #(
    .EQN("~(C*~(D*~(B*~A)))"),
    .INIT(16'hbf0f))
    _al_u7176 (
    .a(_al_u6969_o),
    .b(_al_u6981_o),
    .c(_al_u7175_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgziu6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hcohu6 ));
  AL_MAP_LUT4 #(
    .EQN("~(C*~((D*B))*~(A)+C*(D*B)*~(A)+~(C)*(D*B)*A+C*(D*B)*A)"),
    .INIT(16'h27af))
    _al_u7177 (
    .a(_al_u4289_o),
    .b(_al_u4290_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[8] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [8]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gdjow6 ));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*~(D*B))"),
    .INIT(16'h1050))
    _al_u7178 (
    .a(_al_u7060_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Egziu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gdjow6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [10]),
    .o(_al_u7178_o));
  AL_MAP_LUT4 #(
    .EQN("~(C*~(D*~(B*~A)))"),
    .INIT(16'hbf0f))
    _al_u7179 (
    .a(_al_u6969_o),
    .b(_al_u6989_o),
    .c(_al_u7178_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgziu6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cdohu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u718 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X7now6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Panow6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[12] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[12] ),
    .o(_al_u718_o));
  AL_MAP_LUT4 #(
    .EQN("~(C*~((D*B))*~(A)+C*(D*B)*~(A)+~(C)*(D*B)*A+C*(D*B)*A)"),
    .INIT(16'h27af))
    _al_u7180 (
    .a(_al_u4289_o),
    .b(_al_u4290_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[10] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [10]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eriow6 ));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*~(D*B))"),
    .INIT(16'h1050))
    _al_u7181 (
    .a(_al_u7060_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Egziu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eriow6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [12]),
    .o(_al_u7181_o));
  AL_MAP_LUT4 #(
    .EQN("~(C*~(D*~(B*~A)))"),
    .INIT(16'hbf0f))
    _al_u7182 (
    .a(_al_u6969_o),
    .b(_al_u6994_o),
    .c(_al_u7181_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgziu6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jdohu6 ));
  AL_MAP_LUT4 #(
    .EQN("~(C*~((D*B))*~(A)+C*(D*B)*~(A)+~(C)*(D*B)*A+C*(D*B)*A)"),
    .INIT(16'h27af))
    _al_u7183 (
    .a(_al_u4289_o),
    .b(_al_u4290_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[7] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [7]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jvdow6 ));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*~(D*B))"),
    .INIT(16'h1050))
    _al_u7184 (
    .a(_al_u7060_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Egziu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jvdow6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [9]),
    .o(_al_u7184_o));
  AL_MAP_LUT4 #(
    .EQN("~(C*~(D*~(B*~A)))"),
    .INIT(16'hbf0f))
    _al_u7185 (
    .a(_al_u6969_o),
    .b(_al_u6998_o),
    .c(_al_u7184_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgziu6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xkohu6 ));
  AL_MAP_LUT4 #(
    .EQN("~(C*~((D*B))*~(A)+C*(D*B)*~(A)+~(C)*(D*B)*A+C*(D*B)*A)"),
    .INIT(16'h27af))
    _al_u7186 (
    .a(_al_u4289_o),
    .b(_al_u4290_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[11] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [11]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Prdow6 ));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*~(D*B))"),
    .INIT(16'h1050))
    _al_u7187 (
    .a(_al_u7060_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Egziu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Prdow6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [13]),
    .o(_al_u7187_o));
  AL_MAP_LUT4 #(
    .EQN("~(C*~(D*~(B*~A)))"),
    .INIT(16'hbf0f))
    _al_u7188 (
    .a(_al_u6969_o),
    .b(_al_u7002_o),
    .c(_al_u7187_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgziu6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Elohu6 ));
  AL_MAP_LUT4 #(
    .EQN("~(C*~((D*B))*~(A)+C*(D*B)*~(A)+~(C)*(D*B)*A+C*(D*B)*A)"),
    .INIT(16'h27af))
    _al_u7189 (
    .a(_al_u4289_o),
    .b(_al_u4290_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[12] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [12]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hndow6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u719 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V6now6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wanow6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[12] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[12] ),
    .o(_al_u719_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*~(D*B))"),
    .INIT(16'h1050))
    _al_u7190 (
    .a(_al_u7060_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Egziu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hndow6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [14]),
    .o(_al_u7190_o));
  AL_MAP_LUT4 #(
    .EQN("~(C*~(D*~(B*~A)))"),
    .INIT(16'hbf0f))
    _al_u7191 (
    .a(_al_u6969_o),
    .b(_al_u7006_o),
    .c(_al_u7190_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgziu6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Llohu6 ));
  AL_MAP_LUT4 #(
    .EQN("~(C*~((D*B))*~(A)+C*(D*B)*~(A)+~(C)*(D*B)*A+C*(D*B)*A)"),
    .INIT(16'h27af))
    _al_u7192 (
    .a(_al_u4289_o),
    .b(_al_u4290_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[13] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [13]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eidow6 ));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*~(D*B))"),
    .INIT(16'h1050))
    _al_u7193 (
    .a(_al_u7060_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Egziu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eidow6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [15]),
    .o(_al_u7193_o));
  AL_MAP_LUT4 #(
    .EQN("~(C*~(D*~(B*~A)))"),
    .INIT(16'hbf0f))
    _al_u7194 (
    .a(_al_u6969_o),
    .b(_al_u7010_o),
    .c(_al_u7193_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgziu6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Slohu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*~A)*~(C)*~(B)+~(~D*~A)*C*~(B)+~(~(~D*~A))*C*B+~(~D*~A)*C*B)"),
    .INIT(16'hf3e2))
    _al_u7195 (
    .a(_al_u6236_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ph8iu6_lutinv ),
    .c(_al_u2429_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yi8iu6_lutinv ),
    .o(_al_u7195_o));
  AL_MAP_LUT4 #(
    .EQN("~(C*~(D*~(B*~A)))"),
    .INIT(16'hbf0f))
    _al_u7196 (
    .a(_al_u7092_o),
    .b(_al_u7097_o),
    .c(_al_u7195_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yi8iu6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sf8iu6 ));
  AL_MAP_LUT4 #(
    .EQN("~(C*~((D*B))*~(A)+C*(D*B)*~(A)+~(C)*(D*B)*A+C*(D*B)*A)"),
    .INIT(16'h27af))
    _al_u7197 (
    .a(_al_u4289_o),
    .b(_al_u4290_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[5] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [5]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dkeow6 ));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*~(D*B))"),
    .INIT(16'h1050))
    _al_u7198 (
    .a(_al_u7060_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Egziu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dkeow6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [7]),
    .o(_al_u7198_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C*~A))"),
    .INIT(8'h73))
    _al_u7199 (
    .a(_al_u7049_o),
    .b(_al_u7198_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgziu6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qkohu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u720 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9now6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E8now6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[12] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[12] ),
    .o(_al_u720_o));
  AL_MAP_LUT4 #(
    .EQN("~(C*~((D*B))*~(A)+C*(D*B)*~(A)+~(C)*(D*B)*A+C*(D*B)*A)"),
    .INIT(16'h27af))
    _al_u7200 (
    .a(_al_u4289_o),
    .b(_al_u4290_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[6] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [6]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W48ow6 ));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*~(D*B))"),
    .INIT(16'h1050))
    _al_u7201 (
    .a(_al_u7060_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Egziu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W48ow6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [8]),
    .o(_al_u7201_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C*~A))"),
    .INIT(8'h73))
    _al_u7202 (
    .a(_al_u7053_o),
    .b(_al_u7201_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgziu6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Esohu6 ));
  AL_MAP_LUT4 #(
    .EQN("~(C*~((D*B))*~(A)+C*(D*B)*~(A)+~(C)*(D*B)*A+C*(D*B)*A)"),
    .INIT(16'h27af))
    _al_u7203 (
    .a(_al_u4289_o),
    .b(_al_u4290_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[28] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [28]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cfziu6 ));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*~(D*B))"),
    .INIT(16'h1050))
    _al_u7204 (
    .a(_al_u7060_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Egziu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cfziu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [30]),
    .o(_al_u7204_o));
  AL_MAP_LUT4 #(
    .EQN("~(C*~(D*~(B*~A)))"),
    .INIT(16'hbf0f))
    _al_u7205 (
    .a(_al_u7092_o),
    .b(_al_u7097_o),
    .c(_al_u7204_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgziu6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hxohu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*C)*~(~B*A))"),
    .INIT(16'h0ddd))
    _al_u7206 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jjoiu6 ),
    .b(_al_u1299_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Et8iu6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [1]),
    .o(_al_u7206_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(~D*~(B*~A)))"),
    .INIT(16'hf040))
    _al_u7207 (
    .a(_al_u7013_o),
    .b(_al_u7027_o),
    .c(_al_u7206_o),
    .d(_al_u4172_o),
    .o(_al_u7207_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u7208 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jjoiu6 ),
    .b(_al_u1299_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgkbx6 ),
    .o(_al_u7208_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(B*~(D*~A)))"),
    .INIT(16'h0703))
    _al_u7209 (
    .a(_al_u7101_o),
    .b(_al_u7207_o),
    .c(_al_u7208_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yi8iu6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gn8iu6 ));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u721 (
    .a(_al_u717_o),
    .b(_al_u718_o),
    .c(_al_u719_o),
    .d(_al_u720_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ib0iu6 ));
  AL_MAP_LUT4 #(
    .EQN("~(C*~((D*B))*~(A)+C*(D*B)*~(A)+~(C)*(D*B)*A+C*(D*B)*A)"),
    .INIT(16'h27af))
    _al_u7210 (
    .a(_al_u4289_o),
    .b(_al_u4290_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[23] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [23]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lqcow6 ));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*~(D*B))"),
    .INIT(16'h1050))
    _al_u7211 (
    .a(_al_u7060_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Egziu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lqcow6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [25]),
    .o(_al_u7211_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C*~A))"),
    .INIT(8'h73))
    _al_u7212 (
    .a(_al_u7101_o),
    .b(_al_u7211_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgziu6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pnohu6 ));
  AL_MAP_LUT4 #(
    .EQN("~(C*~((D*B))*~(A)+C*(D*B)*~(A)+~(C)*(D*B)*A+C*(D*B)*A)"),
    .INIT(16'h27af))
    _al_u7213 (
    .a(_al_u4289_o),
    .b(_al_u4290_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[24] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [24]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rmcow6 ));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*~(D*B))"),
    .INIT(16'h1050))
    _al_u7214 (
    .a(_al_u7060_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Egziu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rmcow6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [26]),
    .o(_al_u7214_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C*~A))"),
    .INIT(8'h73))
    _al_u7215 (
    .a(_al_u7105_o),
    .b(_al_u7214_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgziu6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wnohu6 ));
  AL_MAP_LUT4 #(
    .EQN("~(C*~((D*B))*~(A)+C*(D*B)*~(A)+~(C)*(D*B)*A+C*(D*B)*A)"),
    .INIT(16'h27af))
    _al_u7216 (
    .a(_al_u4289_o),
    .b(_al_u4290_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[25] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [25]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vhcow6 ));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*~(D*B))"),
    .INIT(16'h1050))
    _al_u7217 (
    .a(_al_u7060_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Egziu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vhcow6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [27]),
    .o(_al_u7217_o));
  AL_MAP_LUT4 #(
    .EQN("~(C*~(D*~(B*~A)))"),
    .INIT(16'hbf0f))
    _al_u7218 (
    .a(_al_u7092_o),
    .b(_al_u7109_o),
    .c(_al_u7217_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgziu6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Doohu6 ));
  AL_MAP_LUT4 #(
    .EQN("~(C*~((D*B))*~(A)+C*(D*B)*~(A)+~(C)*(D*B)*A+C*(D*B)*A)"),
    .INIT(16'h27af))
    _al_u7219 (
    .a(_al_u4289_o),
    .b(_al_u4290_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[26] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [26]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zccow6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u722 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ib0iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mifpw6 [12]));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*~(D*B))"),
    .INIT(16'h1050))
    _al_u7220 (
    .a(_al_u7060_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Egziu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zccow6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [28]),
    .o(_al_u7220_o));
  AL_MAP_LUT4 #(
    .EQN("~(C*~(D*~(B*~A)))"),
    .INIT(16'hbf0f))
    _al_u7221 (
    .a(_al_u7092_o),
    .b(_al_u7113_o),
    .c(_al_u7220_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgziu6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Koohu6 ));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(B*A))"),
    .INIT(8'h07))
    _al_u7222 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ug8iu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P9niu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ),
    .o(_al_u7222_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*~B))"),
    .INIT(8'h8a))
    _al_u7223 (
    .a(_al_u7222_o),
    .b(_al_u2420_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ph8iu6_lutinv ),
    .o(_al_u7223_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*~B))"),
    .INIT(8'h8a))
    _al_u7224 (
    .a(_al_u7223_o),
    .b(_al_u6242_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ug8iu6_lutinv ),
    .o(_al_u7224_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u7225 (
    .a(_al_u7222_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_apsr_o[0] ),
    .o(_al_u7225_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(B*~(D*~A)))"),
    .INIT(16'h0703))
    _al_u7226 (
    .a(_al_u7122_o),
    .b(_al_u7224_o),
    .c(_al_u7225_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yi8iu6_lutinv ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Glphu6 ));
  AL_MAP_LUT1 #(
    .EQN("(~A)"),
    .INIT(2'h1))
    _al_u7227 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n11 ));
  AL_MAP_LUT1 #(
    .EQN("(~A)"),
    .INIT(2'h1))
    _al_u7228 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tu4iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fd7iu6 ));
  AL_MAP_LUT1 #(
    .EQN("(~A)"),
    .INIT(2'h1))
    _al_u7229 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Etmiu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Afkiu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u723 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X7now6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N9now6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[13] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[13] ),
    .o(_al_u723_o));
  AL_MAP_LUT1 #(
    .EQN("(~A)"),
    .INIT(2'h1))
    _al_u7230 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztmiu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pckiu6 ));
  AL_MAP_LUT1 #(
    .EQN("(~A)"),
    .INIT(2'h1))
    _al_u7231 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jsmiu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rdkiu6 ));
  AL_MAP_LUT1 #(
    .EQN("(~A)"),
    .INIT(2'h1))
    _al_u7232 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qsmiu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ddkiu6 ));
  AL_MAP_LUT1 #(
    .EQN("(~A)"),
    .INIT(2'h1))
    _al_u7233 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gumiu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mx8iu6 ));
  AL_MAP_LUT1 #(
    .EQN("(~A)"),
    .INIT(2'h1))
    _al_u7234 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ltmiu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ofkiu6 ));
  AL_MAP_LUT1 #(
    .EQN("(~A)"),
    .INIT(2'h1))
    _al_u7235 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xsmiu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wckiu6 ));
  AL_MAP_LUT1 #(
    .EQN("(~A)"),
    .INIT(2'h1))
    _al_u7236 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Csmiu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tekiu6 ));
  AL_MAP_LUT1 #(
    .EQN("(~A)"),
    .INIT(2'h1))
    _al_u7237 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Numiu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lf8iu6 ));
  AL_MAP_LUT1 #(
    .EQN("(~A)"),
    .INIT(2'h1))
    _al_u7238 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Stmiu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vfkiu6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u724 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V6now6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C7now6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[13] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[13] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A59pw6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u725 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9now6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Panow6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[13] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[13] ),
    .o(_al_u725_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u726 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wanow6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E8now6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[13] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[13] ),
    .o(_al_u726_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u727 (
    .a(_al_u723_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A59pw6 ),
    .c(_al_u725_o),
    .d(_al_u726_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bb0iu6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u728 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bb0iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mifpw6 [13]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u729 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X7now6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N9now6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[14] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[14] ),
    .o(_al_u729_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u730 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V6now6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C7now6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[14] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[14] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wv8pw6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u731 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9now6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wanow6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[14] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[14] ),
    .o(_al_u731_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u732 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Panow6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E8now6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[14] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[14] ),
    .o(_al_u732_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u733 (
    .a(_al_u729_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wv8pw6 ),
    .c(_al_u731_o),
    .d(_al_u732_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ua0iu6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u734 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ua0iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mifpw6 [14]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u735 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N9now6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C7now6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[15] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[15] ),
    .o(_al_u735_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u736 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X7now6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wanow6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[15] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[15] ),
    .o(_al_u736_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u737 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V6now6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Panow6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[15] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[15] ),
    .o(_al_u737_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u738 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9now6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E8now6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[15] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[15] ),
    .o(_al_u738_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u739 (
    .a(_al_u735_o),
    .b(_al_u736_o),
    .c(_al_u737_o),
    .d(_al_u738_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Na0iu6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u740 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Na0iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mifpw6 [15]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u741 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X7now6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wanow6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[16] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[16] ),
    .o(_al_u741_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u742 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N9now6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Panow6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[16] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[16] ),
    .o(_al_u742_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u743 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V6now6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C7now6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[16] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[16] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ad8pw6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u744 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9now6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E8now6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[16] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[16] ),
    .o(_al_u744_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u745 (
    .a(_al_u741_o),
    .b(_al_u742_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ad8pw6 ),
    .d(_al_u744_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ga0iu6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u746 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ga0iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mifpw6 [16]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u747 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X7now6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N9now6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[17] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[17] ),
    .o(_al_u747_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u748 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V6now6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C7now6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[17] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[17] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W38pw6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u749 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9now6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Panow6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[17] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[17] ),
    .o(_al_u749_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u750 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wanow6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E8now6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[17] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[17] ),
    .o(_al_u750_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u751 (
    .a(_al_u747_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W38pw6 ),
    .c(_al_u749_o),
    .d(_al_u750_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z90iu6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u752 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z90iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mifpw6 [17]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u753 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N9now6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C7now6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[18] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[18] ),
    .o(_al_u753_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u754 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X7now6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Panow6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[18] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[18] ),
    .o(_al_u754_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u755 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V6now6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wanow6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[18] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[18] ),
    .o(_al_u755_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u756 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9now6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E8now6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[18] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[18] ),
    .o(_al_u756_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u757 (
    .a(_al_u753_o),
    .b(_al_u754_o),
    .c(_al_u755_o),
    .d(_al_u756_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S90iu6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u758 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S90iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mifpw6 [18]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u759 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X7now6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9now6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[19] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[19] ),
    .o(_al_u759_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u760 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N9now6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C7now6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[19] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[19] ),
    .o(_al_u760_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u761 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Panow6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E8now6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[19] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[19] ),
    .o(_al_u761_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u762 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V6now6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wanow6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[19] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[19] ),
    .o(_al_u762_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u763 (
    .a(_al_u759_o),
    .b(_al_u760_o),
    .c(_al_u761_o),
    .d(_al_u762_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L90iu6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u764 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L90iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mifpw6 [19]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u765 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X7now6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9now6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[1] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[1] ),
    .o(_al_u765_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u766 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N9now6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C7now6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[1] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[1] ),
    .o(_al_u766_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u767 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Panow6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E8now6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[1] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[1] ),
    .o(_al_u767_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u768 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V6now6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wanow6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[1] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[1] ),
    .o(_al_u768_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u769 (
    .a(_al_u765_o),
    .b(_al_u766_o),
    .c(_al_u767_o),
    .d(_al_u768_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E90iu6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u770 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E90iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mifpw6 [1]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u771 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X7now6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N9now6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[20] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[20] ),
    .o(_al_u771_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u772 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9now6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wanow6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[20] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[20] ),
    .o(_al_u772_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u773 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V6now6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C7now6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[20] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[20] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L27pw6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u774 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Panow6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E8now6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[20] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[20] ),
    .o(_al_u774_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u775 (
    .a(_al_u771_o),
    .b(_al_u772_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L27pw6 ),
    .d(_al_u774_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X80iu6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u776 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X80iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mifpw6 [20]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u777 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N9now6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C7now6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[21] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[21] ),
    .o(_al_u777_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u778 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X7now6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Panow6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[21] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[21] ),
    .o(_al_u778_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u779 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V6now6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wanow6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[21] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[21] ),
    .o(_al_u779_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u780 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9now6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E8now6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[21] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[21] ),
    .o(_al_u780_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u781 (
    .a(_al_u777_o),
    .b(_al_u778_o),
    .c(_al_u779_o),
    .d(_al_u780_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q80iu6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u782 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q80iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mifpw6 [21]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u783 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X7now6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N9now6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[22] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[22] ),
    .o(_al_u783_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u784 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Panow6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wanow6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[22] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[22] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ml6pw6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u785 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V6now6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C7now6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[22] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[22] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dk6pw6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u786 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9now6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E8now6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[22] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[22] ),
    .o(_al_u786_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u787 (
    .a(_al_u783_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ml6pw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dk6pw6 ),
    .d(_al_u786_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J80iu6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u788 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J80iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mifpw6 [22]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u789 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N9now6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E8now6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[23] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[23] ),
    .o(_al_u789_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u790 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X7now6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wanow6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[23] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[23] ),
    .o(_al_u790_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u791 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V6now6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C7now6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[23] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[23] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Za6pw6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u792 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9now6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Panow6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[23] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[23] ),
    .o(_al_u792_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u793 (
    .a(_al_u789_o),
    .b(_al_u790_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Za6pw6 ),
    .d(_al_u792_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C80iu6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u794 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C80iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mifpw6 [23]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u795 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N9now6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C7now6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[24] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[24] ),
    .o(_al_u795_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u796 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X7now6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wanow6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[24] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[24] ),
    .o(_al_u796_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u797 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V6now6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Panow6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[24] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[24] ),
    .o(_al_u797_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u798 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9now6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E8now6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[24] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[24] ),
    .o(_al_u798_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u799 (
    .a(_al_u795_o),
    .b(_al_u796_o),
    .c(_al_u797_o),
    .d(_al_u798_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V70iu6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u800 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V70iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mifpw6 [24]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u801 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X7now6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N9now6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[25] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[25] ),
    .o(_al_u801_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u802 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9now6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Panow6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[25] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[25] ),
    .o(_al_u802_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u803 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V6now6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C7now6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[25] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[25] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rs5pw6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u804 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wanow6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E8now6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[25] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[25] ),
    .o(_al_u804_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u805 (
    .a(_al_u801_o),
    .b(_al_u802_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rs5pw6 ),
    .d(_al_u804_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O70iu6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u806 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O70iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mifpw6 [25]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u807 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X7now6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9now6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[26] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[26] ),
    .o(_al_u807_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u808 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N9now6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C7now6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[26] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[26] ),
    .o(_al_u808_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u809 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V6now6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E8now6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[26] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[26] ),
    .o(_al_u809_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u810 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Panow6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wanow6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[26] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[26] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wk5pw6 ));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u811 (
    .a(_al_u807_o),
    .b(_al_u808_o),
    .c(_al_u809_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wk5pw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H70iu6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u812 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H70iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mifpw6 [26]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u813 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N9now6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C7now6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[27] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[27] ),
    .o(_al_u813_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u814 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X7now6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Panow6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[27] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[27] ),
    .o(_al_u814_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u815 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V6now6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wanow6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[27] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[27] ),
    .o(_al_u815_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u816 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9now6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E8now6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[27] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[27] ),
    .o(_al_u816_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u817 (
    .a(_al_u813_o),
    .b(_al_u814_o),
    .c(_al_u815_o),
    .d(_al_u816_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A70iu6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u818 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A70iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mifpw6 [27]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u819 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X7now6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N9now6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[28] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[28] ),
    .o(_al_u819_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u820 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V6now6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C7now6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[28] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[28] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F15pw6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u821 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9now6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wanow6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[28] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[28] ),
    .o(_al_u821_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u822 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Panow6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E8now6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[28] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[28] ),
    .o(_al_u822_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u823 (
    .a(_al_u819_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F15pw6 ),
    .c(_al_u821_o),
    .d(_al_u822_o),
    .o(_al_u823_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u824 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 ),
    .b(_al_u823_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mifpw6 [28]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u825 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X7now6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wanow6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[29] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[29] ),
    .o(_al_u825_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u826 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N9now6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9now6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[29] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[29] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rt4pw6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u827 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V6now6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C7now6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[29] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[29] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bs4pw6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u828 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Panow6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E8now6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[29] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[29] ),
    .o(_al_u828_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u829 (
    .a(_al_u825_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rt4pw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bs4pw6 ),
    .d(_al_u828_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M60iu6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u830 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M60iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mifpw6 [29]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u831 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X7now6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9now6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[30] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[30] ),
    .o(_al_u831_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u832 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N9now6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C7now6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[30] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[30] ),
    .o(_al_u832_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u833 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V6now6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E8now6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[30] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[30] ),
    .o(_al_u833_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u834 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Panow6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wanow6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[30] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[30] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gk4pw6 ));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u835 (
    .a(_al_u831_o),
    .b(_al_u832_o),
    .c(_al_u833_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gk4pw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y50iu6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u836 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y50iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mifpw6 [30]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u837 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X7now6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N9now6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[6] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[6] ),
    .o(_al_u837_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u838 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V6now6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C7now6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[6] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[6] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ha4pw6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u839 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9now6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wanow6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[6] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[6] ),
    .o(_al_u839_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u840 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Panow6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E8now6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[6] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[6] ),
    .o(_al_u840_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u841 (
    .a(_al_u837_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ha4pw6 ),
    .c(_al_u839_o),
    .d(_al_u840_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P40iu6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u842 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P40iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mifpw6 [6]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u843 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X7now6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N9now6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[9] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[9] ),
    .o(_al_u843_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u844 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9now6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wanow6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[9] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[9] ),
    .o(_al_u844_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u845 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V6now6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C7now6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[9] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[9] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D14pw6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u846 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Panow6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E8now6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[9] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[9] ),
    .o(_al_u846_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u847 (
    .a(_al_u843_o),
    .b(_al_u844_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D14pw6 ),
    .d(_al_u846_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U30iu6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u848 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U30iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mifpw6 [9]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u849 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N9now6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C7now6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[31] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[31] ),
    .o(_al_u849_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u850 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X7now6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Panow6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[31] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[31] ),
    .o(_al_u850_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u851 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V6now6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wanow6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[31] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[31] ),
    .o(_al_u851_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u852 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9now6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E8now6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[31] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[31] ),
    .o(_al_u852_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u853 (
    .a(_al_u849_o),
    .b(_al_u850_o),
    .c(_al_u851_o),
    .d(_al_u852_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R50iu6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u854 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R50iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mifpw6 [31]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u855 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X7now6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N9now6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[4] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[4] ),
    .o(_al_u855_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u856 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Panow6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wanow6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[4] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[4] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J5pow6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u857 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V6now6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C7now6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[4] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[4] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A4pow6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u858 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9now6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E8now6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[4] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[4] ),
    .o(_al_u858_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u859 (
    .a(_al_u855_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J5pow6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A4pow6 ),
    .d(_al_u858_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D50iu6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u860 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D50iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mifpw6 [4]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u861 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N9now6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E8now6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[2] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[2] ),
    .o(_al_u861_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u862 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X7now6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wanow6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[2] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[2] ),
    .o(_al_u862_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u863 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V6now6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C7now6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[2] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[2] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G0pow6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u864 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9now6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Panow6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[2] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[2] ),
    .o(_al_u864_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u865 (
    .a(_al_u861_o),
    .b(_al_u862_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G0pow6 ),
    .d(_al_u864_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F60iu6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u866 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F60iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mifpw6 [2]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u867 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X7now6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wanow6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[3] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[3] ),
    .o(_al_u867_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u868 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N9now6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C7now6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[3] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[3] ),
    .o(_al_u868_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u869 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9now6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E8now6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[3] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[3] ),
    .o(_al_u869_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u870 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V6now6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Panow6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[3] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[3] ),
    .o(_al_u870_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u871 (
    .a(_al_u867_o),
    .b(_al_u868_o),
    .c(_al_u869_o),
    .d(_al_u870_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K50iu6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u872 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K50iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mifpw6 [3]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u873 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X7now6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9now6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[5] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[5] ),
    .o(_al_u873_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u874 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N9now6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C7now6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[5] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[5] ),
    .o(_al_u874_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u875 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Panow6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E8now6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[5] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[5] ),
    .o(_al_u875_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u876 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V6now6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wanow6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[5] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[5] ),
    .o(_al_u876_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u877 (
    .a(_al_u873_o),
    .b(_al_u874_o),
    .c(_al_u875_o),
    .d(_al_u876_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W40iu6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u878 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W40iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mifpw6 [5]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u879 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X7now6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Panow6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[8] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[8] ),
    .o(_al_u879_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u880 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N9now6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wanow6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[8] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[8] ),
    .o(_al_u880_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u881 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V6now6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C7now6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[8] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[8] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rhoow6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u882 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9now6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E8now6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[8] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[8] ),
    .o(_al_u882_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u883 (
    .a(_al_u879_o),
    .b(_al_u880_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rhoow6 ),
    .d(_al_u882_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B40iu6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u884 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B40iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mifpw6 [8]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u885 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N9now6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C7now6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[7] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[7] ),
    .o(_al_u885_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u886 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X7now6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9now6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[7] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[7] ),
    .o(_al_u886_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u887 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V6now6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Panow6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[7] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[7] ),
    .o(_al_u887_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u888 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wanow6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E8now6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[7] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[7] ),
    .o(_al_u888_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u889 (
    .a(_al_u885_o),
    .b(_al_u886_o),
    .c(_al_u887_o),
    .d(_al_u888_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I40iu6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u890 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I40iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mifpw6 [7]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u891 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N9now6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E8now6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[10] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[10] ),
    .o(_al_u891_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u892 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X7now6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wanow6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[10] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[10] ),
    .o(_al_u892_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u893 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V6now6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C7now6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[10] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[10] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cenow6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u894 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9now6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Panow6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[10] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[10] ),
    .o(_al_u894_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u895 (
    .a(_al_u891_o),
    .b(_al_u892_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cenow6 ),
    .d(_al_u894_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wb0iu6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u896 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wb0iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mifpw6 [10]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u897 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X7now6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Panow6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[11] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[11] ),
    .o(_al_u897_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u898 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N9now6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C7now6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[11] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[11] ),
    .o(_al_u898_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u899 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9now6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E8now6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[11] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[11] ),
    .o(_al_u899_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u900 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V6now6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wanow6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[11] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[11] ),
    .o(_al_u900_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u901 (
    .a(_al_u897_o),
    .b(_al_u898_o),
    .c(_al_u899_o),
    .d(_al_u900_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pb0iu6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u902 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pb0iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mifpw6 [11]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u903 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 ),
    .o(_al_u903_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u904 (
    .a(_al_u903_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 ),
    .o(_al_u904_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u905 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D6kiu6_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u906 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D6kiu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 ),
    .o(_al_u906_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u907 (
    .a(_al_u904_o),
    .b(_al_u906_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F85iu6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u908 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D6kiu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ),
    .o(_al_u908_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u909 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 ),
    .o(_al_u909_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u910 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F85iu6 ),
    .b(_al_u908_o),
    .c(_al_u909_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gpyiu6 ));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u911 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P14qw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nbkiu6_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u912 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nbkiu6_lutinv ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Skjax6 ),
    .o(_al_u912_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u913 (
    .a(_al_u912_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 ),
    .o(_al_u913_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u914 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 ),
    .o(_al_u914_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u915 (
    .a(_al_u914_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L45iu6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u916 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iekax6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lgkax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oikax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rkkax6 ),
    .o(_al_u916_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(B*~(C*A)))"),
    .INIT(16'hb300))
    _al_u917 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P14qw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Skjax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K75iu6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*C)*~(B*A))"),
    .INIT(16'h0777))
    _al_u918 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L45iu6_lutinv ),
    .b(_al_u916_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K75iu6_lutinv ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jckax6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aj1ju6 ));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u919 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P14qw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A95iu6_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u920 (
    .a(_al_u696_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A95iu6_lutinv ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Irmpw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oikax6 ),
    .o(_al_u920_o));
  AL_MAP_LUT4 #(
    .EQN("~(D*C*~B*A)"),
    .INIT(16'hdfff))
    _al_u921 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gpyiu6 ),
    .b(_al_u913_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aj1ju6 ),
    .d(_al_u920_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fi1ju6 ));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u922 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K84iu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R84iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y84iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F94iu6 ),
    .o(_al_u922_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    _al_u923 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ra2qw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Urgbx6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yzqpw6 ),
    .o(_al_u923_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    _al_u924 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dg2qw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gwwpw6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H0ebx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jvkpw6 ),
    .o(_al_u924_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u925 (
    .a(_al_u923_o),
    .b(_al_u924_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahdbx6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cfvpw6 ),
    .o(_al_u925_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u926 (
    .a(_al_u922_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G64iu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P74iu6 ),
    .d(_al_u925_o),
    .o(_al_u926_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u927 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vuciu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fnwiu6 ),
    .o(_al_u927_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u928 (
    .a(_al_u926_o),
    .b(_al_u927_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M94iu6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z54iu6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tu4iu6 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u929 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qyniu6_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u930 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ),
    .o(_al_u930_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u931 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qyniu6_lutinv ),
    .b(_al_u930_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 ),
    .o(_al_u931_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u932 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 ),
    .o(_al_u932_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u933 (
    .a(_al_u931_o),
    .b(_al_u932_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 ),
    .o(_al_u933_o));
  AL_MAP_LUT4 #(
    .EQN("~(~B*~(D*~(~C*A)))"),
    .INIT(16'hfdcc))
    _al_u934 (
    .a(_al_u927_o),
    .b(_al_u933_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dg2qw6 ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nj2qw6 ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E7vhu6 ));
  AL_MAP_LUT4 #(
    .EQN("(A*(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C))"),
    .INIT(16'ha808))
    _al_u935 (
    .a(_al_u470_o),
    .b(b_pad_gpio_porta_pad[7]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_ddr [7]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_dr [7]),
    .o(_al_u935_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*(A*~(D)*~(C)+A*D*~(C)+~(A)*D*C+A*D*C))"),
    .INIT(16'h3202))
    _al_u936 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/gpio_ext_porta_int [7]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_ddr [7]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_ls_sync ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/int_pre_in [7]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/ls_int_in [7]));
  AL_MAP_LUT4 #(
    .EQN("(B*(A*~(D)*~(C)+A*D*~(C)+~(A)*D*C+A*D*C))"),
    .INIT(16'hc808))
    _al_u937 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/ls_int_in [7]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inten [7]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inttype_level [7]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/gpio_intr_ed_pm [7]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_raw_intstatus [7]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~(~B*A))"),
    .INIT(16'h000d))
    _al_u938 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_intmask [7]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[4] ),
    .o(_al_u938_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u939 (
    .a(_al_u935_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_raw_intstatus [7]),
    .c(_al_u938_o),
    .o(_al_u939_o));
  EG_PHY_PAD #(
    //.LOCATION("T4"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u94 (
    .ipad(NRST),
    .di(NRST_pad));  // ../RTL/M0demo.v(7)
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h3ff5))
    _al_u940 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inten [7]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_int_polarity [7]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] ),
    .o(_al_u940_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf35f))
    _al_u941 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_intmask [7]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inttype_level [7]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] ),
    .o(_al_u941_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u942 (
    .a(_al_u940_o),
    .b(_al_u941_o),
    .o(_al_u942_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'h00ac))
    _al_u943 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_ddr [7]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_dr [7]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/sel0_b7/B1_0 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+A*~(B)*C*D+A*B*C*D)"),
    .INIT(16'haff3))
    _al_u944 (
    .a(_al_u942_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/sel0_b7/B1_0 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[4] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[5] ),
    .o(_al_u944_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u945 (
    .a(_al_u467_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[4] ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[5] ),
    .o(_al_u945_o));
  AL_MAP_LUT4 #(
    .EQN("~(~A*~((C*B))*~(D)+~A*(C*B)*~(D)+~(~A)*(C*B)*D+~A*(C*B)*D)"),
    .INIT(16'h3faa))
    _al_u946 (
    .a(_al_u944_o),
    .b(_al_u945_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/int_gpio_ls_sync [7]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[6] ),
    .o(_al_u946_o));
  AL_MAP_LUT4 #(
    .EQN("~(B*~(D*~C*~A))"),
    .INIT(16'h3733))
    _al_u947 (
    .a(_al_u939_o),
    .b(_al_u946_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[5] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[6] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n81 [7]));
  AL_MAP_LUT4 #(
    .EQN("(A*(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C))"),
    .INIT(16'ha808))
    _al_u948 (
    .a(_al_u470_o),
    .b(b_pad_gpio_porta_pad[6]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_ddr [6]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_dr [6]),
    .o(_al_u948_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*(A*~(D)*~(C)+A*D*~(C)+~(A)*D*C+A*D*C))"),
    .INIT(16'h3202))
    _al_u949 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/gpio_ext_porta_int [6]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_ddr [6]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_ls_sync ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/int_pre_in [6]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/ls_int_in [6]));
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("INV"))
    _al_u95 (
    .do({open_n451,open_n452,open_n453,\u_cmsdk_mcu/p0_out [15]}),
    .ts(\u_cmsdk_mcu/p0_outen [15]),
    .opad(P0[15]));  // ../RTL/cmsdk_mcu_pin_mux.v(141)
  AL_MAP_LUT4 #(
    .EQN("(B*(A*~(D)*~(C)+A*D*~(C)+~(A)*D*C+A*D*C))"),
    .INIT(16'hc808))
    _al_u950 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/ls_int_in [6]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inten [6]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inttype_level [6]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/gpio_intr_ed_pm [6]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_raw_intstatus [6]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~(~B*A))"),
    .INIT(16'h000d))
    _al_u951 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_intmask [6]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[4] ),
    .o(_al_u951_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(~A*~(C*B)))"),
    .INIT(16'h00ea))
    _al_u952 (
    .a(_al_u948_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_raw_intstatus [6]),
    .c(_al_u951_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[5] ),
    .o(_al_u952_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~A*~(C*B))"),
    .INIT(16'h1500))
    _al_u953 (
    .a(_al_u952_o),
    .b(_al_u945_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/int_gpio_ls_sync [6]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[6] ),
    .o(_al_u953_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h3ff5))
    _al_u954 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inten [6]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_int_polarity [6]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] ),
    .o(_al_u954_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf35f))
    _al_u955 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_intmask [6]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inttype_level [6]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] ),
    .o(_al_u955_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u956 (
    .a(_al_u566_o),
    .b(_al_u954_o),
    .c(_al_u955_o),
    .o(_al_u956_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'h00ac))
    _al_u957 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_ddr [6]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_dr [6]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/sel0_b6/B1_0 ));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(~C*~B*A))"),
    .INIT(16'h00fd))
    _al_u958 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/sel0_b6/B1_0 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[4] ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[5] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[6] ),
    .o(_al_u958_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u959 (
    .a(_al_u953_o),
    .b(_al_u956_o),
    .c(_al_u958_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n81 [6]));
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("INV"))
    _al_u96 (
    .do({open_n467,open_n468,open_n469,\u_cmsdk_mcu/p0_out [14]}),
    .ts(\u_cmsdk_mcu/p0_outen [14]),
    .opad(P0[14]));  // ../RTL/cmsdk_mcu_pin_mux.v(140)
  AL_MAP_LUT4 #(
    .EQN("(A*(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C))"),
    .INIT(16'ha808))
    _al_u960 (
    .a(_al_u470_o),
    .b(b_pad_gpio_porta_pad[5]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_ddr [5]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_dr [5]),
    .o(_al_u960_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*(A*~(D)*~(C)+A*D*~(C)+~(A)*D*C+A*D*C))"),
    .INIT(16'h3202))
    _al_u961 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/gpio_ext_porta_int [5]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_ddr [5]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_ls_sync ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/int_pre_in [5]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/ls_int_in [5]));
  AL_MAP_LUT4 #(
    .EQN("(B*(A*~(D)*~(C)+A*D*~(C)+~(A)*D*C+A*D*C))"),
    .INIT(16'hc808))
    _al_u962 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/ls_int_in [5]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inten [5]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inttype_level [5]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/gpio_intr_ed_pm [5]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_raw_intstatus [5]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~(~B*A))"),
    .INIT(16'h000d))
    _al_u963 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_intmask [5]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[4] ),
    .o(_al_u963_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(~A*~(C*B)))"),
    .INIT(16'h00ea))
    _al_u964 (
    .a(_al_u960_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_raw_intstatus [5]),
    .c(_al_u963_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[5] ),
    .o(_al_u964_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~A*~(C*B))"),
    .INIT(16'h1500))
    _al_u965 (
    .a(_al_u964_o),
    .b(_al_u945_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/int_gpio_ls_sync [5]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[6] ),
    .o(_al_u965_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h3ff5))
    _al_u966 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inten [5]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_int_polarity [5]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] ),
    .o(_al_u966_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf35f))
    _al_u967 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_intmask [5]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inttype_level [5]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] ),
    .o(_al_u967_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u968 (
    .a(_al_u566_o),
    .b(_al_u966_o),
    .c(_al_u967_o),
    .o(_al_u968_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'h00ac))
    _al_u969 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_ddr [5]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_dr [5]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/sel0_b5/B1_0 ));
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("INV"))
    _al_u97 (
    .do({open_n483,open_n484,open_n485,\u_cmsdk_mcu/p0_out [13]}),
    .ts(\u_cmsdk_mcu/p0_outen [13]),
    .opad(P0[13]));  // ../RTL/cmsdk_mcu_pin_mux.v(139)
  AL_MAP_LUT4 #(
    .EQN("(~D*~(~C*~B*A))"),
    .INIT(16'h00fd))
    _al_u970 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/sel0_b5/B1_0 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[4] ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[5] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[6] ),
    .o(_al_u970_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u971 (
    .a(_al_u965_o),
    .b(_al_u968_o),
    .c(_al_u970_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n81 [5]));
  AL_MAP_LUT4 #(
    .EQN("(A*(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C))"),
    .INIT(16'ha808))
    _al_u972 (
    .a(_al_u470_o),
    .b(b_pad_gpio_porta_pad[4]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_ddr [4]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_dr [4]),
    .o(_al_u972_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*(A*~(D)*~(C)+A*D*~(C)+~(A)*D*C+A*D*C))"),
    .INIT(16'h3202))
    _al_u973 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/gpio_ext_porta_int [4]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_ddr [4]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_ls_sync ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/int_pre_in [4]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/ls_int_in [4]));
  AL_MAP_LUT4 #(
    .EQN("(B*(A*~(D)*~(C)+A*D*~(C)+~(A)*D*C+A*D*C))"),
    .INIT(16'hc808))
    _al_u974 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/ls_int_in [4]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inten [4]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inttype_level [4]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/gpio_intr_ed_pm [4]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_raw_intstatus [4]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~(~B*A))"),
    .INIT(16'h000d))
    _al_u975 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_intmask [4]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[4] ),
    .o(_al_u975_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(~A*~(C*B)))"),
    .INIT(16'h00ea))
    _al_u976 (
    .a(_al_u972_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_raw_intstatus [4]),
    .c(_al_u975_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[5] ),
    .o(_al_u976_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~A*~(C*B))"),
    .INIT(16'h1500))
    _al_u977 (
    .a(_al_u976_o),
    .b(_al_u945_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/int_gpio_ls_sync [4]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[6] ),
    .o(_al_u977_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h3ff5))
    _al_u978 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inten [4]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_int_polarity [4]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] ),
    .o(_al_u978_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf35f))
    _al_u979 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_intmask [4]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inttype_level [4]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] ),
    .o(_al_u979_o));
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("INV"))
    _al_u98 (
    .do({open_n499,open_n500,open_n501,\u_cmsdk_mcu/p0_out [12]}),
    .ts(\u_cmsdk_mcu/p0_outen [12]),
    .opad(P0[12]));  // ../RTL/cmsdk_mcu_pin_mux.v(138)
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u980 (
    .a(_al_u566_o),
    .b(_al_u978_o),
    .c(_al_u979_o),
    .o(_al_u980_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'h00ac))
    _al_u981 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_ddr [4]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_dr [4]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/sel0_b4/B1_0 ));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(~C*~B*A))"),
    .INIT(16'h00fd))
    _al_u982 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/sel0_b4/B1_0 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[4] ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[5] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[6] ),
    .o(_al_u982_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u983 (
    .a(_al_u977_o),
    .b(_al_u980_o),
    .c(_al_u982_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n81 [4]));
  AL_MAP_LUT4 #(
    .EQN("(A*(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C))"),
    .INIT(16'ha808))
    _al_u984 (
    .a(_al_u470_o),
    .b(b_pad_gpio_porta_pad[3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_ddr [3]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_dr [3]),
    .o(_al_u984_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*(A*~(D)*~(C)+A*D*~(C)+~(A)*D*C+A*D*C))"),
    .INIT(16'h3202))
    _al_u985 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/gpio_ext_porta_int [3]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_ddr [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_ls_sync ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/int_pre_in [3]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/ls_int_in [3]));
  AL_MAP_LUT4 #(
    .EQN("(B*(A*~(D)*~(C)+A*D*~(C)+~(A)*D*C+A*D*C))"),
    .INIT(16'hc808))
    _al_u986 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/ls_int_in [3]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inten [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inttype_level [3]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/gpio_intr_ed_pm [3]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_raw_intstatus [3]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~(~B*A))"),
    .INIT(16'h000d))
    _al_u987 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_intmask [3]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[4] ),
    .o(_al_u987_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(~A*~(C*B)))"),
    .INIT(16'h00ea))
    _al_u988 (
    .a(_al_u984_o),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_raw_intstatus [3]),
    .c(_al_u987_o),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[5] ),
    .o(_al_u988_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~A*~(C*B))"),
    .INIT(16'h1500))
    _al_u989 (
    .a(_al_u988_o),
    .b(_al_u945_o),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/int_gpio_ls_sync [3]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[6] ),
    .o(_al_u989_o));
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("INV"))
    _al_u99 (
    .do({open_n515,open_n516,open_n517,\u_cmsdk_mcu/p0_out [11]}),
    .ts(\u_cmsdk_mcu/p0_outen [11]),
    .opad(P0[11]));  // ../RTL/cmsdk_mcu_pin_mux.v(137)
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h3ff5))
    _al_u990 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inten [3]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_int_polarity [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] ),
    .o(_al_u990_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf35f))
    _al_u991 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_intmask [3]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inttype_level [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] ),
    .o(_al_u991_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u992 (
    .a(_al_u566_o),
    .b(_al_u990_o),
    .c(_al_u991_o),
    .o(_al_u992_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'h00ac))
    _al_u993 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_ddr [3]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_dr [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/sel0_b3/B1_0 ));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(~C*~B*A))"),
    .INIT(16'h00fd))
    _al_u994 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/sel0_b3/B1_0 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[4] ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[5] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[6] ),
    .o(_al_u994_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u995 (
    .a(_al_u989_o),
    .b(_al_u992_o),
    .c(_al_u994_o),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n81 [3]));
  AL_MAP_LUT4 #(
    .EQN("(A*(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C))"),
    .INIT(16'ha808))
    _al_u996 (
    .a(_al_u470_o),
    .b(b_pad_gpio_porta_pad[2]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_ddr [2]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_dr [2]),
    .o(_al_u996_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*(A*~(D)*~(C)+A*D*~(C)+~(A)*D*C+A*D*C))"),
    .INIT(16'h3202))
    _al_u997 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/gpio_ext_porta_int [2]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_ddr [2]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_ls_sync ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/int_pre_in [2]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/ls_int_in [2]));
  AL_MAP_LUT4 #(
    .EQN("(B*(A*~(D)*~(C)+A*D*~(C)+~(A)*D*C+A*D*C))"),
    .INIT(16'hc808))
    _al_u998 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/ls_int_in [2]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inten [2]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inttype_level [2]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/gpio_intr_ed_pm [2]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_raw_intstatus [2]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~(~B*A))"),
    .INIT(16'h000d))
    _al_u999 (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_intmask [2]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[4] ),
    .o(_al_u999_o));
  EG_PHY_CONFIG #(
    .DONE_PERSISTN("ENABLE"),
    .INIT_PERSISTN("ENABLE"),
    .JTAG_PERSISTN("DISABLE"),
    .PROGRAMN_PERSISTN("DISABLE"))
    config_inst ();
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u1/u0  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_1_0_0 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_1_0 ),
    .c(\u1/c0 ),
    .o({\u1/c1 ,n0[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u1/u1  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_1_0_1 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_1_1 ),
    .c(\u1/c1 ),
    .o({\u1/c2 ,n0[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u1/u10  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_1_0_10 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_1_10 ),
    .c(\u1/c10 ),
    .o({\u1/c11 ,n0[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u1/u11  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_1_0_11 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_1_11 ),
    .c(\u1/c11 ),
    .o({\u1/c12 ,n0[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u1/u12  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_1_0_12 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_1_12 ),
    .c(\u1/c12 ),
    .o({\u1/c13 ,n0[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u1/u13  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_1_0_13 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_1_13 ),
    .c(\u1/c13 ),
    .o({open_n577,n0[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u1/u2  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_1_0_2 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_1_2 ),
    .c(\u1/c2 ),
    .o({\u1/c3 ,n0[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u1/u3  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_1_0_3 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_1_3 ),
    .c(\u1/c3 ),
    .o({\u1/c4 ,n0[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u1/u4  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_1_0_4 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_1_4 ),
    .c(\u1/c4 ),
    .o({\u1/c5 ,n0[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u1/u5  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_1_0_5 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_1_5 ),
    .c(\u1/c5 ),
    .o({\u1/c6 ,n0[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u1/u6  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_1_0_6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_1_6 ),
    .c(\u1/c6 ),
    .o({\u1/c7 ,n0[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u1/u7  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_1_0_7 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_1_7 ),
    .c(\u1/c7 ),
    .o({\u1/c8 ,n0[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u1/u8  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_1_0_8 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_1_8 ),
    .c(\u1/c8 ),
    .o({\u1/c9 ,n0[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u1/u9  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_1_0_9 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_1_9 ),
    .c(\u1/c9 ),
    .o({\u1/c10 ,n0[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u1/ucin  (
    .a(1'b0),
    .o({\u1/c0 ,open_n580}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2/u0  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_18 ),
    .b(n0[0]),
    .c(\u2/c0 ),
    .o({\u2/c1 ,n1[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2/u1  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_19 ),
    .b(n0[1]),
    .c(\u2/c1 ),
    .o({\u2/c2 ,n1[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2/u10  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_28 ),
    .b(n0[10]),
    .c(\u2/c10 ),
    .o({\u2/c11 ,n1[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2/u11  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_29 ),
    .b(n0[11]),
    .c(\u2/c11 ),
    .o({\u2/c12 ,n1[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2/u12  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_30 ),
    .b(n0[12]),
    .c(\u2/c12 ),
    .o({\u2/c13 ,n1[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2/u13  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_31 ),
    .b(n0[13]),
    .c(\u2/c13 ),
    .o({open_n581,n1[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2/u2  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_20 ),
    .b(n0[2]),
    .c(\u2/c2 ),
    .o({\u2/c3 ,n1[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2/u3  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_21 ),
    .b(n0[3]),
    .c(\u2/c3 ),
    .o({\u2/c4 ,n1[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2/u4  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_22 ),
    .b(n0[4]),
    .c(\u2/c4 ),
    .o({\u2/c5 ,n1[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2/u5  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_23 ),
    .b(n0[5]),
    .c(\u2/c5 ),
    .o({\u2/c6 ,n1[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2/u6  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_24 ),
    .b(n0[6]),
    .c(\u2/c6 ),
    .o({\u2/c7 ,n1[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2/u7  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_25 ),
    .b(n0[7]),
    .c(\u2/c7 ),
    .o({\u2/c8 ,n1[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2/u8  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_26 ),
    .b(n0[8]),
    .c(\u2/c8 ),
    .o({\u2/c9 ,n1[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2/u9  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_27 ),
    .b(n0[9]),
    .c(\u2/c9 ),
    .o({\u2/c10 ,n1[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2/ucin  (
    .a(1'b0),
    .o({\u2/c0 ,open_n584}));
  EG_PHY_GCLK \u_M0clkpll/bufg_feedback  (
    .clki(\u_M0clkpll/clk0_buf ),
    .clko(XTAL1_wire));  // al_ip/M0clkpll.v(36)
  EG_PHY_PLL #(
    .CLKC0_CPHASE(124),
    .CLKC0_DIV(125),
    .CLKC0_DIV2_ENABLE("DISABLE"),
    .CLKC0_ENABLE("ENABLE"),
    .CLKC0_FPHASE(0),
    .CLKC1_CPHASE(1),
    .CLKC1_DIV(1),
    .CLKC1_DIV2_ENABLE("DISABLE"),
    .CLKC1_ENABLE("DISABLE"),
    .CLKC1_FPHASE(0),
    .CLKC2_CPHASE(1),
    .CLKC2_DIV(1),
    .CLKC2_DIV2_ENABLE("DISABLE"),
    .CLKC2_ENABLE("DISABLE"),
    .CLKC2_FPHASE(0),
    .CLKC3_CPHASE(1),
    .CLKC3_DIV(1),
    .CLKC3_DIV2_ENABLE("DISABLE"),
    .CLKC3_ENABLE("DISABLE"),
    .CLKC3_FPHASE(0),
    .CLKC4_CPHASE(1),
    .CLKC4_DIV(1),
    .CLKC4_DIV2_ENABLE("DISABLE"),
    .CLKC4_ENABLE("DISABLE"),
    .CLKC4_FPHASE(0),
    .DERIVE_PLL_CLOCKS("DISABLE"),
    .DPHASE_SOURCE("DISABLE"),
    .DYNCFG("DISABLE"),
    .FBCLK_DIV(1),
    .FEEDBK_MODE("NORMAL"),
    .FEEDBK_PATH("CLKC0_EXT"),
    .FIN("24.000"),
    .FREQ_LOCK_ACCURACY(2),
    .GEN_BASIC_CLOCK("DISABLE"),
    .GMC_GAIN(6),
    .GMC_TEST(14),
    .ICP_CURRENT(3),
    .IF_ESCLKSTSW("DISABLE"),
    .INTFB_WAKE("DISABLE"),
    .KVCO(6),
    .LPF_CAPACITOR(3),
    .LPF_RESISTOR(2),
    .NORESET("DISABLE"),
    .ODIV_MUXC0("DIV"),
    .ODIV_MUXC1("DIV"),
    .ODIV_MUXC2("DIV"),
    .ODIV_MUXC3("DIV"),
    .ODIV_MUXC4("DIV"),
    .PLLC2RST_ENA("DISABLE"),
    .PLLC34RST_ENA("DISABLE"),
    .PLLMRST_ENA("DISABLE"),
    .PLLRST_ENA("ENABLE"),
    .PLL_LOCK_MODE(0),
    .PREDIV_MUXC0("VCO"),
    .PREDIV_MUXC1("VCO"),
    .PREDIV_MUXC2("VCO"),
    .PREDIV_MUXC3("VCO"),
    .PREDIV_MUXC4("VCO"),
    .REFCLK_DIV(3),
    .REFCLK_SEL("INTERNAL"),
    .STDBY_ENABLE("ENABLE"),
    .STDBY_VCO_ENA("DISABLE"),
    .SYNC_ENABLE("DISABLE"),
    .VCO_NORESET("DISABLE"))
    \u_M0clkpll/pll_inst  (
    .daddr(6'b000000),
    .dclk(1'b0),
    .dcs(1'b0),
    .di(8'b00000000),
    .dwe(1'b0),
    .fbclk(XTAL1_wire),
    .psclk(1'b0),
    .psclksel(3'b000),
    .psdown(1'b0),
    .psstep(1'b0),
    .refclk(XTAL1_pad),
    .reset(1'b0),
    .stdby(1'b0),
    .clkc({open_n585,open_n586,open_n587,open_n588,\u_M0clkpll/clk0_buf }));  // al_ip/M0clkpll.v(59)
  // address_offset=0;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=32;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("1"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("1"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("ASYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("READBEFOREWRITE"))
    \u_cmsdk_mcu/u_ahb_ram/ram_memory0_1024x32_sub_000000_000  (
    .addra({\u_cmsdk_mcu/HADDR [11:2],3'b111}),
    .addrb({\u_cmsdk_mcu/u_ahb_ram/buf_hwaddr [11:2],3'b111}),
    .clka(XTAL1_wire),
    .clkb(XTAL1_wire),
    .dia(9'b000000000),
    .dib(\u_cmsdk_mcu/u_ahb_ram/n13 [8:0]),
    .web(\u_cmsdk_mcu/u_ahb_ram/n16 ),
    .doa(\u_cmsdk_mcu/sram_hrdata [8:0]));
  // address_offset=0;data_offset=9;depth=1024;width=9;num_section=1;width_per_section=9;section_size=32;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("1"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("1"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("ASYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("READBEFOREWRITE"))
    \u_cmsdk_mcu/u_ahb_ram/ram_memory0_1024x32_sub_000000_009  (
    .addra({\u_cmsdk_mcu/HADDR [11:2],3'b111}),
    .addrb({\u_cmsdk_mcu/u_ahb_ram/buf_hwaddr [11:2],3'b111}),
    .clka(XTAL1_wire),
    .clkb(XTAL1_wire),
    .dia(9'b000000000),
    .dib(\u_cmsdk_mcu/u_ahb_ram/n13 [17:9]),
    .web(\u_cmsdk_mcu/u_ahb_ram/n16 ),
    .doa(\u_cmsdk_mcu/sram_hrdata [17:9]));
  // address_offset=0;data_offset=18;depth=1024;width=9;num_section=1;width_per_section=9;section_size=32;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("1"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("1"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("ASYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("READBEFOREWRITE"))
    \u_cmsdk_mcu/u_ahb_ram/ram_memory0_1024x32_sub_000000_018  (
    .addra({\u_cmsdk_mcu/HADDR [11:2],3'b111}),
    .addrb({\u_cmsdk_mcu/u_ahb_ram/buf_hwaddr [11:2],3'b111}),
    .clka(XTAL1_wire),
    .clkb(XTAL1_wire),
    .dia(9'b000000000),
    .dib(\u_cmsdk_mcu/u_ahb_ram/n13 [26:18]),
    .web(\u_cmsdk_mcu/u_ahb_ram/n16 ),
    .doa(\u_cmsdk_mcu/sram_hrdata [26:18]));
  // address_offset=0;data_offset=27;depth=1024;width=5;num_section=1;width_per_section=5;section_size=32;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("1"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("1"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("ASYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("READBEFOREWRITE"))
    \u_cmsdk_mcu/u_ahb_ram/ram_memory0_1024x32_sub_000000_027  (
    .addra({\u_cmsdk_mcu/HADDR [11:2],3'b111}),
    .addrb({\u_cmsdk_mcu/u_ahb_ram/buf_hwaddr [11:2],3'b111}),
    .clka(XTAL1_wire),
    .clkb(XTAL1_wire),
    .dia({open_n673,open_n674,open_n675,open_n676,5'b00000}),
    .dib({open_n677,open_n678,open_n679,open_n680,\u_cmsdk_mcu/u_ahb_ram/n13 [31:27]}),
    .web(\u_cmsdk_mcu/u_ahb_ram/n16 ),
    .doa({open_n686,open_n687,open_n688,open_n689,\u_cmsdk_mcu/sram_hrdata [31:27]}));
  reg_ar_as_w1 \u_cmsdk_mcu/u_ahb_ram/reg0_b10  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HADDR [10]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n11 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_ahb_ram/buf_hwaddr [10]));  // ../RTL/AHB2MEM.v(51)
  reg_ar_as_w1 \u_cmsdk_mcu/u_ahb_ram/reg0_b11  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HADDR [11]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n11 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_ahb_ram/buf_hwaddr [11]));  // ../RTL/AHB2MEM.v(51)
  reg_ar_as_w1 \u_cmsdk_mcu/u_ahb_ram/reg0_b12  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HADDR [12]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n11 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_ahb_ram/buf_hwaddr [12]));  // ../RTL/AHB2MEM.v(51)
  reg_ar_as_w1 \u_cmsdk_mcu/u_ahb_ram/reg0_b2  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HADDR [2]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n11 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_ahb_ram/buf_hwaddr [2]));  // ../RTL/AHB2MEM.v(51)
  reg_ar_as_w1 \u_cmsdk_mcu/u_ahb_ram/reg0_b3  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HADDR [3]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n11 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_ahb_ram/buf_hwaddr [3]));  // ../RTL/AHB2MEM.v(51)
  reg_ar_as_w1 \u_cmsdk_mcu/u_ahb_ram/reg0_b4  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HADDR [4]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n11 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_ahb_ram/buf_hwaddr [4]));  // ../RTL/AHB2MEM.v(51)
  reg_ar_as_w1 \u_cmsdk_mcu/u_ahb_ram/reg0_b5  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HADDR [5]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n11 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_ahb_ram/buf_hwaddr [5]));  // ../RTL/AHB2MEM.v(51)
  reg_ar_as_w1 \u_cmsdk_mcu/u_ahb_ram/reg0_b6  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HADDR [6]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n11 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_ahb_ram/buf_hwaddr [6]));  // ../RTL/AHB2MEM.v(51)
  reg_ar_as_w1 \u_cmsdk_mcu/u_ahb_ram/reg0_b7  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HADDR [7]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n11 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_ahb_ram/buf_hwaddr [7]));  // ../RTL/AHB2MEM.v(51)
  reg_ar_as_w1 \u_cmsdk_mcu/u_ahb_ram/reg0_b8  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HADDR [8]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n11 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_ahb_ram/buf_hwaddr [8]));  // ../RTL/AHB2MEM.v(51)
  reg_ar_as_w1 \u_cmsdk_mcu/u_ahb_ram/reg0_b9  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HADDR [9]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n11 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_ahb_ram/buf_hwaddr [9]));  // ../RTL/AHB2MEM.v(51)
  reg_ar_as_w1 \u_cmsdk_mcu/u_ahb_ram/reg1_b0  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_ahb_ram/n5 [0]),
    .en(\u_cmsdk_mcu/u_ahb_ram/mux3_b0_sel_is_2_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [0]));  // ../RTL/AHB2MEM.v(51)
  reg_ar_as_w1 \u_cmsdk_mcu/u_ahb_ram/reg1_b10  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_ahb_ram/n5 [10]),
    .en(\u_cmsdk_mcu/u_ahb_ram/mux3_b0_sel_is_2_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [10]));  // ../RTL/AHB2MEM.v(51)
  reg_ar_as_w1 \u_cmsdk_mcu/u_ahb_ram/reg1_b16  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_ahb_ram/n5 [16]),
    .en(\u_cmsdk_mcu/u_ahb_ram/mux3_b0_sel_is_2_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [16]));  // ../RTL/AHB2MEM.v(51)
  reg_ar_as_w1 \u_cmsdk_mcu/u_ahb_ram/reg1_b24  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_ahb_ram/n5 [24]),
    .en(\u_cmsdk_mcu/u_ahb_ram/mux3_b0_sel_is_2_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [24]));  // ../RTL/AHB2MEM.v(51)
  reg_ar_as_w1 \u_cmsdk_mcu/u_ahb_ram/we_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_ahb_ram/n2 ),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n11 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_ahb_ram/we ));  // ../RTL/AHB2MEM.v(51)
  // address_offset=0;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=32;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("1"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("1"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("ASYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("READBEFOREWRITE"))
    \u_cmsdk_mcu/u_ahb_rom/ram_memory0_1024x32_sub_000000_000  (
    .addra({\u_cmsdk_mcu/HADDR [11:2],3'b111}),
    .addrb({\u_cmsdk_mcu/u_ahb_ram/buf_hwaddr [11:2],3'b111}),
    .clka(XTAL1_wire),
    .clkb(XTAL1_wire),
    .dia(9'b000000000),
    .dib(\u_cmsdk_mcu/u_ahb_rom/n13 [8:0]),
    .web(\u_cmsdk_mcu/u_ahb_rom/n16 ),
    .doa(\u_cmsdk_mcu/flash_hrdata [8:0]));
  // address_offset=0;data_offset=9;depth=1024;width=9;num_section=1;width_per_section=9;section_size=32;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("1"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("1"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("ASYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("READBEFOREWRITE"))
    \u_cmsdk_mcu/u_ahb_rom/ram_memory0_1024x32_sub_000000_009  (
    .addra({\u_cmsdk_mcu/HADDR [11:2],3'b111}),
    .addrb({\u_cmsdk_mcu/u_ahb_ram/buf_hwaddr [11:2],3'b111}),
    .clka(XTAL1_wire),
    .clkb(XTAL1_wire),
    .dia(9'b000000000),
    .dib(\u_cmsdk_mcu/u_ahb_rom/n13 [17:9]),
    .web(\u_cmsdk_mcu/u_ahb_rom/n16 ),
    .doa(\u_cmsdk_mcu/flash_hrdata [17:9]));
  // address_offset=0;data_offset=18;depth=1024;width=9;num_section=1;width_per_section=9;section_size=32;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("1"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("1"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("ASYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("READBEFOREWRITE"))
    \u_cmsdk_mcu/u_ahb_rom/ram_memory0_1024x32_sub_000000_018  (
    .addra({\u_cmsdk_mcu/HADDR [11:2],3'b111}),
    .addrb({\u_cmsdk_mcu/u_ahb_ram/buf_hwaddr [11:2],3'b111}),
    .clka(XTAL1_wire),
    .clkb(XTAL1_wire),
    .dia(9'b000000000),
    .dib(\u_cmsdk_mcu/u_ahb_rom/n13 [26:18]),
    .web(\u_cmsdk_mcu/u_ahb_rom/n16 ),
    .doa(\u_cmsdk_mcu/flash_hrdata [26:18]));
  // address_offset=0;data_offset=27;depth=1024;width=5;num_section=1;width_per_section=5;section_size=32;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("1"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("1"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("ASYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("READBEFOREWRITE"))
    \u_cmsdk_mcu/u_ahb_rom/ram_memory0_1024x32_sub_000000_027  (
    .addra({\u_cmsdk_mcu/HADDR [11:2],3'b111}),
    .addrb({\u_cmsdk_mcu/u_ahb_ram/buf_hwaddr [11:2],3'b111}),
    .clka(XTAL1_wire),
    .clkb(XTAL1_wire),
    .dia({open_n773,open_n774,open_n775,open_n776,5'b00000}),
    .dib({open_n777,open_n778,open_n779,open_n780,\u_cmsdk_mcu/u_ahb_rom/n13 [31:27]}),
    .web(\u_cmsdk_mcu/u_ahb_rom/n16 ),
    .doa({open_n786,open_n787,open_n788,open_n789,\u_cmsdk_mcu/flash_hrdata [31:27]}));
  reg_ar_as_w1 \u_cmsdk_mcu/u_ahb_rom/we_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_ahb_rom/n2 ),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n11 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_ahb_rom/we ));  // ../RTL/AHB2MEM.v(51)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/dbgrst_reg_reg  (
    .clk(XTAL1_wire),
    .d(1'b1),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/reset_sync_reg [2]),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/dbgrst_reg ));  // ../RTL/cmsdk_mcu_clkctrl.v(108)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/nxt_hrst ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/reset_sync_reg [2]),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ));  // ../RTL/cmsdk_mcu_clkctrl.v(119)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/reg0_b0  (
    .clk(XTAL1_wire),
    .d(1'b1),
    .en(1'b1),
    .reset(~NRST_pad),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/reset_sync_reg [0]));  // ../RTL/cmsdk_mcu_clkctrl.v(86)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/reg0_b1  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/reset_sync_reg [0]),
    .en(1'b1),
    .reset(~NRST_pad),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/reset_sync_reg [1]));  // ../RTL/cmsdk_mcu_clkctrl.v(86)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/reg0_b2  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/reset_sync_reg [1]),
    .en(1'b1),
    .reset(~NRST_pad),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/reset_sync_reg [2]));  // ../RTL/cmsdk_mcu_clkctrl.v(86)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_ahb_to_gpio/IOSEL_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_ahb_to_gpio/n0 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOSEL ));  // ../RTL/cmsdk_ahb_to_iop.v(69)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_ahb_to_gpio/IOTRANS_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HTRANS [1]),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOTRANS ));  // ../RTL/cmsdk_ahb_to_iop.v(105)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_ahb_to_gpio/IOWRITE_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWRITE ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOWRITE ));  // ../RTL/cmsdk_ahb_to_iop.v(87)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_ahb_to_gpio/reg0_b0  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HADDR [0]),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [0]));  // ../RTL/cmsdk_ahb_to_iop.v(78)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_ahb_to_gpio/reg0_b1  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HADDR [1]),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [1]));  // ../RTL/cmsdk_ahb_to_iop.v(78)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_ahb_to_gpio/reg0_b10  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HADDR [10]),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [10]));  // ../RTL/cmsdk_ahb_to_iop.v(78)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_ahb_to_gpio/reg0_b11  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HADDR [11]),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [11]));  // ../RTL/cmsdk_ahb_to_iop.v(78)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_ahb_to_gpio/reg0_b2  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HADDR [2]),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]));  // ../RTL/cmsdk_ahb_to_iop.v(78)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_ahb_to_gpio/reg0_b3  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HADDR [3]),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]));  // ../RTL/cmsdk_ahb_to_iop.v(78)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_ahb_to_gpio/reg0_b4  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HADDR [4]),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4]));  // ../RTL/cmsdk_ahb_to_iop.v(78)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_ahb_to_gpio/reg0_b5  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HADDR [5]),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [5]));  // ../RTL/cmsdk_ahb_to_iop.v(78)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_ahb_to_gpio/reg0_b6  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HADDR [6]),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [6]));  // ../RTL/cmsdk_ahb_to_iop.v(78)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_ahb_to_gpio/reg0_b7  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HADDR [7]),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [7]));  // ../RTL/cmsdk_ahb_to_iop.v(78)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_ahb_to_gpio/reg0_b8  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HADDR [8]),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [8]));  // ../RTL/cmsdk_ahb_to_iop.v(78)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_ahb_to_gpio/reg0_b9  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HADDR [9]),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [9]));  // ../RTL/cmsdk_ahb_to_iop.v(78)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_ahb_to_gpio/reg1_b0  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HSIZE [0]),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOSIZE [0]));  // ../RTL/cmsdk_ahb_to_iop.v(96)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_ahb_to_gpio/reg1_b1  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HSIZE [1]),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOSIZE [1]));  // ../RTL/cmsdk_ahb_to_iop.v(96)
  AL_MAP_LUT4 #(
    .EQN("(~A*B*~C*D+~A*~B*C*D+~A*B*C*D+A*B*C*D)"),
    .INIT(16'b1101010000000000))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/mux2_b0_rom0  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [5]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n13 [0]));
  AL_MAP_LUT4 #(
    .EQN("(~A*~B*C*~D+~A*~B*C*D+~A*B*C*D)"),
    .INIT(16'b0101000000010000))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/mux2_b2_rom0  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [5]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n13 [2]));
  AL_MAP_LUT4 #(
    .EQN("(A*~B*~C*D+~A*B*~C*D+~A*~B*C*D)"),
    .INIT(16'b0001011000000000))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/mux2_b3_rom0  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [5]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n13 [3]));
  AL_MAP_LUT4 #(
    .EQN("(A*~B*~C*D+~A*B*~C*D+A*~B*C*D+A*B*C*D)"),
    .INIT(16'b1010011000000000))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/mux2_b4_rom0  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [5]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n13 [4]));
  AL_MAP_LUT4 #(
    .EQN("(~A*~B*~C*D+A*~B*~C*D+A*~B*C*D+A*B*C*D)"),
    .INIT(16'b1010001100000000))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/mux2_b5_rom0  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [5]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n13 [5]));
  AL_MAP_LUT4 #(
    .EQN("(A*~B*~C*D+A*~B*C*D+A*B*C*D)"),
    .INIT(16'b1010001000000000))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/mux2_b7_rom0  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [5]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n13 [7]));
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg1_b0  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/nxt_dout_padded [0]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n34 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/p0_out [0]));  // ../RTL/cmsdk_iop_gpio.v(309)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg1_b1  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/nxt_dout_padded [1]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n34 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/p0_out [1]));  // ../RTL/cmsdk_iop_gpio.v(309)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg1_b10  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/nxt_dout_padded [10]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n39 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/p0_out [10]));  // ../RTL/cmsdk_iop_gpio.v(309)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg1_b11  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/nxt_dout_padded [11]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n39 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/p0_out [11]));  // ../RTL/cmsdk_iop_gpio.v(309)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg1_b12  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/nxt_dout_padded [12]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n39 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/p0_out [12]));  // ../RTL/cmsdk_iop_gpio.v(309)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg1_b13  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/nxt_dout_padded [13]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n39 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/p0_out [13]));  // ../RTL/cmsdk_iop_gpio.v(309)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg1_b14  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/nxt_dout_padded [14]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n39 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/p0_out [14]));  // ../RTL/cmsdk_iop_gpio.v(309)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg1_b15  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/nxt_dout_padded [15]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n39 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/p0_out [15]));  // ../RTL/cmsdk_iop_gpio.v(309)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg1_b2  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/nxt_dout_padded [2]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n34 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/p0_out [2]));  // ../RTL/cmsdk_iop_gpio.v(309)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg1_b3  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/nxt_dout_padded [3]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n34 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/p0_out [3]));  // ../RTL/cmsdk_iop_gpio.v(309)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg1_b4  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/nxt_dout_padded [4]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n34 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/p0_out [4]));  // ../RTL/cmsdk_iop_gpio.v(309)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg1_b5  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/nxt_dout_padded [5]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n34 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/p0_out [5]));  // ../RTL/cmsdk_iop_gpio.v(309)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg1_b6  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/nxt_dout_padded [6]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n34 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/p0_out [6]));  // ../RTL/cmsdk_iop_gpio.v(309)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg1_b7  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/nxt_dout_padded [7]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n34 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/p0_out [7]));  // ../RTL/cmsdk_iop_gpio.v(309)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg1_b8  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/nxt_dout_padded [8]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n39 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/p0_out [8]));  // ../RTL/cmsdk_iop_gpio.v(309)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg1_b9  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/nxt_dout_padded [9]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n39 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/p0_out [9]));  // ../RTL/cmsdk_iop_gpio.v(309)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg2_b0  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_doutenset [0]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n54 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/p0_outen [0]));  // ../RTL/cmsdk_iop_gpio.v(348)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg2_b1  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_doutenset [1]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n56 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/p0_outen [1]));  // ../RTL/cmsdk_iop_gpio.v(348)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg2_b10  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_doutenset [10]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n74 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/p0_outen [10]));  // ../RTL/cmsdk_iop_gpio.v(348)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg2_b11  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_doutenset [11]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n76 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/p0_outen [11]));  // ../RTL/cmsdk_iop_gpio.v(348)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg2_b12  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_doutenset [12]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n78 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/p0_outen [12]));  // ../RTL/cmsdk_iop_gpio.v(348)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg2_b13  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_doutenset [13]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n80 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/p0_outen [13]));  // ../RTL/cmsdk_iop_gpio.v(348)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg2_b14  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_doutenset [14]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n82 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/p0_outen [14]));  // ../RTL/cmsdk_iop_gpio.v(348)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg2_b15  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_doutenset [15]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n84 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/p0_outen [15]));  // ../RTL/cmsdk_iop_gpio.v(348)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg2_b2  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_doutenset [2]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n58 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/p0_outen [2]));  // ../RTL/cmsdk_iop_gpio.v(348)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg2_b3  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_doutenset [3]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n60 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/p0_outen [3]));  // ../RTL/cmsdk_iop_gpio.v(348)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg2_b4  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_doutenset [4]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n62 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/p0_outen [4]));  // ../RTL/cmsdk_iop_gpio.v(348)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg2_b5  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_doutenset [5]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n64 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/p0_outen [5]));  // ../RTL/cmsdk_iop_gpio.v(348)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg2_b6  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_doutenset [6]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n66 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/p0_outen [6]));  // ../RTL/cmsdk_iop_gpio.v(348)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg2_b7  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_doutenset [7]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n68 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/p0_outen [7]));  // ../RTL/cmsdk_iop_gpio.v(348)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg2_b8  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_doutenset [8]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n70 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/p0_outen [8]));  // ../RTL/cmsdk_iop_gpio.v(348)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg2_b9  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_doutenset [9]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n72 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/p0_outen [9]));  // ../RTL/cmsdk_iop_gpio.v(348)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg3_b0  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_altfuncset [0]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n99 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/p0_altfunc [0]));  // ../RTL/cmsdk_iop_gpio.v(387)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg3_b1  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_altfuncset [1]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n101 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/p0_altfunc [1]));  // ../RTL/cmsdk_iop_gpio.v(387)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg3_b10  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_altfuncset [10]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n119 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/p0_altfunc [10]));  // ../RTL/cmsdk_iop_gpio.v(387)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg3_b11  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_altfuncset [11]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n121 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/p0_altfunc [11]));  // ../RTL/cmsdk_iop_gpio.v(387)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg3_b12  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_altfuncset [12]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n123 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/p0_altfunc [12]));  // ../RTL/cmsdk_iop_gpio.v(387)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg3_b13  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_altfuncset [13]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n125 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/p0_altfunc [13]));  // ../RTL/cmsdk_iop_gpio.v(387)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg3_b14  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_altfuncset [14]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n127 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/p0_altfunc [14]));  // ../RTL/cmsdk_iop_gpio.v(387)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg3_b15  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_altfuncset [15]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n129 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/p0_altfunc [15]));  // ../RTL/cmsdk_iop_gpio.v(387)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg3_b2  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_altfuncset [2]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n103 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/p0_altfunc [2]));  // ../RTL/cmsdk_iop_gpio.v(387)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg3_b3  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_altfuncset [3]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n105 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/p0_altfunc [3]));  // ../RTL/cmsdk_iop_gpio.v(387)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg3_b4  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_altfuncset [4]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n107 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/p0_altfunc [4]));  // ../RTL/cmsdk_iop_gpio.v(387)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg3_b5  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_altfuncset [5]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n109 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/p0_altfunc [5]));  // ../RTL/cmsdk_iop_gpio.v(387)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg3_b6  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_altfuncset [6]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n111 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/p0_altfunc [6]));  // ../RTL/cmsdk_iop_gpio.v(387)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg3_b7  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_altfuncset [7]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n113 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/p0_altfunc [7]));  // ../RTL/cmsdk_iop_gpio.v(387)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg3_b8  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_altfuncset [8]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n115 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/p0_altfunc [8]));  // ../RTL/cmsdk_iop_gpio.v(387)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg3_b9  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_altfuncset [9]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n117 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/p0_altfunc [9]));  // ../RTL/cmsdk_iop_gpio.v(387)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg4_b0  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intenset [0]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n144 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inten_padded [0]));  // ../RTL/cmsdk_iop_gpio.v(425)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg4_b1  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intenset [1]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n146 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inten_padded [1]));  // ../RTL/cmsdk_iop_gpio.v(425)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg4_b10  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intenset [10]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n164 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inten_padded [10]));  // ../RTL/cmsdk_iop_gpio.v(425)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg4_b11  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intenset [11]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n166 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inten_padded [11]));  // ../RTL/cmsdk_iop_gpio.v(425)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg4_b12  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intenset [12]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n168 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inten_padded [12]));  // ../RTL/cmsdk_iop_gpio.v(425)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg4_b13  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intenset [13]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n170 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inten_padded [13]));  // ../RTL/cmsdk_iop_gpio.v(425)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg4_b14  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intenset [14]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n172 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inten_padded [14]));  // ../RTL/cmsdk_iop_gpio.v(425)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg4_b15  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intenset [15]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n174 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inten_padded [15]));  // ../RTL/cmsdk_iop_gpio.v(425)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg4_b2  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intenset [2]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n148 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inten_padded [2]));  // ../RTL/cmsdk_iop_gpio.v(425)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg4_b3  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intenset [3]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n150 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inten_padded [3]));  // ../RTL/cmsdk_iop_gpio.v(425)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg4_b4  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intenset [4]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n152 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inten_padded [4]));  // ../RTL/cmsdk_iop_gpio.v(425)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg4_b5  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intenset [5]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n154 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inten_padded [5]));  // ../RTL/cmsdk_iop_gpio.v(425)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg4_b6  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intenset [6]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n156 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inten_padded [6]));  // ../RTL/cmsdk_iop_gpio.v(425)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg4_b7  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intenset [7]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n158 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inten_padded [7]));  // ../RTL/cmsdk_iop_gpio.v(425)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg4_b8  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intenset [8]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n160 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inten_padded [8]));  // ../RTL/cmsdk_iop_gpio.v(425)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg4_b9  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intenset [9]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n162 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inten_padded [9]));  // ../RTL/cmsdk_iop_gpio.v(425)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg5_b0  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttypeset [0]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n189 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttype_padded [0]));  // ../RTL/cmsdk_iop_gpio.v(463)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg5_b1  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttypeset [1]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n191 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttype_padded [1]));  // ../RTL/cmsdk_iop_gpio.v(463)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg5_b10  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttypeset [10]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n209 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttype_padded [10]));  // ../RTL/cmsdk_iop_gpio.v(463)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg5_b11  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttypeset [11]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n211 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttype_padded [11]));  // ../RTL/cmsdk_iop_gpio.v(463)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg5_b12  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttypeset [12]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n213 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttype_padded [12]));  // ../RTL/cmsdk_iop_gpio.v(463)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg5_b13  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttypeset [13]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n215 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttype_padded [13]));  // ../RTL/cmsdk_iop_gpio.v(463)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg5_b14  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttypeset [14]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n217 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttype_padded [14]));  // ../RTL/cmsdk_iop_gpio.v(463)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg5_b15  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttypeset [15]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n219 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttype_padded [15]));  // ../RTL/cmsdk_iop_gpio.v(463)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg5_b2  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttypeset [2]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n193 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttype_padded [2]));  // ../RTL/cmsdk_iop_gpio.v(463)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg5_b3  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttypeset [3]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n195 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttype_padded [3]));  // ../RTL/cmsdk_iop_gpio.v(463)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg5_b4  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttypeset [4]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n197 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttype_padded [4]));  // ../RTL/cmsdk_iop_gpio.v(463)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg5_b5  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttypeset [5]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n199 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttype_padded [5]));  // ../RTL/cmsdk_iop_gpio.v(463)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg5_b6  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttypeset [6]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n201 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttype_padded [6]));  // ../RTL/cmsdk_iop_gpio.v(463)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg5_b7  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttypeset [7]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n203 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttype_padded [7]));  // ../RTL/cmsdk_iop_gpio.v(463)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg5_b8  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttypeset [8]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n205 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttype_padded [8]));  // ../RTL/cmsdk_iop_gpio.v(463)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg5_b9  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttypeset [9]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n207 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttype_padded [9]));  // ../RTL/cmsdk_iop_gpio.v(463)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg6_b0  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpolset [0]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n234 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpol_padded [0]));  // ../RTL/cmsdk_iop_gpio.v(501)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg6_b1  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpolset [1]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n236 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpol_padded [1]));  // ../RTL/cmsdk_iop_gpio.v(501)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg6_b10  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpolset [10]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n254 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpol_padded [10]));  // ../RTL/cmsdk_iop_gpio.v(501)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg6_b11  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpolset [11]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n256 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpol_padded [11]));  // ../RTL/cmsdk_iop_gpio.v(501)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg6_b12  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpolset [12]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n258 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpol_padded [12]));  // ../RTL/cmsdk_iop_gpio.v(501)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg6_b13  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpolset [13]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n260 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpol_padded [13]));  // ../RTL/cmsdk_iop_gpio.v(501)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg6_b14  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpolset [14]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n262 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpol_padded [14]));  // ../RTL/cmsdk_iop_gpio.v(501)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg6_b15  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpolset [15]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n264 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpol_padded [15]));  // ../RTL/cmsdk_iop_gpio.v(501)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg6_b2  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpolset [2]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n238 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpol_padded [2]));  // ../RTL/cmsdk_iop_gpio.v(501)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg6_b3  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpolset [3]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n240 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpol_padded [3]));  // ../RTL/cmsdk_iop_gpio.v(501)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg6_b4  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpolset [4]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n242 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpol_padded [4]));  // ../RTL/cmsdk_iop_gpio.v(501)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg6_b5  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpolset [5]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n244 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpol_padded [5]));  // ../RTL/cmsdk_iop_gpio.v(501)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg6_b6  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpolset [6]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n246 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpol_padded [6]));  // ../RTL/cmsdk_iop_gpio.v(501)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg6_b7  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpolset [7]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n248 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpol_padded [7]));  // ../RTL/cmsdk_iop_gpio.v(501)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg6_b8  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpolset [8]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n250 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpol_padded [8]));  // ../RTL/cmsdk_iop_gpio.v(501)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg6_b9  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpolset [9]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n252 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpol_padded [9]));  // ../RTL/cmsdk_iop_gpio.v(501)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg7_b0  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/new_masked_int [0]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n271 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [0]));  // ../RTL/cmsdk_iop_gpio.v(539)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg7_b1  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/new_masked_int [1]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n273 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [1]));  // ../RTL/cmsdk_iop_gpio.v(539)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg7_b10  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/new_masked_int [10]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n291 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [10]));  // ../RTL/cmsdk_iop_gpio.v(539)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg7_b11  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/new_masked_int [11]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n293 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [11]));  // ../RTL/cmsdk_iop_gpio.v(539)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg7_b12  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/new_masked_int [12]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n295 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [12]));  // ../RTL/cmsdk_iop_gpio.v(539)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg7_b13  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/new_masked_int [13]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n297 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [13]));  // ../RTL/cmsdk_iop_gpio.v(539)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg7_b14  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/new_masked_int [14]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n299 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [14]));  // ../RTL/cmsdk_iop_gpio.v(539)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg7_b15  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/new_masked_int [15]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n301 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [15]));  // ../RTL/cmsdk_iop_gpio.v(539)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg7_b2  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/new_masked_int [2]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n275 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [2]));  // ../RTL/cmsdk_iop_gpio.v(539)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg7_b3  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/new_masked_int [3]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n277 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [3]));  // ../RTL/cmsdk_iop_gpio.v(539)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg7_b4  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/new_masked_int [4]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n279 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [4]));  // ../RTL/cmsdk_iop_gpio.v(539)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg7_b5  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/new_masked_int [5]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n281 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [5]));  // ../RTL/cmsdk_iop_gpio.v(539)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg7_b6  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/new_masked_int [6]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n283 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [6]));  // ../RTL/cmsdk_iop_gpio.v(539)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg7_b7  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/new_masked_int [7]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n285 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [7]));  // ../RTL/cmsdk_iop_gpio.v(539)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg7_b8  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/new_masked_int [8]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n287 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [8]));  // ../RTL/cmsdk_iop_gpio.v(539)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg7_b9  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/new_masked_int [9]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n289 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [9]));  // ../RTL/cmsdk_iop_gpio.v(539)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_ahb_to_gpio/IOSEL_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_ahb_to_gpio/n0 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/IOSEL ));  // ../RTL/cmsdk_ahb_to_iop.v(69)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg0_b0  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync1 [0]),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [0]));  // ../RTL/cmsdk_iop_gpio.v(252)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg0_b1  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync1 [1]),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [1]));  // ../RTL/cmsdk_iop_gpio.v(252)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg0_b10  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync1 [10]),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [10]));  // ../RTL/cmsdk_iop_gpio.v(252)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg0_b11  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync1 [11]),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [11]));  // ../RTL/cmsdk_iop_gpio.v(252)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg0_b12  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync1 [12]),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [12]));  // ../RTL/cmsdk_iop_gpio.v(252)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg0_b13  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync1 [13]),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [13]));  // ../RTL/cmsdk_iop_gpio.v(252)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg0_b14  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync1 [14]),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [14]));  // ../RTL/cmsdk_iop_gpio.v(252)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg0_b15  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync1 [15]),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [15]));  // ../RTL/cmsdk_iop_gpio.v(252)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg0_b2  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync1 [2]),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [2]));  // ../RTL/cmsdk_iop_gpio.v(252)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg0_b3  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync1 [3]),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [3]));  // ../RTL/cmsdk_iop_gpio.v(252)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg0_b4  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync1 [4]),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [4]));  // ../RTL/cmsdk_iop_gpio.v(252)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg0_b5  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync1 [5]),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [5]));  // ../RTL/cmsdk_iop_gpio.v(252)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg0_b6  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync1 [6]),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [6]));  // ../RTL/cmsdk_iop_gpio.v(252)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg0_b7  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync1 [7]),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [7]));  // ../RTL/cmsdk_iop_gpio.v(252)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg0_b8  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync1 [8]),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [8]));  // ../RTL/cmsdk_iop_gpio.v(252)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg0_b9  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync1 [9]),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [9]));  // ../RTL/cmsdk_iop_gpio.v(252)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg1_b0  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/nxt_dout_padded [0]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n34 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/p1_out [0]));  // ../RTL/cmsdk_iop_gpio.v(309)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg1_b1  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/nxt_dout_padded [1]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n34 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/p1_out [1]));  // ../RTL/cmsdk_iop_gpio.v(309)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg1_b10  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/nxt_dout_padded [10]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n39 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/p1_out [10]));  // ../RTL/cmsdk_iop_gpio.v(309)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg1_b11  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/nxt_dout_padded [11]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n39 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/p1_out [11]));  // ../RTL/cmsdk_iop_gpio.v(309)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg1_b12  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/nxt_dout_padded [12]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n39 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/p1_out [12]));  // ../RTL/cmsdk_iop_gpio.v(309)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg1_b13  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/nxt_dout_padded [13]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n39 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/p1_out [13]));  // ../RTL/cmsdk_iop_gpio.v(309)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg1_b14  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/nxt_dout_padded [14]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n39 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/p1_out [14]));  // ../RTL/cmsdk_iop_gpio.v(309)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg1_b15  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/nxt_dout_padded [15]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n39 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/p1_out [15]));  // ../RTL/cmsdk_iop_gpio.v(309)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg1_b2  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/nxt_dout_padded [2]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n34 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/p1_out [2]));  // ../RTL/cmsdk_iop_gpio.v(309)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg1_b3  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/nxt_dout_padded [3]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n34 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/p1_out [3]));  // ../RTL/cmsdk_iop_gpio.v(309)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg1_b4  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/nxt_dout_padded [4]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n34 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/p1_out [4]));  // ../RTL/cmsdk_iop_gpio.v(309)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg1_b5  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/nxt_dout_padded [5]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n34 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/p1_out [5]));  // ../RTL/cmsdk_iop_gpio.v(309)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg1_b6  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/nxt_dout_padded [6]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n34 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/p1_out [6]));  // ../RTL/cmsdk_iop_gpio.v(309)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg1_b7  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/nxt_dout_padded [7]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n34 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/p1_out [7]));  // ../RTL/cmsdk_iop_gpio.v(309)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg1_b8  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/nxt_dout_padded [8]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n39 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/p1_out [8]));  // ../RTL/cmsdk_iop_gpio.v(309)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg1_b9  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/nxt_dout_padded [9]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n39 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/p1_out [9]));  // ../RTL/cmsdk_iop_gpio.v(309)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg2_b0  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_doutenset [0]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n54 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/p1_outen [0]));  // ../RTL/cmsdk_iop_gpio.v(348)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg2_b1  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_doutenset [1]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n56 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/p1_outen [1]));  // ../RTL/cmsdk_iop_gpio.v(348)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg2_b10  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_doutenset [10]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n74 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/p1_outen [10]));  // ../RTL/cmsdk_iop_gpio.v(348)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg2_b11  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_doutenset [11]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n76 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/p1_outen [11]));  // ../RTL/cmsdk_iop_gpio.v(348)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg2_b12  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_doutenset [12]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n78 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/p1_outen [12]));  // ../RTL/cmsdk_iop_gpio.v(348)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg2_b13  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_doutenset [13]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n80 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/p1_outen [13]));  // ../RTL/cmsdk_iop_gpio.v(348)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg2_b14  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_doutenset [14]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n82 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/p1_outen [14]));  // ../RTL/cmsdk_iop_gpio.v(348)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg2_b15  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_doutenset [15]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n84 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/p1_outen [15]));  // ../RTL/cmsdk_iop_gpio.v(348)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg2_b2  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_doutenset [2]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n58 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/p1_outen [2]));  // ../RTL/cmsdk_iop_gpio.v(348)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg2_b3  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_doutenset [3]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n60 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/p1_outen [3]));  // ../RTL/cmsdk_iop_gpio.v(348)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg2_b4  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_doutenset [4]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n62 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/p1_outen [4]));  // ../RTL/cmsdk_iop_gpio.v(348)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg2_b5  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_doutenset [5]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n64 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/p1_outen [5]));  // ../RTL/cmsdk_iop_gpio.v(348)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg2_b6  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_doutenset [6]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n66 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/p1_outen [6]));  // ../RTL/cmsdk_iop_gpio.v(348)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg2_b7  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_doutenset [7]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n68 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/p1_outen [7]));  // ../RTL/cmsdk_iop_gpio.v(348)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg2_b8  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_doutenset [8]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n70 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/p1_outen [8]));  // ../RTL/cmsdk_iop_gpio.v(348)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg2_b9  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_doutenset [9]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n72 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/p1_outen [9]));  // ../RTL/cmsdk_iop_gpio.v(348)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg3_b0  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_altfuncset [0]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n99 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/p1_altfunc [0]));  // ../RTL/cmsdk_iop_gpio.v(387)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg3_b1  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_altfuncset [1]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n101 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/p1_altfunc [1]));  // ../RTL/cmsdk_iop_gpio.v(387)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg3_b10  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_altfuncset [10]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n119 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/p1_altfunc [10]));  // ../RTL/cmsdk_iop_gpio.v(387)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg3_b11  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_altfuncset [11]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n121 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/p1_altfunc [11]));  // ../RTL/cmsdk_iop_gpio.v(387)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg3_b12  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_altfuncset [12]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n123 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/p1_altfunc [12]));  // ../RTL/cmsdk_iop_gpio.v(387)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg3_b13  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_altfuncset [13]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n125 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/p1_altfunc [13]));  // ../RTL/cmsdk_iop_gpio.v(387)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg3_b14  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_altfuncset [14]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n127 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/p1_altfunc [14]));  // ../RTL/cmsdk_iop_gpio.v(387)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg3_b15  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_altfuncset [15]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n129 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/p1_altfunc [15]));  // ../RTL/cmsdk_iop_gpio.v(387)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg3_b2  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_altfuncset [2]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n103 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/p1_altfunc [2]));  // ../RTL/cmsdk_iop_gpio.v(387)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg3_b3  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_altfuncset [3]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n105 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/p1_altfunc [3]));  // ../RTL/cmsdk_iop_gpio.v(387)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg3_b4  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_altfuncset [4]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n107 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/p1_altfunc [4]));  // ../RTL/cmsdk_iop_gpio.v(387)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg3_b5  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_altfuncset [5]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n109 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/p1_altfunc [5]));  // ../RTL/cmsdk_iop_gpio.v(387)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg3_b6  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_altfuncset [6]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n111 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/p1_altfunc [6]));  // ../RTL/cmsdk_iop_gpio.v(387)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg3_b7  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_altfuncset [7]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n113 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/p1_altfunc [7]));  // ../RTL/cmsdk_iop_gpio.v(387)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg3_b8  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_altfuncset [8]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n115 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/p1_altfunc [8]));  // ../RTL/cmsdk_iop_gpio.v(387)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg3_b9  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_altfuncset [9]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n117 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/p1_altfunc [9]));  // ../RTL/cmsdk_iop_gpio.v(387)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg4_b0  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intenset [0]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n144 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inten_padded [0]));  // ../RTL/cmsdk_iop_gpio.v(425)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg4_b1  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intenset [1]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n146 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inten_padded [1]));  // ../RTL/cmsdk_iop_gpio.v(425)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg4_b10  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intenset [10]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n164 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inten_padded [10]));  // ../RTL/cmsdk_iop_gpio.v(425)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg4_b11  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intenset [11]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n166 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inten_padded [11]));  // ../RTL/cmsdk_iop_gpio.v(425)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg4_b12  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intenset [12]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n168 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inten_padded [12]));  // ../RTL/cmsdk_iop_gpio.v(425)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg4_b13  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intenset [13]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n170 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inten_padded [13]));  // ../RTL/cmsdk_iop_gpio.v(425)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg4_b14  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intenset [14]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n172 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inten_padded [14]));  // ../RTL/cmsdk_iop_gpio.v(425)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg4_b15  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intenset [15]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n174 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inten_padded [15]));  // ../RTL/cmsdk_iop_gpio.v(425)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg4_b2  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intenset [2]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n148 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inten_padded [2]));  // ../RTL/cmsdk_iop_gpio.v(425)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg4_b3  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intenset [3]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n150 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inten_padded [3]));  // ../RTL/cmsdk_iop_gpio.v(425)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg4_b4  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intenset [4]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n152 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inten_padded [4]));  // ../RTL/cmsdk_iop_gpio.v(425)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg4_b5  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intenset [5]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n154 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inten_padded [5]));  // ../RTL/cmsdk_iop_gpio.v(425)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg4_b6  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intenset [6]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n156 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inten_padded [6]));  // ../RTL/cmsdk_iop_gpio.v(425)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg4_b7  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intenset [7]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n158 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inten_padded [7]));  // ../RTL/cmsdk_iop_gpio.v(425)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg4_b8  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intenset [8]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n160 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inten_padded [8]));  // ../RTL/cmsdk_iop_gpio.v(425)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg4_b9  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intenset [9]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n162 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inten_padded [9]));  // ../RTL/cmsdk_iop_gpio.v(425)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg5_b0  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttypeset [0]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n189 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [0]));  // ../RTL/cmsdk_iop_gpio.v(463)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg5_b1  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttypeset [1]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n191 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [1]));  // ../RTL/cmsdk_iop_gpio.v(463)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg5_b10  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttypeset [10]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n209 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [10]));  // ../RTL/cmsdk_iop_gpio.v(463)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg5_b11  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttypeset [11]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n211 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [11]));  // ../RTL/cmsdk_iop_gpio.v(463)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg5_b12  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttypeset [12]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n213 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [12]));  // ../RTL/cmsdk_iop_gpio.v(463)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg5_b13  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttypeset [13]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n215 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [13]));  // ../RTL/cmsdk_iop_gpio.v(463)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg5_b14  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttypeset [14]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n217 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [14]));  // ../RTL/cmsdk_iop_gpio.v(463)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg5_b15  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttypeset [15]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n219 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [15]));  // ../RTL/cmsdk_iop_gpio.v(463)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg5_b2  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttypeset [2]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n193 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [2]));  // ../RTL/cmsdk_iop_gpio.v(463)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg5_b3  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttypeset [3]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n195 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [3]));  // ../RTL/cmsdk_iop_gpio.v(463)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg5_b4  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttypeset [4]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n197 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [4]));  // ../RTL/cmsdk_iop_gpio.v(463)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg5_b5  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttypeset [5]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n199 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [5]));  // ../RTL/cmsdk_iop_gpio.v(463)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg5_b6  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttypeset [6]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n201 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [6]));  // ../RTL/cmsdk_iop_gpio.v(463)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg5_b7  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttypeset [7]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n203 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [7]));  // ../RTL/cmsdk_iop_gpio.v(463)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg5_b8  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttypeset [8]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n205 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [8]));  // ../RTL/cmsdk_iop_gpio.v(463)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg5_b9  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttypeset [9]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n207 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [9]));  // ../RTL/cmsdk_iop_gpio.v(463)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg6_b0  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpolset [0]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n234 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpol_padded [0]));  // ../RTL/cmsdk_iop_gpio.v(501)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg6_b1  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpolset [1]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n236 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpol_padded [1]));  // ../RTL/cmsdk_iop_gpio.v(501)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg6_b10  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpolset [10]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n254 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpol_padded [10]));  // ../RTL/cmsdk_iop_gpio.v(501)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg6_b11  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpolset [11]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n256 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpol_padded [11]));  // ../RTL/cmsdk_iop_gpio.v(501)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg6_b12  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpolset [12]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n258 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpol_padded [12]));  // ../RTL/cmsdk_iop_gpio.v(501)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg6_b13  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpolset [13]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n260 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpol_padded [13]));  // ../RTL/cmsdk_iop_gpio.v(501)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg6_b14  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpolset [14]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n262 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpol_padded [14]));  // ../RTL/cmsdk_iop_gpio.v(501)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg6_b15  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpolset [15]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n264 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpol_padded [15]));  // ../RTL/cmsdk_iop_gpio.v(501)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg6_b2  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpolset [2]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n238 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpol_padded [2]));  // ../RTL/cmsdk_iop_gpio.v(501)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg6_b3  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpolset [3]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n240 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpol_padded [3]));  // ../RTL/cmsdk_iop_gpio.v(501)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg6_b4  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpolset [4]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n242 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpol_padded [4]));  // ../RTL/cmsdk_iop_gpio.v(501)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg6_b5  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpolset [5]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n244 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpol_padded [5]));  // ../RTL/cmsdk_iop_gpio.v(501)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg6_b6  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpolset [6]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n246 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpol_padded [6]));  // ../RTL/cmsdk_iop_gpio.v(501)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg6_b7  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpolset [7]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n248 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpol_padded [7]));  // ../RTL/cmsdk_iop_gpio.v(501)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg6_b8  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpolset [8]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n250 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpol_padded [8]));  // ../RTL/cmsdk_iop_gpio.v(501)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg6_b9  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpolset [9]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n252 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpol_padded [9]));  // ../RTL/cmsdk_iop_gpio.v(501)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg7_b0  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_masked_int [0]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n271 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[0] ));  // ../RTL/cmsdk_iop_gpio.v(539)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg7_b1  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_masked_int [1]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n273 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[1] ));  // ../RTL/cmsdk_iop_gpio.v(539)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg7_b10  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_masked_int [10]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n291 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[10] ));  // ../RTL/cmsdk_iop_gpio.v(539)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg7_b11  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_masked_int [11]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n293 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[11] ));  // ../RTL/cmsdk_iop_gpio.v(539)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg7_b12  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_masked_int [12]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n295 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[12] ));  // ../RTL/cmsdk_iop_gpio.v(539)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg7_b13  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_masked_int [13]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n297 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[13] ));  // ../RTL/cmsdk_iop_gpio.v(539)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg7_b14  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_masked_int [14]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n299 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[14] ));  // ../RTL/cmsdk_iop_gpio.v(539)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg7_b15  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_masked_int [15]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n301 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[15] ));  // ../RTL/cmsdk_iop_gpio.v(539)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg7_b2  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_masked_int [2]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n275 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[2] ));  // ../RTL/cmsdk_iop_gpio.v(539)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg7_b3  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_masked_int [3]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n277 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[3] ));  // ../RTL/cmsdk_iop_gpio.v(539)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg7_b4  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_masked_int [4]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n279 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[4] ));  // ../RTL/cmsdk_iop_gpio.v(539)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg7_b5  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_masked_int [5]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n281 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[5] ));  // ../RTL/cmsdk_iop_gpio.v(539)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg7_b6  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_masked_int [6]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n283 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[6] ));  // ../RTL/cmsdk_iop_gpio.v(539)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg7_b7  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_masked_int [7]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n285 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[7] ));  // ../RTL/cmsdk_iop_gpio.v(539)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg7_b8  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_masked_int [8]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n287 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[8] ));  // ../RTL/cmsdk_iop_gpio.v(539)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg7_b9  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_masked_int [9]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n289 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[9] ));  // ../RTL/cmsdk_iop_gpio.v(539)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg8_b0  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [0]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n304 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_last_datain [0]));  // ../RTL/cmsdk_iop_gpio.v(561)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg8_b1  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [1]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n304 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_last_datain [1]));  // ../RTL/cmsdk_iop_gpio.v(561)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg8_b10  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [10]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n304 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_last_datain [10]));  // ../RTL/cmsdk_iop_gpio.v(561)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg8_b11  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [11]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n304 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_last_datain [11]));  // ../RTL/cmsdk_iop_gpio.v(561)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg8_b12  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [12]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n304 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_last_datain [12]));  // ../RTL/cmsdk_iop_gpio.v(561)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg8_b13  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [13]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n304 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_last_datain [13]));  // ../RTL/cmsdk_iop_gpio.v(561)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg8_b14  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [14]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n304 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_last_datain [14]));  // ../RTL/cmsdk_iop_gpio.v(561)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg8_b15  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [15]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n304 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_last_datain [15]));  // ../RTL/cmsdk_iop_gpio.v(561)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg8_b2  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [2]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n304 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_last_datain [2]));  // ../RTL/cmsdk_iop_gpio.v(561)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg8_b3  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [3]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n304 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_last_datain [3]));  // ../RTL/cmsdk_iop_gpio.v(561)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg8_b4  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [4]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n304 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_last_datain [4]));  // ../RTL/cmsdk_iop_gpio.v(561)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg8_b5  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [5]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n304 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_last_datain [5]));  // ../RTL/cmsdk_iop_gpio.v(561)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg8_b6  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [6]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n304 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_last_datain [6]));  // ../RTL/cmsdk_iop_gpio.v(561)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg8_b7  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [7]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n304 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_last_datain [7]));  // ../RTL/cmsdk_iop_gpio.v(561)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg8_b8  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [8]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n304 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_last_datain [8]));  // ../RTL/cmsdk_iop_gpio.v(561)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg8_b9  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [9]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n304 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_last_datain [9]));  // ../RTL/cmsdk_iop_gpio.v(561)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg9_b0  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/p1_in [0]),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync1 [0]));  // ../RTL/cmsdk_iop_gpio.v(252)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg9_b1  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/p1_in [1]),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync1 [1]));  // ../RTL/cmsdk_iop_gpio.v(252)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg9_b10  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/p1_in [10]),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync1 [10]));  // ../RTL/cmsdk_iop_gpio.v(252)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg9_b11  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/p1_in [11]),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync1 [11]));  // ../RTL/cmsdk_iop_gpio.v(252)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg9_b12  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/p1_in [12]),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync1 [12]));  // ../RTL/cmsdk_iop_gpio.v(252)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg9_b13  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/p1_in [13]),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync1 [13]));  // ../RTL/cmsdk_iop_gpio.v(252)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg9_b14  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/p1_in [14]),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync1 [14]));  // ../RTL/cmsdk_iop_gpio.v(252)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg9_b15  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/p1_in [15]),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync1 [15]));  // ../RTL/cmsdk_iop_gpio.v(252)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg9_b2  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/p1_in [2]),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync1 [2]));  // ../RTL/cmsdk_iop_gpio.v(252)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg9_b3  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/p1_in [3]),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync1 [3]));  // ../RTL/cmsdk_iop_gpio.v(252)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg9_b4  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/p1_in [4]),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync1 [4]));  // ../RTL/cmsdk_iop_gpio.v(252)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg9_b5  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/p1_in [5]),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync1 [5]));  // ../RTL/cmsdk_iop_gpio.v(252)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg9_b6  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/p1_in [6]),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync1 [6]));  // ../RTL/cmsdk_iop_gpio.v(252)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg9_b7  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/p1_in [7]),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync1 [7]));  // ../RTL/cmsdk_iop_gpio.v(252)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg9_b8  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/p1_in [8]),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync1 [8]));  // ../RTL/cmsdk_iop_gpio.v(252)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg9_b9  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/p1_in [9]),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync1 [9]));  // ../RTL/cmsdk_iop_gpio.v(252)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg0_b0  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/flash_hsel ),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n11 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [0]));  // ../RTL/cmsdk_ahb_slave_mux.v(115)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg0_b1  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/sram_hsel ),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n11 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [1]));  // ../RTL/cmsdk_ahb_slave_mux.v(115)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg0_b4  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/apbsys_hsel ),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n11 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [4]));  // ../RTL/cmsdk_ahb_slave_mux.v(115)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg0_b5  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_hsel ),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n11 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [5]));  // ../RTL/cmsdk_ahb_slave_mux.v(115)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg0_b6  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio1_hsel ),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n11 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [6]));  // ../RTL/cmsdk_ahb_slave_mux.v(115)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg0_b7  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/sysctrl_hsel ),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n11 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [7]));  // ../RTL/cmsdk_ahb_slave_mux.v(115)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg0_b8  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/sysrom_hsel ),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n11 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [8]));  // ../RTL/cmsdk_ahb_slave_mux.v(115)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg0_b0  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [0]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n43 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_ddr [0]));  // ../RTL/gpio_apbif.v(262)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg0_b1  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [1]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n43 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_ddr [1]));  // ../RTL/gpio_apbif.v(262)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg0_b2  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [2]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n43 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_ddr [2]));  // ../RTL/gpio_apbif.v(262)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg0_b3  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [3]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n43 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_ddr [3]));  // ../RTL/gpio_apbif.v(262)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg0_b4  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [4]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n43 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_ddr [4]));  // ../RTL/gpio_apbif.v(262)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg0_b5  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [5]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n43 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_ddr [5]));  // ../RTL/gpio_apbif.v(262)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg0_b6  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [6]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n43 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_ddr [6]));  // ../RTL/gpio_apbif.v(262)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg0_b7  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [7]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n43 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_ddr [7]));  // ../RTL/gpio_apbif.v(262)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg2_b0  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [0]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n49 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inten [0]));  // ../RTL/gpio_apbif.v(303)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg2_b1  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [1]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n49 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inten [1]));  // ../RTL/gpio_apbif.v(303)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg2_b2  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [2]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n49 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inten [2]));  // ../RTL/gpio_apbif.v(303)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg2_b3  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [3]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n49 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inten [3]));  // ../RTL/gpio_apbif.v(303)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg2_b4  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [4]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n49 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inten [4]));  // ../RTL/gpio_apbif.v(303)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg2_b5  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [5]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n49 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inten [5]));  // ../RTL/gpio_apbif.v(303)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg2_b6  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [6]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n49 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inten [6]));  // ../RTL/gpio_apbif.v(303)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg2_b7  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [7]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n49 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inten [7]));  // ../RTL/gpio_apbif.v(303)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg3_b0  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [0]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n52 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_intmask [0]));  // ../RTL/gpio_apbif.v(323)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg3_b1  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [1]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n52 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_intmask [1]));  // ../RTL/gpio_apbif.v(323)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg3_b2  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [2]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n52 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_intmask [2]));  // ../RTL/gpio_apbif.v(323)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg3_b3  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [3]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n52 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_intmask [3]));  // ../RTL/gpio_apbif.v(323)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg3_b4  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [4]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n52 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_intmask [4]));  // ../RTL/gpio_apbif.v(323)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg3_b5  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [5]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n52 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_intmask [5]));  // ../RTL/gpio_apbif.v(323)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg3_b6  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [6]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n52 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_intmask [6]));  // ../RTL/gpio_apbif.v(323)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg3_b7  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [7]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n52 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_intmask [7]));  // ../RTL/gpio_apbif.v(323)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg4_b0  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [0]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n55 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inttype_level [0]));  // ../RTL/gpio_apbif.v(343)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg4_b1  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [1]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n55 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inttype_level [1]));  // ../RTL/gpio_apbif.v(343)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg4_b2  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [2]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n55 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inttype_level [2]));  // ../RTL/gpio_apbif.v(343)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg4_b3  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [3]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n55 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inttype_level [3]));  // ../RTL/gpio_apbif.v(343)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg4_b4  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [4]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n55 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inttype_level [4]));  // ../RTL/gpio_apbif.v(343)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg4_b5  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [5]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n55 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inttype_level [5]));  // ../RTL/gpio_apbif.v(343)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg4_b6  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [6]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n55 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inttype_level [6]));  // ../RTL/gpio_apbif.v(343)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg4_b7  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [7]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n55 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inttype_level [7]));  // ../RTL/gpio_apbif.v(343)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg5_b0  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [0]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n58 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_int_polarity [0]));  // ../RTL/gpio_apbif.v(363)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg5_b1  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [1]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n58 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_int_polarity [1]));  // ../RTL/gpio_apbif.v(363)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg5_b2  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [2]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n58 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_int_polarity [2]));  // ../RTL/gpio_apbif.v(363)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg5_b3  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [3]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n58 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_int_polarity [3]));  // ../RTL/gpio_apbif.v(363)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg5_b4  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [4]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n58 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_int_polarity [4]));  // ../RTL/gpio_apbif.v(363)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg5_b5  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [5]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n58 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_int_polarity [5]));  // ../RTL/gpio_apbif.v(363)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg5_b6  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [6]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n58 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_int_polarity [6]));  // ../RTL/gpio_apbif.v(363)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg5_b7  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [7]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n58 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_int_polarity [7]));  // ../RTL/gpio_apbif.v(363)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg6_b0  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [0]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n61 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_ls_sync ));  // ../RTL/gpio_apbif.v(383)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg6_b1  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [1]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n61 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/int_gpio_ls_sync [1]));  // ../RTL/gpio_apbif.v(383)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg6_b2  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [2]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n61 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/int_gpio_ls_sync [2]));  // ../RTL/gpio_apbif.v(383)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg6_b3  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [3]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n61 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/int_gpio_ls_sync [3]));  // ../RTL/gpio_apbif.v(383)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg6_b4  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [4]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n61 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/int_gpio_ls_sync [4]));  // ../RTL/gpio_apbif.v(383)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg6_b5  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [5]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n61 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/int_gpio_ls_sync [5]));  // ../RTL/gpio_apbif.v(383)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg6_b6  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [6]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n61 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/int_gpio_ls_sync [6]));  // ../RTL/gpio_apbif.v(383)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg6_b7  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [7]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n61 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/int_gpio_ls_sync [7]));  // ../RTL/gpio_apbif.v(383)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg7_b0  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n81 [0]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n68 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gpio0_prdata [0]));  // ../RTL/gpio_apbif.v(453)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg7_b1  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n81 [1]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n68 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gpio0_prdata [1]));  // ../RTL/gpio_apbif.v(453)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg7_b2  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n81 [2]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n68 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gpio0_prdata [2]));  // ../RTL/gpio_apbif.v(453)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg7_b3  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n81 [3]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n68 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gpio0_prdata [3]));  // ../RTL/gpio_apbif.v(453)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg7_b4  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n81 [4]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n68 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gpio0_prdata [4]));  // ../RTL/gpio_apbif.v(453)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg7_b5  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n81 [5]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n68 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gpio0_prdata [5]));  // ../RTL/gpio_apbif.v(453)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg7_b6  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n81 [6]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n68 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gpio0_prdata [6]));  // ../RTL/gpio_apbif.v(453)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg7_b7  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n81 [7]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n68 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gpio0_prdata [7]));  // ../RTL/gpio_apbif.v(453)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg8_b0  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [0]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n40 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_dr [0]));  // ../RTL/gpio_apbif.v(242)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg8_b1  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [1]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n40 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_dr [1]));  // ../RTL/gpio_apbif.v(242)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg8_b2  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [2]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n40 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_dr [2]));  // ../RTL/gpio_apbif.v(242)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg8_b3  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [3]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n40 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_dr [3]));  // ../RTL/gpio_apbif.v(242)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg8_b4  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [4]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n40 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_dr [4]));  // ../RTL/gpio_apbif.v(242)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg8_b5  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [5]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n40 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_dr [5]));  // ../RTL/gpio_apbif.v(242)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg8_b6  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [6]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n40 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_dr [6]));  // ../RTL/gpio_apbif.v(242)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg8_b7  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [7]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n40 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_dr [7]));  // ../RTL/gpio_apbif.v(242)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/reg0_b0  (
    .clk(1'b1),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/gpio_ext_porta_int [0]),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/int_s1 [0]));  // ../RTL/gpio_ctrl.v(184)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/reg0_b1  (
    .clk(1'b1),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/gpio_ext_porta_int [1]),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/int_s1 [1]));  // ../RTL/gpio_ctrl.v(184)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/reg0_b2  (
    .clk(1'b1),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/gpio_ext_porta_int [2]),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/int_s1 [2]));  // ../RTL/gpio_ctrl.v(184)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/reg0_b3  (
    .clk(1'b1),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/gpio_ext_porta_int [3]),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/int_s1 [3]));  // ../RTL/gpio_ctrl.v(184)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/reg0_b4  (
    .clk(1'b1),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/gpio_ext_porta_int [4]),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/int_s1 [4]));  // ../RTL/gpio_ctrl.v(184)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/reg0_b5  (
    .clk(1'b1),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/gpio_ext_porta_int [5]),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/int_s1 [5]));  // ../RTL/gpio_ctrl.v(184)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/reg0_b6  (
    .clk(1'b1),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/gpio_ext_porta_int [6]),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/int_s1 [6]));  // ../RTL/gpio_ctrl.v(184)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/reg0_b7  (
    .clk(1'b1),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/gpio_ext_porta_int [7]),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/int_s1 [7]));  // ../RTL/gpio_ctrl.v(184)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/reg1_b0  (
    .clk(1'b1),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/int_s1 [0]),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/int_pre_in [0]));  // ../RTL/gpio_ctrl.v(192)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/reg1_b1  (
    .clk(1'b1),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/int_s1 [1]),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/int_pre_in [1]));  // ../RTL/gpio_ctrl.v(192)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/reg1_b2  (
    .clk(1'b1),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/int_s1 [2]),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/int_pre_in [2]));  // ../RTL/gpio_ctrl.v(192)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/reg1_b3  (
    .clk(1'b1),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/int_s1 [3]),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/int_pre_in [3]));  // ../RTL/gpio_ctrl.v(192)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/reg1_b4  (
    .clk(1'b1),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/int_s1 [4]),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/int_pre_in [4]));  // ../RTL/gpio_ctrl.v(192)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/reg1_b5  (
    .clk(1'b1),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/int_s1 [5]),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/int_pre_in [5]));  // ../RTL/gpio_ctrl.v(192)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/reg1_b6  (
    .clk(1'b1),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/int_s1 [6]),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/int_pre_in [6]));  // ../RTL/gpio_ctrl.v(192)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/reg1_b7  (
    .clk(1'b1),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/int_s1 [7]),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/int_pre_in [7]));  // ../RTL/gpio_ctrl.v(192)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/reg2_b0  (
    .clk(1'b1),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/int_pre_in [0]),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/ed_int_d1 [0]));  // ../RTL/gpio_ctrl.v(203)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/reg2_b1  (
    .clk(1'b1),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/int_pre_in [1]),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/ed_int_d1 [1]));  // ../RTL/gpio_ctrl.v(203)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/reg2_b2  (
    .clk(1'b1),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/int_pre_in [2]),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/ed_int_d1 [2]));  // ../RTL/gpio_ctrl.v(203)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/reg2_b3  (
    .clk(1'b1),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/int_pre_in [3]),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/ed_int_d1 [3]));  // ../RTL/gpio_ctrl.v(203)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/reg2_b4  (
    .clk(1'b1),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/int_pre_in [4]),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/ed_int_d1 [4]));  // ../RTL/gpio_ctrl.v(203)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/reg2_b5  (
    .clk(1'b1),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/int_pre_in [5]),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/ed_int_d1 [5]));  // ../RTL/gpio_ctrl.v(203)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/reg2_b6  (
    .clk(1'b1),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/int_pre_in [6]),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/ed_int_d1 [6]));  // ../RTL/gpio_ctrl.v(203)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/reg2_b7  (
    .clk(1'b1),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/int_pre_in [7]),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/ed_int_d1 [7]));  // ../RTL/gpio_ctrl.v(203)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/reg3_b0  (
    .clk(1'b1),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/n28 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/gpio_intr_ed_pm [0]));  // ../RTL/gpio_ctrl.v(248)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/reg3_b1  (
    .clk(1'b1),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/n36 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/gpio_intr_ed_pm [1]));  // ../RTL/gpio_ctrl.v(248)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/reg3_b2  (
    .clk(1'b1),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/n44 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/gpio_intr_ed_pm [2]));  // ../RTL/gpio_ctrl.v(248)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/reg3_b3  (
    .clk(1'b1),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/n52 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/gpio_intr_ed_pm [3]));  // ../RTL/gpio_ctrl.v(248)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/reg3_b4  (
    .clk(1'b1),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/n60 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/gpio_intr_ed_pm [4]));  // ../RTL/gpio_ctrl.v(248)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/reg3_b5  (
    .clk(1'b1),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/n68 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/gpio_intr_ed_pm [5]));  // ../RTL/gpio_ctrl.v(248)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/reg3_b6  (
    .clk(1'b1),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/n76 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/gpio_intr_ed_pm [6]));  // ../RTL/gpio_ctrl.v(248)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/reg3_b7  (
    .clk(1'b1),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/n84 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/gpio_intr_ed_pm [7]));  // ../RTL/gpio_ctrl.v(248)
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add0/u0  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_tick_cnt [0]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/BAUDTICK ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add0/c0 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add0/c1 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n55 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add0/u1  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_tick_cnt [1]),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add0/c1 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add0/c2 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n55 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add0/u2  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_tick_cnt [2]),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add0/c2 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add0/c3 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n55 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add0/u3  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_tick_cnt [3]),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add0/c3 ),
    .o({open_n799,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n55 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add0/ucin  (
    .a(1'b0),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add0/c0 ,open_n802}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add1/u0  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_state [0]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_state_inc ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add1/c0 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add1/c1 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n67 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add1/u1  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_state [1]),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add1/c1 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add1/c2 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n67 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add1/u2  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_state [2]),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add1/c2 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add1/c3 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n67 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add1/u3  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_state [3]),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add1/c3 ),
    .o({open_n803,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n67 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add1/ucin  (
    .a(1'b0),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add1/c0 ,open_n806}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add2/u0  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_tick_cnt [0]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/BAUDTICK ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add2/c0 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add2/c1 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n92 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add2/u1  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_tick_cnt [1]),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add2/c1 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add2/c2 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n92 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add2/u2  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_tick_cnt [2]),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add2/c2 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add2/c3 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n92 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add2/u3  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_tick_cnt [3]),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add2/c3 ),
    .o({open_n807,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n92 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add2/ucin  (
    .a(1'b0),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add2/c0 ,open_n810}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add3/u0  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_state [0]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_state_inc ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add3/c0 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add3/c1 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n102 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add3/u1  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_state [1]),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add3/c1 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add3/c2 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n102 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add3/u2  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_state [2]),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add3/c2 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add3/c3 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n102 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add3/u3  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_state [3]),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add3/c3 ),
    .o({open_n811,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n102 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add3/ucin  (
    .a(1'b0),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add3/c0 ,open_n814}));
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/baud_updated_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/write_enable10 ),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n46 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/baud_updated ));  // ../RTL/cmsdk_apb_uart.v(368)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/lt0_0  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [0]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_f [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/lt0_c0 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/lt0_c1 ,open_n815}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/lt0_1  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [1]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_f [2]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/lt0_c1 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/lt0_c2 ,open_n816}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/lt0_2  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [2]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_f [1]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/lt0_c2 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/lt0_c3 ,open_n817}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/lt0_3  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [3]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_f [0]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/lt0_c3 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/lt0_c4 ,open_n818}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/lt0_cin  (
    .a(1'b1),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/lt0_c0 ,open_n821}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/lt0_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/lt0_c4 ),
    .o({open_n822,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n31 }));
  AL_MAP_LUT4 #(
    .EQN("(~A*~B*~C*D+~A*B*~C*D+~A*~B*C*D+~A*B*C*D+A*B*C*D)"),
    .INIT(16'b1101010100000000))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/mux4_b0_rom0  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[4] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[5] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n28 [0]));
  AL_MAP_LUT4 #(
    .EQN("(~A*~B*C*~D+~A*~B*C*D+~A*B*C*D)"),
    .INIT(16'b0101000000010000))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/mux4_b2_rom0  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[4] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[5] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n28 [2]));
  AL_MAP_LUT4 #(
    .EQN("(A*~B*~C*D+~A*B*~C*D+~A*~B*C*D)"),
    .INIT(16'b0001011000000000))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/mux4_b3_rom0  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[4] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[5] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n28 [3]));
  AL_MAP_LUT4 #(
    .EQN("(A*~B*~C*D+~A*B*~C*D+A*~B*C*D+A*B*C*D)"),
    .INIT(16'b1010011000000000))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/mux4_b4_rom0  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[4] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[5] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n28 [4]));
  AL_MAP_LUT4 #(
    .EQN("(~A*~B*~C*D+A*~B*~C*D+A*~B*C*D+A*B*C*D)"),
    .INIT(16'b1010001100000000))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/mux4_b5_rom0  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[4] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[5] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n28 [5]));
  AL_MAP_LUT4 #(
    .EQN("(A*~B*~C*D+A*~B*C*D+A*B*C*D)"),
    .INIT(16'b1010001000000000))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/mux4_b7_rom0  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[4] ),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[5] ),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n28 [7]));
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg0_b0  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [0]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/write_enable08 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(uart0_txen_pad));  // ../RTL/cmsdk_apb_uart.v(238)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg0_b1  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [1]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/write_enable08 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_ctrl [1]));  // ../RTL/cmsdk_apb_uart.v(238)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg0_b2  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [2]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/write_enable08 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_ctrl [2]));  // ../RTL/cmsdk_apb_uart.v(238)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg0_b3  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [3]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/write_enable08 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_ctrl [3]));  // ../RTL/cmsdk_apb_uart.v(238)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg0_b4  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [4]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/write_enable08 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_ctrl [4]));  // ../RTL/cmsdk_apb_uart.v(238)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg0_b5  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [5]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/write_enable08 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_ctrl [5]));  // ../RTL/cmsdk_apb_uart.v(238)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg0_b6  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [6]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/write_enable08 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_ctrl [6]));  // ../RTL/cmsdk_apb_uart.v(238)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg10_b0  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_rx_state [0]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_state_update ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_state [0]));  // ../RTL/cmsdk_apb_uart.v(583)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg10_b1  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_rx_state [1]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_state_update ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_state [1]));  // ../RTL/cmsdk_apb_uart.v(583)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg10_b2  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_rx_state [2]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_state_update ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_state [2]));  // ../RTL/cmsdk_apb_uart.v(583)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg10_b3  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_rx_state [3]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_state_update ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_state [3]));  // ../RTL/cmsdk_apb_uart.v(583)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg11_b0  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_shift_buf [0]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rxbuf_sample ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_rx_buf [0]));  // ../RTL/cmsdk_apb_uart.v(603)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg11_b1  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_shift_buf [1]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rxbuf_sample ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_rx_buf [1]));  // ../RTL/cmsdk_apb_uart.v(603)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg11_b2  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_shift_buf [2]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rxbuf_sample ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_rx_buf [2]));  // ../RTL/cmsdk_apb_uart.v(603)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg11_b3  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_shift_buf [3]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rxbuf_sample ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_rx_buf [3]));  // ../RTL/cmsdk_apb_uart.v(603)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg11_b4  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_shift_buf [4]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rxbuf_sample ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_rx_buf [4]));  // ../RTL/cmsdk_apb_uart.v(603)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg11_b5  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_shift_buf [5]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rxbuf_sample ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_rx_buf [5]));  // ../RTL/cmsdk_apb_uart.v(603)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg11_b6  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_shift_buf [6]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rxbuf_sample ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_rx_buf [6]));  // ../RTL/cmsdk_apb_uart.v(603)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg11_b7  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_shift_in ),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rxbuf_sample ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_rx_buf [7]));  // ../RTL/cmsdk_apb_uart.v(603)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg12_b0  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_shift_buf [1]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_state_inc ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_shift_buf [0]));  // ../RTL/cmsdk_apb_uart.v(614)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg12_b1  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_shift_buf [2]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_state_inc ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_shift_buf [1]));  // ../RTL/cmsdk_apb_uart.v(614)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg12_b2  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_shift_buf [3]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_state_inc ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_shift_buf [2]));  // ../RTL/cmsdk_apb_uart.v(614)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg12_b3  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_shift_buf [4]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_state_inc ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_shift_buf [3]));  // ../RTL/cmsdk_apb_uart.v(614)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg12_b4  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_shift_buf [5]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_state_inc ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_shift_buf [4]));  // ../RTL/cmsdk_apb_uart.v(614)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg12_b5  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_shift_buf [6]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_state_inc ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_shift_buf [5]));  // ../RTL/cmsdk_apb_uart.v(614)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg12_b6  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_shift_in ),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_state_inc ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_shift_buf [6]));  // ../RTL/cmsdk_apb_uart.v(614)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg13_b0  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [0]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/write_enable00 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_tx_buf [0]));  // ../RTL/cmsdk_apb_uart.v(207)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg13_b1  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [1]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/write_enable00 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_tx_buf [1]));  // ../RTL/cmsdk_apb_uart.v(207)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg13_b2  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [2]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/write_enable00 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_tx_buf [2]));  // ../RTL/cmsdk_apb_uart.v(207)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg13_b3  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [3]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/write_enable00 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_tx_buf [3]));  // ../RTL/cmsdk_apb_uart.v(207)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg13_b4  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [4]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/write_enable00 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_tx_buf [4]));  // ../RTL/cmsdk_apb_uart.v(207)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg13_b5  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [5]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/write_enable00 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_tx_buf [5]));  // ../RTL/cmsdk_apb_uart.v(207)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg13_b6  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [6]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/write_enable00 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_tx_buf [6]));  // ../RTL/cmsdk_apb_uart.v(207)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg13_b7  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [7]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/write_enable00 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_tx_buf [7]));  // ../RTL/cmsdk_apb_uart.v(207)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg1_b0  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [0]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/write_enable10 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [0]));  // ../RTL/cmsdk_apb_uart.v(247)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg1_b1  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [1]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/write_enable10 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [1]));  // ../RTL/cmsdk_apb_uart.v(247)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg1_b10  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [10]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/write_enable10 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [10]));  // ../RTL/cmsdk_apb_uart.v(247)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg1_b11  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [11]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/write_enable10 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [11]));  // ../RTL/cmsdk_apb_uart.v(247)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg1_b12  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [12]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/write_enable10 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [12]));  // ../RTL/cmsdk_apb_uart.v(247)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg1_b13  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [13]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/write_enable10 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [13]));  // ../RTL/cmsdk_apb_uart.v(247)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg1_b14  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [14]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/write_enable10 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [14]));  // ../RTL/cmsdk_apb_uart.v(247)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg1_b15  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [15]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/write_enable10 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [15]));  // ../RTL/cmsdk_apb_uart.v(247)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg1_b16  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [16]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/write_enable10 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [16]));  // ../RTL/cmsdk_apb_uart.v(247)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg1_b17  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [17]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/write_enable10 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [17]));  // ../RTL/cmsdk_apb_uart.v(247)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg1_b18  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [18]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/write_enable10 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [18]));  // ../RTL/cmsdk_apb_uart.v(247)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg1_b19  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [19]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/write_enable10 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [19]));  // ../RTL/cmsdk_apb_uart.v(247)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg1_b2  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [2]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/write_enable10 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [2]));  // ../RTL/cmsdk_apb_uart.v(247)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg1_b3  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [3]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/write_enable10 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [3]));  // ../RTL/cmsdk_apb_uart.v(247)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg1_b4  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [4]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/write_enable10 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [4]));  // ../RTL/cmsdk_apb_uart.v(247)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg1_b5  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [5]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/write_enable10 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [5]));  // ../RTL/cmsdk_apb_uart.v(247)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg1_b6  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [6]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/write_enable10 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [6]));  // ../RTL/cmsdk_apb_uart.v(247)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg1_b7  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [7]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/write_enable10 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [7]));  // ../RTL/cmsdk_apb_uart.v(247)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg1_b8  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [8]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/write_enable10 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [8]));  // ../RTL/cmsdk_apb_uart.v(247)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg1_b9  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [9]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/write_enable10 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [9]));  // ../RTL/cmsdk_apb_uart.v(247)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg2_b0  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/read_mux_byte0 [0]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/read_enable ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/read_mux_byte0_reg [0]));  // ../RTL/cmsdk_apb_uart.v(303)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg2_b1  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/read_mux_byte0 [1]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/read_enable ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/read_mux_byte0_reg [1]));  // ../RTL/cmsdk_apb_uart.v(303)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg2_b2  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/read_mux_byte0 [2]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/read_enable ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/read_mux_byte0_reg [2]));  // ../RTL/cmsdk_apb_uart.v(303)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg2_b3  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/read_mux_byte0 [3]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/read_enable ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/read_mux_byte0_reg [3]));  // ../RTL/cmsdk_apb_uart.v(303)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg2_b4  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/read_mux_byte0 [4]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/read_enable ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/read_mux_byte0_reg [4]));  // ../RTL/cmsdk_apb_uart.v(303)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg2_b5  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/read_mux_byte0 [5]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/read_enable ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/read_mux_byte0_reg [5]));  // ../RTL/cmsdk_apb_uart.v(303)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg2_b6  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/read_mux_byte0 [6]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/read_enable ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/read_mux_byte0_reg [6]));  // ../RTL/cmsdk_apb_uart.v(303)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg2_b7  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/read_mux_byte0 [7]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/read_enable ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/read_mux_byte0_reg [7]));  // ../RTL/cmsdk_apb_uart.v(303)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg3_b0  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_baud_cntr_i [0]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n38 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_i [0]));  // ../RTL/cmsdk_apb_uart.v(341)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg3_b1  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_baud_cntr_i [1]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n38 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_i [1]));  // ../RTL/cmsdk_apb_uart.v(341)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg3_b10  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_baud_cntr_i [10]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n38 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_i [10]));  // ../RTL/cmsdk_apb_uart.v(341)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg3_b11  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_baud_cntr_i [11]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n38 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_i [11]));  // ../RTL/cmsdk_apb_uart.v(341)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg3_b12  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_baud_cntr_i [12]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n38 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_i [12]));  // ../RTL/cmsdk_apb_uart.v(341)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg3_b13  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_baud_cntr_i [13]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n38 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_i [13]));  // ../RTL/cmsdk_apb_uart.v(341)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg3_b14  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_baud_cntr_i [14]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n38 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_i [14]));  // ../RTL/cmsdk_apb_uart.v(341)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg3_b15  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_baud_cntr_i [15]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n38 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_i [15]));  // ../RTL/cmsdk_apb_uart.v(341)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg3_b2  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_baud_cntr_i [2]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n38 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_i [2]));  // ../RTL/cmsdk_apb_uart.v(341)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg3_b3  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_baud_cntr_i [3]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n38 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_i [3]));  // ../RTL/cmsdk_apb_uart.v(341)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg3_b4  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_baud_cntr_i [4]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n38 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_i [4]));  // ../RTL/cmsdk_apb_uart.v(341)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg3_b5  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_baud_cntr_i [5]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n38 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_i [5]));  // ../RTL/cmsdk_apb_uart.v(341)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg3_b6  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_baud_cntr_i [6]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n38 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_i [6]));  // ../RTL/cmsdk_apb_uart.v(341)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg3_b7  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_baud_cntr_i [7]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n38 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_i [7]));  // ../RTL/cmsdk_apb_uart.v(341)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg3_b8  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_baud_cntr_i [8]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n38 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_i [8]));  // ../RTL/cmsdk_apb_uart.v(341)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg3_b9  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_baud_cntr_i [9]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n38 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_i [9]));  // ../RTL/cmsdk_apb_uart.v(341)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg4_b0  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_baud_cntr_f [0]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n44 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_f [0]));  // ../RTL/cmsdk_apb_uart.v(358)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg4_b1  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_baud_cntr_f [1]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n44 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_f [1]));  // ../RTL/cmsdk_apb_uart.v(358)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg4_b2  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_baud_cntr_f [2]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n44 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_f [2]));  // ../RTL/cmsdk_apb_uart.v(358)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg4_b3  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_baud_cntr_f [3]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n44 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_f [3]));  // ../RTL/cmsdk_apb_uart.v(358)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg5_b0  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_tx_tick_cnt [0]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/BAUDTICK ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_tick_cnt [0]));  // ../RTL/cmsdk_apb_uart.v(405)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg5_b1  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_tx_tick_cnt [1]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/BAUDTICK ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_tick_cnt [1]));  // ../RTL/cmsdk_apb_uart.v(405)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg5_b2  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_tx_tick_cnt [2]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/BAUDTICK ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_tick_cnt [2]));  // ../RTL/cmsdk_apb_uart.v(405)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg5_b3  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_tx_tick_cnt [3]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/BAUDTICK ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_tick_cnt [3]));  // ../RTL/cmsdk_apb_uart.v(405)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg6_b0  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_tx_state [0]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_state_update ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_state [0]));  // ../RTL/cmsdk_apb_uart.v(445)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg6_b1  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_tx_state [1]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_state_update ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_state [1]));  // ../RTL/cmsdk_apb_uart.v(445)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg6_b2  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_tx_state [2]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_state_update ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_state [2]));  // ../RTL/cmsdk_apb_uart.v(445)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg6_b3  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_tx_state [3]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_state_update ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_state [3]));  // ../RTL/cmsdk_apb_uart.v(445)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg7_b0  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_tx_shift_buf [0]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n74 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_shift_buf [0]));  // ../RTL/cmsdk_apb_uart.v(461)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg7_b1  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_tx_shift_buf [1]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n74 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_shift_buf [1]));  // ../RTL/cmsdk_apb_uart.v(461)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg7_b2  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_tx_shift_buf [2]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n74 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_shift_buf [2]));  // ../RTL/cmsdk_apb_uart.v(461)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg7_b3  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_tx_shift_buf [3]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n74 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_shift_buf [3]));  // ../RTL/cmsdk_apb_uart.v(461)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg7_b4  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_tx_shift_buf [4]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n74 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_shift_buf [4]));  // ../RTL/cmsdk_apb_uart.v(461)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg7_b5  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_tx_shift_buf [5]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n74 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_shift_buf [5]));  // ../RTL/cmsdk_apb_uart.v(461)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg7_b6  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_tx_shift_buf [6]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n74 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_shift_buf [6]));  // ../RTL/cmsdk_apb_uart.v(461)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg7_b7  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_tx_shift_buf [7]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n74 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_shift_buf [7]));  // ../RTL/cmsdk_apb_uart.v(461)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg8_b0  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rxd_sync_2 ),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/BAUDTICK ),
    .reset(1'b0),
    .set(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rxd_lpf [0]));  // ../RTL/cmsdk_apb_uart.v(512)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg8_b1  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rxd_lpf [0]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/BAUDTICK ),
    .reset(1'b0),
    .set(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rxd_lpf [1]));  // ../RTL/cmsdk_apb_uart.v(512)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg8_b2  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rxd_lpf [1]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/BAUDTICK ),
    .reset(1'b0),
    .set(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rxd_lpf [2]));  // ../RTL/cmsdk_apb_uart.v(512)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg9_b0  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_rx_tick_cnt [0]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/update_rx_tick_cnt ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_tick_cnt [0]));  // ../RTL/cmsdk_apb_uart.v(535)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg9_b1  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_rx_tick_cnt [1]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/update_rx_tick_cnt ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_tick_cnt [1]));  // ../RTL/cmsdk_apb_uart.v(535)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg9_b2  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_rx_tick_cnt [2]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/update_rx_tick_cnt ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_tick_cnt [2]));  // ../RTL/cmsdk_apb_uart.v(535)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg9_b3  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_rx_tick_cnt [3]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/update_rx_tick_cnt ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_tick_cnt [3]));  // ../RTL/cmsdk_apb_uart.v(535)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_tick_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reload_i ),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n48 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/BAUDTICK ));  // ../RTL/cmsdk_apb_uart.v(377)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_rx_overrun_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_rx_overrun ),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n17 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_rx_overrun ));  // ../RTL/cmsdk_apb_uart.v(220)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_rxintr_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/intr_stat_set [1]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n117 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/apbsubsys_interrupt [0]));  // ../RTL/cmsdk_apb_uart.v(642)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_tx_overrun_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_tx_overrun ),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n20 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_tx_overrun ));  // ../RTL/cmsdk_apb_uart.v(229)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_txd_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_txd ),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/update_reg_txd ),
    .reset(1'b0),
    .set(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .q(uart0_txd_pad));  // ../RTL/cmsdk_apb_uart.v(476)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_txintr_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/intr_stat_set [0]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n114 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/apbsubsys_interrupt [1]));  // ../RTL/cmsdk_apb_uart.v(634)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_buf_full_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_rx_buf_full ),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n106 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_buf_full ));  // ../RTL/cmsdk_apb_uart.v(592)
  EG_PHY_PAD #(
    //.CLKSRC("CLK"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IDDRPIPEMODE("NONE"),
    .INCEMUX("CE"),
    .INPCLKMUX("CLK"),
    .INRSTMUX("INV"),
    .IN_DFFMODE("FF"),
    .IN_REGSET("SET"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .SRMODE("ASYNC"),
    .TSMUX("1"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rxd_sync_1_reg_IN  (
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_ctrl [1]),
    .ipad(uart0_rxd),
    .ipclk(XTAL1_wire),
    .rst(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .diq({open_n832,open_n833,open_n834,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rxd_sync_1 }));  // ../RTL/cmsdk_apb_uart.v(501)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rxd_sync_2_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rxd_sync_1 ),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_ctrl [1]),
    .reset(1'b0),
    .set(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rxd_sync_2 ));  // ../RTL/cmsdk_apb_uart.v(501)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/u0  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_i [0]),
    .b(1'b1),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/c0 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/c1 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n37 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/u1  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_i [1]),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/c1 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/c2 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n37 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/u10  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_i [10]),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/c10 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/c11 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n37 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/u11  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_i [11]),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/c11 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/c12 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n37 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/u12  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_i [12]),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/c12 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/c13 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n37 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/u13  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_i [13]),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/c13 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/c14 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n37 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/u14  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_i [14]),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/c14 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/c15 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n37 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/u15  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_i [15]),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/c15 ),
    .o({open_n837,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n37 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/u2  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_i [2]),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/c2 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/c3 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n37 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/u3  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_i [3]),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/c3 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/c4 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n37 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/u4  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_i [4]),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/c4 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/c5 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n37 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/u5  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_i [5]),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/c5 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/c6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n37 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/u6  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_i [6]),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/c6 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/c7 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n37 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/u7  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_i [7]),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/c7 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/c8 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n37 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/u8  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_i [8]),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/c8 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/c9 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n37 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/u9  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_i [9]),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/c9 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/c10 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n37 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/ucin  (
    .a(1'b0),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/c0 ,open_n840}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub1/u0  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_f [0]),
    .b(1'b1),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub1/c0 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub1/c1 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n43 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub1/u1  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_f [1]),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub1/c1 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub1/c2 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n43 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub1/u2  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_f [2]),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub1/c2 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub1/c3 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n43 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub1/u3  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_f [3]),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub1/c3 ),
    .o({open_n841,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n43 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub1/ucin  (
    .a(1'b0),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub1/c0 ,open_n844}));
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_buf_full_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/write_enable00 ),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n50 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_buf_full ));  // ../RTL/cmsdk_apb_uart.v(392)
  AL_MAP_LUT3 #(
    .EQN("(~A*~B*~C+~A*~B*C+~A*B*C)"),
    .INIT(8'b01010001))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/mux11_rom0  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/state_reg [0]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/state_reg [1]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/state_reg [2]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/apbsys_hreadyout ));
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/reg2_b0  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/next_state [0]),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/state_reg [0]));  // ../RTL/cmsdk_ahb_to_apb.v(253)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/reg2_b1  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/next_state [1]),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/state_reg [1]));  // ../RTL/cmsdk_ahb_to_apb.v(253)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/reg2_b2  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/next_state [2]),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/state_reg [2]));  // ../RTL/cmsdk_ahb_to_apb.v(253)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/reg3_b0  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_apb_slave_mux/n118 [0]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/apb_tran_end ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/rwdata_reg [0]));  // ../RTL/cmsdk_ahb_to_apb.v(265)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/reg3_b1  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_apb_slave_mux/n118 [1]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/apb_tran_end ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/rwdata_reg [1]));  // ../RTL/cmsdk_ahb_to_apb.v(265)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/reg3_b10  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_apb_slave_mux/n117 [10]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/apb_tran_end ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/rwdata_reg [10]));  // ../RTL/cmsdk_ahb_to_apb.v(265)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/reg3_b11  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_apb_slave_mux/n117 [11]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/apb_tran_end ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/rwdata_reg [11]));  // ../RTL/cmsdk_ahb_to_apb.v(265)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/reg3_b12  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_apb_slave_mux/n117 [12]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/apb_tran_end ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/rwdata_reg [12]));  // ../RTL/cmsdk_ahb_to_apb.v(265)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/reg3_b13  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_apb_slave_mux/n117 [13]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/apb_tran_end ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/rwdata_reg [13]));  // ../RTL/cmsdk_ahb_to_apb.v(265)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/reg3_b14  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_apb_slave_mux/n117 [14]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/apb_tran_end ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/rwdata_reg [14]));  // ../RTL/cmsdk_ahb_to_apb.v(265)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/reg3_b15  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_apb_slave_mux/n117 [15]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/apb_tran_end ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/rwdata_reg [15]));  // ../RTL/cmsdk_ahb_to_apb.v(265)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/reg3_b16  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_apb_slave_mux/n117 [16]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/apb_tran_end ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/rwdata_reg [16]));  // ../RTL/cmsdk_ahb_to_apb.v(265)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/reg3_b17  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_apb_slave_mux/n117 [17]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/apb_tran_end ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/rwdata_reg [17]));  // ../RTL/cmsdk_ahb_to_apb.v(265)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/reg3_b18  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_apb_slave_mux/n117 [18]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/apb_tran_end ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/rwdata_reg [18]));  // ../RTL/cmsdk_ahb_to_apb.v(265)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/reg3_b19  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_apb_slave_mux/n117 [19]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/apb_tran_end ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/rwdata_reg [19]));  // ../RTL/cmsdk_ahb_to_apb.v(265)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/reg3_b2  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_apb_slave_mux/n118 [2]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/apb_tran_end ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/rwdata_reg [2]));  // ../RTL/cmsdk_ahb_to_apb.v(265)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/reg3_b3  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_apb_slave_mux/n118 [3]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/apb_tran_end ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/rwdata_reg [3]));  // ../RTL/cmsdk_ahb_to_apb.v(265)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/reg3_b4  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_apb_slave_mux/n118 [4]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/apb_tran_end ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/rwdata_reg [4]));  // ../RTL/cmsdk_ahb_to_apb.v(265)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/reg3_b5  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_apb_slave_mux/n118 [5]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/apb_tran_end ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/rwdata_reg [5]));  // ../RTL/cmsdk_ahb_to_apb.v(265)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/reg3_b6  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_apb_slave_mux/n118 [6]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/apb_tran_end ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/rwdata_reg [6]));  // ../RTL/cmsdk_ahb_to_apb.v(265)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/reg3_b7  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_apb_slave_mux/n118 [7]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/apb_tran_end ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/rwdata_reg [7]));  // ../RTL/cmsdk_ahb_to_apb.v(265)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/reg3_b8  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_apb_slave_mux/n117 [8]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/apb_tran_end ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/rwdata_reg [8]));  // ../RTL/cmsdk_ahb_to_apb.v(265)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/reg3_b9  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_apb_slave_mux/n117 [9]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/apb_tran_end ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/rwdata_reg [9]));  // ../RTL/cmsdk_ahb_to_apb.v(265)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/reg4_b0  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HADDR [2]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/n1 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] ));  // ../RTL/cmsdk_ahb_to_apb.v(153)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/reg4_b1  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HADDR [3]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/n1 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] ));  // ../RTL/cmsdk_ahb_to_apb.v(153)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/reg4_b10  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HADDR [12]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/n1 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/i_paddr [12]));  // ../RTL/cmsdk_ahb_to_apb.v(153)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/reg4_b11  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HADDR [13]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/n1 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/i_paddr [13]));  // ../RTL/cmsdk_ahb_to_apb.v(153)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/reg4_b12  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HADDR [14]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/n1 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/i_paddr [14]));  // ../RTL/cmsdk_ahb_to_apb.v(153)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/reg4_b13  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HADDR [15]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/n1 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/i_paddr [15]));  // ../RTL/cmsdk_ahb_to_apb.v(153)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/reg4_b2  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HADDR [4]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/n1 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[4] ));  // ../RTL/cmsdk_ahb_to_apb.v(153)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/reg4_b3  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HADDR [5]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/n1 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[5] ));  // ../RTL/cmsdk_ahb_to_apb.v(153)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/reg4_b4  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HADDR [6]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/n1 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[6] ));  // ../RTL/cmsdk_ahb_to_apb.v(153)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/reg4_b5  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HADDR [7]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/n1 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[7] ));  // ../RTL/cmsdk_ahb_to_apb.v(153)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/reg4_b6  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HADDR [8]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/n1 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[8] ));  // ../RTL/cmsdk_ahb_to_apb.v(153)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/reg4_b7  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HADDR [9]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/n1 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[9] ));  // ../RTL/cmsdk_ahb_to_apb.v(153)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/reg4_b8  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HADDR [10]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/n1 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[10] ));  // ../RTL/cmsdk_ahb_to_apb.v(153)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/reg4_b9  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HADDR [11]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/n1 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[11] ));  // ../RTL/cmsdk_ahb_to_apb.v(153)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/wr_reg_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWRITE ),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/n1 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PWRITE ));  // ../RTL/cmsdk_ahb_to_apb.v(153)
  AL_MAP_LUT4 #(
    .EQN("(~A*B*~C*D+~A*~B*C*D+~A*B*C*D+A*B*C*D)"),
    .INIT(16'b1101010000000000))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/mux4_b0_rom0  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [2]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [4]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [5]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/n19 [0]));
  AL_MAP_LUT4 #(
    .EQN("(~A*~B*~C*D+~A*B*~C*D)"),
    .INIT(16'b0000010100000000))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/mux4_b1_rom0  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [2]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [4]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [5]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/n19 [1]));
  AL_MAP_LUT4 #(
    .EQN("(~A*~B*C*~D+~A*~B*~C*D+~A*~B*C*D+~A*B*C*D)"),
    .INIT(16'b0101000100010000))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/mux4_b2_rom0  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [2]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [4]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [5]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/n19 [2]));
  AL_MAP_LUT4 #(
    .EQN("(A*~B*~C*D+~A*B*~C*D+~A*~B*C*D)"),
    .INIT(16'b0001011000000000))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/mux4_b3_rom0  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [2]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [4]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [5]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/n19 [3]));
  AL_MAP_LUT4 #(
    .EQN("(A*~B*~C*D+~A*B*~C*D+A*~B*C*D+A*B*C*D)"),
    .INIT(16'b1010011000000000))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/mux4_b4_rom0  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [2]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [4]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [5]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/n19 [4]));
  AL_MAP_LUT4 #(
    .EQN("(~A*~B*~C*D+A*~B*~C*D+A*~B*C*D+A*B*C*D)"),
    .INIT(16'b1010001100000000))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/mux4_b5_rom0  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [2]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [4]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [5]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/n19 [5]));
  AL_MAP_LUT4 #(
    .EQN("(A*~B*~C*D+A*~B*C*D+A*B*C*D)"),
    .INIT(16'b1010001000000000))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/mux4_b7_rom0  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [2]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [4]),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [5]),
    .o(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/n19 [7]));
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg0_b0  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HADDR [2]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/ahb_access ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [2]));  // ../RTL/cmsdk_mcu_sysctrl.v(156)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg0_b1  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HADDR [3]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/ahb_access ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [3]));  // ../RTL/cmsdk_mcu_sysctrl.v(156)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg0_b2  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HADDR [4]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/ahb_access ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [4]));  // ../RTL/cmsdk_mcu_sysctrl.v(156)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg0_b3  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HADDR [5]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/ahb_access ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [5]));  // ../RTL/cmsdk_mcu_sysctrl.v(156)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg0_b4  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HADDR [6]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/ahb_access ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [6]));  // ../RTL/cmsdk_mcu_sysctrl.v(156)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg0_b5  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HADDR [7]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/ahb_access ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [7]));  // ../RTL/cmsdk_mcu_sysctrl.v(156)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg0_b6  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HADDR [8]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/ahb_access ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [8]));  // ../RTL/cmsdk_mcu_sysctrl.v(156)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg0_b7  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HADDR [9]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/ahb_access ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [9]));  // ../RTL/cmsdk_mcu_sysctrl.v(156)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg0_b8  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HADDR [10]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/ahb_access ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [10]));  // ../RTL/cmsdk_mcu_sysctrl.v(156)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg0_b9  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HADDR [11]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/ahb_access ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [11]));  // ../RTL/cmsdk_mcu_sysctrl.v(156)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg2_b0  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/nxt_resetinfo [0]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_resetinfo_en ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/reset_sync_reg [2]),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_resetinfo [0]));  // ../RTL/cmsdk_mcu_sysctrl.v(318)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg2_b1  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/n38 [1]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_resetinfo_en ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/reset_sync_reg [2]),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_resetinfo [1]));  // ../RTL/cmsdk_mcu_sysctrl.v(318)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg2_b2  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/nxt_resetinfo [2]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_resetinfo_en ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/reset_sync_reg [2]),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_resetinfo [2]));  // ../RTL/cmsdk_mcu_sysctrl.v(318)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg3_b0  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/nxt_byte_strobe [0]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n11 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_byte_strobe [0]));  // ../RTL/cmsdk_mcu_sysctrl.v(147)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_lockupreset_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [0]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_lockupreset_write ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/LOCKUPRESET ));  // ../RTL/cmsdk_mcu_sysctrl.v(290)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_read_enable_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/ahb_read ),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n11 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_read_enable ));  // ../RTL/cmsdk_mcu_sysctrl.v(147)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_remap_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [0]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_remap_write ),
    .reset(1'b0),
    .set(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/remap_ctrl ));  // ../RTL/cmsdk_mcu_sysctrl.v(250)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_write_enable_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/ahb_write ),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n11 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_write_enable ));  // ../RTL/cmsdk_mcu_sysctrl.v(147)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A1qax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K39iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ickiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[30] ));  // ../RTL/cortexm0ds_logic.v(18823)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A2spw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sokiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mx8iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[6] ));  // ../RTL/cortexm0ds_logic.v(17639)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A32qw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fpohu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[29] ));  // ../RTL/cortexm0ds_logic.v(17961)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A3ipw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lf1iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sf1iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A3ipw6 ));  // ../RTL/cortexm0ds_logic.v(17180)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A3qax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D39iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ickiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[31] ));  // ../RTL/cortexm0ds_logic.v(18824)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A5ipw6_reg  (
    .clk(SWCLKTCK_pad),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nrxhu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kxhpw6 ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A5ipw6 ));  // ../RTL/cortexm0ds_logic.v(17185)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A5qax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tx8iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ickiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[0] ));  // ../RTL/cortexm0ds_logic.v(18825)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A6cbx6_reg  (
    .clk(SWCLKTCK_pad),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J4cbx6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C53iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A6cbx6 ));  // ../RTL/cortexm0ds_logic.v(19945)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A7zpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Drkiu6 ),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[5] ));  // ../RTL/cortexm0ds_logic.v(17899)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aa2bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C5phu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aa2bx6 ));  // ../RTL/cortexm0ds_logic.v(19401)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ab9ax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U64iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zg7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ab9ax6 ));  // ../RTL/cortexm0ds_logic.v(18163)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Acebx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I74iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Td7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Acebx6 ));  // ../RTL/cortexm0ds_logic.v(19991)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Acuax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jgkiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wckiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[3] ));  // ../RTL/cortexm0ds_logic.v(18901)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ad7ax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S54iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n382 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ad7ax6 ));  // ../RTL/cortexm0ds_logic.v(18091)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahdax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ud4iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Td7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahdax6 ));  // ../RTL/cortexm0ds_logic.v(18289)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahdbx6_reg  (
    .clk(SWCLKTCK_pad),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jfdbx6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C53iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahdbx6 ));  // ../RTL/cortexm0ds_logic.v(19975)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahlpw6_reg  (
    .clk(SWCLKTCK_pad),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zehpw6 [6]),
    .en(1'b1),
    .reset(1'b0),
    .set(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kxhpw6 ),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahlpw6 ));  // ../RTL/cortexm0ds_logic.v(17362)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Amupw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iauhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Amupw6 ));  // ../RTL/cortexm0ds_logic.v(17710)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aniax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G1vhu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[2] ));  // ../RTL/cortexm0ds_logic.v(18613)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aoeax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z54iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aoeax6 ));  // ../RTL/cortexm0ds_logic.v(18317)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Apcax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K84iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Md7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Apcax6 ));  // ../RTL/cortexm0ds_logic.v(18269)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aqlax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rkkiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hfkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[5] ));  // ../RTL/cortexm0ds_logic.v(18745)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ar1bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vruhu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ar1bx6 ));  // ../RTL/cortexm0ds_logic.v(19347)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Arnpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rgoiu6 ),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y5liu6 ),
    .reset(1'b0),
    .set(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_apsr_o[3] ));  // ../RTL/cortexm0ds_logic.v(17475)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Asupw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hfshu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Asupw6 ));  // ../RTL/cortexm0ds_logic.v(17718)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/At2bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ipthu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/At2bx6 ));  // ../RTL/cortexm0ds_logic.v(19455)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Axohu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 ));  // ../RTL/cortexm0ds_logic.v(17271)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aurpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Drkiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ddkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[7] ));  // ../RTL/cortexm0ds_logic.v(17630)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Auyax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [23]),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B3fiu6 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Auyax6 ));  // ../RTL/cortexm0ds_logic.v(19041)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Avzax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I4eiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R5eiu6 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Avzax6 ));  // ../RTL/cortexm0ds_logic.v(19149)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aw4bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [30]),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzeiu6 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aw4bx6 ));  // ../RTL/cortexm0ds_logic.v(19671)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Awupw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xrohu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[30] ));  // ../RTL/cortexm0ds_logic.v(17729)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Az3bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fsdiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J0fiu6 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Az3bx6 ));  // ../RTL/cortexm0ds_logic.v(19575)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Azpax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vx9iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ickiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[23] ));  // ../RTL/cortexm0ds_logic.v(18822)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B0spw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sokiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lf8iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[6] ));  // ../RTL/cortexm0ds_logic.v(17638)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B3gbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bvuhu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B3gbx6 ));  // ../RTL/cortexm0ds_logic.v(20037)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B4uax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vx9iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wckiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[23] ));  // ../RTL/cortexm0ds_logic.v(18897)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B5zpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sokiu6 ),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[4] ));  // ../RTL/cortexm0ds_logic.v(17898)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B6uax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K39iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wckiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[30] ));  // ../RTL/cortexm0ds_logic.v(18898)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B79bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q44iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n382 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B79bx6 ));  // ../RTL/cortexm0ds_logic.v(19810)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B7lpw6_reg  (
    .clk(SWCLKTCK_pad),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fwohu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kxhpw6 ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B7lpw6 ));  // ../RTL/cortexm0ds_logic.v(17331)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B8uax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D39iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wckiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[31] ));  // ../RTL/cortexm0ds_logic.v(18899)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B9eax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Df4iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Td7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B9eax6 ));  // ../RTL/cortexm0ds_logic.v(18304)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B9jbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ym4iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B9jbx6 ));  // ../RTL/cortexm0ds_logic.v(20186)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bauax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tx8iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wckiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[0] ));  // ../RTL/cortexm0ds_logic.v(18900)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bbjpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bomiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Afkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[12] ));  // ../RTL/cortexm0ds_logic.v(17232)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bc3bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qyohu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bc3bx6 ));  // ../RTL/cortexm0ds_logic.v(19509)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bcabx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [6]),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B3fiu6 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bcabx6 ));  // ../RTL/cortexm0ds_logic.v(19885)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bccax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gk4iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/He7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bccax6 ));  // ../RTL/cortexm0ds_logic.v(18257)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bcdbx6_reg  (
    .clk(SWCLKTCK_pad),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pzxhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bcdbx6 ));  // ../RTL/cortexm0ds_logic.v(19972)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bcgax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lm1iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Md7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bcgax6 ));  // ../RTL/cortexm0ds_logic.v(18404)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bciax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P2vhu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bciax6 ));  // ../RTL/cortexm0ds_logic.v(18577)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bclpw6_reg  (
    .clk(SWCLKTCK_pad),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zehpw6 [0]),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kxhpw6 ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bclpw6 ));  // ../RTL/cortexm0ds_logic.v(17344)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bdjpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bomiu6 ),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[10] ));  // ../RTL/cortexm0ds_logic.v(17233)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bf3qw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P7xhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bf3qw6 ));  // ../RTL/cortexm0ds_logic.v(18033)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bfjpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R5liu6 ),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y5liu6 ),
    .reset(1'b0),
    .set(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_apsr_o[2] ));  // ../RTL/cortexm0ds_logic.v(17238)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Biaax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X44iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qf7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Biaax6 ));  // ../RTL/cortexm0ds_logic.v(18186)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bk7ax6_reg  (
    .clk(SWCLKTCK_pad),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Li7ax6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C53iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bk7ax6 ));  // ../RTL/cortexm0ds_logic.v(18100)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bngax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F94iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Td7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bngax6 ));  // ../RTL/cortexm0ds_logic.v(18410)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bolax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jgkiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hfkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[3] ));  // ../RTL/cortexm0ds_logic.v(18744)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bp2qw6_reg  (
    .clk(SWCLKTCK_pad),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kn2qw6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C53iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bp2qw6 ));  // ../RTL/cortexm0ds_logic.v(17999)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bq9ax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gk4iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zg7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bq9ax6 ));  // ../RTL/cortexm0ds_logic.v(18171)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bsrpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Drkiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Afkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[7] ));  // ../RTL/cortexm0ds_logic.v(17629)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bt2qw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Df4iu6 ),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tu4iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bt2qw6 ));  // ../RTL/cortexm0ds_logic.v(18006)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Btbbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G64iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Md7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Btbbx6 ));  // ../RTL/cortexm0ds_logic.v(19938)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bu6bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vbphu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bu6bx6 ));  // ../RTL/cortexm0ds_logic.v(19762)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Buabx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L54iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Md7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Buabx6 ));  // ../RTL/cortexm0ds_logic.v(19895)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bvaax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ud4iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qf7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bvaax6 ));  // ../RTL/cortexm0ds_logic.v(18193)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bvfbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P74iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n382 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bvfbx6 ));  // ../RTL/cortexm0ds_logic.v(20019)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bwdax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E54iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Td7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bwdax6 ));  // ../RTL/cortexm0ds_logic.v(18297)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bx2qw6_reg  (
    .clk(SWCLKTCK_pad),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bsxhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bx2qw6 ));  // ../RTL/cortexm0ds_logic.v(18008)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bxbax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U64iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/He7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bxbax6 ));  // ../RTL/cortexm0ds_logic.v(18249)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bxpax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ef8iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ickiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[4] ));  // ../RTL/cortexm0ds_logic.v(18821)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C07bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V3qhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C07bx6 ));  // ../RTL/cortexm0ds_logic.v(19765)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C10bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pouhu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C10bx6 ));  // ../RTL/cortexm0ds_logic.v(19167)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C14bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [23]),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J0fiu6 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C14bx6 ));  // ../RTL/cortexm0ds_logic.v(19581)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C1fax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oh4iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C1fax6 ));  // ../RTL/cortexm0ds_logic.v(18324)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C1wpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hyuhu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C1wpw6 ));  // ../RTL/cortexm0ds_logic.v(17800)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C27bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vrmiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lf8iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[11] ));  // ../RTL/cortexm0ds_logic.v(19766)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C2uax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ef8iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wckiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[4] ));  // ../RTL/cortexm0ds_logic.v(18896)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C2ypw6_reg  (
    .clk(SWCLKTCK_pad),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L0ypw6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C53iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C2ypw6 ));  // ../RTL/cortexm0ds_logic.v(17858)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C30bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wouhu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C30bx6 ));  // ../RTL/cortexm0ds_logic.v(19173)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C37ax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Roohu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[22] ));  // ../RTL/cortexm0ds_logic.v(18085)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C3wpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tbvhu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C3wpw6 ));  // ../RTL/cortexm0ds_logic.v(17806)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C3zpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rkkiu6 ),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[3] ));  // ../RTL/cortexm0ds_logic.v(17897)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C47bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vrmiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mx8iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[11] ));  // ../RTL/cortexm0ds_logic.v(19767)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C4dax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J44iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Md7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C4dax6 ));  // ../RTL/cortexm0ds_logic.v(18277)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C50bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kpuhu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C50bx6 ));  // ../RTL/cortexm0ds_logic.v(19179)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C5gbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [22]),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dv9iu6 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C5gbx6 ));  // ../RTL/cortexm0ds_logic.v(20043)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C5wpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Admiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lf8iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[16] ));  // ../RTL/cortexm0ds_logic.v(17808)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C67bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vrmiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ickiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[11] ));  // ../RTL/cortexm0ds_logic.v(19768)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C72qw6_reg  (
    .clk(SWCLKTCK_pad),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1yhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C72qw6 ));  // ../RTL/cortexm0ds_logic.v(17964)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C7wpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Admiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mx8iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[16] ));  // ../RTL/cortexm0ds_logic.v(17809)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C87bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vrmiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pckiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[11] ));  // ../RTL/cortexm0ds_logic.v(19769)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C9wpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Admiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ofkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[16] ));  // ../RTL/cortexm0ds_logic.v(17810)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ca1bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Snthu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ca1bx6 ));  // ../RTL/cortexm0ds_logic.v(19299)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ca7bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vrmiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vfkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[11] ));  // ../RTL/cortexm0ds_logic.v(19770)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cbwpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Admiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Afkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[16] ));  // ../RTL/cortexm0ds_logic.v(17811)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cc2bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ltuhu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cc2bx6 ));  // ../RTL/cortexm0ds_logic.v(19407)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cc7bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vrmiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ofkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[11] ));  // ../RTL/cortexm0ds_logic.v(19771)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cccbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R84iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qf7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cccbx6 ));  // ../RTL/cortexm0ds_logic.v(19948)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cchax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Umohu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[18] ));  // ../RTL/cortexm0ds_logic.v(18483)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cdwpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Admiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ddkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[16] ));  // ../RTL/cortexm0ds_logic.v(17812)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ce7bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vrmiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hfkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[11] ));  // ../RTL/cortexm0ds_logic.v(19772)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ceabx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ldphu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ceabx6 ));  // ../RTL/cortexm0ds_logic.v(19887)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cfvpw6_reg  (
    .clk(SWCLKTCK_pad),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ldvpw6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C53iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cfvpw6 ));  // ../RTL/cortexm0ds_logic.v(17775)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cfwpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Admiu6 ),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[14] ));  // ../RTL/cortexm0ds_logic.v(17813)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cg7bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vrmiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Afkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[11] ));  // ../RTL/cortexm0ds_logic.v(19773)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cglax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vx9iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hfkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[23] ));  // ../RTL/cortexm0ds_logic.v(18740)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Chwpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sqqhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Chwpw6 ));  // ../RTL/cortexm0ds_logic.v(17814)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ci7bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vrmiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wckiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[11] ));  // ../RTL/cortexm0ds_logic.v(19774)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cilax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K39iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hfkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[30] ));  // ../RTL/cortexm0ds_logic.v(18741)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cjqpw6_reg  (
    .clk(SWCLKTCK_pad),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yfxhu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kxhpw6 ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cjqpw6 ));  // ../RTL/cortexm0ds_logic.v(17566)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cjwpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Maphu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cjwpw6 ));  // ../RTL/cortexm0ds_logic.v(17815)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ck7bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vrmiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ddkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[11] ));  // ../RTL/cortexm0ds_logic.v(19775)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cklax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D39iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hfkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[31] ));  // ../RTL/cortexm0ds_logic.v(18742)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cm7bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vrmiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kdkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[11] ));  // ../RTL/cortexm0ds_logic.v(19776)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cmlax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tx8iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hfkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[0] ));  // ../RTL/cortexm0ds_logic.v(18743)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cncbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U7phu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cncbx6 ));  // ../RTL/cortexm0ds_logic.v(19954)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cndbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B74iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qf7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cndbx6 ));  // ../RTL/cortexm0ds_logic.v(19978)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Co7bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vrmiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rdkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[11] ));  // ../RTL/cortexm0ds_logic.v(19777)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cokbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V2row6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cokbx6 ));  // ../RTL/cortexm0ds_logic.v(20266)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Coupw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S8uhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Coupw6 ));  // ../RTL/cortexm0ds_logic.v(17711)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cq3qw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M94iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n382 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cq3qw6 ));  // ../RTL/cortexm0ds_logic.v(18045)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cq7bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vcohu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[14] ));  // ../RTL/cortexm0ds_logic.v(19782)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cqrpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Drkiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ofkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[7] ));  // ../RTL/cortexm0ds_logic.v(17628)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cs6bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X6niu6 ),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztmiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[8] ));  // ../RTL/cortexm0ds_logic.v(19761)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cvpax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qcaiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ickiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[2] ));  // ../RTL/cortexm0ds_logic.v(18820)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cwyax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [30]),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B3fiu6 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cwyax6 ));  // ../RTL/cortexm0ds_logic.v(19047)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cxcbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y84iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/He7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cxcbx6 ));  // ../RTL/cortexm0ds_logic.v(19964)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cxzax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lmuhu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cxzax6 ));  // ../RTL/cortexm0ds_logic.v(19155)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cy4bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [31]),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzeiu6 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cy4bx6 ));  // ../RTL/cortexm0ds_logic.v(19677)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cydbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K9phu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cydbx6 ));  // ../RTL/cortexm0ds_logic.v(19984)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Czzax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nnuhu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Czzax6 ));  // ../RTL/cortexm0ds_logic.v(19161)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D0uax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qcaiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wckiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[2] ));  // ../RTL/cortexm0ds_logic.v(18895)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D12qw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mpohu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[27] ));  // ../RTL/cortexm0ds_logic.v(17955)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D1aax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T24iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qf7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D1aax6 ));  // ../RTL/cortexm0ds_logic.v(18177)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D1zpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jgkiu6 ),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[1] ));  // ../RTL/cortexm0ds_logic.v(17896)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D2opw6_reg  (
    .clk(SWCLKTCK_pad),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wsxhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D2opw6 ));  // ../RTL/cortexm0ds_logic.v(17492)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D2rpw6_reg  (
    .clk(SWCLKTCK_pad),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nfqpw6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C53iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D2rpw6 ));  // ../RTL/cortexm0ds_logic.v(17596)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D43qw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T2xhu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/dbgrst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D43qw6 ));  // ../RTL/cortexm0ds_logic.v(18021)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D46bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fyliu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pckiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[21] ));  // ../RTL/cortexm0ds_logic.v(19749)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D66bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E1miu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pckiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[20] ));  // ../RTL/cortexm0ds_logic.v(19750)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D70bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rpuhu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D70bx6 ));  // ../RTL/cortexm0ds_logic.v(19185)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D7gbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [22]),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F6eiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D7gbx6 ));  // ../RTL/cortexm0ds_logic.v(20045)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D86bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D4miu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pckiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[19] ));  // ../RTL/cortexm0ds_logic.v(19751)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D99ax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D84iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zg7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D99ax6 ));  // ../RTL/cortexm0ds_logic.v(18162)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Da6bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C7miu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pckiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[18] ));  // ../RTL/cortexm0ds_logic.v(19752)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Daebx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I74iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Daebx6 ));  // ../RTL/cortexm0ds_logic.v(19990)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Daiax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ajohu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Daiax6 ));  // ../RTL/cortexm0ds_logic.v(18571)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dc6bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bamiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pckiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[17] ));  // ../RTL/cortexm0ds_logic.v(19753)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/De6bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Admiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pckiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[16] ));  // ../RTL/cortexm0ds_logic.v(19754)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Delax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ef8iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hfkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[4] ));  // ../RTL/cortexm0ds_logic.v(18739)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dfbax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ud4iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cf7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dfbax6 ));  // ../RTL/cortexm0ds_logic.v(18224)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dg2qw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G6xhu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/dbgrst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dg2qw6 ));  // ../RTL/cortexm0ds_logic.v(17983)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dg6bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rimiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pckiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[14] ));  // ../RTL/cortexm0ds_logic.v(19755)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Di3qw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A3xhu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/dbgrst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Di3qw6 ));  // ../RTL/cortexm0ds_logic.v(18039)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Di6bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jlmiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pckiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[13] ));  // ../RTL/cortexm0ds_logic.v(19756)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dk6bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bomiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pckiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[12] ));  // ../RTL/cortexm0ds_logic.v(19757)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dk9bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xi4iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Td7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dk9bx6 ));  // ../RTL/cortexm0ds_logic.v(19817)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dm6bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K8qhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dm6bx6 ));  // ../RTL/cortexm0ds_logic.v(19758)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dmeax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N64iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dmeax6 ));  // ../RTL/cortexm0ds_logic.v(18316)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dncax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T94iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Md7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dncax6 ));  // ../RTL/cortexm0ds_logic.v(18268)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Do6bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hymiu6 ),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztmiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[10] ));  // ../RTL/cortexm0ds_logic.v(19759)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dorpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Drkiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mx8iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[7] ));  // ../RTL/cortexm0ds_logic.v(17627)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dpwpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z54iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n382 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dpwpw6 ));  // ../RTL/cortexm0ds_logic.v(17818)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dq6bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K3niu6 ),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztmiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[9] ));  // ../RTL/cortexm0ds_logic.v(19760)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dqkbx6_reg  (
    .clk(SWCLKTCK_pad),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I5nhu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kxhpw6 ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/dbg_swdo_en ));  // ../RTL/cortexm0ds_logic.v(20272)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Drcbx6_reg  (
    .clk(SWCLKTCK_pad),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S2cbx6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C53iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Drcbx6 ));  // ../RTL/cortexm0ds_logic.v(19961)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Drhax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qkohu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[5] ));  // ../RTL/cortexm0ds_logic.v(18531)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dt1bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I1phu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dt1bx6 ));  // ../RTL/cortexm0ds_logic.v(19353)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dtpax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X6niu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kdkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[8] ));  // ../RTL/cortexm0ds_logic.v(18819)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dugax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O34iu6 ),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M24iu6 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/dbgrst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dugax6 ));  // ../RTL/cortexm0ds_logic.v(18423)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dv2bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nwdpw6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dv2bx6 ));  // ../RTL/cortexm0ds_logic.v(19461)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gfvhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 ));  // ../RTL/cortexm0ds_logic.v(17793)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dzvpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rnbow6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G81ju6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dzvpw6 ));  // ../RTL/cortexm0ds_logic.v(17795)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E05bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [7]),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z1fiu6 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E05bx6 ));  // ../RTL/cortexm0ds_logic.v(19683)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E1npw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X1liu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lf8iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[27] ));  // ../RTL/cortexm0ds_logic.v(17448)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E34bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [30]),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J0fiu6 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E34bx6 ));  // ../RTL/cortexm0ds_logic.v(19587)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E3npw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P4liu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lf8iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[29] ));  // ../RTL/cortexm0ds_logic.v(17449)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E5npw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fyliu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lf8iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[21] ));  // ../RTL/cortexm0ds_logic.v(17450)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E5pax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hsliu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kdkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[25] ));  // ../RTL/cortexm0ds_logic.v(18807)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E6iax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H5vhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E6iax6 ));  // ../RTL/cortexm0ds_logic.v(18565)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E7npw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E1miu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lf8iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[20] ));  // ../RTL/cortexm0ds_logic.v(17451)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E7pax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fyliu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kdkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[21] ));  // ../RTL/cortexm0ds_logic.v(18808)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E8iax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D3vhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E8iax6 ));  // ../RTL/cortexm0ds_logic.v(18566)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E90bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ypuhu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E90bx6 ));  // ../RTL/cortexm0ds_logic.v(19191)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E97ax6_reg  (
    .clk(SWCLKTCK_pad),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sxxhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E97ax6 ));  // ../RTL/cortexm0ds_logic.v(18089)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E9npw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jlmiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lf8iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[13] ));  // ../RTL/cortexm0ds_logic.v(17452)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E9pax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E1miu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kdkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[20] ));  // ../RTL/cortexm0ds_logic.v(18809)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eafax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T24iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rc7iu6 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/dbgrst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eafax6 ));  // ../RTL/cortexm0ds_logic.v(18343)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eagax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lm1iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Td7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eagax6 ));  // ../RTL/cortexm0ds_logic.v(18403)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ebnpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bomiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lf8iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[12] ));  // ../RTL/cortexm0ds_logic.v(17453)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ebpax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D4miu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kdkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[19] ));  // ../RTL/cortexm0ds_logic.v(18810)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eclax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qcaiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hfkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[2] ));  // ../RTL/cortexm0ds_logic.v(18738)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ectax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hsliu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tekiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[25] ));  // ../RTL/cortexm0ds_logic.v(18883)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ednpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gfniu6 ),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Numiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[28] ));  // ../RTL/cortexm0ds_logic.v(17454)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Edpax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C7miu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kdkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[18] ));  // ../RTL/cortexm0ds_logic.v(18811)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ee3bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q6vhu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ee3bx6 ));  // ../RTL/cortexm0ds_logic.v(19515)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eetax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fyliu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tekiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[21] ));  // ../RTL/cortexm0ds_logic.v(18884)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Efdax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T24iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Md7iu6 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/dbgrst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Efdax6 ));  // ../RTL/cortexm0ds_logic.v(18287)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Efnpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D39iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Afkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[31] ));  // ../RTL/cortexm0ds_logic.v(17455)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Efpax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bamiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kdkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[17] ));  // ../RTL/cortexm0ds_logic.v(18812)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Egaax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E54iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qf7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Egaax6 ));  // ../RTL/cortexm0ds_logic.v(18185)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Egtax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E1miu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tekiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[20] ));  // ../RTL/cortexm0ds_logic.v(18885)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ehnpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D39iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lf8iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[31] ));  // ../RTL/cortexm0ds_logic.v(17456)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ehpax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Admiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kdkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[16] ));  // ../RTL/cortexm0ds_logic.v(18813)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ehqpw6_reg  (
    .clk(SWCLKTCK_pad),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nfqpw6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jq3iu6 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kxhpw6 ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ehqpw6 ));  // ../RTL/cortexm0ds_logic.v(17560)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eitax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D4miu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tekiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[19] ));  // ../RTL/cortexm0ds_logic.v(18886)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ejnpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D39iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mx8iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[31] ));  // ../RTL/cortexm0ds_logic.v(17457)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ejpax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rimiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kdkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[14] ));  // ../RTL/cortexm0ds_logic.v(18814)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ektax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C7miu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tekiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[18] ));  // ../RTL/cortexm0ds_logic.v(18887)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Elgax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F94iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Elgax6 ));  // ../RTL/cortexm0ds_logic.v(18409)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eliax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W2vhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[0] ));  // ../RTL/cortexm0ds_logic.v(18607)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Elnpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [31]),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aqgiu6 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Elnpw6 ));  // ../RTL/cortexm0ds_logic.v(17462)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Elpax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jlmiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kdkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[13] ));  // ../RTL/cortexm0ds_logic.v(18815)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Emrpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Drkiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lf8iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[7] ));  // ../RTL/cortexm0ds_logic.v(17626)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Emtax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bamiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tekiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[17] ));  // ../RTL/cortexm0ds_logic.v(18888)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Enpax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bomiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kdkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[12] ));  // ../RTL/cortexm0ds_logic.v(18816)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eotax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Admiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tekiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[16] ));  // ../RTL/cortexm0ds_logic.v(18889)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eppax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hymiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kdkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[10] ));  // ../RTL/cortexm0ds_logic.v(18817)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eqtax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rimiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tekiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[14] ));  // ../RTL/cortexm0ds_logic.v(18890)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Equpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Esohu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[6] ));  // ../RTL/cortexm0ds_logic.v(17716)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Erbbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G64iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Td7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Erbbx6 ));  // ../RTL/cortexm0ds_logic.v(19937)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Erpax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K3niu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kdkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[9] ));  // ../RTL/cortexm0ds_logic.v(18818)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Esabx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L54iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Td7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Esabx6 ));  // ../RTL/cortexm0ds_logic.v(19894)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Estax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jlmiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tekiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[13] ));  // ../RTL/cortexm0ds_logic.v(18891)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Etfbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P74iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Md7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Etfbx6 ));  // ../RTL/cortexm0ds_logic.v(20018)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eudax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S54iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Td7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eudax6 ));  // ../RTL/cortexm0ds_logic.v(18296)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eutax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bomiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tekiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[12] ));  // ../RTL/cortexm0ds_logic.v(18892)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Evbax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D84iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/He7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Evbax6 ));  // ../RTL/cortexm0ds_logic.v(18248)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Evhpw6_reg  (
    .clk(SWCLKTCK_pad),
    .d(1'b1),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/reset_sync_reg [2]),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Evhpw6 ));  // ../RTL/cortexm0ds_logic.v(17154)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Evypw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D39iu6 ),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[29] ));  // ../RTL/cortexm0ds_logic.v(17893)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ewtax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hymiu6 ),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Csmiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[10] ));  // ../RTL/cortexm0ds_logic.v(18893)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Exypw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K39iu6 ),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[28] ));  // ../RTL/cortexm0ds_logic.v(17894)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eytax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X6niu6 ),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Csmiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[8] ));  // ../RTL/cortexm0ds_logic.v(18894)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eyyax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [31]),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B3fiu6 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eyyax6 ));  // ../RTL/cortexm0ds_logic.v(19053)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ez1qw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K3niu6 ),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jsmiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[9] ));  // ../RTL/cortexm0ds_logic.v(17950)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ezypw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ef8iu6 ),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[2] ));  // ../RTL/cortexm0ds_logic.v(17895)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F17ax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rjthu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F17ax6 ));  // ../RTL/cortexm0ds_logic.v(18079)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F1pax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P4liu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kdkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[29] ));  // ../RTL/cortexm0ds_logic.v(18805)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F26bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Czmiu6 ),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jzmiu6 ),
    .reset(1'b0),
    .set(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F26bx6 ));  // ../RTL/cortexm0ds_logic.v(19747)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F2dax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X44iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Md7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F2dax6 ));  // ../RTL/cortexm0ds_logic.v(18276)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F2tax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zvkiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tekiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[24] ));  // ../RTL/cortexm0ds_logic.v(18878)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F3pax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uoliu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kdkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[1] ));  // ../RTL/cortexm0ds_logic.v(18806)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F4iax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I2vhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F4iax6 ));  // ../RTL/cortexm0ds_logic.v(18564)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F4ibx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uephu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/dbgrst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F4ibx6 ));  // ../RTL/cortexm0ds_logic.v(20159)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F4tax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fzkiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tekiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[26] ));  // ../RTL/cortexm0ds_logic.v(18879)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F59bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q44iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Md7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F59bx6 ));  // ../RTL/cortexm0ds_logic.v(19809)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F6dbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dsrhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F6dbx6 ));  // ../RTL/cortexm0ds_logic.v(19969)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F6tax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X1liu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tekiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[27] ));  // ../RTL/cortexm0ds_logic.v(18880)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F7eax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H34iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Td7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F7eax6 ));  // ../RTL/cortexm0ds_logic.v(18303)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F7jbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ym4iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/He7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F7jbx6 ));  // ../RTL/cortexm0ds_logic.v(20185)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F8cbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W5shu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F8cbx6 ));  // ../RTL/cortexm0ds_logic.v(19946)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F8dbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P8phu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F8dbx6 ));  // ../RTL/cortexm0ds_logic.v(19970)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F8tax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P4liu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tekiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[29] ));  // ../RTL/cortexm0ds_logic.v(18881)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F9gbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z8uhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F9gbx6 ));  // ../RTL/cortexm0ds_logic.v(20046)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F9vpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B0biu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n3685 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F9vpw6 ));  // ../RTL/cortexm0ds_logic.v(17771)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Facax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pl4iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/He7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Facax6 ));  // ../RTL/cortexm0ds_logic.v(18256)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Facbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R84iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zg7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Facbx6 ));  // ../RTL/cortexm0ds_logic.v(19947)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fahax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bnohu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[19] ));  // ../RTL/cortexm0ds_logic.v(18477)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fatax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uoliu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tekiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[1] ));  // ../RTL/cortexm0ds_logic.v(18882)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fb0bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fquhu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fb0bx6 ));  // ../RTL/cortexm0ds_logic.v(19197)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fc1bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F3phu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fc1bx6 ));  // ../RTL/cortexm0ds_logic.v(19305)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fe2bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N0phu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fe2bx6 ));  // ../RTL/cortexm0ds_logic.v(19413)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fj8ax6_reg  (
    .clk(SWCLKTCK_pad),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oh8ax6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C53iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fj8ax6 ));  // ../RTL/cortexm0ds_logic.v(18123)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fjdbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A9rhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fjdbx6 ));  // ../RTL/cortexm0ds_logic.v(19976)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fkrpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssohu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fkrpw6 ));  // ../RTL/cortexm0ds_logic.v(17625)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fl2qw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B8phu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fl2qw6 ));  // ../RTL/cortexm0ds_logic.v(17997)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fldbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B74iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zg7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fldbx6 ));  // ../RTL/cortexm0ds_logic.v(19977)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fm7ax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ud4iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fd7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fm7ax6 ));  // ../RTL/cortexm0ds_logic.v(18101)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fnnpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Puohu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fnnpw6 ));  // ../RTL/cortexm0ds_logic.v(17468)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fo9ax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pl4iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zg7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fo9ax6 ));  // ../RTL/cortexm0ds_logic.v(18170)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fpnpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iuohu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fpnpw6 ));  // ../RTL/cortexm0ds_logic.v(17470)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ftaax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Df4iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qf7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ftaax6 ));  // ../RTL/cortexm0ds_logic.v(18192)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ftypw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qcaiu6 ),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[0] ));  // ../RTL/cortexm0ds_logic.v(17892)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fvcbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y84iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qf7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fvcbx6 ));  // ../RTL/cortexm0ds_logic.v(19963)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fvoax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zvkiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kdkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[24] ));  // ../RTL/cortexm0ds_logic.v(18802)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fx1qw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K3niu6 ),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qsmiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[9] ));  // ../RTL/cortexm0ds_logic.v(17949)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fxoax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fzkiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kdkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[26] ));  // ../RTL/cortexm0ds_logic.v(18803)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fzmpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rkkiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lf8iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[5] ));  // ../RTL/cortexm0ds_logic.v(17447)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fzoax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X1liu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kdkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[27] ));  // ../RTL/cortexm0ds_logic.v(18804)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G0tax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Drkiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tekiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[7] ));  // ../RTL/cortexm0ds_logic.v(18877)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G0zax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I4eiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P3fiu6 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G0zax6 ));  // ../RTL/cortexm0ds_logic.v(19059)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G25bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [14]),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z1fiu6 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G25bx6 ));  // ../RTL/cortexm0ds_logic.v(19689)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G2iax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B2vhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G2iax6 ));  // ../RTL/cortexm0ds_logic.v(18563)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G54bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [31]),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J0fiu6 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G54bx6 ));  // ../RTL/cortexm0ds_logic.v(19593)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G79ax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K84iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zg7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G79ax6 ));  // ../RTL/cortexm0ds_logic.v(18161)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G8ebx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I74iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/He7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G8ebx6 ));  // ../RTL/cortexm0ds_logic.v(19989)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gbvpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R9phu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gbvpw6 ));  // ../RTL/cortexm0ds_logic.v(17773)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gc1qw6_reg  (
    .clk(SWCLKTCK_pad),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qa1qw6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C53iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gc1qw6 ));  // ../RTL/cortexm0ds_logic.v(17938)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gd0bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tquhu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gd0bx6 ));  // ../RTL/cortexm0ds_logic.v(19203)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ggabx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hbphu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ggabx6 ));  // ../RTL/cortexm0ds_logic.v(19888)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gihbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H4phu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gihbx6 ));  // ../RTL/cortexm0ds_logic.v(20118)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gkeax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U64iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gkeax6 ));  // ../RTL/cortexm0ds_logic.v(18315)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gl1qw6_reg  (
    .clk(SWCLKTCK_pad),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qj1qw6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C53iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gl1qw6 ));  // ../RTL/cortexm0ds_logic.v(17943)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gnqpw6_reg  (
    .clk(SWCLKTCK_pad),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Krlpw6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C53iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gnqpw6 ));  // ../RTL/cortexm0ds_logic.v(17574)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Golpw6_reg  (
    .clk(SWCLKTCK_pad),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rilpw6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U03iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Golpw6 ));  // ../RTL/cortexm0ds_logic.v(17382)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gp6ax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vx9iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n1552 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[21] ));  // ../RTL/cortexm0ds_logic.v(18064)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gpqpw6_reg  (
    .clk(SWCLKTCK_pad),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vplpw6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C53iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gpqpw6 ));  // ../RTL/cortexm0ds_logic.v(17575)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gr2qw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T24iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fd7iu6 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/dbgrst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gr2qw6 ));  // ../RTL/cortexm0ds_logic.v(18004)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gr6ax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vx9iu6 ),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[21] ));  // ../RTL/cortexm0ds_logic.v(18065)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gt6ax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vx9iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ddkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[23] ));  // ../RTL/cortexm0ds_logic.v(18066)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gtoax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Drkiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kdkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[7] ));  // ../RTL/cortexm0ds_logic.v(18801)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gv1bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgthu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gv1bx6 ));  // ../RTL/cortexm0ds_logic.v(19359)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gv1qw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K3niu6 ),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Etmiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[9] ));  // ../RTL/cortexm0ds_logic.v(17948)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gv6ax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vx9iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lf8iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[23] ));  // ../RTL/cortexm0ds_logic.v(18067)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gvmpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K39iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lf8iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[30] ));  // ../RTL/cortexm0ds_logic.v(17445)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gw6bx6_reg  (
    .clk(SWCLKTCK_pad),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qwxhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gw6bx6 ));  // ../RTL/cortexm0ds_logic.v(19763)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gwwpw6_reg  (
    .clk(SWCLKTCK_pad),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Puwpw6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C53iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gwwpw6 ));  // ../RTL/cortexm0ds_logic.v(17827)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gwxpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gzphu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gwxpw6 ));  // ../RTL/cortexm0ds_logic.v(17855)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gx2bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wpthu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gx2bx6 ));  // ../RTL/cortexm0ds_logic.v(19467)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gx6ax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vx9iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mx8iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[23] ));  // ../RTL/cortexm0ds_logic.v(18068)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gxmpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jgkiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lf8iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[3] ));  // ../RTL/cortexm0ds_logic.v(17446)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gylpw6_reg  (
    .clk(SWCLKTCK_pad),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mmyhu6 ),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U73iu6 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kxhpw6 ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gylpw6 ));  // ../RTL/cortexm0ds_logic.v(17402)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gyxpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ccphu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gyxpw6 ));  // ../RTL/cortexm0ds_logic.v(17856)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gz6ax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [23]),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aqgiu6 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gz6ax6 ));  // ../RTL/cortexm0ds_logic.v(18073)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gzeax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gk4iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gzeax6 ));  // ../RTL/cortexm0ds_logic.v(18323)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H0ebx6_reg  (
    .clk(SWCLKTCK_pad),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sddbx6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C53iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H0ebx6 ));  // ../RTL/cortexm0ds_logic.v(19985)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H3lpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6phu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H3lpw6 ));  // ../RTL/cortexm0ds_logic.v(17325)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H4bax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T24iu6 ),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oe7iu6 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/dbgrst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H4bax6 ));  // ../RTL/cortexm0ds_logic.v(18217)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H4ypw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J44iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n382 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H4ypw6 ));  // ../RTL/cortexm0ds_logic.v(17859)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H4zax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [7]),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L1fiu6 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H4zax6 ));  // ../RTL/cortexm0ds_logic.v(19071)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H7hbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W74iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n382 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H7hbx6 ));  // ../RTL/cortexm0ds_logic.v(20103)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H8gax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lm1iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H8gax6 ));  // ../RTL/cortexm0ds_logic.v(18402)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Halax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z7vhu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Halax6 ));  // ../RTL/cortexm0ds_logic.v(18736)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hbgbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [22]),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzeiu6 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hbgbx6 ));  // ../RTL/cortexm0ds_logic.v(20051)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hdbax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O34iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cf7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hdbax6 ));  // ../RTL/cortexm0ds_logic.v(18223)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hdfax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J44iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rc7iu6 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/dbgrst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hdfax6 ));  // ../RTL/cortexm0ds_logic.v(18355)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Heaax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S54iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qf7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Heaax6 ));  // ../RTL/cortexm0ds_logic.v(18184)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hf0bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hruhu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hf0bx6 ));  // ../RTL/cortexm0ds_logic.v(19209)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hg3bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cyohu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hg3bx6 ));  // ../RTL/cortexm0ds_logic.v(19521)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hg7ax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gephu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hg7ax6 ));  // ../RTL/cortexm0ds_logic.v(18098)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hgrpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X4xhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hgrpw6 ));  // ../RTL/cortexm0ds_logic.v(17617)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hhvpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [19]),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F6eiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hhvpw6 ));  // ../RTL/cortexm0ds_logic.v(17776)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hi9bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xi4iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hi9bx6 ));  // ../RTL/cortexm0ds_logic.v(19816)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsohu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ));  // ../RTL/cortexm0ds_logic.v(17623)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hjgax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F94iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/He7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hjgax6 ));  // ../RTL/cortexm0ds_logic.v(18408)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hkxpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hymiu6 ),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Numiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[10] ));  // ../RTL/cortexm0ds_logic.v(17849)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hlcax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ud4iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Md7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hlcax6 ));  // ../RTL/cortexm0ds_logic.v(18267)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hlwpw6_reg  (
    .clk(SWCLKTCK_pad),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zxxhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hlwpw6 ));  // ../RTL/cortexm0ds_logic.v(17816)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hmbax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n853 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/dbgrst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hmbax6 ));  // ../RTL/cortexm0ds_logic.v(18237)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hmxpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hymiu6 ),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gumiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[10] ));  // ../RTL/cortexm0ds_logic.v(17850)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hoxpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hymiu6 ),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ltmiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[10] ));  // ../RTL/cortexm0ds_logic.v(17851)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hpbbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G64iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hpbbx6 ));  // ../RTL/cortexm0ds_logic.v(19936)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hpcbx6_reg  (
    .clk(SWCLKTCK_pad),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J4cbx6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jq3iu6 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kxhpw6 ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hpcbx6 ));  // ../RTL/cortexm0ds_logic.v(19959)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hphax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xkohu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[7] ));  // ../RTL/cortexm0ds_logic.v(18525)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hqabx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L54iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hqabx6 ));  // ../RTL/cortexm0ds_logic.v(19893)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hqxpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hymiu6 ),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Etmiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[10] ));  // ../RTL/cortexm0ds_logic.v(17852)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hrfbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P74iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Td7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hrfbx6 ));  // ../RTL/cortexm0ds_logic.v(20017)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hroax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sokiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kdkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[6] ));  // ../RTL/cortexm0ds_logic.v(18800)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hsdax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z54iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Td7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hsdax6 ));  // ../RTL/cortexm0ds_logic.v(18295)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hsxpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hymiu6 ),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qsmiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[10] ));  // ../RTL/cortexm0ds_logic.v(17853)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ht1qw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K3niu6 ),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ltmiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[9] ));  // ../RTL/cortexm0ds_logic.v(17947)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Htbax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K84iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/He7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Htbax6 ));  // ../RTL/cortexm0ds_logic.v(18247)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Htmpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fi1ju6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O25iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Htmpw6 ));  // ../RTL/cortexm0ds_logic.v(17444)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Huxpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hymiu6 ),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[8] ));  // ../RTL/cortexm0ds_logic.v(17854)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hw8ax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y1xhu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/dbgrst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hw8ax6 ));  // ../RTL/cortexm0ds_logic.v(18139)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hwhpw6_reg  (
    .clk(SWCLKTCK_pad),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Evhpw6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/reset_sync_reg [2]),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hwhpw6 ));  // ../RTL/cortexm0ds_logic.v(17160)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hysax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sokiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tekiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[6] ));  // ../RTL/cortexm0ds_logic.v(18876)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hz9ax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O34iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zg7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hz9ax6 ));  // ../RTL/cortexm0ds_logic.v(18176)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I0dax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E54iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Md7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I0dax6 ));  // ../RTL/cortexm0ds_logic.v(18275)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I0opw6_reg  (
    .clk(SWCLKTCK_pad),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q3yhu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kxhpw6 ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I0opw6 ));  // ../RTL/cortexm0ds_logic.v(17490)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I1lpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qdvhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I1lpw6 ));  // ../RTL/cortexm0ds_logic.v(17324)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I1qpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fyliu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mx8iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[21] ));  // ../RTL/cortexm0ds_logic.v(17548)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I2zax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G3eiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P3fiu6 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I2zax6 ));  // ../RTL/cortexm0ds_logic.v(19065)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I3qpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E1miu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mx8iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[20] ));  // ../RTL/cortexm0ds_logic.v(17549)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I45bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fsdiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z1fiu6 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I45bx6 ));  // ../RTL/cortexm0ds_logic.v(19695)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I4rpw6_reg  (
    .clk(SWCLKTCK_pad),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L5lpw6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C53iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I4rpw6 ));  // ../RTL/cortexm0ds_logic.v(17597)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I5qpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jlmiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mx8iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[13] ));  // ../RTL/cortexm0ds_logic.v(17550)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I5xax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hcvhu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I5xax6 ));  // ../RTL/cortexm0ds_logic.v(18956)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I74bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [7]),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N2fiu6 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I74bx6 ));  // ../RTL/cortexm0ds_logic.v(19599)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I7qpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bomiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mx8iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[12] ));  // ../RTL/cortexm0ds_logic.v(17551)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I8hax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Inohu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[20] ));  // ../RTL/cortexm0ds_logic.v(18471)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I8lax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fnpiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I8lax6 ));  // ../RTL/cortexm0ds_logic.v(18730)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I9qpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gfniu6 ),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gumiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[28] ));  // ../RTL/cortexm0ds_logic.v(17552)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ibqpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zkphu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ibqpw6 ));  // ../RTL/cortexm0ds_logic.v(17553)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iddax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Df4iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Md7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iddax6 ));  // ../RTL/cortexm0ds_logic.v(18282)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idqpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G7phu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idqpw6 ));  // ../RTL/cortexm0ds_logic.v(17554)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iekax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W7iiu6 ),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D8iiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iekax6 ));  // ../RTL/cortexm0ds_logic.v(18701)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ig2bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztuhu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ig2bx6 ));  // ../RTL/cortexm0ds_logic.v(19419)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ih0bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oruhu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ih0bx6 ));  // ../RTL/cortexm0ds_logic.v(19215)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iixpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H25iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O25iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iixpw6 ));  // ../RTL/cortexm0ds_logic.v(17848)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ijiax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ctthu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[4] ));  // ../RTL/cortexm0ds_logic.v(18601)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ikhbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gnuhu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ikhbx6 ));  // ../RTL/cortexm0ds_logic.v(20124)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Im9ax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J44iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zg7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Im9ax6 ));  // ../RTL/cortexm0ds_logic.v(18169)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Imhbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [4]),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F6eiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Imhbx6 ));  // ../RTL/cortexm0ds_logic.v(20126)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ipoax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rkkiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kdkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[5] ));  // ../RTL/cortexm0ds_logic.v(18799)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ir1qw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K3niu6 ),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gumiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[9] ));  // ../RTL/cortexm0ds_logic.v(17946)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Irmpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uhthu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Irmpw6 ));  // ../RTL/cortexm0ds_logic.v(17442)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Isjpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dt4iu6 ),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kt4iu6 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/dbgrst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Isjpw6 ));  // ../RTL/cortexm0ds_logic.v(17265)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Itcbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y84iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zg7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Itcbx6 ));  // ../RTL/cortexm0ds_logic.v(19962)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iwsax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rkkiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tekiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[5] ));  // ../RTL/cortexm0ds_logic.v(18875)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ixppw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X1liu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mx8iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[27] ));  // ../RTL/cortexm0ds_logic.v(17546)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Izppw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P4liu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mx8iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[29] ));  // ../RTL/cortexm0ds_logic.v(17547)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J06bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cdohu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[8] ));  // ../RTL/cortexm0ds_logic.v(19741)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J0gax6_reg  (
    .clk(SWCLKTCK_pad),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H43iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C53iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J0gax6 ));  // ../RTL/cortexm0ds_logic.v(18398)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J0iax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hjohu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J0iax6 ));  // ../RTL/cortexm0ds_logic.v(18561)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J39bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q44iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Td7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J39bx6 ));  // ../RTL/cortexm0ds_logic.v(19808)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J3xax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ef8iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pckiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[4] ));  // ../RTL/cortexm0ds_logic.v(18951)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J4cbx6_reg  (
    .clk(SWCLKTCK_pad),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R0yhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J4cbx6 ));  // ../RTL/cortexm0ds_logic.v(19944)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J59ax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T94iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zg7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J59ax6 ));  // ../RTL/cortexm0ds_logic.v(18160)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J5eax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oh4iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Td7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J5eax6 ));  // ../RTL/cortexm0ds_logic.v(18302)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J5jbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ym4iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qf7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J5jbx6 ));  // ../RTL/cortexm0ds_logic.v(20184)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J6ebx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I74iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qf7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J6ebx6 ));  // ../RTL/cortexm0ds_logic.v(19988)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J6zax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [14]),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L1fiu6 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J6zax6 ));  // ../RTL/cortexm0ds_logic.v(19077)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J7xax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [23]),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F6eiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J7xax6 ));  // ../RTL/cortexm0ds_logic.v(18958)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J8cax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J44iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/He7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J8cax6 ));  // ../RTL/cortexm0ds_logic.v(18255)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jckax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pithu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jckax6 ));  // ../RTL/cortexm0ds_logic.v(18699)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jdgbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [22]),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J0fiu6 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jdgbx6 ));  // ../RTL/cortexm0ds_logic.v(20057)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jfdbx6_reg  (
    .clk(SWCLKTCK_pad),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bzxhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jfdbx6 ));  // ../RTL/cortexm0ds_logic.v(19974)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jflpw6_reg  (
    .clk(SWCLKTCK_pad),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zehpw6 [3]),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kxhpw6 ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jflpw6 ));  // ../RTL/cortexm0ds_logic.v(17356)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jgxpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iithu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jgxpw6 ));  // ../RTL/cortexm0ds_logic.v(17846)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jhebx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D9phu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jhebx6 ));  // ../RTL/cortexm0ds_logic.v(19994)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jieax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D84iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jieax6 ));  // ../RTL/cortexm0ds_logic.v(18314)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jj0bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Csuhu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jj0bx6 ));  // ../RTL/cortexm0ds_logic.v(19221)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jjvpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D4miu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lf8iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[19] ));  // ../RTL/cortexm0ds_logic.v(17777)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jl3qw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N64iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n382 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jl3qw6 ));  // ../RTL/cortexm0ds_logic.v(18042)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jlvpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D4miu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mx8iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[19] ));  // ../RTL/cortexm0ds_logic.v(17778)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jnoax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jgkiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kdkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[3] ));  // ../RTL/cortexm0ds_logic.v(18798)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jnvpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D4miu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ofkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[19] ));  // ../RTL/cortexm0ds_logic.v(17779)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Johbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vduhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Johbx6 ));  // ../RTL/cortexm0ds_logic.v(20127)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jp1qw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K3niu6 ),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Numiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[9] ));  // ../RTL/cortexm0ds_logic.v(17945)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jp9bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Osthu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jp9bx6 ));  // ../RTL/cortexm0ds_logic.v(19824)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jpmpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N1vhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jpmpw6 ));  // ../RTL/cortexm0ds_logic.v(17437)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jpvpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D4miu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Afkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[19] ));  // ../RTL/cortexm0ds_logic.v(17780)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jraax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H34iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qf7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jraax6 ));  // ../RTL/cortexm0ds_logic.v(18191)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jrvpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D4miu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ddkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[19] ));  // ../RTL/cortexm0ds_logic.v(17781)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jrypw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cy9iu6 ),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jy9iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jrypw6 ));  // ../RTL/cortexm0ds_logic.v(17891)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jtvpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D4miu6 ),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[17] ));  // ../RTL/cortexm0ds_logic.v(17782)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jusax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jgkiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tekiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[3] ));  // ../RTL/cortexm0ds_logic.v(18874)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jvkpw6_reg  (
    .clk(SWCLKTCK_pad),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Stkpw6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C53iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jvkpw6 ));  // ../RTL/cortexm0ds_logic.v(17311)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jvppw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rkkiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mx8iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[5] ));  // ../RTL/cortexm0ds_logic.v(17545)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jvvpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dhvhu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/dbgrst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jvvpw6 ));  // ../RTL/cortexm0ds_logic.v(17787)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jx1bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P1phu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jx1bx6 ));  // ../RTL/cortexm0ds_logic.v(19365)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jxgax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V3xhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/dbgrst_reg ),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jxgax6 ));  // ../RTL/cortexm0ds_logic.v(18435)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jy5bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hsliu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pckiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[25] ));  // ../RTL/cortexm0ds_logic.v(19736)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jz2bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lzohu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jz2bx6 ));  // ../RTL/cortexm0ds_logic.v(19473)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K1xax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qcaiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pckiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[2] ));  // ../RTL/cortexm0ds_logic.v(18950)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K5hbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W74iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Md7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K5hbx6 ));  // ../RTL/cortexm0ds_logic.v(20102)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K65bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [23]),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z1fiu6 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K65bx6 ));  // ../RTL/cortexm0ds_logic.v(19701)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K6gax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lm1iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/He7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K6gax6 ));  // ../RTL/cortexm0ds_logic.v(18401)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K7vpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vyuhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/dbgrst_reg ),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/DBGRESTARTED ));  // ../RTL/cortexm0ds_logic.v(17765)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K94bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [14]),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N2fiu6 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K94bx6 ));  // ../RTL/cortexm0ds_logic.v(19605)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kadbx6_reg  (
    .clk(SWCLKTCK_pad),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wzxhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kadbx6 ));  // ../RTL/cortexm0ds_logic.v(19971)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kakax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Seohu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kakax6 ));  // ../RTL/cortexm0ds_logic.v(18694)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kalpw6_reg  (
    .clk(SWCLKTCK_pad),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zehpw6 [2]),
    .en(1'b1),
    .reset(1'b0),
    .set(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kxhpw6 ),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kalpw6 ));  // ../RTL/cortexm0ds_logic.v(17338)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kcaax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z54iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qf7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kcaax6 ));  // ../RTL/cortexm0ds_logic.v(18183)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ke1qw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U6xhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ke1qw6 ));  // ../RTL/cortexm0ds_logic.v(17939)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kfoax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vx9iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kdkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[23] ));  // ../RTL/cortexm0ds_logic.v(18794)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Khgax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F94iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qf7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Khgax6 ));  // ../RTL/cortexm0ds_logic.v(18407)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Khoax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K39iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kdkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[30] ));  // ../RTL/cortexm0ds_logic.v(18795)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kjoax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D39iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kdkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[31] ));  // ../RTL/cortexm0ds_logic.v(18796)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kkjpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P4liu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Afkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[29] ));  // ../RTL/cortexm0ds_logic.v(17247)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kl0bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qsuhu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kl0bx6 ));  // ../RTL/cortexm0ds_logic.v(19227)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kl8ax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E54iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n382 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kl8ax6 ));  // ../RTL/cortexm0ds_logic.v(18124)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kloax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tx8iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kdkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[0] ));  // ../RTL/cortexm0ds_logic.v(18797)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kmjpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P4liu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vfkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[29] ));  // ../RTL/cortexm0ds_logic.v(17248)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kmsax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vx9iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tekiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[23] ));  // ../RTL/cortexm0ds_logic.v(18870)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kn1qw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kuphu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kn1qw6 ));  // ../RTL/cortexm0ds_logic.v(17944)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kn2qw6_reg  (
    .clk(SWCLKTCK_pad),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K0yhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kn2qw6 ));  // ../RTL/cortexm0ds_logic.v(17998)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Knbbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G64iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/He7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Knbbx6 ));  // ../RTL/cortexm0ds_logic.v(19935)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Knhax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Elohu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[11] ));  // ../RTL/cortexm0ds_logic.v(18519)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Koabx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L54iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/He7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Koabx6 ));  // ../RTL/cortexm0ds_logic.v(19892)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kojpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mxuhu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kojpw6 ));  // ../RTL/cortexm0ds_logic.v(17253)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kosax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K39iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tekiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[30] ));  // ../RTL/cortexm0ds_logic.v(18871)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kpfbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P74iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kpfbx6 ));  // ../RTL/cortexm0ds_logic.v(20016)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kqdax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N64iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Td7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kqdax6 ));  // ../RTL/cortexm0ds_logic.v(18294)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kqhbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [4]),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P3fiu6 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kqhbx6 ));  // ../RTL/cortexm0ds_logic.v(20132)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kqsax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D39iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tekiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[31] ));  // ../RTL/cortexm0ds_logic.v(18872)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Krbax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T94iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/He7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Krbax6 ));  // ../RTL/cortexm0ds_logic.v(18246)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Krlpw6_reg  (
    .clk(SWCLKTCK_pad),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vplpw6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U03iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Krlpw6 ));  // ../RTL/cortexm0ds_logic.v(17384)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ksgax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F24iu6 ),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M24iu6 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/dbgrst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ksgax6 ));  // ../RTL/cortexm0ds_logic.v(18417)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kssax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tx8iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tekiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[0] ));  // ../RTL/cortexm0ds_logic.v(18873)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kswpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y9phu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kswpw6 ));  // ../RTL/cortexm0ds_logic.v(17825)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ktppw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jgkiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mx8iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[3] ));  // ../RTL/cortexm0ds_logic.v(17544)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kwlpw6_reg  (
    .clk(SWCLKTCK_pad),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L5lpw6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jq3iu6 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kxhpw6 ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kwlpw6 ));  // ../RTL/cortexm0ds_logic.v(17396)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kxeax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pl4iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kxeax6 ));  // ../RTL/cortexm0ds_logic.v(18322)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kxhpw6_reg  (
    .clk(SWCLKTCK_pad),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hwhpw6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/reset_sync_reg [2]),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kxhpw6 ));  // ../RTL/cortexm0ds_logic.v(17166)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kzabx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jeuhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kzabx6 ));  // ../RTL/cortexm0ds_logic.v(19903)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L03qw6_reg  (
    .clk(SWCLKTCK_pad),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bx2qw6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C53iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L03qw6 ));  // ../RTL/cortexm0ds_logic.v(18015)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L0ypw6_reg  (
    .clk(SWCLKTCK_pad),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jwxhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L0ypw6 ));  // ../RTL/cortexm0ds_logic.v(17857)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L1bbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Smuhu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L1bbx6 ));  // ../RTL/cortexm0ds_logic.v(19908)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L2bax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O34iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xf7iu6 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/dbgrst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L2bax6 ));  // ../RTL/cortexm0ds_logic.v(18211)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L4lax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wfphu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L4lax6 ));  // ../RTL/cortexm0ds_logic.v(18718)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L5lpw6_reg  (
    .clk(SWCLKTCK_pad),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zqxhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L5lpw6 ));  // ../RTL/cortexm0ds_logic.v(17326)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6hax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pnohu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[23] ));  // ../RTL/cortexm0ds_logic.v(18465)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6lax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qqiow6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ),
    .reset(1'b0),
    .set(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6lax6 ));  // ../RTL/cortexm0ds_logic.v(18724)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L8kax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zeohu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L8kax6 ));  // ../RTL/cortexm0ds_logic.v(18693)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L8zax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fsdiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L1fiu6 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L8zax6 ));  // ../RTL/cortexm0ds_logic.v(19083)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L9bbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nephu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L9bbx6 ));  // ../RTL/cortexm0ds_logic.v(19928)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L9xax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fsdiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F6eiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L9xax6 ));  // ../RTL/cortexm0ds_logic.v(18959)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lbbax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H34iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lg7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lbbax6 ));  // ../RTL/cortexm0ds_logic.v(18222)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ldoax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ef8iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kdkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[4] ));  // ../RTL/cortexm0ds_logic.v(18793)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ldvpw6_reg  (
    .clk(SWCLKTCK_pad),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uyxhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ldvpw6 ));  // ../RTL/cortexm0ds_logic.v(17774)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ldwax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hsliu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rdkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[25] ));  // ../RTL/cortexm0ds_logic.v(18938)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Le2qw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F2xhu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/dbgrst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Le2qw6 ));  // ../RTL/cortexm0ds_logic.v(17977)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lerpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gtohu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[0] ));  // ../RTL/cortexm0ds_logic.v(17611)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lfgbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [22]),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X0fiu6 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lfgbx6 ));  // ../RTL/cortexm0ds_logic.v(20063)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lfppw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X1liu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ddkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[27] ));  // ../RTL/cortexm0ds_logic.v(17537)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lfwax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fyliu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rdkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[21] ));  // ../RTL/cortexm0ds_logic.v(18939)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lg1bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y2phu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lg1bx6 ));  // ../RTL/cortexm0ds_logic.v(19317)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lg9bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xi4iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/He7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lg9bx6 ));  // ../RTL/cortexm0ds_logic.v(19815)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lgkax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qfthu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lgkax6 ));  // ../RTL/cortexm0ds_logic.v(18702)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lhbbx6_reg  (
    .clk(SWCLKTCK_pad),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufbbx6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C53iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lhbbx6 ));  // ../RTL/cortexm0ds_logic.v(19932)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lhppw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P4liu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ddkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[29] ));  // ../RTL/cortexm0ds_logic.v(17538)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lhwax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E1miu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rdkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[20] ));  // ../RTL/cortexm0ds_logic.v(18940)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Li2bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G0phu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Li2bx6 ));  // ../RTL/cortexm0ds_logic.v(19425)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Li7ax6_reg  (
    .clk(SWCLKTCK_pad),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Urxhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Li7ax6 ));  // ../RTL/cortexm0ds_logic.v(18099)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Liabx6_reg  (
    .clk(SWCLKTCK_pad),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xf8ax6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C53iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Liabx6 ));  // ../RTL/cortexm0ds_logic.v(19889)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljcax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T24iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/He7iu6 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/dbgrst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljcax6 ));  // ../RTL/cortexm0ds_logic.v(18265)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljppw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fyliu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ddkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[21] ));  // ../RTL/cortexm0ds_logic.v(17539)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljwax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D4miu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rdkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[19] ));  // ../RTL/cortexm0ds_logic.v(18941)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lk9ax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X44iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zg7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lk9ax6 ));  // ../RTL/cortexm0ds_logic.v(18168)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lksax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ef8iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tekiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[4] ));  // ../RTL/cortexm0ds_logic.v(18869)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Llppw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E1miu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ddkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[20] ));  // ../RTL/cortexm0ds_logic.v(17540)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Llwax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C7miu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rdkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[18] ));  // ../RTL/cortexm0ds_logic.v(18942)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lmkbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pfphu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/dbgrst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lmkbx6 ));  // ../RTL/cortexm0ds_logic.v(20260)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ln0bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Etuhu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ln0bx6 ));  // ../RTL/cortexm0ds_logic.v(19233)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lnppw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jlmiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ddkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[13] ));  // ../RTL/cortexm0ds_logic.v(17541)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lnwax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bamiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rdkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[17] ));  // ../RTL/cortexm0ds_logic.v(18943)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lpppw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bomiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ddkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[12] ));  // ../RTL/cortexm0ds_logic.v(17542)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lpwax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Admiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rdkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[16] ));  // ../RTL/cortexm0ds_logic.v(18944)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lqjpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hxohu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[28] ));  // ../RTL/cortexm0ds_logic.v(17259)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lr9bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T3phu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lr9bx6 ));  // ../RTL/cortexm0ds_logic.v(19830)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lrppw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ef8iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mx8iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[4] ));  // ../RTL/cortexm0ds_logic.v(17543)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lrwax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rimiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rdkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[14] ));  // ../RTL/cortexm0ds_logic.v(18945)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ltwax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jlmiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rdkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[13] ));  // ../RTL/cortexm0ds_logic.v(18946)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lvwax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bomiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rdkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[12] ));  // ../RTL/cortexm0ds_logic.v(18947)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lx9ax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ud4iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zg7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lx9ax6 ));  // ../RTL/cortexm0ds_logic.v(18175)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lxwax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hymiu6 ),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jsmiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[10] ));  // ../RTL/cortexm0ds_logic.v(18948)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lycax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S54iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Md7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lycax6 ));  // ../RTL/cortexm0ds_logic.v(18274)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lywpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [18]),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F6eiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lywpw6 ));  // ../RTL/cortexm0ds_logic.v(17828)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lzwax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X6niu6 ),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jsmiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[8] ));  // ../RTL/cortexm0ds_logic.v(18949)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M13bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dqthu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M13bx6 ));  // ../RTL/cortexm0ds_logic.v(19479)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M2ebx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pdrhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M2ebx6 ));  // ../RTL/cortexm0ds_logic.v(19986)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M2lax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tx8iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mx8iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[0] ));  // ../RTL/cortexm0ds_logic.v(18713)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M3wax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zvkiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rdkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[24] ));  // ../RTL/cortexm0ds_logic.v(18933)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M4ebx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I74iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zg7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M4ebx6 ));  // ../RTL/cortexm0ds_logic.v(19987)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M5wax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fzkiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rdkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[26] ));  // ../RTL/cortexm0ds_logic.v(18934)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6cax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X44iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/He7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6cax6 ));  // ../RTL/cortexm0ds_logic.v(18254)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6kax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jrhow6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G81ju6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6kax6 ));  // ../RTL/cortexm0ds_logic.v(18692)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6rpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [0]),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F6eiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6rpw6 ));  // ../RTL/cortexm0ds_logic.v(17598)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M7wax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X1liu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rdkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[27] ));  // ../RTL/cortexm0ds_logic.v(18935)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M81qw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qcphu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M81qw6 ));  // ../RTL/cortexm0ds_logic.v(17936)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M85bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [30]),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z1fiu6 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M85bx6 ));  // ../RTL/cortexm0ds_logic.v(19707)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M8fax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Czuhu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/dbgrst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M8fax6 ));  // ../RTL/cortexm0ds_logic.v(18337)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M8ipw6_reg  (
    .clk(SWCLKTCK_pad),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W6ipw6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C53iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M8ipw6 ));  // ../RTL/cortexm0ds_logic.v(17188)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M9wax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P4liu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rdkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[29] ));  // ../RTL/cortexm0ds_logic.v(18936)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mb4bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fsdiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N2fiu6 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mb4bx6 ));  // ../RTL/cortexm0ds_logic.v(19611)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mbdax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H34iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Md7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mbdax6 ));  // ../RTL/cortexm0ds_logic.v(18281)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mboax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qcaiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kdkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[2] ));  // ../RTL/cortexm0ds_logic.v(18792)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mbwax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uoliu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rdkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[1] ));  // ../RTL/cortexm0ds_logic.v(18937)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mdppw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rkkiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ddkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[5] ));  // ../RTL/cortexm0ds_logic.v(17536)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mfyax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [7]),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X0fiu6 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mfyax6 ));  // ../RTL/cortexm0ds_logic.v(18999)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mgeax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K84iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mgeax6 ));  // ../RTL/cortexm0ds_logic.v(18313)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mh1qw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jcphu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mh1qw6 ));  // ../RTL/cortexm0ds_logic.v(17941)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Misax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qcaiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tekiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[2] ));  // ../RTL/cortexm0ds_logic.v(18868)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mjmpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X1liu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Afkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[27] ));  // ../RTL/cortexm0ds_logic.v(17429)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mk3bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A4phu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mk3bx6 ));  // ../RTL/cortexm0ds_logic.v(19533)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mlmpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X1liu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vfkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[27] ));  // ../RTL/cortexm0ds_logic.v(17430)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mnmpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xmthu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mnmpw6 ));  // ../RTL/cortexm0ds_logic.v(17435)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mp0bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Stuhu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mp0bx6 ));  // ../RTL/cortexm0ds_logic.v(19239)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ms5bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iiliu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n1465 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ms5bx6 ));  // ../RTL/cortexm0ds_logic.v(19727)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Muhbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O4phu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Muhbx6 ));  // ../RTL/cortexm0ds_logic.v(20144)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mw5bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jdohu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[10] ));  // ../RTL/cortexm0ds_logic.v(19734)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mz1bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jsuhu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mz1bx6 ));  // ../RTL/cortexm0ds_logic.v(19371)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N0cbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N7phu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N0cbx6 ));  // ../RTL/cortexm0ds_logic.v(19942)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N0lax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tx8iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lf8iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[0] ));  // ../RTL/cortexm0ds_logic.v(18712)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N0xpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bauhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N0xpw6 ));  // ../RTL/cortexm0ds_logic.v(17829)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N19bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q44iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N19bx6 ));  // ../RTL/cortexm0ds_logic.v(19807)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N1oax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rimiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mekiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[14] ));  // ../RTL/cortexm0ds_logic.v(18787)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N1wax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Drkiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rdkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[7] ));  // ../RTL/cortexm0ds_logic.v(18932)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N39ax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T24iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zg7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N39ax6 ));  // ../RTL/cortexm0ds_logic.v(18159)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N3eax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gk4iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Td7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N3eax6 ));  // ../RTL/cortexm0ds_logic.v(18301)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N3hbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W74iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Td7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N3hbx6 ));  // ../RTL/cortexm0ds_logic.v(20101)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N3jbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ym4iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zg7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N3jbx6 ));  // ../RTL/cortexm0ds_logic.v(20183)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N3oax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jlmiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mekiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[13] ));  // ../RTL/cortexm0ds_logic.v(18788)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N4gax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lm1iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qf7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N4gax6 ));  // ../RTL/cortexm0ds_logic.v(18400)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N4kax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Djthu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N4kax6 ));  // ../RTL/cortexm0ds_logic.v(18690)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5bbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V4phu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5bbx6 ));  // ../RTL/cortexm0ds_logic.v(19920)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5oax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bomiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mekiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[12] ));  // ../RTL/cortexm0ds_logic.v(18789)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N61qw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vpphu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N61qw6 ));  // ../RTL/cortexm0ds_logic.v(17935)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N7oax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hymiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mekiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[10] ));  // ../RTL/cortexm0ds_logic.v(18790)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N7ppw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K39iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ddkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[30] ));  // ../RTL/cortexm0ds_logic.v(17533)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N8rpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xeuhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N8rpw6 ));  // ../RTL/cortexm0ds_logic.v(17599)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N9oax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X6niu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mekiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[8] ));  // ../RTL/cortexm0ds_logic.v(18791)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N9ppw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D39iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ddkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[31] ));  // ../RTL/cortexm0ds_logic.v(17534)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Naaax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N64iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qf7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Naaax6 ));  // ../RTL/cortexm0ds_logic.v(18182)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nazax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [23]),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L1fiu6 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nazax6 ));  // ../RTL/cortexm0ds_logic.v(19089)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nbppw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jgkiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ddkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[3] ));  // ../RTL/cortexm0ds_logic.v(17535)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nbxax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wauhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nbxax6 ));  // ../RTL/cortexm0ds_logic.v(18960)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nckbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xcphu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nckbx6 ));  // ../RTL/cortexm0ds_logic.v(20246)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nd3qw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B7xhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nd3qw6 ));  // ../RTL/cortexm0ds_logic.v(18032)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nfgax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F94iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zg7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nfgax6 ));  // ../RTL/cortexm0ds_logic.v(18406)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nfnax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zvkiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mekiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[24] ));  // ../RTL/cortexm0ds_logic.v(18776)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nfqpw6_reg  (
    .clk(SWCLKTCK_pad),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F1yhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nfqpw6 ));  // ../RTL/cortexm0ds_logic.v(17555)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ngsax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X6niu6 ),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Stmiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[8] ));  // ../RTL/cortexm0ds_logic.v(18867)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nhgbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [22]),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L1fiu6 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nhgbx6 ));  // ../RTL/cortexm0ds_logic.v(20069)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nhnax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fzkiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mekiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[26] ));  // ../RTL/cortexm0ds_logic.v(18777)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ni5bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zvkiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pckiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[24] ));  // ../RTL/cortexm0ds_logic.v(19718)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nj2qw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E7vhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/dbgrst_reg ),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nj2qw6 ));  // ../RTL/cortexm0ds_logic.v(17995)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Njnax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X1liu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mekiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[27] ));  // ../RTL/cortexm0ds_logic.v(18778)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nk5bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fzkiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pckiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[26] ));  // ../RTL/cortexm0ds_logic.v(19719)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nlbbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G64iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qf7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nlbbx6 ));  // ../RTL/cortexm0ds_logic.v(19934)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nlcbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R84iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n382 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nlcbx6 ));  // ../RTL/cortexm0ds_logic.v(19953)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nlhax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Llohu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[12] ));  // ../RTL/cortexm0ds_logic.v(18513)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nlnax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P4liu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mekiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[29] ));  // ../RTL/cortexm0ds_logic.v(18779)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nm5bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X1liu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pckiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[27] ));  // ../RTL/cortexm0ds_logic.v(19720)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nmabx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L54iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qf7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nmabx6 ));  // ../RTL/cortexm0ds_logic.v(19891)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nmfax6_reg  (
    .clk(SWCLKTCK_pad),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qq3iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C53iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nmfax6 ));  // ../RTL/cortexm0ds_logic.v(18361)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nnfbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P74iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/He7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nnfbx6 ));  // ../RTL/cortexm0ds_logic.v(20015)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nnnax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hsliu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mekiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[25] ));  // ../RTL/cortexm0ds_logic.v(18780)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/No3qw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D84iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n382 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/No3qw6 ));  // ../RTL/cortexm0ds_logic.v(18044)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/No5bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P4liu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pckiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[29] ));  // ../RTL/cortexm0ds_logic.v(19721)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nodax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U64iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Td7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nodax6 ));  // ../RTL/cortexm0ds_logic.v(18293)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Npaax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oh4iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qf7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Npaax6 ));  // ../RTL/cortexm0ds_logic.v(18190)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Npnax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fyliu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mekiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[21] ));  // ../RTL/cortexm0ds_logic.v(18781)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Npypw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yjliu6 ),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fkliu6 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_control_o ));  // ../RTL/cortexm0ds_logic.v(17889)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nq5bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uoliu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pckiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[1] ));  // ../RTL/cortexm0ds_logic.v(19722)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nr0bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Guuhu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nr0bx6 ));  // ../RTL/cortexm0ds_logic.v(19245)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nr7ax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9uhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nr7ax6 ));  // ../RTL/cortexm0ds_logic.v(18109)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nrkpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I8phu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nrkpw6 ));  // ../RTL/cortexm0ds_logic.v(17309)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nrnax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E1miu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mekiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[20] ));  // ../RTL/cortexm0ds_logic.v(18782)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nrqpw6_reg  (
    .clk(SWCLKTCK_pad),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Golpw6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C53iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nrqpw6 ));  // ../RTL/cortexm0ds_logic.v(17576)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ns8ax6_reg  (
    .clk(SWCLKTCK_pad),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wq8ax6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C53iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ns8ax6 ));  // ../RTL/cortexm0ds_logic.v(18133)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nt9bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bouhu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nt9bx6 ));  // ../RTL/cortexm0ds_logic.v(19836)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ntnax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D4miu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mekiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[19] ));  // ../RTL/cortexm0ds_logic.v(18783)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nu5bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Irrhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nu5bx6 ));  // ../RTL/cortexm0ds_logic.v(19729)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nv3qw6_reg  (
    .clk(SWCLKTCK_pad),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wt3qw6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C53iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nv3qw6 ));  // ../RTL/cortexm0ds_logic.v(18048)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nv9bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [6]),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dv9iu6 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nv9bx6 ));  // ../RTL/cortexm0ds_logic.v(19842)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nvnax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C7miu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mekiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[18] ));  // ../RTL/cortexm0ds_logic.v(18784)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nwbbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Anrhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nwbbx6 ));  // ../RTL/cortexm0ds_logic.v(19940)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nwdbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B74iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n382 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nwdbx6 ));  // ../RTL/cortexm0ds_logic.v(19983)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxabx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ocohu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[21] ));  // ../RTL/cortexm0ds_logic.v(19901)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxnax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bamiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mekiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[17] ));  // ../RTL/cortexm0ds_logic.v(18785)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nybbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H1shu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nybbx6 ));  // ../RTL/cortexm0ds_logic.v(19941)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nyhax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ojohu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[1] ));  // ../RTL/cortexm0ds_logic.v(18555)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nyhpw6_reg  (
    .clk(SWCLKTCK_pad),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/cpu0cdbgpwrupreq ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kxhpw6 ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nyhpw6 ));  // ../RTL/cortexm0ds_logic.v(17172)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nznax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Admiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mekiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[16] ));  // ../RTL/cortexm0ds_logic.v(18786)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O0sax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C7miu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vfkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[18] ));  // ../RTL/cortexm0ds_logic.v(18859)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O1jbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K3niu6 ),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[7] ));  // ../RTL/cortexm0ds_logic.v(20182)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O1mpw6_reg  (
    .clk(SWCLKTCK_pad),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yzlpw6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C53iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O1mpw6 ));  // ../RTL/cortexm0ds_logic.v(17405)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O1ppw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jlmiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ofkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[13] ));  // ../RTL/cortexm0ds_logic.v(17530)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O2kax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nfohu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O2kax6 ));  // ../RTL/cortexm0ds_logic.v(18685)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O2sax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bamiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vfkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[17] ));  // ../RTL/cortexm0ds_logic.v(18860)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O3ppw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bomiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ofkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[12] ));  // ../RTL/cortexm0ds_logic.v(17531)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O41qw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X6niu6 ),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[6] ));  // ../RTL/cortexm0ds_logic.v(17934)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O4hax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wnohu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[24] ));  // ../RTL/cortexm0ds_logic.v(18459)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O4sax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Admiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vfkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[16] ));  // ../RTL/cortexm0ds_logic.v(18861)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O5ppw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ef8iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ddkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[4] ));  // ../RTL/cortexm0ds_logic.v(17532)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O6sax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rimiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vfkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[14] ));  // ../RTL/cortexm0ds_logic.v(18862)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O8sax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jlmiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vfkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[13] ));  // ../RTL/cortexm0ds_logic.v(18863)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oa5bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [31]),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z1fiu6 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oa5bx6 ));  // ../RTL/cortexm0ds_logic.v(19713)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oarpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qeuhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oarpw6 ));  // ../RTL/cortexm0ds_logic.v(17600)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oasax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bomiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vfkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[12] ));  // ../RTL/cortexm0ds_logic.v(18864)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ocsax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hymiu6 ),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Stmiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[10] ));  // ../RTL/cortexm0ds_logic.v(18865)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Od4bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [23]),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N2fiu6 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Od4bx6 ));  // ../RTL/cortexm0ds_logic.v(19617)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Odnax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Drkiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mekiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[7] ));  // ../RTL/cortexm0ds_logic.v(18775)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oesax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K3niu6 ),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Stmiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[9] ));  // ../RTL/cortexm0ds_logic.v(18866)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ofmpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [11]),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F6eiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ofmpw6 ));  // ../RTL/cortexm0ds_logic.v(17422)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Og5bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Drkiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pckiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[7] ));  // ../RTL/cortexm0ds_logic.v(19717)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oh8ax6_reg  (
    .clk(SWCLKTCK_pad),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Exxhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oh8ax6 ));  // ../RTL/cortexm0ds_logic.v(18122)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ohyax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [14]),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X0fiu6 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ohyax6 ));  // ../RTL/cortexm0ds_logic.v(19005)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oi9ax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E54iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zg7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oi9ax6 ));  // ../RTL/cortexm0ds_logic.v(18167)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oikax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jfthu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oikax6 ));  // ../RTL/cortexm0ds_logic.v(18703)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ojebx6_reg  (
    .clk(SWCLKTCK_pad),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bcdbx6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C53iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ojebx6 ));  // ../RTL/cortexm0ds_logic.v(19995)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ok2bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ppthu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ok2bx6 ));  // ../RTL/cortexm0ds_logic.v(19431)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Okfax6_reg  (
    .clk(SWCLKTCK_pad),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ne3iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W13iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Okfax6 ));  // ../RTL/cortexm0ds_logic.v(18360)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Om3bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vsthu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Om3bx6 ));  // ../RTL/cortexm0ds_logic.v(19539)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Onypw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uoliu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mekiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[1] ));  // ../RTL/cortexm0ds_logic.v(17884)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Opbax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ud4iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/He7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Opbax6 ));  // ../RTL/cortexm0ds_logic.v(18245)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Osrax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hsliu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vfkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[25] ));  // ../RTL/cortexm0ds_logic.v(18855)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ot0bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wvuhu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ot0bx6 ));  // ../RTL/cortexm0ds_logic.v(19251)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Otopw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X1liu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ofkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[27] ));  // ../RTL/cortexm0ds_logic.v(17526)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oulpw6_reg  (
    .clk(SWCLKTCK_pad),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L5lpw6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W13iu6 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kxhpw6 ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oulpw6 ));  // ../RTL/cortexm0ds_logic.v(17390)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ourax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fyliu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vfkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[21] ));  // ../RTL/cortexm0ds_logic.v(18856)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oveax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J44iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oveax6 ));  // ../RTL/cortexm0ds_logic.v(18321)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ovopw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P4liu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ofkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[29] ));  // ../RTL/cortexm0ds_logic.v(17527)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Owcax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z54iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Md7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Owcax6 ));  // ../RTL/cortexm0ds_logic.v(18273)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Owhbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zmuhu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Owhbx6 ));  // ../RTL/cortexm0ds_logic.v(20150)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Owrax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E1miu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vfkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[20] ));  // ../RTL/cortexm0ds_logic.v(18857)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ox9bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [6]),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F6eiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ox9bx6 ));  // ../RTL/cortexm0ds_logic.v(19844)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oxkpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dwuhu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oxkpw6 ));  // ../RTL/cortexm0ds_logic.v(17316)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oxopw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fyliu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ofkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[21] ));  // ../RTL/cortexm0ds_logic.v(17528)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oyhbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [3]),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F6eiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oyhbx6 ));  // ../RTL/cortexm0ds_logic.v(20152)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oykax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tx8iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ddkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[0] ));  // ../RTL/cortexm0ds_logic.v(18711)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oyrax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D4miu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vfkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[19] ));  // ../RTL/cortexm0ds_logic.v(18858)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ozopw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E1miu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ofkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[20] ));  // ../RTL/cortexm0ds_logic.v(17529)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ozvax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sokiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rdkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[6] ));  // ../RTL/cortexm0ds_logic.v(18931)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0bax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ud4iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xf7iu6 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/dbgrst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0bax6 ));  // ../RTL/cortexm0ds_logic.v(18205)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0ibx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ceuhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0ibx6 ));  // ../RTL/cortexm0ds_logic.v(20153)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V5vhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 ));  // ../RTL/cortexm0ds_logic.v(18683)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P12bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B1phu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P12bx6 ));  // ../RTL/cortexm0ds_logic.v(19377)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P14qw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wgvhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P14qw6 ));  // ../RTL/cortexm0ds_logic.v(18060)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P21qw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X6niu6 ),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qsmiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[8] ));  // ../RTL/cortexm0ds_logic.v(17933)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P23qw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D8xhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P23qw6 ));  // ../RTL/cortexm0ds_logic.v(18016)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P2xpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C7miu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lf8iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[18] ));  // ../RTL/cortexm0ds_logic.v(17830)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P33bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ezohu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P33bx6 ));  // ../RTL/cortexm0ds_logic.v(19485)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P34qw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vx9iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ofkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[23] ));  // ../RTL/cortexm0ds_logic.v(18062)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P4cax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E54iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/He7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P4cax6 ));  // ../RTL/cortexm0ds_logic.v(18253)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P4xpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C7miu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mx8iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[18] ));  // ../RTL/cortexm0ds_logic.v(17831)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P54qw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vx9iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Afkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[23] ));  // ../RTL/cortexm0ds_logic.v(18063)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oqohu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 ));  // ../RTL/cortexm0ds_logic.v(17759)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P6xpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C7miu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ofkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[18] ));  // ../RTL/cortexm0ds_logic.v(17832)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P7bbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hcohu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[9] ));  // ../RTL/cortexm0ds_logic.v(19926)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P8xpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C7miu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Afkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[18] ));  // ../RTL/cortexm0ds_logic.v(17833)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P93qw6_reg  (
    .clk(SWCLKTCK_pad),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z73qw6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C53iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P93qw6 ));  // ../RTL/cortexm0ds_logic.v(18025)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P9bax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Df4iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lg7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P9bax6 ));  // ../RTL/cortexm0ds_logic.v(18221)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Paxpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C7miu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ddkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[18] ));  // ../RTL/cortexm0ds_logic.v(17834)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pbbbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hvqhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pbbbx6 ));  // ../RTL/cortexm0ds_logic.v(19929)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pbnax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sokiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mekiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[6] ));  // ../RTL/cortexm0ds_logic.v(18774)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pcrpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S0vhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[1] ));  // ../RTL/cortexm0ds_logic.v(17605)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pcxpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C7miu6 ),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[16] ));  // ../RTL/cortexm0ds_logic.v(17835)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pczax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [30]),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L1fiu6 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pczax6 ));  // ../RTL/cortexm0ds_logic.v(19095)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pdbbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Faphu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pdbbx6 ));  // ../RTL/cortexm0ds_logic.v(19930)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pdmpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jgkiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vfkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[3] ));  // ../RTL/cortexm0ds_logic.v(17421)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pdxax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [14]),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F6eiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pdxax6 ));  // ../RTL/cortexm0ds_logic.v(18961)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pdyax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Npghu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pdyax6 ));  // ../RTL/cortexm0ds_logic.v(18993)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pe5bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sokiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pckiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[6] ));  // ../RTL/cortexm0ds_logic.v(19716)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pe7ax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M2xhu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/dbgrst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pe7ax6 ));  // ../RTL/cortexm0ds_logic.v(18096)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pe9bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xi4iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qf7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pe9bx6 ));  // ../RTL/cortexm0ds_logic.v(19814)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Peeax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T94iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Peeax6 ));  // ../RTL/cortexm0ds_logic.v(18312)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pejbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gfniu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n1552 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[26] ));  // ../RTL/cortexm0ds_logic.v(20189)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pexpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Khvhu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/dbgrst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pexpw6 ));  // ../RTL/cortexm0ds_logic.v(17840)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pg3qw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W7xhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pg3qw6 ));  // ../RTL/cortexm0ds_logic.v(18034)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Phcax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Df4iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/He7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Phcax6 ));  // ../RTL/cortexm0ds_logic.v(18260)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pifax6_reg  (
    .clk(SWCLKTCK_pad),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T33iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W13iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pifax6 ));  // ../RTL/cortexm0ds_logic.v(18359)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pjgbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [22]),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z1fiu6 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pjgbx6 ));  // ../RTL/cortexm0ds_logic.v(20075)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pkkbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T24iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lg7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pkkbx6 ));  // ../RTL/cortexm0ds_logic.v(20255)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Plypw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uoliu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ddkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[1] ));  // ../RTL/cortexm0ds_logic.v(17883)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pmlpw6_reg  (
    .clk(SWCLKTCK_pad),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zehpw6 [5]),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kxhpw6 ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pmlpw6 ));  // ../RTL/cortexm0ds_logic.v(17380)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pqrax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uoliu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vfkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[1] ));  // ../RTL/cortexm0ds_logic.v(18854)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Propw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rkkiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ofkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[5] ));  // ../RTL/cortexm0ds_logic.v(17525)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pt7ax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ybuhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pt7ax6 ));  // ../RTL/cortexm0ds_logic.v(18110)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Puwpw6_reg  (
    .clk(SWCLKTCK_pad),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nyxhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Puwpw6 ));  // ../RTL/cortexm0ds_logic.v(17826)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pv0bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kwuhu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pv0bx6 ));  // ../RTL/cortexm0ds_logic.v(19257)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pv9ax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Df4iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zg7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pv9ax6 ));  // ../RTL/cortexm0ds_logic.v(18174)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pwkax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tx8iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Afkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[0] ));  // ../RTL/cortexm0ds_logic.v(18710)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pxvax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rkkiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rdkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[5] ));  // ../RTL/cortexm0ds_logic.v(18930)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pz9bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [6]),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzeiu6 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pz9bx6 ));  // ../RTL/cortexm0ds_logic.v(19849)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pzibx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K3niu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n1552 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[7] ));  // ../RTL/cortexm0ds_logic.v(20181)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pzkpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gn8iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nn8iu6 ),
    .reset(1'b0),
    .set(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_tbit_o ));  // ../RTL/cortexm0ds_logic.v(17322)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q01qw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X6niu6 ),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Etmiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[8] ));  // ../RTL/cortexm0ds_logic.v(17932)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q1hbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W74iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q1hbx6 ));  // ../RTL/cortexm0ds_logic.v(20100)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q2gax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lm1iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zg7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q2gax6 ));  // ../RTL/cortexm0ds_logic.v(18399)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q2ibx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K84iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n382 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q2ibx6 ));  // ../RTL/cortexm0ds_logic.v(20154)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q4dbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y84iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n382 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q4dbx6 ));  // ../RTL/cortexm0ds_logic.v(19968)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q6fax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T24iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae7iu6 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/dbgrst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q6fax6 ));  // ../RTL/cortexm0ds_logic.v(18331)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q89bx6_reg  (
    .clk(SWCLKTCK_pad),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgfax6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C53iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q89bx6 ));  // ../RTL/cortexm0ds_logic.v(19811)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q8aax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U64iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qf7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q8aax6 ));  // ../RTL/cortexm0ds_logic.v(18181)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q9dax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oh4iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Md7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q9dax6 ));  // ../RTL/cortexm0ds_logic.v(18280)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q9nax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rkkiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mekiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[5] ));  // ../RTL/cortexm0ds_logic.v(18773)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qa1qw6_reg  (
    .clk(SWCLKTCK_pad),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vvxhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qa1qw6 ));  // ../RTL/cortexm0ds_logic.v(17937)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qaipw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sgthu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qaipw6 ));  // ../RTL/cortexm0ds_logic.v(17193)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qakbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rqthu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qakbx6 ));  // ../RTL/cortexm0ds_logic.v(20244)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbmpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jgkiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Afkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[3] ));  // ../RTL/cortexm0ds_logic.v(17420)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qc5bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Loshu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qc5bx6 ));  // ../RTL/cortexm0ds_logic.v(19715)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qehbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y8xhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qehbx6 ));  // ../RTL/cortexm0ds_logic.v(20107)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qf4bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [30]),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N2fiu6 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qf4bx6 ));  // ../RTL/cortexm0ds_logic.v(19623)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qhmpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mrthu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[3] ));  // ../RTL/cortexm0ds_logic.v(17427)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qijpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sf8iu6 ),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zf8iu6 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_apsr_o[1] ));  // ../RTL/cortexm0ds_logic.v(17245)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qirax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vx9iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vfkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[23] ));  // ../RTL/cortexm0ds_logic.v(18850)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qj1qw6_reg  (
    .clk(SWCLKTCK_pad),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cwxhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qj1qw6 ));  // ../RTL/cortexm0ds_logic.v(17942)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qjbbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G64iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zg7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qjbbx6 ));  // ../RTL/cortexm0ds_logic.v(19933)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qjcbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R84iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Md7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qjcbx6 ));  // ../RTL/cortexm0ds_logic.v(19952)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qjhax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Slohu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[13] ));  // ../RTL/cortexm0ds_logic.v(18507)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qjyax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fsdiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X0fiu6 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qjyax6 ));  // ../RTL/cortexm0ds_logic.v(19011)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qjypw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uoliu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Afkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[1] ));  // ../RTL/cortexm0ds_logic.v(17882)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qkabx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L54iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zg7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qkabx6 ));  // ../RTL/cortexm0ds_logic.v(19890)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qkrax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K39iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vfkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[30] ));  // ../RTL/cortexm0ds_logic.v(18851)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qlfbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P74iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qf7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qlfbx6 ));  // ../RTL/cortexm0ds_logic.v(20014)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qlopw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K39iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ofkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[30] ));  // ../RTL/cortexm0ds_logic.v(17522)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qmdax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D84iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Td7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qmdax6 ));  // ../RTL/cortexm0ds_logic.v(18292)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qmrax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D39iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vfkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[31] ));  // ../RTL/cortexm0ds_logic.v(18852)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qnopw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D39iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ofkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[31] ));  // ../RTL/cortexm0ds_logic.v(17523)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qo3bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M3phu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qo3bx6 ));  // ../RTL/cortexm0ds_logic.v(19545)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qorax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tx8iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vfkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[0] ));  // ../RTL/cortexm0ds_logic.v(18853)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qpopw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jgkiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ofkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[3] ));  // ../RTL/cortexm0ds_logic.v(17524)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qsfax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxqpw6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n265 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/dbgrst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qsfax6 ));  // ../RTL/cortexm0ds_logic.v(18378)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qudbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B74iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Md7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qudbx6 ));  // ../RTL/cortexm0ds_logic.v(19982)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qufax6_reg  (
    .clk(SWCLKTCK_pad),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qsfax6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kxhpw6 ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qufax6 ));  // ../RTL/cortexm0ds_logic.v(18384)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qukax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tx8iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ofkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[0] ));  // ../RTL/cortexm0ds_logic.v(18709)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qvvax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jgkiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rdkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[3] ));  // ../RTL/cortexm0ds_logic.v(18929)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qwfax6_reg  (
    .clk(SWCLKTCK_pad),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qufax6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kxhpw6 ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qwfax6 ));  // ../RTL/cortexm0ds_logic.v(18390)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qwfbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W8phu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qwfbx6 ));  // ../RTL/cortexm0ds_logic.v(20020)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qx0bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ywuhu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qx0bx6 ));  // ../RTL/cortexm0ds_logic.v(19263)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qxibx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K3niu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mekiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[9] ));  // ../RTL/cortexm0ds_logic.v(20180)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qyjax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufohu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qyjax6 ));  // ../RTL/cortexm0ds_logic.v(18678)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qynpw6_reg  (
    .clk(SWCLKTCK_pad),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I13iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W13iu6 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kxhpw6 ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P13iu6 ));  // ../RTL/cortexm0ds_logic.v(17484)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R19ax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O34iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bs4iu6 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/dbgrst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R19ax6 ));  // ../RTL/cortexm0ds_logic.v(18157)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R1abx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [6]),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J0fiu6 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R1abx6 ));  // ../RTL/cortexm0ds_logic.v(19855)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R1eax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pl4iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Td7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R1eax6 ));  // ../RTL/cortexm0ds_logic.v(18300)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R2hax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Doohu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[25] ));  // ../RTL/cortexm0ds_logic.v(18453)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vqohu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 ));  // ../RTL/cortexm0ds_logic.v(17753)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R7ibx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gfniu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ickiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[28] ));  // ../RTL/cortexm0ds_logic.v(20167)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R7kpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [13]),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F6eiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R7kpw6 ));  // ../RTL/cortexm0ds_logic.v(17289)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R7nax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jgkiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mekiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[3] ));  // ../RTL/cortexm0ds_logic.v(18772)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R9ibx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gfniu6 ),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztmiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[28] ));  // ../RTL/cortexm0ds_logic.v(20168)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R9mpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S5biu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F58iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R9mpw6 ));  // ../RTL/cortexm0ds_logic.v(17419)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R9yax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mbvhu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R9yax6 ));  // ../RTL/cortexm0ds_logic.v(18981)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ra2qw6_reg  (
    .clk(SWCLKTCK_pad),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C72qw6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C53iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ra2qw6 ));  // ../RTL/cortexm0ds_logic.v(17971)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rbibx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gfniu6 ),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Stmiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[28] ));  // ../RTL/cortexm0ds_logic.v(20169)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rdibx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gfniu6 ),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ltmiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[28] ));  // ../RTL/cortexm0ds_logic.v(20170)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rdkpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fyliu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Afkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[21] ));  // ../RTL/cortexm0ds_logic.v(17297)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rekbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yaohu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/SYSRESETREQ ));  // ../RTL/cortexm0ds_logic.v(20251)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rezax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [31]),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L1fiu6 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rezax6 ));  // ../RTL/cortexm0ds_logic.v(19101)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rfibx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gfniu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hfkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[28] ));  // ../RTL/cortexm0ds_logic.v(20171)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rfkpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fyliu6 ),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[19] ));  // ../RTL/cortexm0ds_logic.v(17298)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rfxax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dbuhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rfxax6 ));  // ../RTL/cortexm0ds_logic.v(18962)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rg9ax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S54iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zg7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rg9ax6 ));  // ../RTL/cortexm0ds_logic.v(18166)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rgrax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ef8iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vfkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[4] ));  // ../RTL/cortexm0ds_logic.v(18849)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rhibx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gfniu6 ),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xsmiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[28] ));  // ../RTL/cortexm0ds_logic.v(20172)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rhkpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [21]),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F6eiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rhkpw6 ));  // ../RTL/cortexm0ds_logic.v(17299)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rhypw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uoliu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ofkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[1] ));  // ../RTL/cortexm0ds_logic.v(17881)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rijbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uwdpw6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rijbx6 ));  // ../RTL/cortexm0ds_logic.v(20200)
  EG_PHY_PAD #(
    //.CLKSRC("CLK"),
    //.LOCATION("A7"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IDDRPIPEMODE("NONE"),
    .INCEMUX("INV"),
    .INPCLKMUX("CLK"),
    .INRSTMUX("INV"),
    .IN_DFFMODE("FF"),
    .IN_REGSET("SET"),
    .IOTYPE("LVCMOS25"),
    .MODE("BI"),
    .SRMODE("ASYNC"),
    .TSMUX("INV"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rilpw6_reg_IN  (
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tw2iu6 ),
    .do({open_n845,open_n846,open_n847,\u_cmsdk_mcu/dbg_swdo }),
    .ipclk(SWCLKTCK_pad),
    .rst(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kxhpw6 ),
    .ts(\u_cmsdk_mcu/dbg_swdo_en ),
    .diq({open_n853,open_n854,open_n855,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rilpw6 }),
    .bpad(SWDIOTMS));  // ../RTL/cmsdk_mcu.v(167)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rjibx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gfniu6 ),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qsmiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[28] ));  // ../RTL/cortexm0ds_logic.v(20173)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rjopw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ef8iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ofkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[4] ));  // ../RTL/cortexm0ds_logic.v(17521)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rk1bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K2phu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rk1bx6 ));  // ../RTL/cortexm0ds_logic.v(19329)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rkbax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ifphu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/dbgrst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rkbax6 ));  // ../RTL/cortexm0ds_logic.v(18231)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rkkax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cfthu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rkkax6 ));  // ../RTL/cortexm0ds_logic.v(18704)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rlgbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [22]),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N2fiu6 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rlgbx6 ));  // ../RTL/cortexm0ds_logic.v(20081)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rlibx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gfniu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kdkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[28] ));  // ../RTL/cortexm0ds_logic.v(20174)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rm2bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gwdpw6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rm2bx6 ));  // ../RTL/cortexm0ds_logic.v(19437)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rnaax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gk4iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qf7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rnaax6 ));  // ../RTL/cortexm0ds_logic.v(18189)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rnibx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gfniu6 ),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jsmiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[28] ));  // ../RTL/cortexm0ds_logic.v(20175)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rnvax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vx9iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rdkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[23] ));  // ../RTL/cortexm0ds_logic.v(18925)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ro8ax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Obphu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ro8ax6 ));  // ../RTL/cortexm0ds_logic.v(18131)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rpibx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gfniu6 ),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Csmiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[28] ));  // ../RTL/cortexm0ds_logic.v(20176)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rpvax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K39iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rdkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[30] ));  // ../RTL/cortexm0ds_logic.v(18926)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rq0qw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [8]),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F6eiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rq0qw6 ));  // ../RTL/cortexm0ds_logic.v(17927)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rr3qw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z6phu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rr3qw6 ));  // ../RTL/cortexm0ds_logic.v(18046)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rribx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gfniu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mekiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[28] ));  // ../RTL/cortexm0ds_logic.v(20177)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rrvax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D39iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rdkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[31] ));  // ../RTL/cortexm0ds_logic.v(18927)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rskax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Agjiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F58iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rskax6 ));  // ../RTL/cortexm0ds_logic.v(18708)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rteax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X44iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rteax6 ));  // ../RTL/cortexm0ds_logic.v(18320)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rtibx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gfniu6 ),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[26] ));  // ../RTL/cortexm0ds_logic.v(20178)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rtvax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tx8iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rdkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[0] ));  // ../RTL/cortexm0ds_logic.v(18928)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rucax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N64iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Md7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rucax6 ));  // ../RTL/cortexm0ds_logic.v(18272)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rv7ax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hduhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rv7ax6 ));  // ../RTL/cortexm0ds_logic.v(18111)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rvibx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K3niu6 ),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Csmiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[9] ));  // ../RTL/cortexm0ds_logic.v(20179)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rwhax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vjohu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[2] ));  // ../RTL/cortexm0ds_logic.v(18549)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rwjax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jzuhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rwjax6 ));  // ../RTL/cortexm0ds_logic.v(18676)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ry0qw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X6niu6 ),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ltmiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[8] ));  // ../RTL/cortexm0ds_logic.v(17931)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ry2qw6_reg  (
    .clk(SWCLKTCK_pad),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J3yhu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kxhpw6 ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ry2qw6 ));  // ../RTL/cortexm0ds_logic.v(18013)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ryfax6_reg  (
    .clk(SWCLKTCK_pad),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rtxhu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kxhpw6 ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ryfax6 ));  // ../RTL/cortexm0ds_logic.v(18396)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rz0bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ayuhu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rz0bx6 ));  // ../RTL/cortexm0ds_logic.v(19269)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rz8bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q44iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/He7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rz8bx6 ));  // ../RTL/cortexm0ds_logic.v(19806)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S0kbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Acvhu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S0kbx6 ));  // ../RTL/cortexm0ds_logic.v(20219)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S11bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mivhu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S11bx6 ));  // ../RTL/cortexm0ds_logic.v(19275)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S18ax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rimiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ofkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[14] ));  // ../RTL/cortexm0ds_logic.v(18114)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S1nax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K39iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mekiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[30] ));  // ../RTL/cortexm0ds_logic.v(18769)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S2cax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S54iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/He7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S2cax6 ));  // ../RTL/cortexm0ds_logic.v(18252)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S2cbx6_reg  (
    .clk(SWCLKTCK_pad),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y0yhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S2cbx6 ));  // ../RTL/cortexm0ds_logic.v(19943)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S32bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xsuhu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S32bx6 ));  // ../RTL/cortexm0ds_logic.v(19383)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S38ax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rimiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Afkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[14] ));  // ../RTL/cortexm0ds_logic.v(18115)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S3mpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [7]),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B3fiu6 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S3mpw6 ));  // ../RTL/cortexm0ds_logic.v(17410)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S3nax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D39iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mekiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[31] ));  // ../RTL/cortexm0ds_logic.v(18770)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S4kbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ay8iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n1465 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S4kbx6 ));  // ../RTL/cortexm0ds_logic.v(20231)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S53bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kqthu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S53bx6 ));  // ../RTL/cortexm0ds_logic.v(19491)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S58ax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rimiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ddkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[14] ));  // ../RTL/cortexm0ds_logic.v(18116)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S5kpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rkkiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vfkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[5] ));  // ../RTL/cortexm0ds_logic.v(17288)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S5nax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tx8iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mekiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[0] ));  // ../RTL/cortexm0ds_logic.v(18771)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S78ax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rimiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n1552 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[12] ));  // ../RTL/cortexm0ds_logic.v(18117)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S7mpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nhthu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S7mpw6 ));  // ../RTL/cortexm0ds_logic.v(17417)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S7yax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rkkiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pckiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[5] ));  // ../RTL/cortexm0ds_logic.v(18976)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S98ax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rimiu6 ),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[12] ));  // ../RTL/cortexm0ds_logic.v(18118)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sb8ax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ohqhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sb8ax6 ));  // ../RTL/cortexm0ds_logic.v(18119)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sbfax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D84iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rc7iu6 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/dbgrst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sbfax6 ));  // ../RTL/cortexm0ds_logic.v(18349)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sd8ax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Abphu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sd8ax6 ));  // ../RTL/cortexm0ds_logic.v(18120)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sddbx6_reg  (
    .clk(SWCLKTCK_pad),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Izxhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sddbx6 ));  // ../RTL/cortexm0ds_logic.v(19973)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sdlpw6_reg  (
    .clk(SWCLKTCK_pad),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zehpw6 [1]),
    .en(1'b1),
    .reset(1'b0),
    .set(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kxhpw6 ),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sdlpw6 ));  // ../RTL/cortexm0ds_logic.v(17350)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sejax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Khohu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sejax6 ));  // ../RTL/cortexm0ds_logic.v(18648)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Serax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qcaiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vfkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[2] ));  // ../RTL/cortexm0ds_logic.v(18848)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sfypw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uoliu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mx8iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[1] ));  // ../RTL/cortexm0ds_logic.v(17880)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sgjax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dhohu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sgjax6 ));  // ../RTL/cortexm0ds_logic.v(18649)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sh4bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [31]),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N2fiu6 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sh4bx6 ));  // ../RTL/cortexm0ds_logic.v(19629)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Shopw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zp6ow6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G81ju6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Shopw6 ));  // ../RTL/cortexm0ds_logic.v(17520)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sijax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wgohu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sijax6 ));  // ../RTL/cortexm0ds_logic.v(18650)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Skjax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E0vhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Skjax6 ));  // ../RTL/cortexm0ds_logic.v(18655)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Slvax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ef8iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rdkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[4] ));  // ../RTL/cortexm0ds_logic.v(18924)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Slyax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [23]),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X0fiu6 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Slyax6 ));  // ../RTL/cortexm0ds_logic.v(19017)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Smjax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pgohu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Smjax6 ));  // ../RTL/cortexm0ds_logic.v(18657)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sn4bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [7]),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzeiu6 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sn4bx6 ));  // ../RTL/cortexm0ds_logic.v(19647)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/So0qw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X6niu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n1552 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[6] ));  // ../RTL/cortexm0ds_logic.v(17926)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xzuhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 ));  // ../RTL/cortexm0ds_logic.v(18662)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sq3bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Enthu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sq3bx6 ));  // ../RTL/cortexm0ds_logic.v(19551)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sqfax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pkhpw6 [0]),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/dbgrst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sqfax6 ));  // ../RTL/cortexm0ds_logic.v(18372)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sqjax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Igohu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sqjax6 ));  // ../RTL/cortexm0ds_logic.v(18664)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sqkax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y48iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F58iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sqkax6 ));  // ../RTL/cortexm0ds_logic.v(18707)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sqwpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O3xhu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/dbgrst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sqwpw6 ));  // ../RTL/cortexm0ds_logic.v(17823)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ss0qw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tcuhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ss0qw6 ));  // ../RTL/cortexm0ds_logic.v(17928)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qzuhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6 ));  // ../RTL/cortexm0ds_logic.v(18669)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Stkpw6_reg  (
    .clk(SWCLKTCK_pad),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D0yhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Stkpw6 ));  // ../RTL/cortexm0ds_logic.v(17310)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Su8ax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X44iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n382 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Su8ax6 ));  // ../RTL/cortexm0ds_logic.v(18134)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sujax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bgohu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sujax6 ));  // ../RTL/cortexm0ds_logic.v(18671)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sw0qw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X6niu6 ),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gumiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[8] ));  // ../RTL/cortexm0ds_logic.v(17930)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Swjbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rw8iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qqhiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Swjbx6 ));  // ../RTL/cortexm0ds_logic.v(20213)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sx3qw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufvhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sx3qw6 ));  // ../RTL/cortexm0ds_logic.v(18049)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sx7ax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rimiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lf8iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[14] ));  // ../RTL/cortexm0ds_logic.v(18112)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Syjbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wzqhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Syjbx6 ));  // ../RTL/cortexm0ds_logic.v(20214)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sz3qw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I7cow6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n3436 ),
    .reset(1'b0),
    .set(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sz3qw6 ));  // ../RTL/cortexm0ds_logic.v(18054)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sz7ax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rimiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mx8iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[14] ));  // ../RTL/cortexm0ds_logic.v(18113)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Szmax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vx9iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mekiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[23] ));  // ../RTL/cortexm0ds_logic.v(18768)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T00qw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X1liu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n1552 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[25] ));  // ../RTL/cortexm0ds_logic.v(17914)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T0ipw6_reg  (
    .clk(SWCLKTCK_pad),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nyhpw6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kxhpw6 ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T0ipw6 ));  // ../RTL/cortexm0ds_logic.v(17178)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1fbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zuliu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Afkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[22] ));  // ../RTL/cortexm0ds_logic.v(20004)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Crohu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 ));  // ../RTL/cortexm0ds_logic.v(17747)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T20qw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P4liu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n1552 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[27] ));  // ../RTL/cortexm0ds_logic.v(17915)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T2dbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y84iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Md7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T2dbx6 ));  // ../RTL/cortexm0ds_logic.v(19967)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T2kbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kjthu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T2kbx6 ));  // ../RTL/cortexm0ds_logic.v(20225)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T3abx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [6]),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X0fiu6 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T3abx6 ));  // ../RTL/cortexm0ds_logic.v(19861)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T3fbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zuliu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wckiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[22] ));  // ../RTL/cortexm0ds_logic.v(20005)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T3kpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rkkiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Afkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[5] ));  // ../RTL/cortexm0ds_logic.v(17287)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T3opw6_reg  (
    .clk(SWCLKTCK_pad),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D2opw6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C53iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T3opw6 ));  // ../RTL/cortexm0ds_logic.v(17493)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T40qw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hsliu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n1552 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[23] ));  // ../RTL/cortexm0ds_logic.v(17916)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T5fbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zuliu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ddkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[22] ));  // ../RTL/cortexm0ds_logic.v(20006)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T5mpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z0vhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T5mpw6 ));  // ../RTL/cortexm0ds_logic.v(17412)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T5yax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Htshu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T5yax6 ));  // ../RTL/cortexm0ds_logic.v(18975)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T60qw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fyliu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n1552 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[19] ));  // ../RTL/cortexm0ds_logic.v(17917)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T6aax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D84iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qf7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T6aax6 ));  // ../RTL/cortexm0ds_logic.v(18180)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T6kbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L4rhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T6kbx6 ));  // ../RTL/cortexm0ds_logic.v(20233)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T7bax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ud4iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lg7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T7bax6 ));  // ../RTL/cortexm0ds_logic.v(18220)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T7fbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zuliu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kdkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[22] ));  // ../RTL/cortexm0ds_logic.v(20007)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T80qw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E1miu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n1552 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[18] ));  // ../RTL/cortexm0ds_logic.v(17918)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T82qw6_reg  (
    .clk(SWCLKTCK_pad),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C72qw6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jq3iu6 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kxhpw6 ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T82qw6 ));  // ../RTL/cortexm0ds_logic.v(17969)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T8kbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G8vhu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T8kbx6 ));  // ../RTL/cortexm0ds_logic.v(20238)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T9fbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zuliu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rdkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[22] ));  // ../RTL/cortexm0ds_logic.v(20008)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T9kpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kbuhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T9kpw6 ));  // ../RTL/cortexm0ds_logic.v(17290)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ta0qw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D4miu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n1552 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[17] ));  // ../RTL/cortexm0ds_logic.v(17919)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tajax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wz4iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qqhiu6 ),
    .reset(1'b0),
    .set(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tajax6 ));  // ../RTL/cortexm0ds_logic.v(18645)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tb3qw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H34iu6 ),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M24iu6 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/dbgrst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tb3qw6 ));  // ../RTL/cortexm0ds_logic.v(18030)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tbfbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zuliu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tekiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[22] ));  // ../RTL/cortexm0ds_logic.v(20009)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tc0qw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C7miu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n1552 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[16] ));  // ../RTL/cortexm0ds_logic.v(17920)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tc9bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xi4iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zg7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tc9bx6 ));  // ../RTL/cortexm0ds_logic.v(19813)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tceax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ud4iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tceax6 ));  // ../RTL/cortexm0ds_logic.v(18311)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tchbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M94iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qf7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tchbx6 ));  // ../RTL/cortexm0ds_logic.v(20106)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tcipw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jyohu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tcipw6 ));  // ../RTL/cortexm0ds_logic.v(17199)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tcjax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rhohu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tcjax6 ));  // ../RTL/cortexm0ds_logic.v(18647)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tcjbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ym4iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Md7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tcjbx6 ));  // ../RTL/cortexm0ds_logic.v(20188)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tcrax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X6niu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ickiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[8] ));  // ../RTL/cortexm0ds_logic.v(18847)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tdfbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zuliu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mekiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[22] ));  // ../RTL/cortexm0ds_logic.v(20010)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tdypw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uoliu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lf8iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[1] ));  // ../RTL/cortexm0ds_logic.v(17879)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Te0qw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bamiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n1552 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[15] ));  // ../RTL/cortexm0ds_logic.v(17921)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tfcax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H34iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/He7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tfcax6 ));  // ../RTL/cortexm0ds_logic.v(18259)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tffbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zuliu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n1552 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[20] ));  // ../RTL/cortexm0ds_logic.v(20011)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tg0qw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Admiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n1552 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[14] ));  // ../RTL/cortexm0ds_logic.v(17922)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgkbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lashu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgkbx6 ));  // ../RTL/cortexm0ds_logic.v(20253)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgzax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [31]),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dv9iu6 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgzax6 ));  // ../RTL/cortexm0ds_logic.v(19107)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Thcbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R84iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Td7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Thcbx6 ));  // ../RTL/cortexm0ds_logic.v(19951)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Thfbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zuliu6 ),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[20] ));  // ../RTL/cortexm0ds_logic.v(20012)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Thhax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zlohu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[15] ));  // ../RTL/cortexm0ds_logic.v(18501)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Thiax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Frthu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/dbgrst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Thiax6 ));  // ../RTL/cortexm0ds_logic.v(18595)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Thxax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [7]),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F6eiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Thxax6 ));  // ../RTL/cortexm0ds_logic.v(18963)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ti0qw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jlmiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n1552 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[11] ));  // ../RTL/cortexm0ds_logic.v(17923)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tikbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T24iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cf7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tikbx6 ));  // ../RTL/cortexm0ds_logic.v(20254)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tjfbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P74iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zg7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tjfbx6 ));  // ../RTL/cortexm0ds_logic.v(20013)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tjkpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G9uhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tjkpw6 ));  // ../RTL/cortexm0ds_logic.v(17300)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tjvax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qcaiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rdkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[2] ));  // ../RTL/cortexm0ds_logic.v(18923)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tk0qw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bomiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n1552 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[10] ));  // ../RTL/cortexm0ds_logic.v(17924)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tkdax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K84iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Td7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tkdax6 ));  // ../RTL/cortexm0ds_logic.v(18291)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tkjbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dpuhu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tkjbx6 ));  // ../RTL/cortexm0ds_logic.v(20206)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tl4bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [30]),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mpgiu6 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tl4bx6 ));  // ../RTL/cortexm0ds_logic.v(19641)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tlebx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eirhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tlebx6 ));  // ../RTL/cortexm0ds_logic.v(19996)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tm0qw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hymiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n1552 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[8] ));  // ../RTL/cortexm0ds_logic.v(17925)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tmjbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [9]),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F6eiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tmjbx6 ));  // ../RTL/cortexm0ds_logic.v(20208)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tnebx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zuliu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lf8iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[22] ));  // ../RTL/cortexm0ds_logic.v(19997)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tngbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [22]),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B3fiu6 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tngbx6 ));  // ../RTL/cortexm0ds_logic.v(20087)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tokax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eeohu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tokax6 ));  // ../RTL/cortexm0ds_logic.v(18706)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tpebx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zuliu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mx8iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[22] ));  // ../RTL/cortexm0ds_logic.v(19998)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tptpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [10]),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F6eiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tptpw6 ));  // ../RTL/cortexm0ds_logic.v(17689)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Trebx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zuliu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ickiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[22] ));  // ../RTL/cortexm0ds_logic.v(19999)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tsdbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B74iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Td7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tsdbx6 ));  // ../RTL/cortexm0ds_logic.v(19981)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tt9ax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H34iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zg7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tt9ax6 ));  // ../RTL/cortexm0ds_logic.v(18173)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ttebx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zuliu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pckiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[22] ));  // ../RTL/cortexm0ds_logic.v(20000)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tu0qw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X6niu6 ),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Numiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[8] ));  // ../RTL/cortexm0ds_logic.v(17929)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tujbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mbohu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tujbx6 ));  // ../RTL/cortexm0ds_logic.v(20212)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tvebx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zuliu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vfkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[22] ));  // ../RTL/cortexm0ds_logic.v(20001)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Twzpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zvkiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n1552 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[22] ));  // ../RTL/cortexm0ds_logic.v(17912)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Txebx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zuliu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ofkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[22] ));  // ../RTL/cortexm0ds_logic.v(20002)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Txmax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ef8iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mekiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[4] ));  // ../RTL/cortexm0ds_logic.v(18767)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tyaax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T24iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xf7iu6 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/dbgrst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tyaax6 ));  // ../RTL/cortexm0ds_logic.v(18199)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tyipw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [12]),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F6eiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tyipw6 ));  // ../RTL/cortexm0ds_logic.v(17226)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tyzpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fzkiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n1552 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[24] ));  // ../RTL/cortexm0ds_logic.v(17913)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tzebx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zuliu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hfkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[22] ));  // ../RTL/cortexm0ds_logic.v(20003)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tzgbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W74iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/He7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tzgbx6 ));  // ../RTL/cortexm0ds_logic.v(20099)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U0hax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Koohu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[26] ));  // ../RTL/cortexm0ds_logic.v(18447)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U0rax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Admiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ickiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[16] ));  // ../RTL/cortexm0ds_logic.v(18841)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U1kpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y7jiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F58iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U1kpw6 ));  // ../RTL/cortexm0ds_logic.v(17286)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U2rax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rimiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ickiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[14] ));  // ../RTL/cortexm0ds_logic.v(18842)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U31bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J5phu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U31bx6 ));  // ../RTL/cortexm0ds_logic.v(19281)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U3yax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jgkiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pckiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[3] ));  // ../RTL/cortexm0ds_logic.v(18974)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U4fax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Df4iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U4fax6 ));  // ../RTL/cortexm0ds_logic.v(18326)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U4rax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jlmiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ickiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[13] ));  // ../RTL/cortexm0ds_logic.v(18843)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U6rax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bomiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ickiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[12] ));  // ../RTL/cortexm0ds_logic.v(18844)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U7dax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gk4iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Md7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U7dax6 ));  // ../RTL/cortexm0ds_logic.v(18279)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U8jax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W7cow6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U8jax6 ));  // ../RTL/cortexm0ds_logic.v(18639)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U8rax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hymiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ickiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[10] ));  // ../RTL/cortexm0ds_logic.v(18845)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9ypw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rhvhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9ypw6 ));  // ../RTL/cortexm0ds_logic.v(17876)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ua9bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wjshu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ua9bx6 ));  // ../RTL/cortexm0ds_logic.v(19812)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uarax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K3niu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ickiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[9] ));  // ../RTL/cortexm0ds_logic.v(18846)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ubypw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tpohu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ubypw6 ));  // ../RTL/cortexm0ds_logic.v(17878)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ue9ax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z54iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zg7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ue9ax6 ));  // ../RTL/cortexm0ds_logic.v(18165)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufbbx6_reg  (
    .clk(SWCLKTCK_pad),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gyxhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufbbx6 ));  // ../RTL/cortexm0ds_logic.v(19931)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufebx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I74iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n382 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufebx6 ));  // ../RTL/cortexm0ds_logic.v(19993)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Utohu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 ));  // ../RTL/cortexm0ds_logic.v(17518)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uh2qw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ghthu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/dbgrst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uh2qw6 ));  // ../RTL/cortexm0ds_logic.v(17989)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uhvax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X6niu6 ),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xsmiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[8] ));  // ../RTL/cortexm0ds_logic.v(18922)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uizax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [30]),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dv9iu6 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uizax6 ));  // ../RTL/cortexm0ds_logic.v(19113)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uj4bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [31]),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mpgiu6 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uj4bx6 ));  // ../RTL/cortexm0ds_logic.v(19635)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ujspw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [16]),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F6eiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ujspw6 ));  // ../RTL/cortexm0ds_logic.v(17658)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ujxax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aduhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ujxax6 ));  // ../RTL/cortexm0ds_logic.v(18964)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Umkax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Leohu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Umkax6 ));  // ../RTL/cortexm0ds_logic.v(18705)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Untpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qcaiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mx8iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[2] ));  // ../RTL/cortexm0ds_logic.v(17688)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Unyax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [30]),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X0fiu6 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Unyax6 ));  // ../RTL/cortexm0ds_logic.v(19023)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uo2bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pvuhu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uo2bx6 ));  // ../RTL/cortexm0ds_logic.v(19443)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uofax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pkhpw6 [1]),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/dbgrst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uofax6 ));  // ../RTL/cortexm0ds_logic.v(18366)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uoipw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K39iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Afkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[30] ));  // ../RTL/cortexm0ds_logic.v(17216)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uojbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mcuhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uojbx6 ));  // ../RTL/cortexm0ds_logic.v(20209)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uoqax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hsliu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ickiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[25] ));  // ../RTL/cortexm0ds_logic.v(18835)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Up4bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [14]),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzeiu6 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Up4bx6 ));  // ../RTL/cortexm0ds_logic.v(19653)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uqipw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gfniu6 ),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Etmiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[28] ));  // ../RTL/cortexm0ds_logic.v(17217)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uqqax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fyliu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ickiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[21] ));  // ../RTL/cortexm0ds_logic.v(18836)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ureax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E54iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ureax6 ));  // ../RTL/cortexm0ds_logic.v(18319)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Urgbx6_reg  (
    .clk(SWCLKTCK_pad),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kadbx6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C53iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Urgbx6 ));  // ../RTL/cortexm0ds_logic.v(20095)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Us3bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bxdpw6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Us3bx6 ));  // ../RTL/cortexm0ds_logic.v(19557)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uscax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U64iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Md7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uscax6 ));  // ../RTL/cortexm0ds_logic.v(18271)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Usipw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fxuhu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Usipw6 ));  // ../RTL/cortexm0ds_logic.v(17222)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Usjbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tbohu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Usjbx6 ));  // ../RTL/cortexm0ds_logic.v(20211)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Usnpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dgphu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Usnpw6 ));  // ../RTL/cortexm0ds_logic.v(17477)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Usqax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E1miu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ickiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[20] ));  // ../RTL/cortexm0ds_logic.v(18837)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Utqpw6_reg  (
    .clk(SWCLKTCK_pad),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fuxhu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kxhpw6 ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Utqpw6 ));  // ../RTL/cortexm0ds_logic.v(17581)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uunpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H2yhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uunpw6 ));  // ../RTL/cortexm0ds_logic.v(17478)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uuqax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D4miu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ickiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[19] ));  // ../RTL/cortexm0ds_logic.v(18838)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uuzpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Drkiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n1552 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[5] ));  // ../RTL/cortexm0ds_logic.v(17911)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uvmax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qcaiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mekiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[2] ));  // ../RTL/cortexm0ds_logic.v(18766)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uwipw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ef8iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lf8iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[4] ));  // ../RTL/cortexm0ds_logic.v(17225)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uwqax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C7miu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ickiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[18] ));  // ../RTL/cortexm0ds_logic.v(18839)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ux8bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q44iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qf7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ux8bx6 ));  // ../RTL/cortexm0ds_logic.v(19805)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uyqax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bamiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ickiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[17] ));  // ../RTL/cortexm0ds_logic.v(18840)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V0cax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z54iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/He7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V0cax6 ));  // ../RTL/cortexm0ds_logic.v(18251)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V0jpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rbuhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V0jpw6 ));  // ../RTL/cortexm0ds_logic.v(17227)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V1vax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C7miu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wckiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[18] ));  // ../RTL/cortexm0ds_logic.v(18914)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V1yax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tx8iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pckiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[0] ));  // ../RTL/cortexm0ds_logic.v(18973)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V3vax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bamiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wckiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[17] ));  // ../RTL/cortexm0ds_logic.v(18915)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V52bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U0phu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V52bx6 ));  // ../RTL/cortexm0ds_logic.v(19389)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V53qw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sdphu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V53qw6 ));  // ../RTL/cortexm0ds_logic.v(18023)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V5abx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [6]),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L1fiu6 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V5abx6 ));  // ../RTL/cortexm0ds_logic.v(19867)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V5vax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Admiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wckiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[16] ));  // ../RTL/cortexm0ds_logic.v(18916)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V6jax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Miohu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V6jax6 ));  // ../RTL/cortexm0ds_logic.v(18634)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V73bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xyohu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V73bx6 ));  // ../RTL/cortexm0ds_logic.v(19497)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V7vax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rimiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wckiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[14] ));  // ../RTL/cortexm0ds_logic.v(18917)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V9vax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jlmiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wckiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[13] ));  // ../RTL/cortexm0ds_logic.v(18918)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Va7ax6_reg  (
    .clk(SWCLKTCK_pad),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E97ax6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C53iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Va7ax6 ));  // ../RTL/cortexm0ds_logic.v(18090)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vbkpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C6vhu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[5] ));  // ../RTL/cortexm0ds_logic.v(17295)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vbspw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [14]),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B3fiu6 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vbspw6 ));  // ../RTL/cortexm0ds_logic.v(17648)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vbvax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bomiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wckiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[12] ));  // ../RTL/cortexm0ds_logic.v(18919)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vdvax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hymiu6 ),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xsmiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[10] ));  // ../RTL/cortexm0ds_logic.v(18920)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vefax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Edphu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vefax6 ));  // ../RTL/cortexm0ds_logic.v(18357)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Veqax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zvkiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ickiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[24] ));  // ../RTL/cortexm0ds_logic.v(18830)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vfvax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K3niu6 ),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xsmiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[9] ));  // ../RTL/cortexm0ds_logic.v(18921)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vgjpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oxohu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vgjpw6 ));  // ../RTL/cortexm0ds_logic.v(17240)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vgqax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fzkiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ickiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[26] ));  // ../RTL/cortexm0ds_logic.v(18831)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vhspw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jn7ow6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O25iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vhspw6 ));  // ../RTL/cortexm0ds_logic.v(17657)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vibax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H34iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cf7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vibax6 ));  // ../RTL/cortexm0ds_logic.v(18226)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Viqax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X1liu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ickiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[27] ));  // ../RTL/cortexm0ds_logic.v(18832)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vj3qw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R8xhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vj3qw6 ));  // ../RTL/cortexm0ds_logic.v(18041)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vkqax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P4liu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ickiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[29] ));  // ../RTL/cortexm0ds_logic.v(18833)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vkzax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [23]),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dv9iu6 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vkzax6 ));  // ../RTL/cortexm0ds_logic.v(19119)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vlaax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pl4iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qf7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vlaax6 ));  // ../RTL/cortexm0ds_logic.v(18188)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vlkpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jlmiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Afkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[13] ));  // ../RTL/cortexm0ds_logic.v(17301)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vltpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qcaiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lf8iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[2] ));  // ../RTL/cortexm0ds_logic.v(17687)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vlxax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G3eiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F6eiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vlxax6 ));  // ../RTL/cortexm0ds_logic.v(18965)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vmipw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Flyiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O25iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vmipw6 ));  // ../RTL/cortexm0ds_logic.v(17215)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vmqax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uoliu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ickiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[1] ));  // ../RTL/cortexm0ds_logic.v(18834)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vn9bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I7xhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vn9bx6 ));  // ../RTL/cortexm0ds_logic.v(19819)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vnkpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jlmiu6 ),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[11] ));  // ../RTL/cortexm0ds_logic.v(17302)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vpgbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [22]),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aqgiu6 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vpgbx6 ));  // ../RTL/cortexm0ds_logic.v(20093)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vpkpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bfphu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/dbgrst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vpkpw6 ));  // ../RTL/cortexm0ds_logic.v(17307)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vplpw6_reg  (
    .clk(SWCLKTCK_pad),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Golpw6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U03iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vplpw6 ));  // ../RTL/cortexm0ds_logic.v(17383)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vqgax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F94iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n382 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vqgax6 ));  // ../RTL/cortexm0ds_logic.v(18412)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vqjbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Acohu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vqjbx6 ));  // ../RTL/cortexm0ds_logic.v(20210)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vrtpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fcuhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vrtpw6 ));  // ../RTL/cortexm0ds_logic.v(17690)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vszpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sokiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n1552 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[4] ));  // ../RTL/cortexm0ds_logic.v(17910)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vtmax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X6niu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hfkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[8] ));  // ../RTL/cortexm0ds_logic.v(18765)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vtuax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hsliu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wckiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[25] ));  // ../RTL/cortexm0ds_logic.v(18910)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vuhax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ckohu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[3] ));  // ../RTL/cortexm0ds_logic.v(18543)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vuipw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ef8iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Afkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[4] ));  // ../RTL/cortexm0ds_logic.v(17224)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vvuax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fyliu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wckiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[21] ));  // ../RTL/cortexm0ds_logic.v(18911)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vvxax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vx9iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pckiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[23] ));  // ../RTL/cortexm0ds_logic.v(18970)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vxuax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E1miu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wckiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[20] ));  // ../RTL/cortexm0ds_logic.v(18912)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vxxax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K39iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pckiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[30] ));  // ../RTL/cortexm0ds_logic.v(18971)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vyfbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uuuhu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vyfbx6 ));  // ../RTL/cortexm0ds_logic.v(20025)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vygax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U8vhu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vygax6 ));  // ../RTL/cortexm0ds_logic.v(18441)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vz8ax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ud4iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bs4iu6 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/dbgrst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vz8ax6 ));  // ../RTL/cortexm0ds_logic.v(18151)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzdax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J44iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Td7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzdax6 ));  // ../RTL/cortexm0ds_logic.v(18299)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzjpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fivhu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzjpw6 ));  // ../RTL/cortexm0ds_logic.v(17284)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzuax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D4miu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wckiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[19] ));  // ../RTL/cortexm0ds_logic.v(18913)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jrohu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ));  // ../RTL/cortexm0ds_logic.v(17741)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzxax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D39iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pckiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[31] ));  // ../RTL/cortexm0ds_logic.v(18972)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W0dbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y84iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Td7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W0dbx6 ));  // ../RTL/cortexm0ds_logic.v(19966)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W0jax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T4vhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W0jax6 ));  // ../RTL/cortexm0ds_logic.v(18626)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W2jax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A5vhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W2jax6 ));  // ../RTL/cortexm0ds_logic.v(18627)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4aax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K84iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qf7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4aax6 ));  // ../RTL/cortexm0ds_logic.v(18179)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4jax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Withu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4jax6 ));  // ../RTL/cortexm0ds_logic.v(18632)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W51bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gothu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W51bx6 ));  // ../RTL/cortexm0ds_logic.v(19287)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W5max6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hsliu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hfkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[25] ));  // ../RTL/cortexm0ds_logic.v(18753)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W5ypw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yavhu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W5ypw6 ));  // ../RTL/cortexm0ds_logic.v(17864)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W6ipw6_reg  (
    .clk(SWCLKTCK_pad),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Grxhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W6ipw6 ));  // ../RTL/cortexm0ds_logic.v(17187)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W7max6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fyliu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hfkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[21] ));  // ../RTL/cortexm0ds_logic.v(18754)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W8hbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yhvhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W8hbx6 ));  // ../RTL/cortexm0ds_logic.v(20104)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W9max6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E1miu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hfkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[20] ));  // ../RTL/cortexm0ds_logic.v(18755)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W9spw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sokiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vfkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[6] ));  // ../RTL/cortexm0ds_logic.v(17643)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wahbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M94iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zg7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wahbx6 ));  // ../RTL/cortexm0ds_logic.v(20105)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wbmax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D4miu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hfkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[19] ));  // ../RTL/cortexm0ds_logic.v(18756)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wc2qw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T94iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n382 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wc2qw6 ));  // ../RTL/cortexm0ds_logic.v(17972)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wcqax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Drkiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ickiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[7] ));  // ../RTL/cortexm0ds_logic.v(18829)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wdmax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C7miu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hfkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[18] ));  // ../RTL/cortexm0ds_logic.v(18757)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Weipw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K39iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mx8iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[30] ));  // ../RTL/cortexm0ds_logic.v(17201)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wfcbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R84iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wfcbx6 ));  // ../RTL/cortexm0ds_logic.v(19950)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wfhax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gmohu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[16] ));  // ../RTL/cortexm0ds_logic.v(18495)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wfmax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bamiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hfkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[17] ));  // ../RTL/cortexm0ds_logic.v(18758)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wfspw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S7vhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wfspw6 ));  // ../RTL/cortexm0ds_logic.v(17655)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wgipw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [30]),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aqgiu6 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wgipw6 ));  // ../RTL/cortexm0ds_logic.v(17206)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Whmax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Admiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hfkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[16] ));  // ../RTL/cortexm0ds_logic.v(18759)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Widax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T94iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Td7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Widax6 ));  // ../RTL/cortexm0ds_logic.v(18290)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wjmax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rimiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hfkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[14] ));  // ../RTL/cortexm0ds_logic.v(18760)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wjtpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qcaiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ddkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[2] ));  // ../RTL/cortexm0ds_logic.v(17686)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wjuax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zvkiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wckiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[24] ));  // ../RTL/cortexm0ds_logic.v(18905)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wkipw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bithu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wkipw6 ));  // ../RTL/cortexm0ds_logic.v(17213)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wlmax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jlmiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hfkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[13] ));  // ../RTL/cortexm0ds_logic.v(18761)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wlspw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pauhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wlspw6 ));  // ../RTL/cortexm0ds_logic.v(17659)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wluax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fzkiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wckiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[26] ));  // ../RTL/cortexm0ds_logic.v(18906)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wmzax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fsdiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dv9iu6 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wmzax6 ));  // ../RTL/cortexm0ds_logic.v(19125)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wnmax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bomiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hfkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[12] ));  // ../RTL/cortexm0ds_logic.v(18762)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wnuax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X1liu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wckiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[27] ));  // ../RTL/cortexm0ds_logic.v(18907)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wnxax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I4eiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F6eiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wnxax6 ));  // ../RTL/cortexm0ds_logic.v(18966)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wpmax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hymiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hfkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[10] ));  // ../RTL/cortexm0ds_logic.v(18763)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wpuax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P4liu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wckiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[29] ));  // ../RTL/cortexm0ds_logic.v(18908)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wpyax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [31]),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X0fiu6 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wpyax6 ));  // ../RTL/cortexm0ds_logic.v(19029)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wq8ax6_reg  (
    .clk(SWCLKTCK_pad),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xwxhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wq8ax6 ));  // ../RTL/cortexm0ds_logic.v(18132)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wqdbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B74iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wqdbx6 ));  // ../RTL/cortexm0ds_logic.v(19980)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wqzpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rkkiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n1552 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[3] ));  // ../RTL/cortexm0ds_logic.v(17909)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wr4bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fsdiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzeiu6 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wr4bx6 ));  // ../RTL/cortexm0ds_logic.v(19659)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wrmax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K3niu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hfkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[9] ));  // ../RTL/cortexm0ds_logic.v(18764)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wruax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uoliu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wckiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[1] ));  // ../RTL/cortexm0ds_logic.v(18909)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wt3qw6_reg  (
    .clk(SWCLKTCK_pad),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M1yhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wt3qw6 ));  // ../RTL/cortexm0ds_logic.v(18047)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wtxax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lgthu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wtxax6 ));  // ../RTL/cortexm0ds_logic.v(18969)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wu3bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [7]),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J0fiu6 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wu3bx6 ));  // ../RTL/cortexm0ds_logic.v(19563)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wvgax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xg6iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/dbgrst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wvgax6 ));  // ../RTL/cortexm0ds_logic.v(18429)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wwiax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F4vhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wwiax6 ));  // ../RTL/cortexm0ds_logic.v(18624)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wxgbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W74iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qf7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wxgbx6 ));  // ../RTL/cortexm0ds_logic.v(20098)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wxjpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z71ju6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G81ju6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wxjpw6 ));  // ../RTL/cortexm0ds_logic.v(17279)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wyiax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M4vhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wyiax6 ));  // ../RTL/cortexm0ds_logic.v(18625)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X1max6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P4liu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hfkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[29] ));  // ../RTL/cortexm0ds_logic.v(18751)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X1upw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fzkiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ddkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[26] ));  // ../RTL/cortexm0ds_logic.v(17695)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X2jpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E1miu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Afkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[20] ));  // ../RTL/cortexm0ds_logic.v(17228)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X3max6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uoliu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hfkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[1] ));  // ../RTL/cortexm0ds_logic.v(18752)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X3upw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fzkiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vfkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[26] ));  // ../RTL/cortexm0ds_logic.v(17696)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X42qw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S6phu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X42qw6 ));  // ../RTL/cortexm0ds_logic.v(17963)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X4jpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E1miu6 ),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[18] ));  // ../RTL/cortexm0ds_logic.v(17229)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X5bax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O34iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lg7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X5bax6 ));  // ../RTL/cortexm0ds_logic.v(18219)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X5ibx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Glphu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_apsr_o[0] ));  // ../RTL/cortexm0ds_logic.v(20165)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X5opw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [5]),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F6eiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X5opw6 ));  // ../RTL/cortexm0ds_logic.v(17494)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X5upw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rwuhu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X5upw6 ));  // ../RTL/cortexm0ds_logic.v(17701)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X6jpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [20]),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F6eiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X6jpw6 ));  // ../RTL/cortexm0ds_logic.v(17230)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X7abx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [6]),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z1fiu6 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X7abx6 ));  // ../RTL/cortexm0ds_logic.v(19873)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X7spw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sokiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ddkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[6] ));  // ../RTL/cortexm0ds_logic.v(17642)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X7ypw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L0vhu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X7ypw6 ));  // ../RTL/cortexm0ds_logic.v(17870)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xaeax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T24iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Td7iu6 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/dbgrst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xaeax6 ));  // ../RTL/cortexm0ds_logic.v(18309)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xajbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ym4iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Td7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xajbx6 ));  // ../RTL/cortexm0ds_logic.v(20187)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xaqax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sokiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ickiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[6] ));  // ../RTL/cortexm0ds_logic.v(18828)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xbopw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n689 ),
    .en(1'b1),
    .reset(1'b0),
    .set(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/SLEEPHOLDACKn ));  // ../RTL/cortexm0ds_logic.v(17506)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xc9ax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N64iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zg7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xc9ax6 ));  // ../RTL/cortexm0ds_logic.v(18164)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xdcax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oh4iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/He7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xdcax6 ));  // ../RTL/cortexm0ds_logic.v(18258)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xdebx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I74iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Md7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xdebx6 ));  // ../RTL/cortexm0ds_logic.v(19992)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xdspw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O5vhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xdspw6 ));  // ../RTL/cortexm0ds_logic.v(17650)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xf8ax6_reg  (
    .clk(SWCLKTCK_pad),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lxxhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xf8ax6 ));  // ../RTL/cortexm0ds_logic.v(18121)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xfiax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oy8iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n590 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_primask_o ));  // ../RTL/cortexm0ds_logic.v(18589)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xhtpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qcaiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Afkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[2] ));  // ../RTL/cortexm0ds_logic.v(17685)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xhuax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Drkiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wckiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[7] ));  // ../RTL/cortexm0ds_logic.v(18904)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xiipw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U1vhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xiipw6 ));  // ../RTL/cortexm0ds_logic.v(17208)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xkqpw6_reg  (
    .clk(SWCLKTCK_pad),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cjqpw6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n267 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kxhpw6 ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/cpu0cdbgpwrupreq ));  // ../RTL/cortexm0ds_logic.v(17572)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xn7ax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K8xhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xn7ax6 ));  // ../RTL/cortexm0ds_logic.v(18102)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xnbax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X6vhu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/dbgrst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xnbax6 ));  // ../RTL/cortexm0ds_logic.v(18243)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xo1bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D2phu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xo1bx6 ));  // ../RTL/cortexm0ds_logic.v(19341)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xozax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [14]),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dv9iu6 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xozax6 ));  // ../RTL/cortexm0ds_logic.v(19131)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xozpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jgkiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n1552 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[1] ));  // ../RTL/cortexm0ds_logic.v(17908)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xpeax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S54iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xpeax6 ));  // ../RTL/cortexm0ds_logic.v(18318)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xpxax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zcqhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xpxax6 ));  // ../RTL/cortexm0ds_logic.v(18967)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xq2bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Szohu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xq2bx6 ));  // ../RTL/cortexm0ds_logic.v(19449)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xqcax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D84iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Md7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xqcax6 ));  // ../RTL/cortexm0ds_logic.v(18270)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xr9ax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oh4iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zg7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xr9ax6 ));  // ../RTL/cortexm0ds_logic.v(18172)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xrxax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Egthu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xrxax6 ));  // ../RTL/cortexm0ds_logic.v(18968)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xttpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fzkiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lf8iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[26] ));  // ../RTL/cortexm0ds_logic.v(17691)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xu2qw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zdphu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xu2qw6 ));  // ../RTL/cortexm0ds_logic.v(18007)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuiax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y3vhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuiax6 ));  // ../RTL/cortexm0ds_logic.v(18623)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xv8bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q44iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zg7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xv8bx6 ));  // ../RTL/cortexm0ds_logic.v(19804)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xvlax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zvkiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hfkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[24] ));  // ../RTL/cortexm0ds_logic.v(18748)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xvqpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Utqpw6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/dbgrst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xvqpw6 ));  // ../RTL/cortexm0ds_logic.v(17587)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xvtpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fzkiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mx8iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[26] ));  // ../RTL/cortexm0ds_logic.v(17692)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xwaax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O34iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qf7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xwaax6 ));  // ../RTL/cortexm0ds_logic.v(18194)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xx6bx6_reg  (
    .clk(SWCLKTCK_pad),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gw6bx6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C53iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xx6bx6 ));  // ../RTL/cortexm0ds_logic.v(19764)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxlax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fzkiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hfkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[26] ));  // ../RTL/cortexm0ds_logic.v(18749)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxqpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xvqpw6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/dbgrst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxqpw6 ));  // ../RTL/cortexm0ds_logic.v(17593)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxtpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fzkiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ofkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[26] ));  // ../RTL/cortexm0ds_logic.v(17693)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qrohu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 ));  // ../RTL/cortexm0ds_logic.v(17735)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xzlax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X1liu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hfkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[27] ));  // ../RTL/cortexm0ds_logic.v(18750)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xztpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fzkiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Afkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[26] ));  // ../RTL/cortexm0ds_logic.v(17694)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y0gbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zzohu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y0gbx6 ));  // ../RTL/cortexm0ds_logic.v(20031)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y2fax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H34iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y2fax6 ));  // ../RTL/cortexm0ds_logic.v(18325)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y5dax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pl4iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Md7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y5dax6 ));  // ../RTL/cortexm0ds_logic.v(18278)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y5spw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sokiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Afkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[6] ));  // ../RTL/cortexm0ds_logic.v(17641)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y72bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cmthu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y72bx6 ));  // ../RTL/cortexm0ds_logic.v(19395)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y7opw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oduhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y7opw6 ));  // ../RTL/cortexm0ds_logic.v(17495)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y7upw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bamiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lf8iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[17] ));  // ../RTL/cortexm0ds_logic.v(17703)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y8lpw6_reg  (
    .clk(SWCLKTCK_pad),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rfxhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y8lpw6 ));  // ../RTL/cortexm0ds_logic.v(17333)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y8qax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rkkiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ickiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[5] ));  // ../RTL/cortexm0ds_logic.v(18827)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y93bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J6vhu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y93bx6 ));  // ../RTL/cortexm0ds_logic.v(19503)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y9upw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bamiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mx8iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[17] ));  // ../RTL/cortexm0ds_logic.v(17704)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ybupw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bamiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ofkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[17] ));  // ../RTL/cortexm0ds_logic.v(17705)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydgax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lm1iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n382 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydgax6 ));  // ../RTL/cortexm0ds_logic.v(18405)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Buohu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 ));  // ../RTL/cortexm0ds_logic.v(17512)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydupw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bamiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Afkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[17] ));  // ../RTL/cortexm0ds_logic.v(17706)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yf1qw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N6xhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yf1qw6 ));  // ../RTL/cortexm0ds_logic.v(17940)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yftpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qcaiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ofkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[2] ));  // ../RTL/cortexm0ds_logic.v(17684)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yfuax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sokiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wckiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[6] ));  // ../RTL/cortexm0ds_logic.v(18903)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yfupw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bamiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ddkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[17] ));  // ../RTL/cortexm0ds_logic.v(17707)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yhupw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bamiu6 ),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[15] ));  // ../RTL/cortexm0ds_logic.v(17708)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yizpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D39iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n1552 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[29] ));  // ../RTL/cortexm0ds_logic.v(17905)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yjaax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J44iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qf7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yjaax6 ));  // ../RTL/cortexm0ds_logic.v(18187)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yjupw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [17]),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F6eiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yjupw6 ));  // ../RTL/cortexm0ds_logic.v(17709)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yklpw6_reg  (
    .clk(SWCLKTCK_pad),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zehpw6 [4]),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kxhpw6 ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yklpw6 ));  // ../RTL/cortexm0ds_logic.v(17374)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ykzpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K39iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n1552 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[28] ));  // ../RTL/cortexm0ds_logic.v(17906)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ym3qw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U64iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n382 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ym3qw6 ));  // ../RTL/cortexm0ds_logic.v(18043)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ymwpw6_reg  (
    .clk(SWCLKTCK_pad),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hlwpw6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C53iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ymwpw6 ));  // ../RTL/cortexm0ds_logic.v(17817)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ymzpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ef8iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n1552 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[2] ));  // ../RTL/cortexm0ds_logic.v(17907)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ynspw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zvkiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lf8iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[24] ));  // ../RTL/cortexm0ds_logic.v(17660)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yogax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F94iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Md7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yogax6 ));  // ../RTL/cortexm0ds_logic.v(18411)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ypspw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zvkiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mx8iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[24] ));  // ../RTL/cortexm0ds_logic.v(17661)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yqzax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [7]),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dv9iu6 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yqzax6 ));  // ../RTL/cortexm0ds_logic.v(19137)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yrspw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zvkiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ofkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[24] ));  // ../RTL/cortexm0ds_logic.v(17662)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yryax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fsdiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B3fiu6 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yryax6 ));  // ../RTL/cortexm0ds_logic.v(19035)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ysiax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ysiax6 ));  // ../RTL/cortexm0ds_logic.v(18622)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yt4bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [23]),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzeiu6 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yt4bx6 ));  // ../RTL/cortexm0ds_logic.v(19665)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yt8bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vrmiu6 ),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[9] ));  // ../RTL/cortexm0ds_logic.v(19803)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ytlax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Drkiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hfkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[7] ));  // ../RTL/cortexm0ds_logic.v(18747)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ytspw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zvkiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Afkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[24] ));  // ../RTL/cortexm0ds_logic.v(17663)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yubbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G64iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n382 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yubbx6 ));  // ../RTL/cortexm0ds_logic.v(19939)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvabx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L54iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n382 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvabx6 ));  // ../RTL/cortexm0ds_logic.v(19896)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Twohu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 ));  // ../RTL/cortexm0ds_logic.v(17277)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvspw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zvkiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ddkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[24] ));  // ../RTL/cortexm0ds_logic.v(17664)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yw3bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [14]),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J0fiu6 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yw3bx6 ));  // ../RTL/cortexm0ds_logic.v(19569)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yxdax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X44iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Td7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yxdax6 ));  // ../RTL/cortexm0ds_logic.v(18298)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yxrpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W1phu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yxrpw6 ));  // ../RTL/cortexm0ds_logic.v(17636)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yxspw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zvkiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vfkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[24] ));  // ../RTL/cortexm0ds_logic.v(17665)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yybax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N64iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/He7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yybax6 ));  // ../RTL/cortexm0ds_logic.v(18250)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yzlpw6_reg  (
    .clk(SWCLKTCK_pad),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C3yhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yzlpw6 ));  // ../RTL/cortexm0ds_logic.v(17404)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yzqpw6_reg  (
    .clk(SWCLKTCK_pad),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zwnpw6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C53iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yzqpw6 ));  // ../RTL/cortexm0ds_logic.v(17595)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yzspw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tivhu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yzspw6 ));  // ../RTL/cortexm0ds_logic.v(17670)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z18bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zfmiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ofkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[15] ));  // ../RTL/cortexm0ds_logic.v(19789)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z1tpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hsliu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lf8iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[25] ));  // ../RTL/cortexm0ds_logic.v(17672)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z2aax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T94iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qf7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z2aax6 ));  // ../RTL/cortexm0ds_logic.v(18178)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z38bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zfmiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hfkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[15] ));  // ../RTL/cortexm0ds_logic.v(19790)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z3spw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sokiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ofkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[6] ));  // ../RTL/cortexm0ds_logic.v(17640)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z3tpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hsliu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mx8iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[25] ));  // ../RTL/cortexm0ds_logic.v(17673)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z47ax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dmqhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z47ax6 ));  // ../RTL/cortexm0ds_logic.v(18087)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z58bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zfmiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Afkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[15] ));  // ../RTL/cortexm0ds_logic.v(19791)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z5tpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hsliu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ofkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[25] ));  // ../RTL/cortexm0ds_logic.v(17674)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z67ax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Taphu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z67ax6 ));  // ../RTL/cortexm0ds_logic.v(18088)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z6qax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jgkiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ickiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[3] ));  // ../RTL/cortexm0ds_logic.v(18826)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z71bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R2phu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z71bx6 ));  // ../RTL/cortexm0ds_logic.v(19293)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z73qw6_reg  (
    .clk(SWCLKTCK_pad),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Psxhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z73qw6 ));  // ../RTL/cortexm0ds_logic.v(18024)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z78bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zfmiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wckiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[15] ));  // ../RTL/cortexm0ds_logic.v(19792)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z7tpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hsliu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Afkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[25] ));  // ../RTL/cortexm0ds_logic.v(17675)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z8jpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N9uhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z8jpw6 ));  // ../RTL/cortexm0ds_logic.v(17231)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z8zpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zvkiu6 ),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[22] ));  // ../RTL/cortexm0ds_logic.v(17900)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z98bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zfmiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ddkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[15] ));  // ../RTL/cortexm0ds_logic.v(19793)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z9abx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [6]),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N2fiu6 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z9abx6 ));  // ../RTL/cortexm0ds_logic.v(19879)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z9opw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J4xhu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z9opw6 ));  // ../RTL/cortexm0ds_logic.v(17500)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z9tpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hsliu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ddkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[25] ));  // ../RTL/cortexm0ds_logic.v(17676)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zazpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fzkiu6 ),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[24] ));  // ../RTL/cortexm0ds_logic.v(17901)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zb8bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zfmiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kdkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[15] ));  // ../RTL/cortexm0ds_logic.v(19794)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zbtpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hsliu6 ),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[23] ));  // ../RTL/cortexm0ds_logic.v(17677)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zczpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X1liu6 ),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[25] ));  // ../RTL/cortexm0ds_logic.v(17902)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zd8bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zfmiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rdkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[15] ));  // ../RTL/cortexm0ds_logic.v(19795)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zdcbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R84iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/He7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zdcbx6 ));  // ../RTL/cortexm0ds_logic.v(19949)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zdhax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nmohu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[17] ));  // ../RTL/cortexm0ds_logic.v(18489)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zdiax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mihow6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zdiax6 ));  // ../RTL/cortexm0ds_logic.v(18583)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zdtpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qmthu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zdtpw6 ));  // ../RTL/cortexm0ds_logic.v(17682)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zduax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rkkiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wckiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[5] ));  // ../RTL/cortexm0ds_logic.v(18902)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zezpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P4liu6 ),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[27] ));  // ../RTL/cortexm0ds_logic.v(17903)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zf8bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zfmiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tekiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[15] ));  // ../RTL/cortexm0ds_logic.v(19796)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgbax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Df4iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cf7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgbax6 ));  // ../RTL/cortexm0ds_logic.v(18225)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgfax6_reg  (
    .clk(SWCLKTCK_pad),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dtxhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgfax6 ));  // ../RTL/cortexm0ds_logic.v(18358)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgzpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qcaiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n1552 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[0] ));  // ../RTL/cortexm0ds_logic.v(17904)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zh8bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zfmiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mekiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[15] ));  // ../RTL/cortexm0ds_logic.v(19797)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zj8bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zfmiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n1552 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[13] ));  // ../RTL/cortexm0ds_logic.v(19798)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zl8bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zfmiu6 ),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[13] ));  // ../RTL/cortexm0ds_logic.v(19799)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zl9bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xi4iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Md7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zl9bx6 ));  // ../RTL/cortexm0ds_logic.v(19818)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zm8ax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H3xhu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/dbgrst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zm8ax6 ));  // ../RTL/cortexm0ds_logic.v(18129)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zn8bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vrmiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tekiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[11] ));  // ../RTL/cortexm0ds_logic.v(19800)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zodbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B74iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/He7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zodbx6 ));  // ../RTL/cortexm0ds_logic.v(19979)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zp8bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vrmiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mekiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[11] ));  // ../RTL/cortexm0ds_logic.v(19801)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zqiax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K3vhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zqiax6 ));  // ../RTL/cortexm0ds_logic.v(18621)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zr7bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zfmiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lf8iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[15] ));  // ../RTL/cortexm0ds_logic.v(19784)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zr8bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vrmiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n1552 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[9] ));  // ../RTL/cortexm0ds_logic.v(19802)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zrlax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sokiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hfkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[6] ));  // ../RTL/cortexm0ds_logic.v(18746)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zshax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jkohu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[4] ));  // ../RTL/cortexm0ds_logic.v(18537)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zslpw6_reg  (
    .clk(SWCLKTCK_pad),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Krlpw6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U03iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zslpw6 ));  // ../RTL/cortexm0ds_logic.v(17385)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zszax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [0]),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R5eiu6 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zszax6 ));  // ../RTL/cortexm0ds_logic.v(19143)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zt7bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zfmiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mx8iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[15] ));  // ../RTL/cortexm0ds_logic.v(19785)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztgbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kavhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztgbx6 ));  // ../RTL/cortexm0ds_logic.v(20096)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztupw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fbvhu6 ),
    .en(1'b1),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztupw6 ));  // ../RTL/cortexm0ds_logic.v(17723)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zv7bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zfmiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ickiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[15] ));  // ../RTL/cortexm0ds_logic.v(19786)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zvgbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W74iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zg7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zvgbx6 ));  // ../RTL/cortexm0ds_logic.v(20097)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zvrpw6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Drkiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vfkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[7] ));  // ../RTL/cortexm0ds_logic.v(17631)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zwnpw6_reg  (
    .clk(SWCLKTCK_pad),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A2yhu6 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zwnpw6 ));  // ../RTL/cortexm0ds_logic.v(17479)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zx7bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zfmiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pckiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[15] ));  // ../RTL/cortexm0ds_logic.v(19787)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zx8ax6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T24iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bs4iu6 ),
    .reset(~\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/dbgrst_reg ),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zx8ax6 ));  // ../RTL/cortexm0ds_logic.v(18145)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zycbx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y84iu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae7iu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zycbx6 ));  // ../RTL/cortexm0ds_logic.v(19965)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zz7bx6_reg  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zfmiu6 ),
    .en(~\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vfkiu6 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[15] ));  // ../RTL/cortexm0ds_logic.v(19788)
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add0/u0  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qehbx6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E4yhu6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add0/c0 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add0/c1 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vrkbx6 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add0/u1  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vj3qw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ksgax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add0/c1 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add0/c2 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vrkbx6 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add0/u2  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xn7ax6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dugax6 ),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add0/c2 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add0/c3 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vrkbx6 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add0/u3  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P23qw6 ),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add0/c3 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add0/c4 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vrkbx6 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add0/u4  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pg3qw6 ),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add0/c4 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add0/c5 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vrkbx6 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add0/u5  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bf3qw6 ),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add0/c5 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add0/c6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vrkbx6 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add0/u6  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vn9bx6 ),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add0/c6 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add0/c7 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vrkbx6 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add0/u7  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nd3qw6 ),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add0/c7 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add0/c8 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vrkbx6 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add0/u8  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ke1qw6 ),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add0/c8 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add0/c9 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vrkbx6 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add0/u9  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yf1qw6 ),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add0/c9 ),
    .o({open_n857,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vrkbx6 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add0/ucin  (
    .a(1'b0),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add0/c0 ,open_n860}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/u0  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[0] ),
    .b(1'b1),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c0 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c1 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/u1  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[1] ),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c1 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c2 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/u10  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[10] ),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c10 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c11 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/u11  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[11] ),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c11 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c12 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/u12  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[12] ),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c12 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c13 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/u13  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[13] ),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c13 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c14 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/u14  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[14] ),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c14 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c15 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/u15  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[15] ),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c15 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c16 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/u16  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[16] ),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c16 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c17 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/u17  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[17] ),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c17 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c18 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/u18  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[18] ),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c18 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c19 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/u19  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[19] ),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c19 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c20 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/u2  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[2] ),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c2 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c3 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/u20  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[20] ),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c20 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c21 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/u21  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[21] ),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c21 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c22 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/u22  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[22] ),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c22 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c23 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/u23  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[23] ),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c23 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c24 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/u24  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[24] ),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c24 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c25 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/u25  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[25] ),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c25 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c26 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/u26  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[26] ),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c26 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c27 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/u27  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[27] ),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c27 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c28 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/u28  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[28] ),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c28 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c29 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/u29  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[29] ),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c29 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c30 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/u3  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[3] ),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c3 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c4 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/u30  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[30] ),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c30 ),
    .o({open_n861,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/u4  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[4] ),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c4 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c5 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/u5  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[5] ),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c5 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/u6  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[6] ),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c6 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c7 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/u7  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[7] ),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c7 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c8 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/u8  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[8] ),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c8 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c9 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/u9  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[9] ),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c9 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c10 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/ucin  (
    .a(1'b0),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c0 ,open_n864}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/u0  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R0ghu6 ),
    .b(1'b1),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c0 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c1 ,open_n865}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/u1  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[2] ),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c1 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c2 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/u10  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[11] ),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c10 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c11 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/u11  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[12] ),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c11 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c12 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/u12  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[13] ),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c12 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c13 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/u13  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[14] ),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c13 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c14 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/u14  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[15] ),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c14 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c15 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/u15  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[16] ),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c15 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c16 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/u16  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[17] ),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c16 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c17 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/u17  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[18] ),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c17 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c18 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/u18  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[19] ),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c18 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c19 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/u19  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[20] ),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c19 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c20 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/u2  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[3] ),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c2 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c3 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/u20  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[21] ),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c20 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c21 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/u21  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[22] ),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c21 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c22 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/u22  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[23] ),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c22 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c23 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/u23  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[24] ),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c23 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c24 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/u24  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[25] ),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c24 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c25 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/u25  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[26] ),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c25 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c26 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/u26  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[27] ),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c26 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c27 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/u27  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[28] ),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c27 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c28 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/u28  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[29] ),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c28 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c29 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/u29  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[30] ),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c29 ),
    .o({open_n866,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/u3  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[4] ),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c3 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c4 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/u4  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[5] ),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c4 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c5 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/u5  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[6] ),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c5 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/u6  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[7] ),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c6 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c7 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/u7  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[8] ),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c7 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c8 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/u8  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[9] ),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c8 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c9 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/u9  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[10] ),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c9 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c10 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/ucin  (
    .a(1'b0),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c0 ,open_n869}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/u0  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [0]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [0]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c0 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c1 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/u1  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [1]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [1]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c1 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c2 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/u10  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [10]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [10]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c10 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c11 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/u11  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C1epw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [11]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c11 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c12 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/u12  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J1epw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [12]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c12 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c13 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/u13  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q1epw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [13]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c13 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c14 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/u14  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X1epw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [14]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c14 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c15 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/u15  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L2epw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [15]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c15 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c16 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/u16  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z2epw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [16]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c16 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c17 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/u17  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G3epw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [17]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c17 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c18 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/u18  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N3epw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [18]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c18 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c19 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/u19  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U3epw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [19]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c19 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c20 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/u2  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [2]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [2]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c2 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c3 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/u20  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B4epw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [20]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c20 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c21 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/u21  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I4epw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [21]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c21 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c22 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/u22  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P4epw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [22]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c22 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c23 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/u23  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [23]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [23]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c23 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c24 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/u24  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [24]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [24]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c24 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c25 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/u25  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [25]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [25]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c25 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c26 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/u26  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [26]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [26]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c26 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c27 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/u27  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [27]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [27]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c27 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c28 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/u28  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [28]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [28]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c28 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c29 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/u29  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [29]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [29]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c29 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c30 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/u3  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [3]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [3]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c3 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c4 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/u30  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [30]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [30]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c30 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c31 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/u31  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D5epw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [31]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c31 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c32 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [32]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/u4  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [4]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [4]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c4 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c5 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/u5  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [5]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [5]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c5 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/u6  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E2epw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [6]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c6 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c7 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/u7  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S2epw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [7]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c7 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c8 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/u8  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4epw6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [8]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c8 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c9 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/u9  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q5phu6 ),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [9]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c9 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c10 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/ucin  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dqfhu6 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c0 ,open_n872}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/ucout  (
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c32 ),
    .o({open_n875,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [33]}));
  EG_PHY_MULT18 #(
    .INPUTREGA("DISABLE"),
    .INPUTREGB("DISABLE"),
    .MODE("MULT18X18C"),
    .OUTPUTREG("DISABLE"),
    .SIGNEDAMUX("0"),
    .SIGNEDBMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mifpw6 [17:0]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgfpw6 [17:0]),
    .p({open_n959,open_n960,open_n961,open_n962,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_31 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_30 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_29 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_28 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_27 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_26 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_25 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_24 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_23 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_22 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_21 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_20 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_19 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_18 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_17 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_16 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_15 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_14 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_13 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_12 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_11 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_10 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_9 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_8 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_7 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_5 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_4 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_3 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_2 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_1 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_0 }));
  EG_PHY_MULT18 #(
    .INPUTREGA("DISABLE"),
    .INPUTREGB("DISABLE"),
    .MODE("MULT18X18C"),
    .OUTPUTREG("DISABLE"),
    .SIGNEDAMUX("0"),
    .SIGNEDBMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_1_  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mifpw6 [17:0]),
    .b({4'b0000,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgfpw6 [31:18]}),
    .p({open_n1046,open_n1047,open_n1048,open_n1049,open_n1050,open_n1051,open_n1052,open_n1053,open_n1054,open_n1055,open_n1056,open_n1057,open_n1058,open_n1059,open_n1060,open_n1061,open_n1062,open_n1063,open_n1064,open_n1065,open_n1066,open_n1067,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_1_13 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_1_12 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_1_11 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_1_10 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_1_9 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_1_8 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_1_7 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_1_6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_1_5 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_1_4 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_1_3 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_1_2 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_1_1 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_1_0 }));
  EG_PHY_MULT18 #(
    .INPUTREGA("DISABLE"),
    .INPUTREGB("DISABLE"),
    .MODE("MULT18X18C"),
    .OUTPUTREG("DISABLE"),
    .SIGNEDAMUX("0"),
    .SIGNEDBMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_1_0_  (
    .a({4'b0000,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mifpw6 [31:18]}),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgfpw6 [17:0]),
    .p({open_n1151,open_n1152,open_n1153,open_n1154,open_n1155,open_n1156,open_n1157,open_n1158,open_n1159,open_n1160,open_n1161,open_n1162,open_n1163,open_n1164,open_n1165,open_n1166,open_n1167,open_n1168,open_n1169,open_n1170,open_n1171,open_n1172,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_1_0_13 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_1_0_12 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_1_0_11 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_1_0_10 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_1_0_9 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_1_0_8 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_1_0_7 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_1_0_6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_1_0_5 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_1_0_4 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_1_0_3 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_1_0_2 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_1_0_1 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_1_0_0 }));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/u0  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N8rpw6 ),
    .b(1'b1),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/c0 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/c1 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6gpw6 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/u1  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oarpw6 ),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/c1 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/c2 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6gpw6 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/u10  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vrtpw6 ),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/c10 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/c11 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6gpw6 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/u11  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pt7ax6 ),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/c11 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/c12 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6gpw6 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/u12  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V0jpw6 ),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/c12 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/c13 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6gpw6 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/u13  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T9kpw6 ),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/c13 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/c14 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6gpw6 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/u14  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rfxax6 ),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/c14 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/c15 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6gpw6 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/u15  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nbxax6 ),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/c15 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/c16 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6gpw6 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/u16  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wlspw6 ),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/c16 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/c17 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6gpw6 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/u17  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Amupw6 ),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/c17 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/c18 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6gpw6 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/u18  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N0xpw6 ),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/c18 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/c19 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6gpw6 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/u19  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nr7ax6 ),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/c19 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/c20 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6gpw6 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/u2  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kzabx6 ),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/c2 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/c3 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6gpw6 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/u20  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z8jpw6 ),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/c20 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/c21 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6gpw6 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/u21  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tjkpw6 ),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/c21 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/c22 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6gpw6 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/u22  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F9gbx6 ),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/c22 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/c23 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6gpw6 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/u23  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Coupw6 ),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/c23 ),
    .o({open_n1173,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6gpw6 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/u3  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0ibx6 ),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/c3 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/c4 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6gpw6 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/u4  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Johbx6 ),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/c4 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/c5 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6gpw6 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/u5  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y7opw6 ),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/c5 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/c6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6gpw6 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/u6  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rv7ax6 ),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/c6 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/c7 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6gpw6 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/u7  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ujxax6 ),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/c7 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/c8 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6gpw6 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/u8  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ss0qw6 ),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/c8 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/c9 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6gpw6 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/u9  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uojbx6 ),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/c9 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/c10 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6gpw6 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/ucin  (
    .a(1'b0),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/c0 ,open_n1176}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub1/u0  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X5phu6 ),
    .b(1'b1),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub1/c0 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub1/c1 ,open_n1177}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub1/u1  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vnfpw6 [0]),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub1/c1 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub1/c2 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xlfpw6 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub1/u2  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vnfpw6 [1]),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub1/c2 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub1/c3 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xlfpw6 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub1/u3  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vnfpw6 [2]),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub1/c3 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub1/c4 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xlfpw6 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub1/u4  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vnfpw6 [3]),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub1/c4 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub1/c5 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xlfpw6 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub1/u5  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vnfpw6 [4]),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub1/c5 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub1/c6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xlfpw6 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub1/u6  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vnfpw6 [5]),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub1/c6 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub1/c7 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xlfpw6 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub1/u7  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vnfpw6 [6]),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub1/c7 ),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub1/c8 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xlfpw6 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub1/u8  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vnfpw6 [7]),
    .b(1'b0),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub1/c8 ),
    .o({open_n1178,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xlfpw6 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub1/ucin  (
    .a(1'b0),
    .o({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub1/c0 ,open_n1181}));
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/reg0_b0  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HADDR [2]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/trans_valid ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/haddr_reg [0]));  // ../RTL/cmsdk_ahb_cs_rom_table.v(161)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/reg0_b1  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HADDR [3]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/trans_valid ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/haddr_reg [1]));  // ../RTL/cmsdk_ahb_cs_rom_table.v(161)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/reg0_b2  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HADDR [4]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/trans_valid ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/haddr_reg [2]));  // ../RTL/cmsdk_ahb_cs_rom_table.v(161)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/reg0_b3  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HADDR [5]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/trans_valid ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/haddr_reg [3]));  // ../RTL/cmsdk_ahb_cs_rom_table.v(161)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/reg0_b4  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HADDR [6]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/trans_valid ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/haddr_reg [4]));  // ../RTL/cmsdk_ahb_cs_rom_table.v(161)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/reg0_b5  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HADDR [7]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/trans_valid ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/haddr_reg [5]));  // ../RTL/cmsdk_ahb_cs_rom_table.v(161)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/reg0_b6  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HADDR [8]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/trans_valid ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/haddr_reg [6]));  // ../RTL/cmsdk_ahb_cs_rom_table.v(161)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/reg0_b7  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HADDR [9]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/trans_valid ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/haddr_reg [7]));  // ../RTL/cmsdk_ahb_cs_rom_table.v(161)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/reg0_b8  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HADDR [10]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/trans_valid ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/haddr_reg [8]));  // ../RTL/cmsdk_ahb_cs_rom_table.v(161)
  reg_ar_as_w1 \u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/reg0_b9  (
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HADDR [11]),
    .en(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/trans_valid ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/haddr_reg [9]));  // ../RTL/cmsdk_ahb_cs_rom_table.v(161)

endmodule 

module reg_ar_as_w1
  (
  clk,
  d,
  en,
  reset,
  set,
  q
  );

  input clk;
  input d;
  input en;
  input reset;
  input set;
  output q;

  parameter REGSET = "RESET";
  wire enout;

  AL_MUX u_en0 (
    .i0(q),
    .i1(d),
    .sel(en),
    .o(enout));
  AL_DFF #(
    .INI((REGSET == "SET") ? 1'b1 : 1'b0))
    u_seq0 (
    .clk(clk),
    .d(enout),
    .reset(reset),
    .set(set),
    .q(q));

endmodule 

module AL_MUX
  (
  input i0,
  input i1,
  input sel,
  output o
  );

  wire not_sel, sel_i0, sel_i1;
  not u0 (not_sel, sel);
  and u1 (sel_i1, sel, i1);
  and u2 (sel_i0, not_sel, i0);
  or u3 (o, sel_i1, sel_i0);

endmodule

module AL_DFF
  (
  input reset,
  input set,
  input clk,
  input d,
  output reg q
  );

  parameter INI = 1'b0;

  always @(posedge reset or posedge set or posedge clk)
  begin
    if (reset)
      q <= 1'b0;
    else if (set)
      q <= 1'b1;
    else
      q <= d;
  end

endmodule

