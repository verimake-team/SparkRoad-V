// Verilog netlist created by TD v4.6.12906
// Thu Aug  8 15:19:06 2019

`timescale 1ns / 1ps
module VGA_Demo  // source/rtl/VGA_Demo.v(2)
  (
  clk_24m,
  rst_n,
  vga_b,
  vga_clk,
  vga_de,
  vga_g,
  vga_hs,
  vga_r,
  vga_vs
  );

  input clk_24m;  // source/rtl/VGA_Demo.v(4)
  input rst_n;  // source/rtl/VGA_Demo.v(5)
  output [7:0] vga_b;  // source/rtl/VGA_Demo.v(16)
  output vga_clk;  // source/rtl/VGA_Demo.v(8)
  output vga_de;  // source/rtl/VGA_Demo.v(12)
  output [7:0] vga_g;  // source/rtl/VGA_Demo.v(15)
  output vga_hs;  // source/rtl/VGA_Demo.v(9)
  output [7:0] vga_r;  // source/rtl/VGA_Demo.v(14)
  output vga_vs;  // source/rtl/VGA_Demo.v(10)

  wire [23:0] lcd_data;  // source/rtl/VGA_Demo.v(22)
  wire [11:0] lcd_xpos;  // source/rtl/VGA_Demo.v(20)
  wire [11:0] lcd_ypos;  // source/rtl/VGA_Demo.v(21)
  wire [23:0] \u2_Display/n1 ;
  wire clk_vga;  // source/rtl/VGA_Demo.v(19)

  Clk_div u0_PLL (
    .clk(clk_24m),
    .rst_n(rst_n),
    .clk_div(clk_vga));  // source/rtl/VGA_Demo.v(25)
  Driver u1_Driver (
    .clk(clk_vga),
    .lcd_data(lcd_data),
    .rst_n(rst_n),
    .lcd_dclk(vga_clk),
    .lcd_en(vga_de),
    .lcd_hs(vga_hs),
    .lcd_rgb({vga_r,vga_g,vga_b}),
    .lcd_vs(vga_vs),
    .lcd_xpos(lcd_xpos),
    .lcd_ypos(lcd_ypos));  // source/rtl/VGA_Demo.v(34)
  mult_u12_u12_o24 \u2_Display/mult0  (
    .i0(lcd_xpos),
    .i1(lcd_ypos),
    .o(\u2_Display/n1 ));  // source/rtl/Display.v(93)
  reg_ar_as_w1 \u2_Display/reg0_b0  (
    .clk(clk_vga),
    .d(\u2_Display/n1 [0]),
    .en(1'b1),
    .reset(~rst_n),
    .set(1'b0),
    .q(lcd_data[0]));  // source/rtl/Display.v(93)
  reg_ar_as_w1 \u2_Display/reg0_b1  (
    .clk(clk_vga),
    .d(\u2_Display/n1 [1]),
    .en(1'b1),
    .reset(~rst_n),
    .set(1'b0),
    .q(lcd_data[1]));  // source/rtl/Display.v(93)
  reg_ar_as_w1 \u2_Display/reg0_b10  (
    .clk(clk_vga),
    .d(\u2_Display/n1 [10]),
    .en(1'b1),
    .reset(~rst_n),
    .set(1'b0),
    .q(lcd_data[10]));  // source/rtl/Display.v(93)
  reg_ar_as_w1 \u2_Display/reg0_b11  (
    .clk(clk_vga),
    .d(\u2_Display/n1 [11]),
    .en(1'b1),
    .reset(~rst_n),
    .set(1'b0),
    .q(lcd_data[11]));  // source/rtl/Display.v(93)
  reg_ar_as_w1 \u2_Display/reg0_b12  (
    .clk(clk_vga),
    .d(\u2_Display/n1 [12]),
    .en(1'b1),
    .reset(~rst_n),
    .set(1'b0),
    .q(lcd_data[12]));  // source/rtl/Display.v(93)
  reg_ar_as_w1 \u2_Display/reg0_b13  (
    .clk(clk_vga),
    .d(\u2_Display/n1 [13]),
    .en(1'b1),
    .reset(~rst_n),
    .set(1'b0),
    .q(lcd_data[13]));  // source/rtl/Display.v(93)
  reg_ar_as_w1 \u2_Display/reg0_b14  (
    .clk(clk_vga),
    .d(\u2_Display/n1 [14]),
    .en(1'b1),
    .reset(~rst_n),
    .set(1'b0),
    .q(lcd_data[14]));  // source/rtl/Display.v(93)
  reg_ar_as_w1 \u2_Display/reg0_b15  (
    .clk(clk_vga),
    .d(\u2_Display/n1 [15]),
    .en(1'b1),
    .reset(~rst_n),
    .set(1'b0),
    .q(lcd_data[15]));  // source/rtl/Display.v(93)
  reg_ar_as_w1 \u2_Display/reg0_b16  (
    .clk(clk_vga),
    .d(\u2_Display/n1 [16]),
    .en(1'b1),
    .reset(~rst_n),
    .set(1'b0),
    .q(lcd_data[16]));  // source/rtl/Display.v(93)
  reg_ar_as_w1 \u2_Display/reg0_b17  (
    .clk(clk_vga),
    .d(\u2_Display/n1 [17]),
    .en(1'b1),
    .reset(~rst_n),
    .set(1'b0),
    .q(lcd_data[17]));  // source/rtl/Display.v(93)
  reg_ar_as_w1 \u2_Display/reg0_b18  (
    .clk(clk_vga),
    .d(\u2_Display/n1 [18]),
    .en(1'b1),
    .reset(~rst_n),
    .set(1'b0),
    .q(lcd_data[18]));  // source/rtl/Display.v(93)
  reg_ar_as_w1 \u2_Display/reg0_b19  (
    .clk(clk_vga),
    .d(\u2_Display/n1 [19]),
    .en(1'b1),
    .reset(~rst_n),
    .set(1'b0),
    .q(lcd_data[19]));  // source/rtl/Display.v(93)
  reg_ar_as_w1 \u2_Display/reg0_b2  (
    .clk(clk_vga),
    .d(\u2_Display/n1 [2]),
    .en(1'b1),
    .reset(~rst_n),
    .set(1'b0),
    .q(lcd_data[2]));  // source/rtl/Display.v(93)
  reg_ar_as_w1 \u2_Display/reg0_b20  (
    .clk(clk_vga),
    .d(\u2_Display/n1 [20]),
    .en(1'b1),
    .reset(~rst_n),
    .set(1'b0),
    .q(lcd_data[20]));  // source/rtl/Display.v(93)
  reg_ar_as_w1 \u2_Display/reg0_b21  (
    .clk(clk_vga),
    .d(\u2_Display/n1 [21]),
    .en(1'b1),
    .reset(~rst_n),
    .set(1'b0),
    .q(lcd_data[21]));  // source/rtl/Display.v(93)
  reg_ar_as_w1 \u2_Display/reg0_b22  (
    .clk(clk_vga),
    .d(\u2_Display/n1 [22]),
    .en(1'b1),
    .reset(~rst_n),
    .set(1'b0),
    .q(lcd_data[22]));  // source/rtl/Display.v(93)
  reg_ar_as_w1 \u2_Display/reg0_b23  (
    .clk(clk_vga),
    .d(\u2_Display/n1 [23]),
    .en(1'b1),
    .reset(~rst_n),
    .set(1'b0),
    .q(lcd_data[23]));  // source/rtl/Display.v(93)
  reg_ar_as_w1 \u2_Display/reg0_b3  (
    .clk(clk_vga),
    .d(\u2_Display/n1 [3]),
    .en(1'b1),
    .reset(~rst_n),
    .set(1'b0),
    .q(lcd_data[3]));  // source/rtl/Display.v(93)
  reg_ar_as_w1 \u2_Display/reg0_b4  (
    .clk(clk_vga),
    .d(\u2_Display/n1 [4]),
    .en(1'b1),
    .reset(~rst_n),
    .set(1'b0),
    .q(lcd_data[4]));  // source/rtl/Display.v(93)
  reg_ar_as_w1 \u2_Display/reg0_b5  (
    .clk(clk_vga),
    .d(\u2_Display/n1 [5]),
    .en(1'b1),
    .reset(~rst_n),
    .set(1'b0),
    .q(lcd_data[5]));  // source/rtl/Display.v(93)
  reg_ar_as_w1 \u2_Display/reg0_b6  (
    .clk(clk_vga),
    .d(\u2_Display/n1 [6]),
    .en(1'b1),
    .reset(~rst_n),
    .set(1'b0),
    .q(lcd_data[6]));  // source/rtl/Display.v(93)
  reg_ar_as_w1 \u2_Display/reg0_b7  (
    .clk(clk_vga),
    .d(\u2_Display/n1 [7]),
    .en(1'b1),
    .reset(~rst_n),
    .set(1'b0),
    .q(lcd_data[7]));  // source/rtl/Display.v(93)
  reg_ar_as_w1 \u2_Display/reg0_b8  (
    .clk(clk_vga),
    .d(\u2_Display/n1 [8]),
    .en(1'b1),
    .reset(~rst_n),
    .set(1'b0),
    .q(lcd_data[8]));  // source/rtl/Display.v(93)
  reg_ar_as_w1 \u2_Display/reg0_b9  (
    .clk(clk_vga),
    .d(\u2_Display/n1 [9]),
    .en(1'b1),
    .reset(~rst_n),
    .set(1'b0),
    .q(lcd_data[9]));  // source/rtl/Display.v(93)

endmodule 

module Clk_div  // source/rtl/Clk_div.v(2)
  (
  clk,
  rst_n,
  clk_div
  );

  input clk;  // source/rtl/Clk_div.v(4)
  input rst_n;  // source/rtl/Clk_div.v(5)
  output clk_div;  // source/rtl/Clk_div.v(7)

  wire n0;

  not u0 (n0, rst_n);  // source/rtl/Clk_div.v(15)
  PLL uut (
    .refclk(clk),
    .reset(n0),
    .clk0_out(clk_div));  // source/rtl/Clk_div.v(12)

endmodule 

module Driver  // source/rtl/Driver.v(11)
  (
  clk,
  lcd_data,
  rst_n,
  lcd_dclk,
  lcd_en,
  lcd_hs,
  lcd_rgb,
  lcd_vs,
  lcd_xpos,
  lcd_ypos
  );

  input clk;  // source/rtl/Driver.v(26)
  input [23:0] lcd_data;  // source/rtl/Driver.v(28)
  input rst_n;  // source/rtl/Driver.v(27)
  output lcd_dclk;  // source/rtl/Driver.v(31)
  output lcd_en;  // source/rtl/Driver.v(34)
  output lcd_hs;  // source/rtl/Driver.v(32)
  output [23:0] lcd_rgb;  // source/rtl/Driver.v(35)
  output lcd_vs;  // source/rtl/Driver.v(33)
  output [11:0] lcd_xpos;  // source/rtl/Driver.v(38)
  output [11:0] lcd_ypos;  // source/rtl/Driver.v(39)

  parameter H_BACK = 248;
  parameter H_DISP = 1280;
  parameter H_FRONT = 48;
  parameter H_SYNC = 112;
  parameter H_TOTAL = 1688;
  parameter V_BACK = 38;
  parameter V_DISP = 1024;
  parameter V_FRONT = 1;
  parameter V_SYNC = 3;
  parameter V_TOTAL = 1066;
  // localparam H_AHEAD = 12'b000000000001;
  wire [11:0] hcnt;  // source/rtl/Driver.v(44)
  wire [11:0] n2;
  wire [12:0] n20;
  wire [12:0] n21;
  wire [11:0] n3;
  wire [11:0] n7;
  wire [11:0] n8;
  wire [11:0] vcnt;  // source/rtl/Driver.v(45)
  wire lcd_request;  // source/rtl/Driver.v(46)
  wire n1;
  wire n10;
  wire n11;
  wire n12;
  wire n13;
  wire n14;
  wire n15;
  wire n16;
  wire n17;
  wire n18;
  wire n19;
  wire n4;
  wire n5;
  wire n6;

  add_pu12_pu12_o12 add0 (
    .i0(hcnt),
    .i1(12'b000000000001),
    .o(n2));  // source/rtl/Driver.v(59)
  add_pu12_pu12_o12 add1 (
    .i0(vcnt),
    .i1(12'b000000000001),
    .o(n7));  // source/rtl/Driver.v(77)
  eq_w12 eq0 (
    .i0(hcnt),
    .i1(12'b011010010111),
    .o(n5));  // source/rtl/Driver.v(72)
  eq_w12 eq1 (
    .i0(vcnt),
    .i1(12'b010000101001),
    .o(n6));  // source/rtl/Driver.v(74)
  lt_u12_u12 lt0 (
    .ci(1'b0),
    .i0(hcnt),
    .i1(12'b011010010111),
    .o(n1));  // source/rtl/Driver.v(58)
  lt_u12_u12 lt1 (
    .ci(1'b1),
    .i0(hcnt),
    .i1(12'b000001101111),
    .o(n4));  // source/rtl/Driver.v(65)
  lt_u12_u12 lt2 (
    .ci(1'b1),
    .i0(vcnt),
    .i1(12'b000000000010),
    .o(n10));  // source/rtl/Driver.v(81)
  lt_u12_u12 lt3 (
    .ci(1'b1),
    .i0(12'b000101101000),
    .i1(hcnt),
    .o(n11));  // source/rtl/Driver.v(87)
  lt_u12_u12 lt4 (
    .ci(1'b0),
    .i0(hcnt),
    .i1(12'b011001101000),
    .o(n12));  // source/rtl/Driver.v(87)
  lt_u12_u12 lt5 (
    .ci(1'b1),
    .i0(12'b000000101001),
    .i1(vcnt),
    .o(n14));  // source/rtl/Driver.v(88)
  lt_u12_u12 lt6 (
    .ci(1'b0),
    .i0(vcnt),
    .i1(12'b010000101001),
    .o(n15));  // source/rtl/Driver.v(88)
  lt_u12_u12 lt7 (
    .ci(1'b1),
    .i0(12'b000101100111),
    .i1(hcnt),
    .o(n17));  // source/rtl/Driver.v(94)
  lt_u12_u12 lt8 (
    .ci(1'b0),
    .i0(hcnt),
    .i1(12'b011001100111),
    .o(n18));  // source/rtl/Driver.v(94)
  binary_mux_s1_w1 mux0_b0 (
    .i0(1'b0),
    .i1(n2[0]),
    .sel(n1),
    .o(n3[0]));  // source/rtl/Driver.v(61)
  binary_mux_s1_w1 mux0_b1 (
    .i0(1'b0),
    .i1(n2[1]),
    .sel(n1),
    .o(n3[1]));  // source/rtl/Driver.v(61)
  binary_mux_s1_w1 mux0_b10 (
    .i0(1'b0),
    .i1(n2[10]),
    .sel(n1),
    .o(n3[10]));  // source/rtl/Driver.v(61)
  binary_mux_s1_w1 mux0_b11 (
    .i0(1'b0),
    .i1(n2[11]),
    .sel(n1),
    .o(n3[11]));  // source/rtl/Driver.v(61)
  binary_mux_s1_w1 mux0_b2 (
    .i0(1'b0),
    .i1(n2[2]),
    .sel(n1),
    .o(n3[2]));  // source/rtl/Driver.v(61)
  binary_mux_s1_w1 mux0_b3 (
    .i0(1'b0),
    .i1(n2[3]),
    .sel(n1),
    .o(n3[3]));  // source/rtl/Driver.v(61)
  binary_mux_s1_w1 mux0_b4 (
    .i0(1'b0),
    .i1(n2[4]),
    .sel(n1),
    .o(n3[4]));  // source/rtl/Driver.v(61)
  binary_mux_s1_w1 mux0_b5 (
    .i0(1'b0),
    .i1(n2[5]),
    .sel(n1),
    .o(n3[5]));  // source/rtl/Driver.v(61)
  binary_mux_s1_w1 mux0_b6 (
    .i0(1'b0),
    .i1(n2[6]),
    .sel(n1),
    .o(n3[6]));  // source/rtl/Driver.v(61)
  binary_mux_s1_w1 mux0_b7 (
    .i0(1'b0),
    .i1(n2[7]),
    .sel(n1),
    .o(n3[7]));  // source/rtl/Driver.v(61)
  binary_mux_s1_w1 mux0_b8 (
    .i0(1'b0),
    .i1(n2[8]),
    .sel(n1),
    .o(n3[8]));  // source/rtl/Driver.v(61)
  binary_mux_s1_w1 mux0_b9 (
    .i0(1'b0),
    .i1(n2[9]),
    .sel(n1),
    .o(n3[9]));  // source/rtl/Driver.v(61)
  binary_mux_s1_w1 mux1_b0 (
    .i0(n7[0]),
    .i1(1'b0),
    .sel(n6),
    .o(n8[0]));  // source/rtl/Driver.v(77)
  binary_mux_s1_w1 mux1_b1 (
    .i0(n7[1]),
    .i1(1'b0),
    .sel(n6),
    .o(n8[1]));  // source/rtl/Driver.v(77)
  binary_mux_s1_w1 mux1_b10 (
    .i0(n7[10]),
    .i1(1'b0),
    .sel(n6),
    .o(n8[10]));  // source/rtl/Driver.v(77)
  binary_mux_s1_w1 mux1_b11 (
    .i0(n7[11]),
    .i1(1'b0),
    .sel(n6),
    .o(n8[11]));  // source/rtl/Driver.v(77)
  binary_mux_s1_w1 mux1_b2 (
    .i0(n7[2]),
    .i1(1'b0),
    .sel(n6),
    .o(n8[2]));  // source/rtl/Driver.v(77)
  binary_mux_s1_w1 mux1_b3 (
    .i0(n7[3]),
    .i1(1'b0),
    .sel(n6),
    .o(n8[3]));  // source/rtl/Driver.v(77)
  binary_mux_s1_w1 mux1_b4 (
    .i0(n7[4]),
    .i1(1'b0),
    .sel(n6),
    .o(n8[4]));  // source/rtl/Driver.v(77)
  binary_mux_s1_w1 mux1_b5 (
    .i0(n7[5]),
    .i1(1'b0),
    .sel(n6),
    .o(n8[5]));  // source/rtl/Driver.v(77)
  binary_mux_s1_w1 mux1_b6 (
    .i0(n7[6]),
    .i1(1'b0),
    .sel(n6),
    .o(n8[6]));  // source/rtl/Driver.v(77)
  binary_mux_s1_w1 mux1_b7 (
    .i0(n7[7]),
    .i1(1'b0),
    .sel(n6),
    .o(n8[7]));  // source/rtl/Driver.v(77)
  binary_mux_s1_w1 mux1_b8 (
    .i0(n7[8]),
    .i1(1'b0),
    .sel(n6),
    .o(n8[8]));  // source/rtl/Driver.v(77)
  binary_mux_s1_w1 mux1_b9 (
    .i0(n7[9]),
    .i1(1'b0),
    .sel(n6),
    .o(n8[9]));  // source/rtl/Driver.v(77)
  binary_mux_s1_w1 mux3_b0 (
    .i0(1'b0),
    .i1(lcd_data[0]),
    .sel(lcd_en),
    .o(lcd_rgb[0]));  // source/rtl/Driver.v(91)
  binary_mux_s1_w1 mux3_b1 (
    .i0(1'b0),
    .i1(lcd_data[1]),
    .sel(lcd_en),
    .o(lcd_rgb[1]));  // source/rtl/Driver.v(91)
  binary_mux_s1_w1 mux3_b10 (
    .i0(1'b0),
    .i1(lcd_data[10]),
    .sel(lcd_en),
    .o(lcd_rgb[10]));  // source/rtl/Driver.v(91)
  binary_mux_s1_w1 mux3_b11 (
    .i0(1'b0),
    .i1(lcd_data[11]),
    .sel(lcd_en),
    .o(lcd_rgb[11]));  // source/rtl/Driver.v(91)
  binary_mux_s1_w1 mux3_b12 (
    .i0(1'b0),
    .i1(lcd_data[12]),
    .sel(lcd_en),
    .o(lcd_rgb[12]));  // source/rtl/Driver.v(91)
  binary_mux_s1_w1 mux3_b13 (
    .i0(1'b0),
    .i1(lcd_data[13]),
    .sel(lcd_en),
    .o(lcd_rgb[13]));  // source/rtl/Driver.v(91)
  binary_mux_s1_w1 mux3_b14 (
    .i0(1'b0),
    .i1(lcd_data[14]),
    .sel(lcd_en),
    .o(lcd_rgb[14]));  // source/rtl/Driver.v(91)
  binary_mux_s1_w1 mux3_b15 (
    .i0(1'b0),
    .i1(lcd_data[15]),
    .sel(lcd_en),
    .o(lcd_rgb[15]));  // source/rtl/Driver.v(91)
  binary_mux_s1_w1 mux3_b16 (
    .i0(1'b0),
    .i1(lcd_data[16]),
    .sel(lcd_en),
    .o(lcd_rgb[16]));  // source/rtl/Driver.v(91)
  binary_mux_s1_w1 mux3_b17 (
    .i0(1'b0),
    .i1(lcd_data[17]),
    .sel(lcd_en),
    .o(lcd_rgb[17]));  // source/rtl/Driver.v(91)
  binary_mux_s1_w1 mux3_b18 (
    .i0(1'b0),
    .i1(lcd_data[18]),
    .sel(lcd_en),
    .o(lcd_rgb[18]));  // source/rtl/Driver.v(91)
  binary_mux_s1_w1 mux3_b19 (
    .i0(1'b0),
    .i1(lcd_data[19]),
    .sel(lcd_en),
    .o(lcd_rgb[19]));  // source/rtl/Driver.v(91)
  binary_mux_s1_w1 mux3_b2 (
    .i0(1'b0),
    .i1(lcd_data[2]),
    .sel(lcd_en),
    .o(lcd_rgb[2]));  // source/rtl/Driver.v(91)
  binary_mux_s1_w1 mux3_b20 (
    .i0(1'b0),
    .i1(lcd_data[20]),
    .sel(lcd_en),
    .o(lcd_rgb[20]));  // source/rtl/Driver.v(91)
  binary_mux_s1_w1 mux3_b21 (
    .i0(1'b0),
    .i1(lcd_data[21]),
    .sel(lcd_en),
    .o(lcd_rgb[21]));  // source/rtl/Driver.v(91)
  binary_mux_s1_w1 mux3_b22 (
    .i0(1'b0),
    .i1(lcd_data[22]),
    .sel(lcd_en),
    .o(lcd_rgb[22]));  // source/rtl/Driver.v(91)
  binary_mux_s1_w1 mux3_b23 (
    .i0(1'b0),
    .i1(lcd_data[23]),
    .sel(lcd_en),
    .o(lcd_rgb[23]));  // source/rtl/Driver.v(91)
  binary_mux_s1_w1 mux3_b3 (
    .i0(1'b0),
    .i1(lcd_data[3]),
    .sel(lcd_en),
    .o(lcd_rgb[3]));  // source/rtl/Driver.v(91)
  binary_mux_s1_w1 mux3_b4 (
    .i0(1'b0),
    .i1(lcd_data[4]),
    .sel(lcd_en),
    .o(lcd_rgb[4]));  // source/rtl/Driver.v(91)
  binary_mux_s1_w1 mux3_b5 (
    .i0(1'b0),
    .i1(lcd_data[5]),
    .sel(lcd_en),
    .o(lcd_rgb[5]));  // source/rtl/Driver.v(91)
  binary_mux_s1_w1 mux3_b6 (
    .i0(1'b0),
    .i1(lcd_data[6]),
    .sel(lcd_en),
    .o(lcd_rgb[6]));  // source/rtl/Driver.v(91)
  binary_mux_s1_w1 mux3_b7 (
    .i0(1'b0),
    .i1(lcd_data[7]),
    .sel(lcd_en),
    .o(lcd_rgb[7]));  // source/rtl/Driver.v(91)
  binary_mux_s1_w1 mux3_b8 (
    .i0(1'b0),
    .i1(lcd_data[8]),
    .sel(lcd_en),
    .o(lcd_rgb[8]));  // source/rtl/Driver.v(91)
  binary_mux_s1_w1 mux3_b9 (
    .i0(1'b0),
    .i1(lcd_data[9]),
    .sel(lcd_en),
    .o(lcd_rgb[9]));  // source/rtl/Driver.v(91)
  binary_mux_s1_w1 mux4_b0 (
    .i0(1'b0),
    .i1(n20[0]),
    .sel(lcd_request),
    .o(lcd_xpos[0]));  // source/rtl/Driver.v(98)
  binary_mux_s1_w1 mux4_b1 (
    .i0(1'b0),
    .i1(n20[1]),
    .sel(lcd_request),
    .o(lcd_xpos[1]));  // source/rtl/Driver.v(98)
  binary_mux_s1_w1 mux4_b10 (
    .i0(1'b0),
    .i1(n20[10]),
    .sel(lcd_request),
    .o(lcd_xpos[10]));  // source/rtl/Driver.v(98)
  binary_mux_s1_w1 mux4_b11 (
    .i0(1'b0),
    .i1(n20[11]),
    .sel(lcd_request),
    .o(lcd_xpos[11]));  // source/rtl/Driver.v(98)
  binary_mux_s1_w1 mux4_b2 (
    .i0(1'b0),
    .i1(n20[2]),
    .sel(lcd_request),
    .o(lcd_xpos[2]));  // source/rtl/Driver.v(98)
  binary_mux_s1_w1 mux4_b3 (
    .i0(1'b0),
    .i1(n20[3]),
    .sel(lcd_request),
    .o(lcd_xpos[3]));  // source/rtl/Driver.v(98)
  binary_mux_s1_w1 mux4_b4 (
    .i0(1'b0),
    .i1(n20[4]),
    .sel(lcd_request),
    .o(lcd_xpos[4]));  // source/rtl/Driver.v(98)
  binary_mux_s1_w1 mux4_b5 (
    .i0(1'b0),
    .i1(n20[5]),
    .sel(lcd_request),
    .o(lcd_xpos[5]));  // source/rtl/Driver.v(98)
  binary_mux_s1_w1 mux4_b6 (
    .i0(1'b0),
    .i1(n20[6]),
    .sel(lcd_request),
    .o(lcd_xpos[6]));  // source/rtl/Driver.v(98)
  binary_mux_s1_w1 mux4_b7 (
    .i0(1'b0),
    .i1(n20[7]),
    .sel(lcd_request),
    .o(lcd_xpos[7]));  // source/rtl/Driver.v(98)
  binary_mux_s1_w1 mux4_b8 (
    .i0(1'b0),
    .i1(n20[8]),
    .sel(lcd_request),
    .o(lcd_xpos[8]));  // source/rtl/Driver.v(98)
  binary_mux_s1_w1 mux4_b9 (
    .i0(1'b0),
    .i1(n20[9]),
    .sel(lcd_request),
    .o(lcd_xpos[9]));  // source/rtl/Driver.v(98)
  binary_mux_s1_w1 mux5_b0 (
    .i0(1'b0),
    .i1(n21[0]),
    .sel(lcd_request),
    .o(lcd_ypos[0]));  // source/rtl/Driver.v(99)
  binary_mux_s1_w1 mux5_b1 (
    .i0(1'b0),
    .i1(n21[1]),
    .sel(lcd_request),
    .o(lcd_ypos[1]));  // source/rtl/Driver.v(99)
  binary_mux_s1_w1 mux5_b10 (
    .i0(1'b0),
    .i1(n21[10]),
    .sel(lcd_request),
    .o(lcd_ypos[10]));  // source/rtl/Driver.v(99)
  binary_mux_s1_w1 mux5_b11 (
    .i0(1'b0),
    .i1(n21[11]),
    .sel(lcd_request),
    .o(lcd_ypos[11]));  // source/rtl/Driver.v(99)
  binary_mux_s1_w1 mux5_b2 (
    .i0(1'b0),
    .i1(n21[2]),
    .sel(lcd_request),
    .o(lcd_ypos[2]));  // source/rtl/Driver.v(99)
  binary_mux_s1_w1 mux5_b3 (
    .i0(1'b0),
    .i1(n21[3]),
    .sel(lcd_request),
    .o(lcd_ypos[3]));  // source/rtl/Driver.v(99)
  binary_mux_s1_w1 mux5_b4 (
    .i0(1'b0),
    .i1(n21[4]),
    .sel(lcd_request),
    .o(lcd_ypos[4]));  // source/rtl/Driver.v(99)
  binary_mux_s1_w1 mux5_b5 (
    .i0(1'b0),
    .i1(n21[5]),
    .sel(lcd_request),
    .o(lcd_ypos[5]));  // source/rtl/Driver.v(99)
  binary_mux_s1_w1 mux5_b6 (
    .i0(1'b0),
    .i1(n21[6]),
    .sel(lcd_request),
    .o(lcd_ypos[6]));  // source/rtl/Driver.v(99)
  binary_mux_s1_w1 mux5_b7 (
    .i0(1'b0),
    .i1(n21[7]),
    .sel(lcd_request),
    .o(lcd_ypos[7]));  // source/rtl/Driver.v(99)
  binary_mux_s1_w1 mux5_b8 (
    .i0(1'b0),
    .i1(n21[8]),
    .sel(lcd_request),
    .o(lcd_ypos[8]));  // source/rtl/Driver.v(99)
  binary_mux_s1_w1 mux5_b9 (
    .i0(1'b0),
    .i1(n21[9]),
    .sel(lcd_request),
    .o(lcd_ypos[9]));  // source/rtl/Driver.v(99)
  reg_ar_as_w1 reg0_b0 (
    .clk(clk),
    .d(n8[0]),
    .en(n5),
    .reset(~rst_n),
    .set(1'b0),
    .q(vcnt[0]));  // source/rtl/Driver.v(78)
  reg_ar_as_w1 reg0_b1 (
    .clk(clk),
    .d(n8[1]),
    .en(n5),
    .reset(~rst_n),
    .set(1'b0),
    .q(vcnt[1]));  // source/rtl/Driver.v(78)
  reg_ar_as_w1 reg0_b10 (
    .clk(clk),
    .d(n8[10]),
    .en(n5),
    .reset(~rst_n),
    .set(1'b0),
    .q(vcnt[10]));  // source/rtl/Driver.v(78)
  reg_ar_as_w1 reg0_b11 (
    .clk(clk),
    .d(n8[11]),
    .en(n5),
    .reset(~rst_n),
    .set(1'b0),
    .q(vcnt[11]));  // source/rtl/Driver.v(78)
  reg_ar_as_w1 reg0_b2 (
    .clk(clk),
    .d(n8[2]),
    .en(n5),
    .reset(~rst_n),
    .set(1'b0),
    .q(vcnt[2]));  // source/rtl/Driver.v(78)
  reg_ar_as_w1 reg0_b3 (
    .clk(clk),
    .d(n8[3]),
    .en(n5),
    .reset(~rst_n),
    .set(1'b0),
    .q(vcnt[3]));  // source/rtl/Driver.v(78)
  reg_ar_as_w1 reg0_b4 (
    .clk(clk),
    .d(n8[4]),
    .en(n5),
    .reset(~rst_n),
    .set(1'b0),
    .q(vcnt[4]));  // source/rtl/Driver.v(78)
  reg_ar_as_w1 reg0_b5 (
    .clk(clk),
    .d(n8[5]),
    .en(n5),
    .reset(~rst_n),
    .set(1'b0),
    .q(vcnt[5]));  // source/rtl/Driver.v(78)
  reg_ar_as_w1 reg0_b6 (
    .clk(clk),
    .d(n8[6]),
    .en(n5),
    .reset(~rst_n),
    .set(1'b0),
    .q(vcnt[6]));  // source/rtl/Driver.v(78)
  reg_ar_as_w1 reg0_b7 (
    .clk(clk),
    .d(n8[7]),
    .en(n5),
    .reset(~rst_n),
    .set(1'b0),
    .q(vcnt[7]));  // source/rtl/Driver.v(78)
  reg_ar_as_w1 reg0_b8 (
    .clk(clk),
    .d(n8[8]),
    .en(n5),
    .reset(~rst_n),
    .set(1'b0),
    .q(vcnt[8]));  // source/rtl/Driver.v(78)
  reg_ar_as_w1 reg0_b9 (
    .clk(clk),
    .d(n8[9]),
    .en(n5),
    .reset(~rst_n),
    .set(1'b0),
    .q(vcnt[9]));  // source/rtl/Driver.v(78)
  reg_ar_as_w1 reg1_b0 (
    .clk(clk),
    .d(n3[0]),
    .en(1'b1),
    .reset(~rst_n),
    .set(1'b0),
    .q(hcnt[0]));  // source/rtl/Driver.v(62)
  reg_ar_as_w1 reg1_b1 (
    .clk(clk),
    .d(n3[1]),
    .en(1'b1),
    .reset(~rst_n),
    .set(1'b0),
    .q(hcnt[1]));  // source/rtl/Driver.v(62)
  reg_ar_as_w1 reg1_b10 (
    .clk(clk),
    .d(n3[10]),
    .en(1'b1),
    .reset(~rst_n),
    .set(1'b0),
    .q(hcnt[10]));  // source/rtl/Driver.v(62)
  reg_ar_as_w1 reg1_b11 (
    .clk(clk),
    .d(n3[11]),
    .en(1'b1),
    .reset(~rst_n),
    .set(1'b0),
    .q(hcnt[11]));  // source/rtl/Driver.v(62)
  reg_ar_as_w1 reg1_b2 (
    .clk(clk),
    .d(n3[2]),
    .en(1'b1),
    .reset(~rst_n),
    .set(1'b0),
    .q(hcnt[2]));  // source/rtl/Driver.v(62)
  reg_ar_as_w1 reg1_b3 (
    .clk(clk),
    .d(n3[3]),
    .en(1'b1),
    .reset(~rst_n),
    .set(1'b0),
    .q(hcnt[3]));  // source/rtl/Driver.v(62)
  reg_ar_as_w1 reg1_b4 (
    .clk(clk),
    .d(n3[4]),
    .en(1'b1),
    .reset(~rst_n),
    .set(1'b0),
    .q(hcnt[4]));  // source/rtl/Driver.v(62)
  reg_ar_as_w1 reg1_b5 (
    .clk(clk),
    .d(n3[5]),
    .en(1'b1),
    .reset(~rst_n),
    .set(1'b0),
    .q(hcnt[5]));  // source/rtl/Driver.v(62)
  reg_ar_as_w1 reg1_b6 (
    .clk(clk),
    .d(n3[6]),
    .en(1'b1),
    .reset(~rst_n),
    .set(1'b0),
    .q(hcnt[6]));  // source/rtl/Driver.v(62)
  reg_ar_as_w1 reg1_b7 (
    .clk(clk),
    .d(n3[7]),
    .en(1'b1),
    .reset(~rst_n),
    .set(1'b0),
    .q(hcnt[7]));  // source/rtl/Driver.v(62)
  reg_ar_as_w1 reg1_b8 (
    .clk(clk),
    .d(n3[8]),
    .en(1'b1),
    .reset(~rst_n),
    .set(1'b0),
    .q(hcnt[8]));  // source/rtl/Driver.v(62)
  reg_ar_as_w1 reg1_b9 (
    .clk(clk),
    .d(n3[9]),
    .en(1'b1),
    .reset(~rst_n),
    .set(1'b0),
    .q(hcnt[9]));  // source/rtl/Driver.v(62)
  add_pu12_mu12_o12 sub0 (
    .i0(hcnt),
    .i1(12'b000101100111),
    .o(n20[11:0]));  // source/rtl/Driver.v(98)
  add_pu12_mu12_o12 sub1 (
    .i0(vcnt),
    .i1(12'b000000101001),
    .o(n21[11:0]));  // source/rtl/Driver.v(99)
  and u10 (lcd_request, n19, n16);  // source/rtl/Driver.v(95)
  not u3 (lcd_hs, n4);  // source/rtl/Driver.v(65)
  not u4 (lcd_vs, n10);  // source/rtl/Driver.v(81)
  not u5 (lcd_dclk, clk);  // source/rtl/Driver.v(84)
  and u6 (n13, n11, n12);  // source/rtl/Driver.v(87)
  and u7 (n16, n14, n15);  // source/rtl/Driver.v(88)
  and u8 (lcd_en, n13, n16);  // source/rtl/Driver.v(88)
  and u9 (n19, n17, n18);  // source/rtl/Driver.v(94)

endmodule 

module mult_u12_u12_o24
  (
  i0,
  i1,
  o
  );

  input [11:0] i0;
  input [11:0] i1;
  output [23:0] o;

  wire a0;
  wire a1;
  wire a10;
  wire a11;
  wire a2;
  wire a3;
  wire a4;
  wire a5;
  wire a6;
  wire a7;
  wire a8;
  wire a9;
  wire b0;
  wire b1;
  wire b10;
  wire b11;
  wire b2;
  wire b3;
  wire b4;
  wire b5;
  wire b6;
  wire b7;
  wire b8;
  wire b9;
  wire net_and_a0_b0;
  wire net_and_a0_b1;
  wire net_and_a0_b10;
  wire net_and_a0_b11;
  wire net_and_a0_b2;
  wire net_and_a0_b3;
  wire net_and_a0_b4;
  wire net_and_a0_b5;
  wire net_and_a0_b6;
  wire net_and_a0_b7;
  wire net_and_a0_b8;
  wire net_and_a0_b9;
  wire net_and_a10_b0;
  wire net_and_a10_b1;
  wire net_and_a10_b10;
  wire net_and_a10_b11;
  wire net_and_a10_b2;
  wire net_and_a10_b3;
  wire net_and_a10_b4;
  wire net_and_a10_b5;
  wire net_and_a10_b6;
  wire net_and_a10_b7;
  wire net_and_a10_b8;
  wire net_and_a10_b9;
  wire net_and_a11_b0;
  wire net_and_a11_b1;
  wire net_and_a11_b10;
  wire net_and_a11_b11;
  wire net_and_a11_b2;
  wire net_and_a11_b3;
  wire net_and_a11_b4;
  wire net_and_a11_b5;
  wire net_and_a11_b6;
  wire net_and_a11_b7;
  wire net_and_a11_b8;
  wire net_and_a11_b9;
  wire net_and_a1_b0;
  wire net_and_a1_b1;
  wire net_and_a1_b10;
  wire net_and_a1_b11;
  wire net_and_a1_b2;
  wire net_and_a1_b3;
  wire net_and_a1_b4;
  wire net_and_a1_b5;
  wire net_and_a1_b6;
  wire net_and_a1_b7;
  wire net_and_a1_b8;
  wire net_and_a1_b9;
  wire net_and_a2_b0;
  wire net_and_a2_b1;
  wire net_and_a2_b10;
  wire net_and_a2_b11;
  wire net_and_a2_b2;
  wire net_and_a2_b3;
  wire net_and_a2_b4;
  wire net_and_a2_b5;
  wire net_and_a2_b6;
  wire net_and_a2_b7;
  wire net_and_a2_b8;
  wire net_and_a2_b9;
  wire net_and_a3_b0;
  wire net_and_a3_b1;
  wire net_and_a3_b10;
  wire net_and_a3_b11;
  wire net_and_a3_b2;
  wire net_and_a3_b3;
  wire net_and_a3_b4;
  wire net_and_a3_b5;
  wire net_and_a3_b6;
  wire net_and_a3_b7;
  wire net_and_a3_b8;
  wire net_and_a3_b9;
  wire net_and_a4_b0;
  wire net_and_a4_b1;
  wire net_and_a4_b10;
  wire net_and_a4_b11;
  wire net_and_a4_b2;
  wire net_and_a4_b3;
  wire net_and_a4_b4;
  wire net_and_a4_b5;
  wire net_and_a4_b6;
  wire net_and_a4_b7;
  wire net_and_a4_b8;
  wire net_and_a4_b9;
  wire net_and_a5_b0;
  wire net_and_a5_b1;
  wire net_and_a5_b10;
  wire net_and_a5_b11;
  wire net_and_a5_b2;
  wire net_and_a5_b3;
  wire net_and_a5_b4;
  wire net_and_a5_b5;
  wire net_and_a5_b6;
  wire net_and_a5_b7;
  wire net_and_a5_b8;
  wire net_and_a5_b9;
  wire net_and_a6_b0;
  wire net_and_a6_b1;
  wire net_and_a6_b10;
  wire net_and_a6_b11;
  wire net_and_a6_b2;
  wire net_and_a6_b3;
  wire net_and_a6_b4;
  wire net_and_a6_b5;
  wire net_and_a6_b6;
  wire net_and_a6_b7;
  wire net_and_a6_b8;
  wire net_and_a6_b9;
  wire net_and_a7_b0;
  wire net_and_a7_b1;
  wire net_and_a7_b10;
  wire net_and_a7_b11;
  wire net_and_a7_b2;
  wire net_and_a7_b3;
  wire net_and_a7_b4;
  wire net_and_a7_b5;
  wire net_and_a7_b6;
  wire net_and_a7_b7;
  wire net_and_a7_b8;
  wire net_and_a7_b9;
  wire net_and_a8_b0;
  wire net_and_a8_b1;
  wire net_and_a8_b10;
  wire net_and_a8_b11;
  wire net_and_a8_b2;
  wire net_and_a8_b3;
  wire net_and_a8_b4;
  wire net_and_a8_b5;
  wire net_and_a8_b6;
  wire net_and_a8_b7;
  wire net_and_a8_b8;
  wire net_and_a8_b9;
  wire net_and_a9_b0;
  wire net_and_a9_b1;
  wire net_and_a9_b10;
  wire net_and_a9_b11;
  wire net_and_a9_b2;
  wire net_and_a9_b3;
  wire net_and_a9_b4;
  wire net_and_a9_b5;
  wire net_and_a9_b6;
  wire net_and_a9_b7;
  wire net_and_a9_b8;
  wire net_and_a9_b9;
  wire o_0;
  wire o_1;
  wire o_10;
  wire o_11;
  wire o_12;
  wire o_13;
  wire o_14;
  wire o_15;
  wire o_16;
  wire o_17;
  wire o_18;
  wire o_19;
  wire o_2;
  wire o_20;
  wire o_21;
  wire o_22;
  wire o_23;
  wire o_3;
  wire o_4;
  wire o_5;
  wire o_6;
  wire o_7;
  wire o_8;
  wire o_9;

  assign a11 = i0[11];
  assign a10 = i0[10];
  assign a9 = i0[9];
  assign a8 = i0[8];
  assign a7 = i0[7];
  assign a6 = i0[6];
  assign a5 = i0[5];
  assign a4 = i0[4];
  assign a3 = i0[3];
  assign a2 = i0[2];
  assign a1 = i0[1];
  assign a0 = i0[0];
  assign b11 = i1[11];
  assign b10 = i1[10];
  assign b9 = i1[9];
  assign b8 = i1[8];
  assign b7 = i1[7];
  assign b6 = i1[6];
  assign b5 = i1[5];
  assign b4 = i1[4];
  assign b3 = i1[3];
  assign b2 = i1[2];
  assign b1 = i1[1];
  assign b0 = i1[0];
  assign o[23] = o_23;
  assign o[22] = o_22;
  assign o[21] = o_21;
  assign o[20] = o_20;
  assign o[19] = o_19;
  assign o[18] = o_18;
  assign o[17] = o_17;
  assign o[16] = o_16;
  assign o[15] = o_15;
  assign o[14] = o_14;
  assign o[13] = o_13;
  assign o[12] = o_12;
  assign o[11] = o_11;
  assign o[10] = o_10;
  assign o[9] = o_9;
  assign o[8] = o_8;
  assign o[7] = o_7;
  assign o[6] = o_6;
  assign o[5] = o_5;
  assign o[4] = o_4;
  assign o[3] = o_3;
  assign o[2] = o_2;
  assign o[1] = o_1;
  assign o[0] = o_0;
  and and_a0_b0 (net_and_a0_b0, a0, b0);
  and and_a0_b1 (net_and_a0_b1, a0, b1);
  and and_a0_b10 (net_and_a0_b10, a0, b10);
  and and_a0_b11 (net_and_a0_b11, a0, b11);
  and and_a0_b2 (net_and_a0_b2, a0, b2);
  and and_a0_b3 (net_and_a0_b3, a0, b3);
  and and_a0_b4 (net_and_a0_b4, a0, b4);
  and and_a0_b5 (net_and_a0_b5, a0, b5);
  and and_a0_b6 (net_and_a0_b6, a0, b6);
  and and_a0_b7 (net_and_a0_b7, a0, b7);
  and and_a0_b8 (net_and_a0_b8, a0, b8);
  and and_a0_b9 (net_and_a0_b9, a0, b9);
  and and_a10_b0 (net_and_a10_b0, a10, b0);
  and and_a10_b1 (net_and_a10_b1, a10, b1);
  and and_a10_b10 (net_and_a10_b10, a10, b10);
  and and_a10_b11 (net_and_a10_b11, a10, b11);
  and and_a10_b2 (net_and_a10_b2, a10, b2);
  and and_a10_b3 (net_and_a10_b3, a10, b3);
  and and_a10_b4 (net_and_a10_b4, a10, b4);
  and and_a10_b5 (net_and_a10_b5, a10, b5);
  and and_a10_b6 (net_and_a10_b6, a10, b6);
  and and_a10_b7 (net_and_a10_b7, a10, b7);
  and and_a10_b8 (net_and_a10_b8, a10, b8);
  and and_a10_b9 (net_and_a10_b9, a10, b9);
  and and_a11_b0 (net_and_a11_b0, a11, b0);
  and and_a11_b1 (net_and_a11_b1, a11, b1);
  and and_a11_b10 (net_and_a11_b10, a11, b10);
  and and_a11_b11 (net_and_a11_b11, a11, b11);
  and and_a11_b2 (net_and_a11_b2, a11, b2);
  and and_a11_b3 (net_and_a11_b3, a11, b3);
  and and_a11_b4 (net_and_a11_b4, a11, b4);
  and and_a11_b5 (net_and_a11_b5, a11, b5);
  and and_a11_b6 (net_and_a11_b6, a11, b6);
  and and_a11_b7 (net_and_a11_b7, a11, b7);
  and and_a11_b8 (net_and_a11_b8, a11, b8);
  and and_a11_b9 (net_and_a11_b9, a11, b9);
  and and_a1_b0 (net_and_a1_b0, a1, b0);
  and and_a1_b1 (net_and_a1_b1, a1, b1);
  and and_a1_b10 (net_and_a1_b10, a1, b10);
  and and_a1_b11 (net_and_a1_b11, a1, b11);
  and and_a1_b2 (net_and_a1_b2, a1, b2);
  and and_a1_b3 (net_and_a1_b3, a1, b3);
  and and_a1_b4 (net_and_a1_b4, a1, b4);
  and and_a1_b5 (net_and_a1_b5, a1, b5);
  and and_a1_b6 (net_and_a1_b6, a1, b6);
  and and_a1_b7 (net_and_a1_b7, a1, b7);
  and and_a1_b8 (net_and_a1_b8, a1, b8);
  and and_a1_b9 (net_and_a1_b9, a1, b9);
  and and_a2_b0 (net_and_a2_b0, a2, b0);
  and and_a2_b1 (net_and_a2_b1, a2, b1);
  and and_a2_b10 (net_and_a2_b10, a2, b10);
  and and_a2_b11 (net_and_a2_b11, a2, b11);
  and and_a2_b2 (net_and_a2_b2, a2, b2);
  and and_a2_b3 (net_and_a2_b3, a2, b3);
  and and_a2_b4 (net_and_a2_b4, a2, b4);
  and and_a2_b5 (net_and_a2_b5, a2, b5);
  and and_a2_b6 (net_and_a2_b6, a2, b6);
  and and_a2_b7 (net_and_a2_b7, a2, b7);
  and and_a2_b8 (net_and_a2_b8, a2, b8);
  and and_a2_b9 (net_and_a2_b9, a2, b9);
  and and_a3_b0 (net_and_a3_b0, a3, b0);
  and and_a3_b1 (net_and_a3_b1, a3, b1);
  and and_a3_b10 (net_and_a3_b10, a3, b10);
  and and_a3_b11 (net_and_a3_b11, a3, b11);
  and and_a3_b2 (net_and_a3_b2, a3, b2);
  and and_a3_b3 (net_and_a3_b3, a3, b3);
  and and_a3_b4 (net_and_a3_b4, a3, b4);
  and and_a3_b5 (net_and_a3_b5, a3, b5);
  and and_a3_b6 (net_and_a3_b6, a3, b6);
  and and_a3_b7 (net_and_a3_b7, a3, b7);
  and and_a3_b8 (net_and_a3_b8, a3, b8);
  and and_a3_b9 (net_and_a3_b9, a3, b9);
  and and_a4_b0 (net_and_a4_b0, a4, b0);
  and and_a4_b1 (net_and_a4_b1, a4, b1);
  and and_a4_b10 (net_and_a4_b10, a4, b10);
  and and_a4_b11 (net_and_a4_b11, a4, b11);
  and and_a4_b2 (net_and_a4_b2, a4, b2);
  and and_a4_b3 (net_and_a4_b3, a4, b3);
  and and_a4_b4 (net_and_a4_b4, a4, b4);
  and and_a4_b5 (net_and_a4_b5, a4, b5);
  and and_a4_b6 (net_and_a4_b6, a4, b6);
  and and_a4_b7 (net_and_a4_b7, a4, b7);
  and and_a4_b8 (net_and_a4_b8, a4, b8);
  and and_a4_b9 (net_and_a4_b9, a4, b9);
  and and_a5_b0 (net_and_a5_b0, a5, b0);
  and and_a5_b1 (net_and_a5_b1, a5, b1);
  and and_a5_b10 (net_and_a5_b10, a5, b10);
  and and_a5_b11 (net_and_a5_b11, a5, b11);
  and and_a5_b2 (net_and_a5_b2, a5, b2);
  and and_a5_b3 (net_and_a5_b3, a5, b3);
  and and_a5_b4 (net_and_a5_b4, a5, b4);
  and and_a5_b5 (net_and_a5_b5, a5, b5);
  and and_a5_b6 (net_and_a5_b6, a5, b6);
  and and_a5_b7 (net_and_a5_b7, a5, b7);
  and and_a5_b8 (net_and_a5_b8, a5, b8);
  and and_a5_b9 (net_and_a5_b9, a5, b9);
  and and_a6_b0 (net_and_a6_b0, a6, b0);
  and and_a6_b1 (net_and_a6_b1, a6, b1);
  and and_a6_b10 (net_and_a6_b10, a6, b10);
  and and_a6_b11 (net_and_a6_b11, a6, b11);
  and and_a6_b2 (net_and_a6_b2, a6, b2);
  and and_a6_b3 (net_and_a6_b3, a6, b3);
  and and_a6_b4 (net_and_a6_b4, a6, b4);
  and and_a6_b5 (net_and_a6_b5, a6, b5);
  and and_a6_b6 (net_and_a6_b6, a6, b6);
  and and_a6_b7 (net_and_a6_b7, a6, b7);
  and and_a6_b8 (net_and_a6_b8, a6, b8);
  and and_a6_b9 (net_and_a6_b9, a6, b9);
  and and_a7_b0 (net_and_a7_b0, a7, b0);
  and and_a7_b1 (net_and_a7_b1, a7, b1);
  and and_a7_b10 (net_and_a7_b10, a7, b10);
  and and_a7_b11 (net_and_a7_b11, a7, b11);
  and and_a7_b2 (net_and_a7_b2, a7, b2);
  and and_a7_b3 (net_and_a7_b3, a7, b3);
  and and_a7_b4 (net_and_a7_b4, a7, b4);
  and and_a7_b5 (net_and_a7_b5, a7, b5);
  and and_a7_b6 (net_and_a7_b6, a7, b6);
  and and_a7_b7 (net_and_a7_b7, a7, b7);
  and and_a7_b8 (net_and_a7_b8, a7, b8);
  and and_a7_b9 (net_and_a7_b9, a7, b9);
  and and_a8_b0 (net_and_a8_b0, a8, b0);
  and and_a8_b1 (net_and_a8_b1, a8, b1);
  and and_a8_b10 (net_and_a8_b10, a8, b10);
  and and_a8_b11 (net_and_a8_b11, a8, b11);
  and and_a8_b2 (net_and_a8_b2, a8, b2);
  and and_a8_b3 (net_and_a8_b3, a8, b3);
  and and_a8_b4 (net_and_a8_b4, a8, b4);
  and and_a8_b5 (net_and_a8_b5, a8, b5);
  and and_a8_b6 (net_and_a8_b6, a8, b6);
  and and_a8_b7 (net_and_a8_b7, a8, b7);
  and and_a8_b8 (net_and_a8_b8, a8, b8);
  and and_a8_b9 (net_and_a8_b9, a8, b9);
  and and_a9_b0 (net_and_a9_b0, a9, b0);
  and and_a9_b1 (net_and_a9_b1, a9, b1);
  and and_a9_b10 (net_and_a9_b10, a9, b10);
  and and_a9_b11 (net_and_a9_b11, a9, b11);
  and and_a9_b2 (net_and_a9_b2, a9, b2);
  and and_a9_b3 (net_and_a9_b3, a9, b3);
  and and_a9_b4 (net_and_a9_b4, a9, b4);
  and and_a9_b5 (net_and_a9_b5, a9, b5);
  and and_a9_b6 (net_and_a9_b6, a9, b6);
  and and_a9_b7 (net_and_a9_b7, a9, b7);
  and and_a9_b8 (net_and_a9_b8, a9, b8);
  and and_a9_b9 (net_and_a9_b9, a9, b9);
  add_pu23_pu22_pu21_pu20_pu19_pu18_pu17_pu16_pu15_pu14_pu13_pu12_o24 sum (
    .i0({net_and_a11_b11,net_and_a11_b10,net_and_a11_b9,net_and_a11_b8,net_and_a11_b7,net_and_a11_b6,net_and_a11_b5,net_and_a11_b4,net_and_a11_b3,net_and_a11_b2,net_and_a11_b1,net_and_a11_b0,net_and_a10_b0,net_and_a9_b0,net_and_a8_b0,net_and_a7_b0,net_and_a6_b0,net_and_a5_b0,net_and_a4_b0,net_and_a3_b0,net_and_a2_b0,net_and_a1_b0,net_and_a0_b0}),
    .i1({net_and_a10_b11,net_and_a10_b10,net_and_a10_b9,net_and_a10_b8,net_and_a10_b7,net_and_a10_b6,net_and_a10_b5,net_and_a10_b4,net_and_a10_b3,net_and_a10_b2,net_and_a10_b1,net_and_a9_b1,net_and_a8_b1,net_and_a7_b1,net_and_a6_b1,net_and_a5_b1,net_and_a4_b1,net_and_a3_b1,net_and_a2_b1,net_and_a1_b1,net_and_a0_b1,1'b0}),
    .i10({net_and_a1_b11,net_and_a1_b10,net_and_a0_b10,10'b0000000000}),
    .i11({net_and_a0_b11,11'b00000000000}),
    .i2({net_and_a9_b11,net_and_a9_b10,net_and_a9_b9,net_and_a9_b8,net_and_a9_b7,net_and_a9_b6,net_and_a9_b5,net_and_a9_b4,net_and_a9_b3,net_and_a9_b2,net_and_a8_b2,net_and_a7_b2,net_and_a6_b2,net_and_a5_b2,net_and_a4_b2,net_and_a3_b2,net_and_a2_b2,net_and_a1_b2,net_and_a0_b2,2'b00}),
    .i3({net_and_a8_b11,net_and_a8_b10,net_and_a8_b9,net_and_a8_b8,net_and_a8_b7,net_and_a8_b6,net_and_a8_b5,net_and_a8_b4,net_and_a8_b3,net_and_a7_b3,net_and_a6_b3,net_and_a5_b3,net_and_a4_b3,net_and_a3_b3,net_and_a2_b3,net_and_a1_b3,net_and_a0_b3,3'b000}),
    .i4({net_and_a7_b11,net_and_a7_b10,net_and_a7_b9,net_and_a7_b8,net_and_a7_b7,net_and_a7_b6,net_and_a7_b5,net_and_a7_b4,net_and_a6_b4,net_and_a5_b4,net_and_a4_b4,net_and_a3_b4,net_and_a2_b4,net_and_a1_b4,net_and_a0_b4,4'b0000}),
    .i5({net_and_a6_b11,net_and_a6_b10,net_and_a6_b9,net_and_a6_b8,net_and_a6_b7,net_and_a6_b6,net_and_a6_b5,net_and_a5_b5,net_and_a4_b5,net_and_a3_b5,net_and_a2_b5,net_and_a1_b5,net_and_a0_b5,5'b00000}),
    .i6({net_and_a5_b11,net_and_a5_b10,net_and_a5_b9,net_and_a5_b8,net_and_a5_b7,net_and_a5_b6,net_and_a4_b6,net_and_a3_b6,net_and_a2_b6,net_and_a1_b6,net_and_a0_b6,6'b000000}),
    .i7({net_and_a4_b11,net_and_a4_b10,net_and_a4_b9,net_and_a4_b8,net_and_a4_b7,net_and_a3_b7,net_and_a2_b7,net_and_a1_b7,net_and_a0_b7,7'b0000000}),
    .i8({net_and_a3_b11,net_and_a3_b10,net_and_a3_b9,net_and_a3_b8,net_and_a2_b8,net_and_a1_b8,net_and_a0_b8,8'b00000000}),
    .i9({net_and_a2_b11,net_and_a2_b10,net_and_a2_b9,net_and_a1_b9,net_and_a0_b9,9'b000000000}),
    .o({o_23,o_22,o_21,o_20,o_19,o_18,o_17,o_16,o_15,o_14,o_13,o_12,o_11,o_10,o_9,o_8,o_7,o_6,o_5,o_4,o_3,o_2,o_1,o_0}));

endmodule 

module reg_ar_as_w1
  (
  clk,
  d,
  en,
  reset,
  set,
  q
  );

  input clk;
  input d;
  input en;
  input reset;
  input set;
  output q;

  parameter REGSET = "RESET";
  wire enout;

  AL_MUX u_en0 (
    .i0(q),
    .i1(d),
    .sel(en),
    .o(enout));
  AL_DFF #(
    .INI((REGSET == "SET") ? 1'b1 : 1'b0))
    u_seq0 (
    .clk(clk),
    .d(enout),
    .reset(reset),
    .set(set),
    .q(q));

endmodule 

module PLL  // al_ip/PLL.v(22)
  (
  refclk,
  reset,
  clk0_out,
  extlock
  );

  input refclk;  // al_ip/PLL.v(27)
  input reset;  // al_ip/PLL.v(28)
  output clk0_out;  // al_ip/PLL.v(30)
  output extlock;  // al_ip/PLL.v(29)

  wire clk0_buf;  // al_ip/PLL.v(32)

  EG_LOGIC_BUFG bufg_feedback (
    .i(clk0_buf),
    .o(clk0_out));  // al_ip/PLL.v(34)
  EG_PHY_PLL #(
    .CLKC0_CPHASE(8),
    .CLKC0_DIV(9),
    .CLKC0_DIV2_ENABLE("DISABLE"),
    .CLKC0_ENABLE("ENABLE"),
    .CLKC0_FPHASE(0),
    .CLKC1_CPHASE(1),
    .CLKC1_DIV(1),
    .CLKC1_DIV2_ENABLE("DISABLE"),
    .CLKC1_ENABLE("DISABLE"),
    .CLKC1_FPHASE(0),
    .CLKC2_CPHASE(1),
    .CLKC2_DIV(1),
    .CLKC2_DIV2_ENABLE("DISABLE"),
    .CLKC2_ENABLE("DISABLE"),
    .CLKC2_FPHASE(0),
    .CLKC3_CPHASE(1),
    .CLKC3_DIV(1),
    .CLKC3_DIV2_ENABLE("DISABLE"),
    .CLKC3_ENABLE("DISABLE"),
    .CLKC3_FPHASE(0),
    .CLKC4_CPHASE(1),
    .CLKC4_DIV(1),
    .CLKC4_DIV2_ENABLE("DISABLE"),
    .CLKC4_ENABLE("DISABLE"),
    .CLKC4_FPHASE(0),
    .DERIVE_PLL_CLOCKS("DISABLE"),
    .DPHASE_SOURCE("DISABLE"),
    .DYNCFG("DISABLE"),
    .FBCLK_DIV(9),
    .FEEDBK_MODE("NORMAL"),
    .FEEDBK_PATH("CLKC0_EXT"),
    .FIN("24.000"),
    .FREQ_LOCK_ACCURACY(2),
    .GEN_BASIC_CLOCK("DISABLE"),
    .GMC_GAIN(6),
    .GMC_TEST(14),
    .ICP_CURRENT(3),
    .IF_ESCLKSTSW("DISABLE"),
    .INTFB_WAKE("DISABLE"),
    .KVCO(6),
    .LPF_CAPACITOR(3),
    .LPF_RESISTOR(2),
    .NORESET("DISABLE"),
    .ODIV_MUXC0("DIV"),
    .ODIV_MUXC1("DIV"),
    .ODIV_MUXC2("DIV"),
    .ODIV_MUXC3("DIV"),
    .ODIV_MUXC4("DIV"),
    .PLLC2RST_ENA("DISABLE"),
    .PLLC34RST_ENA("DISABLE"),
    .PLLMRST_ENA("DISABLE"),
    .PLLRST_ENA("ENABLE"),
    .PLL_LOCK_MODE(0),
    .PREDIV_MUXC0("VCO"),
    .PREDIV_MUXC1("VCO"),
    .PREDIV_MUXC2("VCO"),
    .PREDIV_MUXC3("VCO"),
    .PREDIV_MUXC4("VCO"),
    .REFCLK_DIV(2),
    .REFCLK_SEL("INTERNAL"),
    .STDBY_ENABLE("DISABLE"),
    .STDBY_VCO_ENA("DISABLE"),
    .SYNC_ENABLE("DISABLE"),
    .VCO_NORESET("DISABLE"))
    pll_inst (
    .daddr(6'b000000),
    .dclk(1'b0),
    .dcs(1'b0),
    .di(8'b00000000),
    .dwe(1'b0),
    .fbclk(clk0_out),
    .psclk(1'b0),
    .psclksel(3'b000),
    .psdown(1'b0),
    .psstep(1'b0),
    .refclk(refclk),
    .reset(reset),
    .stdby(1'b0),
    .clkc({open_n0,open_n1,open_n2,open_n3,clk0_buf}),
    .extlock(extlock));  // al_ip/PLL.v(57)

endmodule 

module add_pu12_pu12_o12
  (
  i0,
  i1,
  o
  );

  input [11:0] i0;
  input [11:0] i1;
  output [11:0] o;

  wire net_a0;
  wire net_a1;
  wire net_a10;
  wire net_a11;
  wire net_a2;
  wire net_a3;
  wire net_a4;
  wire net_a5;
  wire net_a6;
  wire net_a7;
  wire net_a8;
  wire net_a9;
  wire net_b0;
  wire net_b1;
  wire net_b10;
  wire net_b11;
  wire net_b2;
  wire net_b3;
  wire net_b4;
  wire net_b5;
  wire net_b6;
  wire net_b7;
  wire net_b8;
  wire net_b9;
  wire net_cout0;
  wire net_cout1;
  wire net_cout10;
  wire net_cout11;
  wire net_cout2;
  wire net_cout3;
  wire net_cout4;
  wire net_cout5;
  wire net_cout6;
  wire net_cout7;
  wire net_cout8;
  wire net_cout9;
  wire net_sum0;
  wire net_sum1;
  wire net_sum10;
  wire net_sum11;
  wire net_sum2;
  wire net_sum3;
  wire net_sum4;
  wire net_sum5;
  wire net_sum6;
  wire net_sum7;
  wire net_sum8;
  wire net_sum9;

  assign net_a11 = i0[11];
  assign net_a10 = i0[10];
  assign net_a9 = i0[9];
  assign net_a8 = i0[8];
  assign net_a7 = i0[7];
  assign net_a6 = i0[6];
  assign net_a5 = i0[5];
  assign net_a4 = i0[4];
  assign net_a3 = i0[3];
  assign net_a2 = i0[2];
  assign net_a1 = i0[1];
  assign net_a0 = i0[0];
  assign net_b11 = i1[11];
  assign net_b10 = i1[10];
  assign net_b9 = i1[9];
  assign net_b8 = i1[8];
  assign net_b7 = i1[7];
  assign net_b6 = i1[6];
  assign net_b5 = i1[5];
  assign net_b4 = i1[4];
  assign net_b3 = i1[3];
  assign net_b2 = i1[2];
  assign net_b1 = i1[1];
  assign net_b0 = i1[0];
  assign o[11] = net_sum11;
  assign o[10] = net_sum10;
  assign o[9] = net_sum9;
  assign o[8] = net_sum8;
  assign o[7] = net_sum7;
  assign o[6] = net_sum6;
  assign o[5] = net_sum5;
  assign o[4] = net_sum4;
  assign o[3] = net_sum3;
  assign o[2] = net_sum2;
  assign o[1] = net_sum1;
  assign o[0] = net_sum0;
  AL_FADD comp_0 (
    .a(net_a0),
    .b(net_b0),
    .c(1'b0),
    .cout(net_cout0),
    .sum(net_sum0));
  AL_FADD comp_1 (
    .a(net_a1),
    .b(net_b1),
    .c(net_cout0),
    .cout(net_cout1),
    .sum(net_sum1));
  AL_FADD comp_10 (
    .a(net_a10),
    .b(net_b10),
    .c(net_cout9),
    .cout(net_cout10),
    .sum(net_sum10));
  AL_FADD comp_11 (
    .a(net_a11),
    .b(net_b11),
    .c(net_cout10),
    .cout(net_cout11),
    .sum(net_sum11));
  AL_FADD comp_2 (
    .a(net_a2),
    .b(net_b2),
    .c(net_cout1),
    .cout(net_cout2),
    .sum(net_sum2));
  AL_FADD comp_3 (
    .a(net_a3),
    .b(net_b3),
    .c(net_cout2),
    .cout(net_cout3),
    .sum(net_sum3));
  AL_FADD comp_4 (
    .a(net_a4),
    .b(net_b4),
    .c(net_cout3),
    .cout(net_cout4),
    .sum(net_sum4));
  AL_FADD comp_5 (
    .a(net_a5),
    .b(net_b5),
    .c(net_cout4),
    .cout(net_cout5),
    .sum(net_sum5));
  AL_FADD comp_6 (
    .a(net_a6),
    .b(net_b6),
    .c(net_cout5),
    .cout(net_cout6),
    .sum(net_sum6));
  AL_FADD comp_7 (
    .a(net_a7),
    .b(net_b7),
    .c(net_cout6),
    .cout(net_cout7),
    .sum(net_sum7));
  AL_FADD comp_8 (
    .a(net_a8),
    .b(net_b8),
    .c(net_cout7),
    .cout(net_cout8),
    .sum(net_sum8));
  AL_FADD comp_9 (
    .a(net_a9),
    .b(net_b9),
    .c(net_cout8),
    .cout(net_cout9),
    .sum(net_sum9));

endmodule 

module eq_w12
  (
  i0,
  i1,
  o
  );

  input [11:0] i0;
  input [11:0] i1;
  output o;

  wire \or_or_or_xor_i0[0]_i_o ;
  wire \or_or_xor_i0[0]_i1[0_o ;
  wire \or_or_xor_i0[6]_i1[6_o ;
  wire \or_xor_i0[0]_i1[0]_o_o ;
  wire \or_xor_i0[10]_i1[10]_o ;
  wire \or_xor_i0[1]_i1[1]_o_o ;
  wire \or_xor_i0[3]_i1[3]_o_o ;
  wire \or_xor_i0[4]_i1[4]_o_o ;
  wire \or_xor_i0[6]_i1[6]_o_o ;
  wire \or_xor_i0[7]_i1[7]_o_o ;
  wire \or_xor_i0[9]_i1[9]_o_o ;
  wire \xor_i0[0]_i1[0]_o ;
  wire \xor_i0[10]_i1[10]_o ;
  wire \xor_i0[11]_i1[11]_o ;
  wire \xor_i0[1]_i1[1]_o ;
  wire \xor_i0[2]_i1[2]_o ;
  wire \xor_i0[3]_i1[3]_o ;
  wire \xor_i0[4]_i1[4]_o ;
  wire \xor_i0[5]_i1[5]_o ;
  wire \xor_i0[6]_i1[6]_o ;
  wire \xor_i0[7]_i1[7]_o ;
  wire \xor_i0[8]_i1[8]_o ;
  wire \xor_i0[9]_i1[9]_o ;

  not none_diff (o, \or_or_or_xor_i0[0]_i_o );
  or \or_or_or_xor_i0[0]_i  (\or_or_or_xor_i0[0]_i_o , \or_or_xor_i0[0]_i1[0_o , \or_or_xor_i0[6]_i1[6_o );
  or \or_or_xor_i0[0]_i1[0  (\or_or_xor_i0[0]_i1[0_o , \or_xor_i0[0]_i1[0]_o_o , \or_xor_i0[3]_i1[3]_o_o );
  or \or_or_xor_i0[6]_i1[6  (\or_or_xor_i0[6]_i1[6_o , \or_xor_i0[6]_i1[6]_o_o , \or_xor_i0[9]_i1[9]_o_o );
  or \or_xor_i0[0]_i1[0]_o  (\or_xor_i0[0]_i1[0]_o_o , \xor_i0[0]_i1[0]_o , \or_xor_i0[1]_i1[1]_o_o );
  or \or_xor_i0[10]_i1[10]  (\or_xor_i0[10]_i1[10]_o , \xor_i0[10]_i1[10]_o , \xor_i0[11]_i1[11]_o );
  or \or_xor_i0[1]_i1[1]_o  (\or_xor_i0[1]_i1[1]_o_o , \xor_i0[1]_i1[1]_o , \xor_i0[2]_i1[2]_o );
  or \or_xor_i0[3]_i1[3]_o  (\or_xor_i0[3]_i1[3]_o_o , \xor_i0[3]_i1[3]_o , \or_xor_i0[4]_i1[4]_o_o );
  or \or_xor_i0[4]_i1[4]_o  (\or_xor_i0[4]_i1[4]_o_o , \xor_i0[4]_i1[4]_o , \xor_i0[5]_i1[5]_o );
  or \or_xor_i0[6]_i1[6]_o  (\or_xor_i0[6]_i1[6]_o_o , \xor_i0[6]_i1[6]_o , \or_xor_i0[7]_i1[7]_o_o );
  or \or_xor_i0[7]_i1[7]_o  (\or_xor_i0[7]_i1[7]_o_o , \xor_i0[7]_i1[7]_o , \xor_i0[8]_i1[8]_o );
  or \or_xor_i0[9]_i1[9]_o  (\or_xor_i0[9]_i1[9]_o_o , \xor_i0[9]_i1[9]_o , \or_xor_i0[10]_i1[10]_o );
  xor \xor_i0[0]_i1[0]  (\xor_i0[0]_i1[0]_o , i0[0], i1[0]);
  xor \xor_i0[10]_i1[10]  (\xor_i0[10]_i1[10]_o , i0[10], i1[10]);
  xor \xor_i0[11]_i1[11]  (\xor_i0[11]_i1[11]_o , i0[11], i1[11]);
  xor \xor_i0[1]_i1[1]  (\xor_i0[1]_i1[1]_o , i0[1], i1[1]);
  xor \xor_i0[2]_i1[2]  (\xor_i0[2]_i1[2]_o , i0[2], i1[2]);
  xor \xor_i0[3]_i1[3]  (\xor_i0[3]_i1[3]_o , i0[3], i1[3]);
  xor \xor_i0[4]_i1[4]  (\xor_i0[4]_i1[4]_o , i0[4], i1[4]);
  xor \xor_i0[5]_i1[5]  (\xor_i0[5]_i1[5]_o , i0[5], i1[5]);
  xor \xor_i0[6]_i1[6]  (\xor_i0[6]_i1[6]_o , i0[6], i1[6]);
  xor \xor_i0[7]_i1[7]  (\xor_i0[7]_i1[7]_o , i0[7], i1[7]);
  xor \xor_i0[8]_i1[8]  (\xor_i0[8]_i1[8]_o , i0[8], i1[8]);
  xor \xor_i0[9]_i1[9]  (\xor_i0[9]_i1[9]_o , i0[9], i1[9]);

endmodule 

module lt_u12_u12
  (
  ci,
  i0,
  i1,
  o
  );

  input ci;
  input [11:0] i0;
  input [11:0] i1;
  output o;

  wire [11:0] diff;
  wire diff_6_11;
  wire less_6_11;
  wire \less_6_11_inst/diff_0 ;
  wire \less_6_11_inst/diff_1 ;
  wire \less_6_11_inst/diff_2 ;
  wire \less_6_11_inst/diff_3 ;
  wire \less_6_11_inst/diff_4 ;
  wire \less_6_11_inst/diff_5 ;
  wire \less_6_11_inst/o_0 ;
  wire \less_6_11_inst/o_1 ;
  wire \less_6_11_inst/o_2 ;
  wire \less_6_11_inst/o_3 ;
  wire \less_6_11_inst/o_4 ;
  wire o_0;
  wire o_1;
  wire o_2;
  wire o_3;
  wire o_4;
  wire o_5;

  or any_diff_6_11 (diff_6_11, diff[6], diff[7], diff[8], diff[9], diff[10], diff[11]);
  xor diff_0 (diff[0], i0[0], i1[0]);
  xor diff_1 (diff[1], i0[1], i1[1]);
  xor diff_10 (diff[10], i0[10], i1[10]);
  xor diff_11 (diff[11], i0[11], i1[11]);
  xor diff_2 (diff[2], i0[2], i1[2]);
  xor diff_3 (diff[3], i0[3], i1[3]);
  xor diff_4 (diff[4], i0[4], i1[4]);
  xor diff_5 (diff[5], i0[5], i1[5]);
  xor diff_6 (diff[6], i0[6], i1[6]);
  xor diff_7 (diff[7], i0[7], i1[7]);
  xor diff_8 (diff[8], i0[8], i1[8]);
  xor diff_9 (diff[9], i0[9], i1[9]);
  AL_MUX \less_6_11_inst/mux_0  (
    .i0(1'b0),
    .i1(i1[6]),
    .sel(\less_6_11_inst/diff_0 ),
    .o(\less_6_11_inst/o_0 ));
  AL_MUX \less_6_11_inst/mux_1  (
    .i0(\less_6_11_inst/o_0 ),
    .i1(i1[7]),
    .sel(\less_6_11_inst/diff_1 ),
    .o(\less_6_11_inst/o_1 ));
  AL_MUX \less_6_11_inst/mux_2  (
    .i0(\less_6_11_inst/o_1 ),
    .i1(i1[8]),
    .sel(\less_6_11_inst/diff_2 ),
    .o(\less_6_11_inst/o_2 ));
  AL_MUX \less_6_11_inst/mux_3  (
    .i0(\less_6_11_inst/o_2 ),
    .i1(i1[9]),
    .sel(\less_6_11_inst/diff_3 ),
    .o(\less_6_11_inst/o_3 ));
  AL_MUX \less_6_11_inst/mux_4  (
    .i0(\less_6_11_inst/o_3 ),
    .i1(i1[10]),
    .sel(\less_6_11_inst/diff_4 ),
    .o(\less_6_11_inst/o_4 ));
  AL_MUX \less_6_11_inst/mux_5  (
    .i0(\less_6_11_inst/o_4 ),
    .i1(i1[11]),
    .sel(\less_6_11_inst/diff_5 ),
    .o(less_6_11));
  xor \less_6_11_inst/xor_0  (\less_6_11_inst/diff_0 , i0[6], i1[6]);
  xor \less_6_11_inst/xor_1  (\less_6_11_inst/diff_1 , i0[7], i1[7]);
  xor \less_6_11_inst/xor_2  (\less_6_11_inst/diff_2 , i0[8], i1[8]);
  xor \less_6_11_inst/xor_3  (\less_6_11_inst/diff_3 , i0[9], i1[9]);
  xor \less_6_11_inst/xor_4  (\less_6_11_inst/diff_4 , i0[10], i1[10]);
  xor \less_6_11_inst/xor_5  (\less_6_11_inst/diff_5 , i0[11], i1[11]);
  AL_MUX mux_0 (
    .i0(ci),
    .i1(i1[0]),
    .sel(diff[0]),
    .o(o_0));
  AL_MUX mux_1 (
    .i0(o_0),
    .i1(i1[1]),
    .sel(diff[1]),
    .o(o_1));
  AL_MUX mux_2 (
    .i0(o_1),
    .i1(i1[2]),
    .sel(diff[2]),
    .o(o_2));
  AL_MUX mux_3 (
    .i0(o_2),
    .i1(i1[3]),
    .sel(diff[3]),
    .o(o_3));
  AL_MUX mux_4 (
    .i0(o_3),
    .i1(i1[4]),
    .sel(diff[4]),
    .o(o_4));
  AL_MUX mux_5 (
    .i0(o_4),
    .i1(i1[5]),
    .sel(diff[5]),
    .o(o_5));
  AL_MUX mux_6 (
    .i0(o_5),
    .i1(less_6_11),
    .sel(diff_6_11),
    .o(o));

endmodule 

module binary_mux_s1_w1
  (
  i0,
  i1,
  sel,
  o
  );

  input i0;
  input i1;
  input sel;
  output o;


  AL_MUX al_mux_b0_0_0 (
    .i0(i0),
    .i1(i1),
    .sel(sel),
    .o(o));

endmodule 

module add_pu12_mu12_o12
  (
  i0,
  i1,
  o
  );

  input [11:0] i0;
  input [11:0] i1;
  output [11:0] o;

  wire net_a0;
  wire net_a1;
  wire net_a10;
  wire net_a11;
  wire net_a2;
  wire net_a3;
  wire net_a4;
  wire net_a5;
  wire net_a6;
  wire net_a7;
  wire net_a8;
  wire net_a9;
  wire net_b0;
  wire net_b1;
  wire net_b10;
  wire net_b11;
  wire net_b2;
  wire net_b3;
  wire net_b4;
  wire net_b5;
  wire net_b6;
  wire net_b7;
  wire net_b8;
  wire net_b9;
  wire net_cout0;
  wire net_cout1;
  wire net_cout10;
  wire net_cout11;
  wire net_cout2;
  wire net_cout3;
  wire net_cout4;
  wire net_cout5;
  wire net_cout6;
  wire net_cout7;
  wire net_cout8;
  wire net_cout9;
  wire net_nb0;
  wire net_nb1;
  wire net_nb10;
  wire net_nb11;
  wire net_nb2;
  wire net_nb3;
  wire net_nb4;
  wire net_nb5;
  wire net_nb6;
  wire net_nb7;
  wire net_nb8;
  wire net_nb9;
  wire net_sum0;
  wire net_sum1;
  wire net_sum10;
  wire net_sum11;
  wire net_sum2;
  wire net_sum3;
  wire net_sum4;
  wire net_sum5;
  wire net_sum6;
  wire net_sum7;
  wire net_sum8;
  wire net_sum9;

  assign net_a11 = i0[11];
  assign net_a10 = i0[10];
  assign net_a9 = i0[9];
  assign net_a8 = i0[8];
  assign net_a7 = i0[7];
  assign net_a6 = i0[6];
  assign net_a5 = i0[5];
  assign net_a4 = i0[4];
  assign net_a3 = i0[3];
  assign net_a2 = i0[2];
  assign net_a1 = i0[1];
  assign net_a0 = i0[0];
  assign net_b11 = i1[11];
  assign net_b10 = i1[10];
  assign net_b9 = i1[9];
  assign net_b8 = i1[8];
  assign net_b7 = i1[7];
  assign net_b6 = i1[6];
  assign net_b5 = i1[5];
  assign net_b4 = i1[4];
  assign net_b3 = i1[3];
  assign net_b2 = i1[2];
  assign net_b1 = i1[1];
  assign net_b0 = i1[0];
  assign o[11] = net_sum11;
  assign o[10] = net_sum10;
  assign o[9] = net_sum9;
  assign o[8] = net_sum8;
  assign o[7] = net_sum7;
  assign o[6] = net_sum6;
  assign o[5] = net_sum5;
  assign o[4] = net_sum4;
  assign o[3] = net_sum3;
  assign o[2] = net_sum2;
  assign o[1] = net_sum1;
  assign o[0] = net_sum0;
  AL_FADD comp_0 (
    .a(net_a0),
    .b(net_nb0),
    .c(1'b1),
    .cout(net_cout0),
    .sum(net_sum0));
  AL_FADD comp_1 (
    .a(net_a1),
    .b(net_nb1),
    .c(net_cout0),
    .cout(net_cout1),
    .sum(net_sum1));
  AL_FADD comp_10 (
    .a(net_a10),
    .b(net_nb10),
    .c(net_cout9),
    .cout(net_cout10),
    .sum(net_sum10));
  AL_FADD comp_11 (
    .a(net_a11),
    .b(net_nb11),
    .c(net_cout10),
    .cout(net_cout11),
    .sum(net_sum11));
  AL_FADD comp_2 (
    .a(net_a2),
    .b(net_nb2),
    .c(net_cout1),
    .cout(net_cout2),
    .sum(net_sum2));
  AL_FADD comp_3 (
    .a(net_a3),
    .b(net_nb3),
    .c(net_cout2),
    .cout(net_cout3),
    .sum(net_sum3));
  AL_FADD comp_4 (
    .a(net_a4),
    .b(net_nb4),
    .c(net_cout3),
    .cout(net_cout4),
    .sum(net_sum4));
  AL_FADD comp_5 (
    .a(net_a5),
    .b(net_nb5),
    .c(net_cout4),
    .cout(net_cout5),
    .sum(net_sum5));
  AL_FADD comp_6 (
    .a(net_a6),
    .b(net_nb6),
    .c(net_cout5),
    .cout(net_cout6),
    .sum(net_sum6));
  AL_FADD comp_7 (
    .a(net_a7),
    .b(net_nb7),
    .c(net_cout6),
    .cout(net_cout7),
    .sum(net_sum7));
  AL_FADD comp_8 (
    .a(net_a8),
    .b(net_nb8),
    .c(net_cout7),
    .cout(net_cout8),
    .sum(net_sum8));
  AL_FADD comp_9 (
    .a(net_a9),
    .b(net_nb9),
    .c(net_cout8),
    .cout(net_cout9),
    .sum(net_sum9));
  not inv_b0 (net_nb0, net_b0);
  not inv_b1 (net_nb1, net_b1);
  not inv_b10 (net_nb10, net_b10);
  not inv_b11 (net_nb11, net_b11);
  not inv_b2 (net_nb2, net_b2);
  not inv_b3 (net_nb3, net_b3);
  not inv_b4 (net_nb4, net_b4);
  not inv_b5 (net_nb5, net_b5);
  not inv_b6 (net_nb6, net_b6);
  not inv_b7 (net_nb7, net_b7);
  not inv_b8 (net_nb8, net_b8);
  not inv_b9 (net_nb9, net_b9);

endmodule 

module add_pu23_pu22_pu21_pu20_pu19_pu18_pu17_pu16_pu15_pu14_pu13_pu12_o24
  (
  i0,
  i1,
  i10,
  i11,
  i2,
  i3,
  i4,
  i5,
  i6,
  i7,
  i8,
  i9,
  o
  );

  input [22:0] i0;
  input [21:0] i1;
  input [12:0] i10;
  input [11:0] i11;
  input [20:0] i2;
  input [19:0] i3;
  input [18:0] i4;
  input [17:0] i5;
  input [16:0] i6;
  input [15:0] i7;
  input [14:0] i8;
  input [13:0] i9;
  output [23:0] o;

  wire net_a0_0;
  wire net_a0_1;
  wire net_a0_10;
  wire net_a0_11;
  wire net_a0_12;
  wire net_a0_13;
  wire net_a0_14;
  wire net_a0_15;
  wire net_a0_16;
  wire net_a0_17;
  wire net_a0_18;
  wire net_a0_19;
  wire net_a0_2;
  wire net_a0_20;
  wire net_a0_21;
  wire net_a0_22;
  wire net_a0_3;
  wire net_a0_4;
  wire net_a0_5;
  wire net_a0_6;
  wire net_a0_7;
  wire net_a0_8;
  wire net_a0_9;
  wire net_a10_0;
  wire net_a10_1;
  wire net_a10_10;
  wire net_a10_11;
  wire net_a10_12;
  wire net_a10_2;
  wire net_a10_3;
  wire net_a10_4;
  wire net_a10_5;
  wire net_a10_6;
  wire net_a10_7;
  wire net_a10_8;
  wire net_a10_9;
  wire net_a11_0;
  wire net_a11_1;
  wire net_a11_10;
  wire net_a11_11;
  wire net_a11_2;
  wire net_a11_3;
  wire net_a11_4;
  wire net_a11_5;
  wire net_a11_6;
  wire net_a11_7;
  wire net_a11_8;
  wire net_a11_9;
  wire net_a1_0;
  wire net_a1_1;
  wire net_a1_10;
  wire net_a1_11;
  wire net_a1_12;
  wire net_a1_13;
  wire net_a1_14;
  wire net_a1_15;
  wire net_a1_16;
  wire net_a1_17;
  wire net_a1_18;
  wire net_a1_19;
  wire net_a1_2;
  wire net_a1_20;
  wire net_a1_21;
  wire net_a1_3;
  wire net_a1_4;
  wire net_a1_5;
  wire net_a1_6;
  wire net_a1_7;
  wire net_a1_8;
  wire net_a1_9;
  wire net_a2_0;
  wire net_a2_1;
  wire net_a2_10;
  wire net_a2_11;
  wire net_a2_12;
  wire net_a2_13;
  wire net_a2_14;
  wire net_a2_15;
  wire net_a2_16;
  wire net_a2_17;
  wire net_a2_18;
  wire net_a2_19;
  wire net_a2_2;
  wire net_a2_20;
  wire net_a2_3;
  wire net_a2_4;
  wire net_a2_5;
  wire net_a2_6;
  wire net_a2_7;
  wire net_a2_8;
  wire net_a2_9;
  wire net_a3_0;
  wire net_a3_1;
  wire net_a3_10;
  wire net_a3_11;
  wire net_a3_12;
  wire net_a3_13;
  wire net_a3_14;
  wire net_a3_15;
  wire net_a3_16;
  wire net_a3_17;
  wire net_a3_18;
  wire net_a3_19;
  wire net_a3_2;
  wire net_a3_3;
  wire net_a3_4;
  wire net_a3_5;
  wire net_a3_6;
  wire net_a3_7;
  wire net_a3_8;
  wire net_a3_9;
  wire net_a4_0;
  wire net_a4_1;
  wire net_a4_10;
  wire net_a4_11;
  wire net_a4_12;
  wire net_a4_13;
  wire net_a4_14;
  wire net_a4_15;
  wire net_a4_16;
  wire net_a4_17;
  wire net_a4_18;
  wire net_a4_2;
  wire net_a4_3;
  wire net_a4_4;
  wire net_a4_5;
  wire net_a4_6;
  wire net_a4_7;
  wire net_a4_8;
  wire net_a4_9;
  wire net_a5_0;
  wire net_a5_1;
  wire net_a5_10;
  wire net_a5_11;
  wire net_a5_12;
  wire net_a5_13;
  wire net_a5_14;
  wire net_a5_15;
  wire net_a5_16;
  wire net_a5_17;
  wire net_a5_2;
  wire net_a5_3;
  wire net_a5_4;
  wire net_a5_5;
  wire net_a5_6;
  wire net_a5_7;
  wire net_a5_8;
  wire net_a5_9;
  wire net_a6_0;
  wire net_a6_1;
  wire net_a6_10;
  wire net_a6_11;
  wire net_a6_12;
  wire net_a6_13;
  wire net_a6_14;
  wire net_a6_15;
  wire net_a6_16;
  wire net_a6_2;
  wire net_a6_3;
  wire net_a6_4;
  wire net_a6_5;
  wire net_a6_6;
  wire net_a6_7;
  wire net_a6_8;
  wire net_a6_9;
  wire net_a7_0;
  wire net_a7_1;
  wire net_a7_10;
  wire net_a7_11;
  wire net_a7_12;
  wire net_a7_13;
  wire net_a7_14;
  wire net_a7_15;
  wire net_a7_2;
  wire net_a7_3;
  wire net_a7_4;
  wire net_a7_5;
  wire net_a7_6;
  wire net_a7_7;
  wire net_a7_8;
  wire net_a7_9;
  wire net_a8_0;
  wire net_a8_1;
  wire net_a8_10;
  wire net_a8_11;
  wire net_a8_12;
  wire net_a8_13;
  wire net_a8_14;
  wire net_a8_2;
  wire net_a8_3;
  wire net_a8_4;
  wire net_a8_5;
  wire net_a8_6;
  wire net_a8_7;
  wire net_a8_8;
  wire net_a8_9;
  wire net_a9_0;
  wire net_a9_1;
  wire net_a9_10;
  wire net_a9_11;
  wire net_a9_12;
  wire net_a9_13;
  wire net_a9_2;
  wire net_a9_3;
  wire net_a9_4;
  wire net_a9_5;
  wire net_a9_6;
  wire net_a9_7;
  wire net_a9_8;
  wire net_a9_9;
  wire net_cout10_0;
  wire net_cout10_1;
  wire net_cout10_10;
  wire net_cout10_11;
  wire net_cout10_12;
  wire net_cout10_13;
  wire net_cout10_14;
  wire net_cout10_15;
  wire net_cout10_16;
  wire net_cout10_17;
  wire net_cout10_18;
  wire net_cout10_19;
  wire net_cout10_2;
  wire net_cout10_20;
  wire net_cout10_21;
  wire net_cout10_22;
  wire net_cout10_23;
  wire net_cout10_3;
  wire net_cout10_4;
  wire net_cout10_5;
  wire net_cout10_6;
  wire net_cout10_7;
  wire net_cout10_8;
  wire net_cout10_9;
  wire net_cout11_0;
  wire net_cout11_1;
  wire net_cout11_10;
  wire net_cout11_11;
  wire net_cout11_12;
  wire net_cout11_13;
  wire net_cout11_14;
  wire net_cout11_15;
  wire net_cout11_16;
  wire net_cout11_17;
  wire net_cout11_18;
  wire net_cout11_19;
  wire net_cout11_2;
  wire net_cout11_20;
  wire net_cout11_21;
  wire net_cout11_22;
  wire net_cout11_23;
  wire net_cout11_3;
  wire net_cout11_4;
  wire net_cout11_5;
  wire net_cout11_6;
  wire net_cout11_7;
  wire net_cout11_8;
  wire net_cout11_9;
  wire net_cout1_0;
  wire net_cout1_1;
  wire net_cout1_10;
  wire net_cout1_11;
  wire net_cout1_12;
  wire net_cout1_13;
  wire net_cout1_14;
  wire net_cout1_15;
  wire net_cout1_16;
  wire net_cout1_17;
  wire net_cout1_18;
  wire net_cout1_19;
  wire net_cout1_2;
  wire net_cout1_20;
  wire net_cout1_21;
  wire net_cout1_22;
  wire net_cout1_3;
  wire net_cout1_4;
  wire net_cout1_5;
  wire net_cout1_6;
  wire net_cout1_7;
  wire net_cout1_8;
  wire net_cout1_9;
  wire net_cout2_0;
  wire net_cout2_1;
  wire net_cout2_10;
  wire net_cout2_11;
  wire net_cout2_12;
  wire net_cout2_13;
  wire net_cout2_14;
  wire net_cout2_15;
  wire net_cout2_16;
  wire net_cout2_17;
  wire net_cout2_18;
  wire net_cout2_19;
  wire net_cout2_2;
  wire net_cout2_20;
  wire net_cout2_21;
  wire net_cout2_22;
  wire net_cout2_23;
  wire net_cout2_3;
  wire net_cout2_4;
  wire net_cout2_5;
  wire net_cout2_6;
  wire net_cout2_7;
  wire net_cout2_8;
  wire net_cout2_9;
  wire net_cout3_0;
  wire net_cout3_1;
  wire net_cout3_10;
  wire net_cout3_11;
  wire net_cout3_12;
  wire net_cout3_13;
  wire net_cout3_14;
  wire net_cout3_15;
  wire net_cout3_16;
  wire net_cout3_17;
  wire net_cout3_18;
  wire net_cout3_19;
  wire net_cout3_2;
  wire net_cout3_20;
  wire net_cout3_21;
  wire net_cout3_22;
  wire net_cout3_23;
  wire net_cout3_3;
  wire net_cout3_4;
  wire net_cout3_5;
  wire net_cout3_6;
  wire net_cout3_7;
  wire net_cout3_8;
  wire net_cout3_9;
  wire net_cout4_0;
  wire net_cout4_1;
  wire net_cout4_10;
  wire net_cout4_11;
  wire net_cout4_12;
  wire net_cout4_13;
  wire net_cout4_14;
  wire net_cout4_15;
  wire net_cout4_16;
  wire net_cout4_17;
  wire net_cout4_18;
  wire net_cout4_19;
  wire net_cout4_2;
  wire net_cout4_20;
  wire net_cout4_21;
  wire net_cout4_22;
  wire net_cout4_23;
  wire net_cout4_3;
  wire net_cout4_4;
  wire net_cout4_5;
  wire net_cout4_6;
  wire net_cout4_7;
  wire net_cout4_8;
  wire net_cout4_9;
  wire net_cout5_0;
  wire net_cout5_1;
  wire net_cout5_10;
  wire net_cout5_11;
  wire net_cout5_12;
  wire net_cout5_13;
  wire net_cout5_14;
  wire net_cout5_15;
  wire net_cout5_16;
  wire net_cout5_17;
  wire net_cout5_18;
  wire net_cout5_19;
  wire net_cout5_2;
  wire net_cout5_20;
  wire net_cout5_21;
  wire net_cout5_22;
  wire net_cout5_23;
  wire net_cout5_3;
  wire net_cout5_4;
  wire net_cout5_5;
  wire net_cout5_6;
  wire net_cout5_7;
  wire net_cout5_8;
  wire net_cout5_9;
  wire net_cout6_0;
  wire net_cout6_1;
  wire net_cout6_10;
  wire net_cout6_11;
  wire net_cout6_12;
  wire net_cout6_13;
  wire net_cout6_14;
  wire net_cout6_15;
  wire net_cout6_16;
  wire net_cout6_17;
  wire net_cout6_18;
  wire net_cout6_19;
  wire net_cout6_2;
  wire net_cout6_20;
  wire net_cout6_21;
  wire net_cout6_22;
  wire net_cout6_23;
  wire net_cout6_3;
  wire net_cout6_4;
  wire net_cout6_5;
  wire net_cout6_6;
  wire net_cout6_7;
  wire net_cout6_8;
  wire net_cout6_9;
  wire net_cout7_0;
  wire net_cout7_1;
  wire net_cout7_10;
  wire net_cout7_11;
  wire net_cout7_12;
  wire net_cout7_13;
  wire net_cout7_14;
  wire net_cout7_15;
  wire net_cout7_16;
  wire net_cout7_17;
  wire net_cout7_18;
  wire net_cout7_19;
  wire net_cout7_2;
  wire net_cout7_20;
  wire net_cout7_21;
  wire net_cout7_22;
  wire net_cout7_23;
  wire net_cout7_3;
  wire net_cout7_4;
  wire net_cout7_5;
  wire net_cout7_6;
  wire net_cout7_7;
  wire net_cout7_8;
  wire net_cout7_9;
  wire net_cout8_0;
  wire net_cout8_1;
  wire net_cout8_10;
  wire net_cout8_11;
  wire net_cout8_12;
  wire net_cout8_13;
  wire net_cout8_14;
  wire net_cout8_15;
  wire net_cout8_16;
  wire net_cout8_17;
  wire net_cout8_18;
  wire net_cout8_19;
  wire net_cout8_2;
  wire net_cout8_20;
  wire net_cout8_21;
  wire net_cout8_22;
  wire net_cout8_23;
  wire net_cout8_3;
  wire net_cout8_4;
  wire net_cout8_5;
  wire net_cout8_6;
  wire net_cout8_7;
  wire net_cout8_8;
  wire net_cout8_9;
  wire net_cout9_0;
  wire net_cout9_1;
  wire net_cout9_10;
  wire net_cout9_11;
  wire net_cout9_12;
  wire net_cout9_13;
  wire net_cout9_14;
  wire net_cout9_15;
  wire net_cout9_16;
  wire net_cout9_17;
  wire net_cout9_18;
  wire net_cout9_19;
  wire net_cout9_2;
  wire net_cout9_20;
  wire net_cout9_21;
  wire net_cout9_22;
  wire net_cout9_23;
  wire net_cout9_3;
  wire net_cout9_4;
  wire net_cout9_5;
  wire net_cout9_6;
  wire net_cout9_7;
  wire net_cout9_8;
  wire net_cout9_9;
  wire net_sum10_0;
  wire net_sum10_1;
  wire net_sum10_10;
  wire net_sum10_11;
  wire net_sum10_12;
  wire net_sum10_13;
  wire net_sum10_14;
  wire net_sum10_15;
  wire net_sum10_16;
  wire net_sum10_17;
  wire net_sum10_18;
  wire net_sum10_19;
  wire net_sum10_2;
  wire net_sum10_20;
  wire net_sum10_21;
  wire net_sum10_22;
  wire net_sum10_23;
  wire net_sum10_3;
  wire net_sum10_4;
  wire net_sum10_5;
  wire net_sum10_6;
  wire net_sum10_7;
  wire net_sum10_8;
  wire net_sum10_9;
  wire net_sum11_0;
  wire net_sum11_1;
  wire net_sum11_10;
  wire net_sum11_11;
  wire net_sum11_12;
  wire net_sum11_13;
  wire net_sum11_14;
  wire net_sum11_15;
  wire net_sum11_16;
  wire net_sum11_17;
  wire net_sum11_18;
  wire net_sum11_19;
  wire net_sum11_2;
  wire net_sum11_20;
  wire net_sum11_21;
  wire net_sum11_22;
  wire net_sum11_23;
  wire net_sum11_3;
  wire net_sum11_4;
  wire net_sum11_5;
  wire net_sum11_6;
  wire net_sum11_7;
  wire net_sum11_8;
  wire net_sum11_9;
  wire net_sum1_0;
  wire net_sum1_1;
  wire net_sum1_10;
  wire net_sum1_11;
  wire net_sum1_12;
  wire net_sum1_13;
  wire net_sum1_14;
  wire net_sum1_15;
  wire net_sum1_16;
  wire net_sum1_17;
  wire net_sum1_18;
  wire net_sum1_19;
  wire net_sum1_2;
  wire net_sum1_20;
  wire net_sum1_21;
  wire net_sum1_22;
  wire net_sum1_3;
  wire net_sum1_4;
  wire net_sum1_5;
  wire net_sum1_6;
  wire net_sum1_7;
  wire net_sum1_8;
  wire net_sum1_9;
  wire net_sum2_0;
  wire net_sum2_1;
  wire net_sum2_10;
  wire net_sum2_11;
  wire net_sum2_12;
  wire net_sum2_13;
  wire net_sum2_14;
  wire net_sum2_15;
  wire net_sum2_16;
  wire net_sum2_17;
  wire net_sum2_18;
  wire net_sum2_19;
  wire net_sum2_2;
  wire net_sum2_20;
  wire net_sum2_21;
  wire net_sum2_22;
  wire net_sum2_23;
  wire net_sum2_3;
  wire net_sum2_4;
  wire net_sum2_5;
  wire net_sum2_6;
  wire net_sum2_7;
  wire net_sum2_8;
  wire net_sum2_9;
  wire net_sum3_0;
  wire net_sum3_1;
  wire net_sum3_10;
  wire net_sum3_11;
  wire net_sum3_12;
  wire net_sum3_13;
  wire net_sum3_14;
  wire net_sum3_15;
  wire net_sum3_16;
  wire net_sum3_17;
  wire net_sum3_18;
  wire net_sum3_19;
  wire net_sum3_2;
  wire net_sum3_20;
  wire net_sum3_21;
  wire net_sum3_22;
  wire net_sum3_23;
  wire net_sum3_3;
  wire net_sum3_4;
  wire net_sum3_5;
  wire net_sum3_6;
  wire net_sum3_7;
  wire net_sum3_8;
  wire net_sum3_9;
  wire net_sum4_0;
  wire net_sum4_1;
  wire net_sum4_10;
  wire net_sum4_11;
  wire net_sum4_12;
  wire net_sum4_13;
  wire net_sum4_14;
  wire net_sum4_15;
  wire net_sum4_16;
  wire net_sum4_17;
  wire net_sum4_18;
  wire net_sum4_19;
  wire net_sum4_2;
  wire net_sum4_20;
  wire net_sum4_21;
  wire net_sum4_22;
  wire net_sum4_23;
  wire net_sum4_3;
  wire net_sum4_4;
  wire net_sum4_5;
  wire net_sum4_6;
  wire net_sum4_7;
  wire net_sum4_8;
  wire net_sum4_9;
  wire net_sum5_0;
  wire net_sum5_1;
  wire net_sum5_10;
  wire net_sum5_11;
  wire net_sum5_12;
  wire net_sum5_13;
  wire net_sum5_14;
  wire net_sum5_15;
  wire net_sum5_16;
  wire net_sum5_17;
  wire net_sum5_18;
  wire net_sum5_19;
  wire net_sum5_2;
  wire net_sum5_20;
  wire net_sum5_21;
  wire net_sum5_22;
  wire net_sum5_23;
  wire net_sum5_3;
  wire net_sum5_4;
  wire net_sum5_5;
  wire net_sum5_6;
  wire net_sum5_7;
  wire net_sum5_8;
  wire net_sum5_9;
  wire net_sum6_0;
  wire net_sum6_1;
  wire net_sum6_10;
  wire net_sum6_11;
  wire net_sum6_12;
  wire net_sum6_13;
  wire net_sum6_14;
  wire net_sum6_15;
  wire net_sum6_16;
  wire net_sum6_17;
  wire net_sum6_18;
  wire net_sum6_19;
  wire net_sum6_2;
  wire net_sum6_20;
  wire net_sum6_21;
  wire net_sum6_22;
  wire net_sum6_23;
  wire net_sum6_3;
  wire net_sum6_4;
  wire net_sum6_5;
  wire net_sum6_6;
  wire net_sum6_7;
  wire net_sum6_8;
  wire net_sum6_9;
  wire net_sum7_0;
  wire net_sum7_1;
  wire net_sum7_10;
  wire net_sum7_11;
  wire net_sum7_12;
  wire net_sum7_13;
  wire net_sum7_14;
  wire net_sum7_15;
  wire net_sum7_16;
  wire net_sum7_17;
  wire net_sum7_18;
  wire net_sum7_19;
  wire net_sum7_2;
  wire net_sum7_20;
  wire net_sum7_21;
  wire net_sum7_22;
  wire net_sum7_23;
  wire net_sum7_3;
  wire net_sum7_4;
  wire net_sum7_5;
  wire net_sum7_6;
  wire net_sum7_7;
  wire net_sum7_8;
  wire net_sum7_9;
  wire net_sum8_0;
  wire net_sum8_1;
  wire net_sum8_10;
  wire net_sum8_11;
  wire net_sum8_12;
  wire net_sum8_13;
  wire net_sum8_14;
  wire net_sum8_15;
  wire net_sum8_16;
  wire net_sum8_17;
  wire net_sum8_18;
  wire net_sum8_19;
  wire net_sum8_2;
  wire net_sum8_20;
  wire net_sum8_21;
  wire net_sum8_22;
  wire net_sum8_23;
  wire net_sum8_3;
  wire net_sum8_4;
  wire net_sum8_5;
  wire net_sum8_6;
  wire net_sum8_7;
  wire net_sum8_8;
  wire net_sum8_9;
  wire net_sum9_0;
  wire net_sum9_1;
  wire net_sum9_10;
  wire net_sum9_11;
  wire net_sum9_12;
  wire net_sum9_13;
  wire net_sum9_14;
  wire net_sum9_15;
  wire net_sum9_16;
  wire net_sum9_17;
  wire net_sum9_18;
  wire net_sum9_19;
  wire net_sum9_2;
  wire net_sum9_20;
  wire net_sum9_21;
  wire net_sum9_22;
  wire net_sum9_23;
  wire net_sum9_3;
  wire net_sum9_4;
  wire net_sum9_5;
  wire net_sum9_6;
  wire net_sum9_7;
  wire net_sum9_8;
  wire net_sum9_9;

  assign net_a0_22 = i0[22];
  assign net_a0_21 = i0[21];
  assign net_a0_20 = i0[20];
  assign net_a0_19 = i0[19];
  assign net_a0_18 = i0[18];
  assign net_a0_17 = i0[17];
  assign net_a0_16 = i0[16];
  assign net_a0_15 = i0[15];
  assign net_a0_14 = i0[14];
  assign net_a0_13 = i0[13];
  assign net_a0_12 = i0[12];
  assign net_a0_11 = i0[11];
  assign net_a0_10 = i0[10];
  assign net_a0_9 = i0[9];
  assign net_a0_8 = i0[8];
  assign net_a0_7 = i0[7];
  assign net_a0_6 = i0[6];
  assign net_a0_5 = i0[5];
  assign net_a0_4 = i0[4];
  assign net_a0_3 = i0[3];
  assign net_a0_2 = i0[2];
  assign net_a0_1 = i0[1];
  assign net_a0_0 = i0[0];
  assign net_a1_21 = i1[21];
  assign net_a1_20 = i1[20];
  assign net_a1_19 = i1[19];
  assign net_a1_18 = i1[18];
  assign net_a1_17 = i1[17];
  assign net_a1_16 = i1[16];
  assign net_a1_15 = i1[15];
  assign net_a1_14 = i1[14];
  assign net_a1_13 = i1[13];
  assign net_a1_12 = i1[12];
  assign net_a1_11 = i1[11];
  assign net_a1_10 = i1[10];
  assign net_a1_9 = i1[9];
  assign net_a1_8 = i1[8];
  assign net_a1_7 = i1[7];
  assign net_a1_6 = i1[6];
  assign net_a1_5 = i1[5];
  assign net_a1_4 = i1[4];
  assign net_a1_3 = i1[3];
  assign net_a1_2 = i1[2];
  assign net_a1_1 = i1[1];
  assign net_a1_0 = i1[0];
  assign net_a10_12 = i10[12];
  assign net_a10_11 = i10[11];
  assign net_a10_10 = i10[10];
  assign net_a10_9 = i10[9];
  assign net_a10_8 = i10[8];
  assign net_a10_7 = i10[7];
  assign net_a10_6 = i10[6];
  assign net_a10_5 = i10[5];
  assign net_a10_4 = i10[4];
  assign net_a10_3 = i10[3];
  assign net_a10_2 = i10[2];
  assign net_a10_1 = i10[1];
  assign net_a10_0 = i10[0];
  assign net_a11_11 = i11[11];
  assign net_a11_10 = i11[10];
  assign net_a11_9 = i11[9];
  assign net_a11_8 = i11[8];
  assign net_a11_7 = i11[7];
  assign net_a11_6 = i11[6];
  assign net_a11_5 = i11[5];
  assign net_a11_4 = i11[4];
  assign net_a11_3 = i11[3];
  assign net_a11_2 = i11[2];
  assign net_a11_1 = i11[1];
  assign net_a11_0 = i11[0];
  assign net_a2_20 = i2[20];
  assign net_a2_19 = i2[19];
  assign net_a2_18 = i2[18];
  assign net_a2_17 = i2[17];
  assign net_a2_16 = i2[16];
  assign net_a2_15 = i2[15];
  assign net_a2_14 = i2[14];
  assign net_a2_13 = i2[13];
  assign net_a2_12 = i2[12];
  assign net_a2_11 = i2[11];
  assign net_a2_10 = i2[10];
  assign net_a2_9 = i2[9];
  assign net_a2_8 = i2[8];
  assign net_a2_7 = i2[7];
  assign net_a2_6 = i2[6];
  assign net_a2_5 = i2[5];
  assign net_a2_4 = i2[4];
  assign net_a2_3 = i2[3];
  assign net_a2_2 = i2[2];
  assign net_a2_1 = i2[1];
  assign net_a2_0 = i2[0];
  assign net_a3_19 = i3[19];
  assign net_a3_18 = i3[18];
  assign net_a3_17 = i3[17];
  assign net_a3_16 = i3[16];
  assign net_a3_15 = i3[15];
  assign net_a3_14 = i3[14];
  assign net_a3_13 = i3[13];
  assign net_a3_12 = i3[12];
  assign net_a3_11 = i3[11];
  assign net_a3_10 = i3[10];
  assign net_a3_9 = i3[9];
  assign net_a3_8 = i3[8];
  assign net_a3_7 = i3[7];
  assign net_a3_6 = i3[6];
  assign net_a3_5 = i3[5];
  assign net_a3_4 = i3[4];
  assign net_a3_3 = i3[3];
  assign net_a3_2 = i3[2];
  assign net_a3_1 = i3[1];
  assign net_a3_0 = i3[0];
  assign net_a4_18 = i4[18];
  assign net_a4_17 = i4[17];
  assign net_a4_16 = i4[16];
  assign net_a4_15 = i4[15];
  assign net_a4_14 = i4[14];
  assign net_a4_13 = i4[13];
  assign net_a4_12 = i4[12];
  assign net_a4_11 = i4[11];
  assign net_a4_10 = i4[10];
  assign net_a4_9 = i4[9];
  assign net_a4_8 = i4[8];
  assign net_a4_7 = i4[7];
  assign net_a4_6 = i4[6];
  assign net_a4_5 = i4[5];
  assign net_a4_4 = i4[4];
  assign net_a4_3 = i4[3];
  assign net_a4_2 = i4[2];
  assign net_a4_1 = i4[1];
  assign net_a4_0 = i4[0];
  assign net_a5_17 = i5[17];
  assign net_a5_16 = i5[16];
  assign net_a5_15 = i5[15];
  assign net_a5_14 = i5[14];
  assign net_a5_13 = i5[13];
  assign net_a5_12 = i5[12];
  assign net_a5_11 = i5[11];
  assign net_a5_10 = i5[10];
  assign net_a5_9 = i5[9];
  assign net_a5_8 = i5[8];
  assign net_a5_7 = i5[7];
  assign net_a5_6 = i5[6];
  assign net_a5_5 = i5[5];
  assign net_a5_4 = i5[4];
  assign net_a5_3 = i5[3];
  assign net_a5_2 = i5[2];
  assign net_a5_1 = i5[1];
  assign net_a5_0 = i5[0];
  assign net_a6_16 = i6[16];
  assign net_a6_15 = i6[15];
  assign net_a6_14 = i6[14];
  assign net_a6_13 = i6[13];
  assign net_a6_12 = i6[12];
  assign net_a6_11 = i6[11];
  assign net_a6_10 = i6[10];
  assign net_a6_9 = i6[9];
  assign net_a6_8 = i6[8];
  assign net_a6_7 = i6[7];
  assign net_a6_6 = i6[6];
  assign net_a6_5 = i6[5];
  assign net_a6_4 = i6[4];
  assign net_a6_3 = i6[3];
  assign net_a6_2 = i6[2];
  assign net_a6_1 = i6[1];
  assign net_a6_0 = i6[0];
  assign net_a7_15 = i7[15];
  assign net_a7_14 = i7[14];
  assign net_a7_13 = i7[13];
  assign net_a7_12 = i7[12];
  assign net_a7_11 = i7[11];
  assign net_a7_10 = i7[10];
  assign net_a7_9 = i7[9];
  assign net_a7_8 = i7[8];
  assign net_a7_7 = i7[7];
  assign net_a7_6 = i7[6];
  assign net_a7_5 = i7[5];
  assign net_a7_4 = i7[4];
  assign net_a7_3 = i7[3];
  assign net_a7_2 = i7[2];
  assign net_a7_1 = i7[1];
  assign net_a7_0 = i7[0];
  assign net_a8_14 = i8[14];
  assign net_a8_13 = i8[13];
  assign net_a8_12 = i8[12];
  assign net_a8_11 = i8[11];
  assign net_a8_10 = i8[10];
  assign net_a8_9 = i8[9];
  assign net_a8_8 = i8[8];
  assign net_a8_7 = i8[7];
  assign net_a8_6 = i8[6];
  assign net_a8_5 = i8[5];
  assign net_a8_4 = i8[4];
  assign net_a8_3 = i8[3];
  assign net_a8_2 = i8[2];
  assign net_a8_1 = i8[1];
  assign net_a8_0 = i8[0];
  assign net_a9_13 = i9[13];
  assign net_a9_12 = i9[12];
  assign net_a9_11 = i9[11];
  assign net_a9_10 = i9[10];
  assign net_a9_9 = i9[9];
  assign net_a9_8 = i9[8];
  assign net_a9_7 = i9[7];
  assign net_a9_6 = i9[6];
  assign net_a9_5 = i9[5];
  assign net_a9_4 = i9[4];
  assign net_a9_3 = i9[3];
  assign net_a9_2 = i9[2];
  assign net_a9_1 = i9[1];
  assign net_a9_0 = i9[0];
  assign o[23] = net_sum11_23;
  assign o[22] = net_sum11_22;
  assign o[21] = net_sum11_21;
  assign o[20] = net_sum11_20;
  assign o[19] = net_sum11_19;
  assign o[18] = net_sum11_18;
  assign o[17] = net_sum11_17;
  assign o[16] = net_sum11_16;
  assign o[15] = net_sum11_15;
  assign o[14] = net_sum11_14;
  assign o[13] = net_sum11_13;
  assign o[12] = net_sum11_12;
  assign o[11] = net_sum11_11;
  assign o[10] = net_sum11_10;
  assign o[9] = net_sum11_9;
  assign o[8] = net_sum11_8;
  assign o[7] = net_sum11_7;
  assign o[6] = net_sum11_6;
  assign o[5] = net_sum11_5;
  assign o[4] = net_sum11_4;
  assign o[3] = net_sum11_3;
  assign o[2] = net_sum11_2;
  assign o[1] = net_sum11_1;
  assign o[0] = net_sum11_0;
  AL_FADD comp10_0 (
    .a(net_a10_0),
    .b(net_sum9_0),
    .c(1'b0),
    .cout(net_cout10_0),
    .sum(net_sum10_0));
  AL_FADD comp10_1 (
    .a(net_a10_1),
    .b(net_sum9_1),
    .c(net_cout10_0),
    .cout(net_cout10_1),
    .sum(net_sum10_1));
  AL_FADD comp10_10 (
    .a(net_a10_10),
    .b(net_sum9_10),
    .c(net_cout10_9),
    .cout(net_cout10_10),
    .sum(net_sum10_10));
  AL_FADD comp10_11 (
    .a(net_a10_11),
    .b(net_sum9_11),
    .c(net_cout10_10),
    .cout(net_cout10_11),
    .sum(net_sum10_11));
  AL_FADD comp10_12 (
    .a(net_a10_12),
    .b(net_sum9_12),
    .c(net_cout10_11),
    .cout(net_cout10_12),
    .sum(net_sum10_12));
  AL_FADD comp10_13 (
    .a(1'b0),
    .b(net_sum9_13),
    .c(net_cout10_12),
    .cout(net_cout10_13),
    .sum(net_sum10_13));
  AL_FADD comp10_14 (
    .a(1'b0),
    .b(net_sum9_14),
    .c(net_cout10_13),
    .cout(net_cout10_14),
    .sum(net_sum10_14));
  AL_FADD comp10_15 (
    .a(1'b0),
    .b(net_sum9_15),
    .c(net_cout10_14),
    .cout(net_cout10_15),
    .sum(net_sum10_15));
  AL_FADD comp10_16 (
    .a(1'b0),
    .b(net_sum9_16),
    .c(net_cout10_15),
    .cout(net_cout10_16),
    .sum(net_sum10_16));
  AL_FADD comp10_17 (
    .a(1'b0),
    .b(net_sum9_17),
    .c(net_cout10_16),
    .cout(net_cout10_17),
    .sum(net_sum10_17));
  AL_FADD comp10_18 (
    .a(1'b0),
    .b(net_sum9_18),
    .c(net_cout10_17),
    .cout(net_cout10_18),
    .sum(net_sum10_18));
  AL_FADD comp10_19 (
    .a(1'b0),
    .b(net_sum9_19),
    .c(net_cout10_18),
    .cout(net_cout10_19),
    .sum(net_sum10_19));
  AL_FADD comp10_2 (
    .a(net_a10_2),
    .b(net_sum9_2),
    .c(net_cout10_1),
    .cout(net_cout10_2),
    .sum(net_sum10_2));
  AL_FADD comp10_20 (
    .a(1'b0),
    .b(net_sum9_20),
    .c(net_cout10_19),
    .cout(net_cout10_20),
    .sum(net_sum10_20));
  AL_FADD comp10_21 (
    .a(1'b0),
    .b(net_sum9_21),
    .c(net_cout10_20),
    .cout(net_cout10_21),
    .sum(net_sum10_21));
  AL_FADD comp10_22 (
    .a(1'b0),
    .b(net_sum9_22),
    .c(net_cout10_21),
    .cout(net_cout10_22),
    .sum(net_sum10_22));
  AL_FADD comp10_23 (
    .a(1'b0),
    .b(net_sum9_23),
    .c(net_cout10_22),
    .cout(net_cout10_23),
    .sum(net_sum10_23));
  AL_FADD comp10_3 (
    .a(net_a10_3),
    .b(net_sum9_3),
    .c(net_cout10_2),
    .cout(net_cout10_3),
    .sum(net_sum10_3));
  AL_FADD comp10_4 (
    .a(net_a10_4),
    .b(net_sum9_4),
    .c(net_cout10_3),
    .cout(net_cout10_4),
    .sum(net_sum10_4));
  AL_FADD comp10_5 (
    .a(net_a10_5),
    .b(net_sum9_5),
    .c(net_cout10_4),
    .cout(net_cout10_5),
    .sum(net_sum10_5));
  AL_FADD comp10_6 (
    .a(net_a10_6),
    .b(net_sum9_6),
    .c(net_cout10_5),
    .cout(net_cout10_6),
    .sum(net_sum10_6));
  AL_FADD comp10_7 (
    .a(net_a10_7),
    .b(net_sum9_7),
    .c(net_cout10_6),
    .cout(net_cout10_7),
    .sum(net_sum10_7));
  AL_FADD comp10_8 (
    .a(net_a10_8),
    .b(net_sum9_8),
    .c(net_cout10_7),
    .cout(net_cout10_8),
    .sum(net_sum10_8));
  AL_FADD comp10_9 (
    .a(net_a10_9),
    .b(net_sum9_9),
    .c(net_cout10_8),
    .cout(net_cout10_9),
    .sum(net_sum10_9));
  AL_FADD comp11_0 (
    .a(net_a11_0),
    .b(net_sum10_0),
    .c(1'b0),
    .cout(net_cout11_0),
    .sum(net_sum11_0));
  AL_FADD comp11_1 (
    .a(net_a11_1),
    .b(net_sum10_1),
    .c(net_cout11_0),
    .cout(net_cout11_1),
    .sum(net_sum11_1));
  AL_FADD comp11_10 (
    .a(net_a11_10),
    .b(net_sum10_10),
    .c(net_cout11_9),
    .cout(net_cout11_10),
    .sum(net_sum11_10));
  AL_FADD comp11_11 (
    .a(net_a11_11),
    .b(net_sum10_11),
    .c(net_cout11_10),
    .cout(net_cout11_11),
    .sum(net_sum11_11));
  AL_FADD comp11_12 (
    .a(1'b0),
    .b(net_sum10_12),
    .c(net_cout11_11),
    .cout(net_cout11_12),
    .sum(net_sum11_12));
  AL_FADD comp11_13 (
    .a(1'b0),
    .b(net_sum10_13),
    .c(net_cout11_12),
    .cout(net_cout11_13),
    .sum(net_sum11_13));
  AL_FADD comp11_14 (
    .a(1'b0),
    .b(net_sum10_14),
    .c(net_cout11_13),
    .cout(net_cout11_14),
    .sum(net_sum11_14));
  AL_FADD comp11_15 (
    .a(1'b0),
    .b(net_sum10_15),
    .c(net_cout11_14),
    .cout(net_cout11_15),
    .sum(net_sum11_15));
  AL_FADD comp11_16 (
    .a(1'b0),
    .b(net_sum10_16),
    .c(net_cout11_15),
    .cout(net_cout11_16),
    .sum(net_sum11_16));
  AL_FADD comp11_17 (
    .a(1'b0),
    .b(net_sum10_17),
    .c(net_cout11_16),
    .cout(net_cout11_17),
    .sum(net_sum11_17));
  AL_FADD comp11_18 (
    .a(1'b0),
    .b(net_sum10_18),
    .c(net_cout11_17),
    .cout(net_cout11_18),
    .sum(net_sum11_18));
  AL_FADD comp11_19 (
    .a(1'b0),
    .b(net_sum10_19),
    .c(net_cout11_18),
    .cout(net_cout11_19),
    .sum(net_sum11_19));
  AL_FADD comp11_2 (
    .a(net_a11_2),
    .b(net_sum10_2),
    .c(net_cout11_1),
    .cout(net_cout11_2),
    .sum(net_sum11_2));
  AL_FADD comp11_20 (
    .a(1'b0),
    .b(net_sum10_20),
    .c(net_cout11_19),
    .cout(net_cout11_20),
    .sum(net_sum11_20));
  AL_FADD comp11_21 (
    .a(1'b0),
    .b(net_sum10_21),
    .c(net_cout11_20),
    .cout(net_cout11_21),
    .sum(net_sum11_21));
  AL_FADD comp11_22 (
    .a(1'b0),
    .b(net_sum10_22),
    .c(net_cout11_21),
    .cout(net_cout11_22),
    .sum(net_sum11_22));
  AL_FADD comp11_23 (
    .a(1'b0),
    .b(net_sum10_23),
    .c(net_cout11_22),
    .cout(net_cout11_23),
    .sum(net_sum11_23));
  AL_FADD comp11_3 (
    .a(net_a11_3),
    .b(net_sum10_3),
    .c(net_cout11_2),
    .cout(net_cout11_3),
    .sum(net_sum11_3));
  AL_FADD comp11_4 (
    .a(net_a11_4),
    .b(net_sum10_4),
    .c(net_cout11_3),
    .cout(net_cout11_4),
    .sum(net_sum11_4));
  AL_FADD comp11_5 (
    .a(net_a11_5),
    .b(net_sum10_5),
    .c(net_cout11_4),
    .cout(net_cout11_5),
    .sum(net_sum11_5));
  AL_FADD comp11_6 (
    .a(net_a11_6),
    .b(net_sum10_6),
    .c(net_cout11_5),
    .cout(net_cout11_6),
    .sum(net_sum11_6));
  AL_FADD comp11_7 (
    .a(net_a11_7),
    .b(net_sum10_7),
    .c(net_cout11_6),
    .cout(net_cout11_7),
    .sum(net_sum11_7));
  AL_FADD comp11_8 (
    .a(net_a11_8),
    .b(net_sum10_8),
    .c(net_cout11_7),
    .cout(net_cout11_8),
    .sum(net_sum11_8));
  AL_FADD comp11_9 (
    .a(net_a11_9),
    .b(net_sum10_9),
    .c(net_cout11_8),
    .cout(net_cout11_9),
    .sum(net_sum11_9));
  AL_FADD comp1_0 (
    .a(net_a1_0),
    .b(net_a0_0),
    .c(1'b0),
    .cout(net_cout1_0),
    .sum(net_sum1_0));
  AL_FADD comp1_1 (
    .a(net_a1_1),
    .b(net_a0_1),
    .c(net_cout1_0),
    .cout(net_cout1_1),
    .sum(net_sum1_1));
  AL_FADD comp1_10 (
    .a(net_a1_10),
    .b(net_a0_10),
    .c(net_cout1_9),
    .cout(net_cout1_10),
    .sum(net_sum1_10));
  AL_FADD comp1_11 (
    .a(net_a1_11),
    .b(net_a0_11),
    .c(net_cout1_10),
    .cout(net_cout1_11),
    .sum(net_sum1_11));
  AL_FADD comp1_12 (
    .a(net_a1_12),
    .b(net_a0_12),
    .c(net_cout1_11),
    .cout(net_cout1_12),
    .sum(net_sum1_12));
  AL_FADD comp1_13 (
    .a(net_a1_13),
    .b(net_a0_13),
    .c(net_cout1_12),
    .cout(net_cout1_13),
    .sum(net_sum1_13));
  AL_FADD comp1_14 (
    .a(net_a1_14),
    .b(net_a0_14),
    .c(net_cout1_13),
    .cout(net_cout1_14),
    .sum(net_sum1_14));
  AL_FADD comp1_15 (
    .a(net_a1_15),
    .b(net_a0_15),
    .c(net_cout1_14),
    .cout(net_cout1_15),
    .sum(net_sum1_15));
  AL_FADD comp1_16 (
    .a(net_a1_16),
    .b(net_a0_16),
    .c(net_cout1_15),
    .cout(net_cout1_16),
    .sum(net_sum1_16));
  AL_FADD comp1_17 (
    .a(net_a1_17),
    .b(net_a0_17),
    .c(net_cout1_16),
    .cout(net_cout1_17),
    .sum(net_sum1_17));
  AL_FADD comp1_18 (
    .a(net_a1_18),
    .b(net_a0_18),
    .c(net_cout1_17),
    .cout(net_cout1_18),
    .sum(net_sum1_18));
  AL_FADD comp1_19 (
    .a(net_a1_19),
    .b(net_a0_19),
    .c(net_cout1_18),
    .cout(net_cout1_19),
    .sum(net_sum1_19));
  AL_FADD comp1_2 (
    .a(net_a1_2),
    .b(net_a0_2),
    .c(net_cout1_1),
    .cout(net_cout1_2),
    .sum(net_sum1_2));
  AL_FADD comp1_20 (
    .a(net_a1_20),
    .b(net_a0_20),
    .c(net_cout1_19),
    .cout(net_cout1_20),
    .sum(net_sum1_20));
  AL_FADD comp1_21 (
    .a(net_a1_21),
    .b(net_a0_21),
    .c(net_cout1_20),
    .cout(net_cout1_21),
    .sum(net_sum1_21));
  AL_FADD comp1_22 (
    .a(1'b0),
    .b(net_a0_22),
    .c(net_cout1_21),
    .cout(net_cout1_22),
    .sum(net_sum1_22));
  AL_FADD comp1_3 (
    .a(net_a1_3),
    .b(net_a0_3),
    .c(net_cout1_2),
    .cout(net_cout1_3),
    .sum(net_sum1_3));
  AL_FADD comp1_4 (
    .a(net_a1_4),
    .b(net_a0_4),
    .c(net_cout1_3),
    .cout(net_cout1_4),
    .sum(net_sum1_4));
  AL_FADD comp1_5 (
    .a(net_a1_5),
    .b(net_a0_5),
    .c(net_cout1_4),
    .cout(net_cout1_5),
    .sum(net_sum1_5));
  AL_FADD comp1_6 (
    .a(net_a1_6),
    .b(net_a0_6),
    .c(net_cout1_5),
    .cout(net_cout1_6),
    .sum(net_sum1_6));
  AL_FADD comp1_7 (
    .a(net_a1_7),
    .b(net_a0_7),
    .c(net_cout1_6),
    .cout(net_cout1_7),
    .sum(net_sum1_7));
  AL_FADD comp1_8 (
    .a(net_a1_8),
    .b(net_a0_8),
    .c(net_cout1_7),
    .cout(net_cout1_8),
    .sum(net_sum1_8));
  AL_FADD comp1_9 (
    .a(net_a1_9),
    .b(net_a0_9),
    .c(net_cout1_8),
    .cout(net_cout1_9),
    .sum(net_sum1_9));
  AL_FADD comp2_0 (
    .a(net_a2_0),
    .b(net_sum1_0),
    .c(1'b0),
    .cout(net_cout2_0),
    .sum(net_sum2_0));
  AL_FADD comp2_1 (
    .a(net_a2_1),
    .b(net_sum1_1),
    .c(net_cout2_0),
    .cout(net_cout2_1),
    .sum(net_sum2_1));
  AL_FADD comp2_10 (
    .a(net_a2_10),
    .b(net_sum1_10),
    .c(net_cout2_9),
    .cout(net_cout2_10),
    .sum(net_sum2_10));
  AL_FADD comp2_11 (
    .a(net_a2_11),
    .b(net_sum1_11),
    .c(net_cout2_10),
    .cout(net_cout2_11),
    .sum(net_sum2_11));
  AL_FADD comp2_12 (
    .a(net_a2_12),
    .b(net_sum1_12),
    .c(net_cout2_11),
    .cout(net_cout2_12),
    .sum(net_sum2_12));
  AL_FADD comp2_13 (
    .a(net_a2_13),
    .b(net_sum1_13),
    .c(net_cout2_12),
    .cout(net_cout2_13),
    .sum(net_sum2_13));
  AL_FADD comp2_14 (
    .a(net_a2_14),
    .b(net_sum1_14),
    .c(net_cout2_13),
    .cout(net_cout2_14),
    .sum(net_sum2_14));
  AL_FADD comp2_15 (
    .a(net_a2_15),
    .b(net_sum1_15),
    .c(net_cout2_14),
    .cout(net_cout2_15),
    .sum(net_sum2_15));
  AL_FADD comp2_16 (
    .a(net_a2_16),
    .b(net_sum1_16),
    .c(net_cout2_15),
    .cout(net_cout2_16),
    .sum(net_sum2_16));
  AL_FADD comp2_17 (
    .a(net_a2_17),
    .b(net_sum1_17),
    .c(net_cout2_16),
    .cout(net_cout2_17),
    .sum(net_sum2_17));
  AL_FADD comp2_18 (
    .a(net_a2_18),
    .b(net_sum1_18),
    .c(net_cout2_17),
    .cout(net_cout2_18),
    .sum(net_sum2_18));
  AL_FADD comp2_19 (
    .a(net_a2_19),
    .b(net_sum1_19),
    .c(net_cout2_18),
    .cout(net_cout2_19),
    .sum(net_sum2_19));
  AL_FADD comp2_2 (
    .a(net_a2_2),
    .b(net_sum1_2),
    .c(net_cout2_1),
    .cout(net_cout2_2),
    .sum(net_sum2_2));
  AL_FADD comp2_20 (
    .a(net_a2_20),
    .b(net_sum1_20),
    .c(net_cout2_19),
    .cout(net_cout2_20),
    .sum(net_sum2_20));
  AL_FADD comp2_21 (
    .a(1'b0),
    .b(net_sum1_21),
    .c(net_cout2_20),
    .cout(net_cout2_21),
    .sum(net_sum2_21));
  AL_FADD comp2_22 (
    .a(1'b0),
    .b(net_sum1_22),
    .c(net_cout2_21),
    .cout(net_cout2_22),
    .sum(net_sum2_22));
  AL_FADD comp2_23 (
    .a(1'b0),
    .b(net_cout1_22),
    .c(net_cout2_22),
    .cout(net_cout2_23),
    .sum(net_sum2_23));
  AL_FADD comp2_3 (
    .a(net_a2_3),
    .b(net_sum1_3),
    .c(net_cout2_2),
    .cout(net_cout2_3),
    .sum(net_sum2_3));
  AL_FADD comp2_4 (
    .a(net_a2_4),
    .b(net_sum1_4),
    .c(net_cout2_3),
    .cout(net_cout2_4),
    .sum(net_sum2_4));
  AL_FADD comp2_5 (
    .a(net_a2_5),
    .b(net_sum1_5),
    .c(net_cout2_4),
    .cout(net_cout2_5),
    .sum(net_sum2_5));
  AL_FADD comp2_6 (
    .a(net_a2_6),
    .b(net_sum1_6),
    .c(net_cout2_5),
    .cout(net_cout2_6),
    .sum(net_sum2_6));
  AL_FADD comp2_7 (
    .a(net_a2_7),
    .b(net_sum1_7),
    .c(net_cout2_6),
    .cout(net_cout2_7),
    .sum(net_sum2_7));
  AL_FADD comp2_8 (
    .a(net_a2_8),
    .b(net_sum1_8),
    .c(net_cout2_7),
    .cout(net_cout2_8),
    .sum(net_sum2_8));
  AL_FADD comp2_9 (
    .a(net_a2_9),
    .b(net_sum1_9),
    .c(net_cout2_8),
    .cout(net_cout2_9),
    .sum(net_sum2_9));
  AL_FADD comp3_0 (
    .a(net_a3_0),
    .b(net_sum2_0),
    .c(1'b0),
    .cout(net_cout3_0),
    .sum(net_sum3_0));
  AL_FADD comp3_1 (
    .a(net_a3_1),
    .b(net_sum2_1),
    .c(net_cout3_0),
    .cout(net_cout3_1),
    .sum(net_sum3_1));
  AL_FADD comp3_10 (
    .a(net_a3_10),
    .b(net_sum2_10),
    .c(net_cout3_9),
    .cout(net_cout3_10),
    .sum(net_sum3_10));
  AL_FADD comp3_11 (
    .a(net_a3_11),
    .b(net_sum2_11),
    .c(net_cout3_10),
    .cout(net_cout3_11),
    .sum(net_sum3_11));
  AL_FADD comp3_12 (
    .a(net_a3_12),
    .b(net_sum2_12),
    .c(net_cout3_11),
    .cout(net_cout3_12),
    .sum(net_sum3_12));
  AL_FADD comp3_13 (
    .a(net_a3_13),
    .b(net_sum2_13),
    .c(net_cout3_12),
    .cout(net_cout3_13),
    .sum(net_sum3_13));
  AL_FADD comp3_14 (
    .a(net_a3_14),
    .b(net_sum2_14),
    .c(net_cout3_13),
    .cout(net_cout3_14),
    .sum(net_sum3_14));
  AL_FADD comp3_15 (
    .a(net_a3_15),
    .b(net_sum2_15),
    .c(net_cout3_14),
    .cout(net_cout3_15),
    .sum(net_sum3_15));
  AL_FADD comp3_16 (
    .a(net_a3_16),
    .b(net_sum2_16),
    .c(net_cout3_15),
    .cout(net_cout3_16),
    .sum(net_sum3_16));
  AL_FADD comp3_17 (
    .a(net_a3_17),
    .b(net_sum2_17),
    .c(net_cout3_16),
    .cout(net_cout3_17),
    .sum(net_sum3_17));
  AL_FADD comp3_18 (
    .a(net_a3_18),
    .b(net_sum2_18),
    .c(net_cout3_17),
    .cout(net_cout3_18),
    .sum(net_sum3_18));
  AL_FADD comp3_19 (
    .a(net_a3_19),
    .b(net_sum2_19),
    .c(net_cout3_18),
    .cout(net_cout3_19),
    .sum(net_sum3_19));
  AL_FADD comp3_2 (
    .a(net_a3_2),
    .b(net_sum2_2),
    .c(net_cout3_1),
    .cout(net_cout3_2),
    .sum(net_sum3_2));
  AL_FADD comp3_20 (
    .a(1'b0),
    .b(net_sum2_20),
    .c(net_cout3_19),
    .cout(net_cout3_20),
    .sum(net_sum3_20));
  AL_FADD comp3_21 (
    .a(1'b0),
    .b(net_sum2_21),
    .c(net_cout3_20),
    .cout(net_cout3_21),
    .sum(net_sum3_21));
  AL_FADD comp3_22 (
    .a(1'b0),
    .b(net_sum2_22),
    .c(net_cout3_21),
    .cout(net_cout3_22),
    .sum(net_sum3_22));
  AL_FADD comp3_23 (
    .a(1'b0),
    .b(net_sum2_23),
    .c(net_cout3_22),
    .cout(net_cout3_23),
    .sum(net_sum3_23));
  AL_FADD comp3_3 (
    .a(net_a3_3),
    .b(net_sum2_3),
    .c(net_cout3_2),
    .cout(net_cout3_3),
    .sum(net_sum3_3));
  AL_FADD comp3_4 (
    .a(net_a3_4),
    .b(net_sum2_4),
    .c(net_cout3_3),
    .cout(net_cout3_4),
    .sum(net_sum3_4));
  AL_FADD comp3_5 (
    .a(net_a3_5),
    .b(net_sum2_5),
    .c(net_cout3_4),
    .cout(net_cout3_5),
    .sum(net_sum3_5));
  AL_FADD comp3_6 (
    .a(net_a3_6),
    .b(net_sum2_6),
    .c(net_cout3_5),
    .cout(net_cout3_6),
    .sum(net_sum3_6));
  AL_FADD comp3_7 (
    .a(net_a3_7),
    .b(net_sum2_7),
    .c(net_cout3_6),
    .cout(net_cout3_7),
    .sum(net_sum3_7));
  AL_FADD comp3_8 (
    .a(net_a3_8),
    .b(net_sum2_8),
    .c(net_cout3_7),
    .cout(net_cout3_8),
    .sum(net_sum3_8));
  AL_FADD comp3_9 (
    .a(net_a3_9),
    .b(net_sum2_9),
    .c(net_cout3_8),
    .cout(net_cout3_9),
    .sum(net_sum3_9));
  AL_FADD comp4_0 (
    .a(net_a4_0),
    .b(net_sum3_0),
    .c(1'b0),
    .cout(net_cout4_0),
    .sum(net_sum4_0));
  AL_FADD comp4_1 (
    .a(net_a4_1),
    .b(net_sum3_1),
    .c(net_cout4_0),
    .cout(net_cout4_1),
    .sum(net_sum4_1));
  AL_FADD comp4_10 (
    .a(net_a4_10),
    .b(net_sum3_10),
    .c(net_cout4_9),
    .cout(net_cout4_10),
    .sum(net_sum4_10));
  AL_FADD comp4_11 (
    .a(net_a4_11),
    .b(net_sum3_11),
    .c(net_cout4_10),
    .cout(net_cout4_11),
    .sum(net_sum4_11));
  AL_FADD comp4_12 (
    .a(net_a4_12),
    .b(net_sum3_12),
    .c(net_cout4_11),
    .cout(net_cout4_12),
    .sum(net_sum4_12));
  AL_FADD comp4_13 (
    .a(net_a4_13),
    .b(net_sum3_13),
    .c(net_cout4_12),
    .cout(net_cout4_13),
    .sum(net_sum4_13));
  AL_FADD comp4_14 (
    .a(net_a4_14),
    .b(net_sum3_14),
    .c(net_cout4_13),
    .cout(net_cout4_14),
    .sum(net_sum4_14));
  AL_FADD comp4_15 (
    .a(net_a4_15),
    .b(net_sum3_15),
    .c(net_cout4_14),
    .cout(net_cout4_15),
    .sum(net_sum4_15));
  AL_FADD comp4_16 (
    .a(net_a4_16),
    .b(net_sum3_16),
    .c(net_cout4_15),
    .cout(net_cout4_16),
    .sum(net_sum4_16));
  AL_FADD comp4_17 (
    .a(net_a4_17),
    .b(net_sum3_17),
    .c(net_cout4_16),
    .cout(net_cout4_17),
    .sum(net_sum4_17));
  AL_FADD comp4_18 (
    .a(net_a4_18),
    .b(net_sum3_18),
    .c(net_cout4_17),
    .cout(net_cout4_18),
    .sum(net_sum4_18));
  AL_FADD comp4_19 (
    .a(1'b0),
    .b(net_sum3_19),
    .c(net_cout4_18),
    .cout(net_cout4_19),
    .sum(net_sum4_19));
  AL_FADD comp4_2 (
    .a(net_a4_2),
    .b(net_sum3_2),
    .c(net_cout4_1),
    .cout(net_cout4_2),
    .sum(net_sum4_2));
  AL_FADD comp4_20 (
    .a(1'b0),
    .b(net_sum3_20),
    .c(net_cout4_19),
    .cout(net_cout4_20),
    .sum(net_sum4_20));
  AL_FADD comp4_21 (
    .a(1'b0),
    .b(net_sum3_21),
    .c(net_cout4_20),
    .cout(net_cout4_21),
    .sum(net_sum4_21));
  AL_FADD comp4_22 (
    .a(1'b0),
    .b(net_sum3_22),
    .c(net_cout4_21),
    .cout(net_cout4_22),
    .sum(net_sum4_22));
  AL_FADD comp4_23 (
    .a(1'b0),
    .b(net_sum3_23),
    .c(net_cout4_22),
    .cout(net_cout4_23),
    .sum(net_sum4_23));
  AL_FADD comp4_3 (
    .a(net_a4_3),
    .b(net_sum3_3),
    .c(net_cout4_2),
    .cout(net_cout4_3),
    .sum(net_sum4_3));
  AL_FADD comp4_4 (
    .a(net_a4_4),
    .b(net_sum3_4),
    .c(net_cout4_3),
    .cout(net_cout4_4),
    .sum(net_sum4_4));
  AL_FADD comp4_5 (
    .a(net_a4_5),
    .b(net_sum3_5),
    .c(net_cout4_4),
    .cout(net_cout4_5),
    .sum(net_sum4_5));
  AL_FADD comp4_6 (
    .a(net_a4_6),
    .b(net_sum3_6),
    .c(net_cout4_5),
    .cout(net_cout4_6),
    .sum(net_sum4_6));
  AL_FADD comp4_7 (
    .a(net_a4_7),
    .b(net_sum3_7),
    .c(net_cout4_6),
    .cout(net_cout4_7),
    .sum(net_sum4_7));
  AL_FADD comp4_8 (
    .a(net_a4_8),
    .b(net_sum3_8),
    .c(net_cout4_7),
    .cout(net_cout4_8),
    .sum(net_sum4_8));
  AL_FADD comp4_9 (
    .a(net_a4_9),
    .b(net_sum3_9),
    .c(net_cout4_8),
    .cout(net_cout4_9),
    .sum(net_sum4_9));
  AL_FADD comp5_0 (
    .a(net_a5_0),
    .b(net_sum4_0),
    .c(1'b0),
    .cout(net_cout5_0),
    .sum(net_sum5_0));
  AL_FADD comp5_1 (
    .a(net_a5_1),
    .b(net_sum4_1),
    .c(net_cout5_0),
    .cout(net_cout5_1),
    .sum(net_sum5_1));
  AL_FADD comp5_10 (
    .a(net_a5_10),
    .b(net_sum4_10),
    .c(net_cout5_9),
    .cout(net_cout5_10),
    .sum(net_sum5_10));
  AL_FADD comp5_11 (
    .a(net_a5_11),
    .b(net_sum4_11),
    .c(net_cout5_10),
    .cout(net_cout5_11),
    .sum(net_sum5_11));
  AL_FADD comp5_12 (
    .a(net_a5_12),
    .b(net_sum4_12),
    .c(net_cout5_11),
    .cout(net_cout5_12),
    .sum(net_sum5_12));
  AL_FADD comp5_13 (
    .a(net_a5_13),
    .b(net_sum4_13),
    .c(net_cout5_12),
    .cout(net_cout5_13),
    .sum(net_sum5_13));
  AL_FADD comp5_14 (
    .a(net_a5_14),
    .b(net_sum4_14),
    .c(net_cout5_13),
    .cout(net_cout5_14),
    .sum(net_sum5_14));
  AL_FADD comp5_15 (
    .a(net_a5_15),
    .b(net_sum4_15),
    .c(net_cout5_14),
    .cout(net_cout5_15),
    .sum(net_sum5_15));
  AL_FADD comp5_16 (
    .a(net_a5_16),
    .b(net_sum4_16),
    .c(net_cout5_15),
    .cout(net_cout5_16),
    .sum(net_sum5_16));
  AL_FADD comp5_17 (
    .a(net_a5_17),
    .b(net_sum4_17),
    .c(net_cout5_16),
    .cout(net_cout5_17),
    .sum(net_sum5_17));
  AL_FADD comp5_18 (
    .a(1'b0),
    .b(net_sum4_18),
    .c(net_cout5_17),
    .cout(net_cout5_18),
    .sum(net_sum5_18));
  AL_FADD comp5_19 (
    .a(1'b0),
    .b(net_sum4_19),
    .c(net_cout5_18),
    .cout(net_cout5_19),
    .sum(net_sum5_19));
  AL_FADD comp5_2 (
    .a(net_a5_2),
    .b(net_sum4_2),
    .c(net_cout5_1),
    .cout(net_cout5_2),
    .sum(net_sum5_2));
  AL_FADD comp5_20 (
    .a(1'b0),
    .b(net_sum4_20),
    .c(net_cout5_19),
    .cout(net_cout5_20),
    .sum(net_sum5_20));
  AL_FADD comp5_21 (
    .a(1'b0),
    .b(net_sum4_21),
    .c(net_cout5_20),
    .cout(net_cout5_21),
    .sum(net_sum5_21));
  AL_FADD comp5_22 (
    .a(1'b0),
    .b(net_sum4_22),
    .c(net_cout5_21),
    .cout(net_cout5_22),
    .sum(net_sum5_22));
  AL_FADD comp5_23 (
    .a(1'b0),
    .b(net_sum4_23),
    .c(net_cout5_22),
    .cout(net_cout5_23),
    .sum(net_sum5_23));
  AL_FADD comp5_3 (
    .a(net_a5_3),
    .b(net_sum4_3),
    .c(net_cout5_2),
    .cout(net_cout5_3),
    .sum(net_sum5_3));
  AL_FADD comp5_4 (
    .a(net_a5_4),
    .b(net_sum4_4),
    .c(net_cout5_3),
    .cout(net_cout5_4),
    .sum(net_sum5_4));
  AL_FADD comp5_5 (
    .a(net_a5_5),
    .b(net_sum4_5),
    .c(net_cout5_4),
    .cout(net_cout5_5),
    .sum(net_sum5_5));
  AL_FADD comp5_6 (
    .a(net_a5_6),
    .b(net_sum4_6),
    .c(net_cout5_5),
    .cout(net_cout5_6),
    .sum(net_sum5_6));
  AL_FADD comp5_7 (
    .a(net_a5_7),
    .b(net_sum4_7),
    .c(net_cout5_6),
    .cout(net_cout5_7),
    .sum(net_sum5_7));
  AL_FADD comp5_8 (
    .a(net_a5_8),
    .b(net_sum4_8),
    .c(net_cout5_7),
    .cout(net_cout5_8),
    .sum(net_sum5_8));
  AL_FADD comp5_9 (
    .a(net_a5_9),
    .b(net_sum4_9),
    .c(net_cout5_8),
    .cout(net_cout5_9),
    .sum(net_sum5_9));
  AL_FADD comp6_0 (
    .a(net_a6_0),
    .b(net_sum5_0),
    .c(1'b0),
    .cout(net_cout6_0),
    .sum(net_sum6_0));
  AL_FADD comp6_1 (
    .a(net_a6_1),
    .b(net_sum5_1),
    .c(net_cout6_0),
    .cout(net_cout6_1),
    .sum(net_sum6_1));
  AL_FADD comp6_10 (
    .a(net_a6_10),
    .b(net_sum5_10),
    .c(net_cout6_9),
    .cout(net_cout6_10),
    .sum(net_sum6_10));
  AL_FADD comp6_11 (
    .a(net_a6_11),
    .b(net_sum5_11),
    .c(net_cout6_10),
    .cout(net_cout6_11),
    .sum(net_sum6_11));
  AL_FADD comp6_12 (
    .a(net_a6_12),
    .b(net_sum5_12),
    .c(net_cout6_11),
    .cout(net_cout6_12),
    .sum(net_sum6_12));
  AL_FADD comp6_13 (
    .a(net_a6_13),
    .b(net_sum5_13),
    .c(net_cout6_12),
    .cout(net_cout6_13),
    .sum(net_sum6_13));
  AL_FADD comp6_14 (
    .a(net_a6_14),
    .b(net_sum5_14),
    .c(net_cout6_13),
    .cout(net_cout6_14),
    .sum(net_sum6_14));
  AL_FADD comp6_15 (
    .a(net_a6_15),
    .b(net_sum5_15),
    .c(net_cout6_14),
    .cout(net_cout6_15),
    .sum(net_sum6_15));
  AL_FADD comp6_16 (
    .a(net_a6_16),
    .b(net_sum5_16),
    .c(net_cout6_15),
    .cout(net_cout6_16),
    .sum(net_sum6_16));
  AL_FADD comp6_17 (
    .a(1'b0),
    .b(net_sum5_17),
    .c(net_cout6_16),
    .cout(net_cout6_17),
    .sum(net_sum6_17));
  AL_FADD comp6_18 (
    .a(1'b0),
    .b(net_sum5_18),
    .c(net_cout6_17),
    .cout(net_cout6_18),
    .sum(net_sum6_18));
  AL_FADD comp6_19 (
    .a(1'b0),
    .b(net_sum5_19),
    .c(net_cout6_18),
    .cout(net_cout6_19),
    .sum(net_sum6_19));
  AL_FADD comp6_2 (
    .a(net_a6_2),
    .b(net_sum5_2),
    .c(net_cout6_1),
    .cout(net_cout6_2),
    .sum(net_sum6_2));
  AL_FADD comp6_20 (
    .a(1'b0),
    .b(net_sum5_20),
    .c(net_cout6_19),
    .cout(net_cout6_20),
    .sum(net_sum6_20));
  AL_FADD comp6_21 (
    .a(1'b0),
    .b(net_sum5_21),
    .c(net_cout6_20),
    .cout(net_cout6_21),
    .sum(net_sum6_21));
  AL_FADD comp6_22 (
    .a(1'b0),
    .b(net_sum5_22),
    .c(net_cout6_21),
    .cout(net_cout6_22),
    .sum(net_sum6_22));
  AL_FADD comp6_23 (
    .a(1'b0),
    .b(net_sum5_23),
    .c(net_cout6_22),
    .cout(net_cout6_23),
    .sum(net_sum6_23));
  AL_FADD comp6_3 (
    .a(net_a6_3),
    .b(net_sum5_3),
    .c(net_cout6_2),
    .cout(net_cout6_3),
    .sum(net_sum6_3));
  AL_FADD comp6_4 (
    .a(net_a6_4),
    .b(net_sum5_4),
    .c(net_cout6_3),
    .cout(net_cout6_4),
    .sum(net_sum6_4));
  AL_FADD comp6_5 (
    .a(net_a6_5),
    .b(net_sum5_5),
    .c(net_cout6_4),
    .cout(net_cout6_5),
    .sum(net_sum6_5));
  AL_FADD comp6_6 (
    .a(net_a6_6),
    .b(net_sum5_6),
    .c(net_cout6_5),
    .cout(net_cout6_6),
    .sum(net_sum6_6));
  AL_FADD comp6_7 (
    .a(net_a6_7),
    .b(net_sum5_7),
    .c(net_cout6_6),
    .cout(net_cout6_7),
    .sum(net_sum6_7));
  AL_FADD comp6_8 (
    .a(net_a6_8),
    .b(net_sum5_8),
    .c(net_cout6_7),
    .cout(net_cout6_8),
    .sum(net_sum6_8));
  AL_FADD comp6_9 (
    .a(net_a6_9),
    .b(net_sum5_9),
    .c(net_cout6_8),
    .cout(net_cout6_9),
    .sum(net_sum6_9));
  AL_FADD comp7_0 (
    .a(net_a7_0),
    .b(net_sum6_0),
    .c(1'b0),
    .cout(net_cout7_0),
    .sum(net_sum7_0));
  AL_FADD comp7_1 (
    .a(net_a7_1),
    .b(net_sum6_1),
    .c(net_cout7_0),
    .cout(net_cout7_1),
    .sum(net_sum7_1));
  AL_FADD comp7_10 (
    .a(net_a7_10),
    .b(net_sum6_10),
    .c(net_cout7_9),
    .cout(net_cout7_10),
    .sum(net_sum7_10));
  AL_FADD comp7_11 (
    .a(net_a7_11),
    .b(net_sum6_11),
    .c(net_cout7_10),
    .cout(net_cout7_11),
    .sum(net_sum7_11));
  AL_FADD comp7_12 (
    .a(net_a7_12),
    .b(net_sum6_12),
    .c(net_cout7_11),
    .cout(net_cout7_12),
    .sum(net_sum7_12));
  AL_FADD comp7_13 (
    .a(net_a7_13),
    .b(net_sum6_13),
    .c(net_cout7_12),
    .cout(net_cout7_13),
    .sum(net_sum7_13));
  AL_FADD comp7_14 (
    .a(net_a7_14),
    .b(net_sum6_14),
    .c(net_cout7_13),
    .cout(net_cout7_14),
    .sum(net_sum7_14));
  AL_FADD comp7_15 (
    .a(net_a7_15),
    .b(net_sum6_15),
    .c(net_cout7_14),
    .cout(net_cout7_15),
    .sum(net_sum7_15));
  AL_FADD comp7_16 (
    .a(1'b0),
    .b(net_sum6_16),
    .c(net_cout7_15),
    .cout(net_cout7_16),
    .sum(net_sum7_16));
  AL_FADD comp7_17 (
    .a(1'b0),
    .b(net_sum6_17),
    .c(net_cout7_16),
    .cout(net_cout7_17),
    .sum(net_sum7_17));
  AL_FADD comp7_18 (
    .a(1'b0),
    .b(net_sum6_18),
    .c(net_cout7_17),
    .cout(net_cout7_18),
    .sum(net_sum7_18));
  AL_FADD comp7_19 (
    .a(1'b0),
    .b(net_sum6_19),
    .c(net_cout7_18),
    .cout(net_cout7_19),
    .sum(net_sum7_19));
  AL_FADD comp7_2 (
    .a(net_a7_2),
    .b(net_sum6_2),
    .c(net_cout7_1),
    .cout(net_cout7_2),
    .sum(net_sum7_2));
  AL_FADD comp7_20 (
    .a(1'b0),
    .b(net_sum6_20),
    .c(net_cout7_19),
    .cout(net_cout7_20),
    .sum(net_sum7_20));
  AL_FADD comp7_21 (
    .a(1'b0),
    .b(net_sum6_21),
    .c(net_cout7_20),
    .cout(net_cout7_21),
    .sum(net_sum7_21));
  AL_FADD comp7_22 (
    .a(1'b0),
    .b(net_sum6_22),
    .c(net_cout7_21),
    .cout(net_cout7_22),
    .sum(net_sum7_22));
  AL_FADD comp7_23 (
    .a(1'b0),
    .b(net_sum6_23),
    .c(net_cout7_22),
    .cout(net_cout7_23),
    .sum(net_sum7_23));
  AL_FADD comp7_3 (
    .a(net_a7_3),
    .b(net_sum6_3),
    .c(net_cout7_2),
    .cout(net_cout7_3),
    .sum(net_sum7_3));
  AL_FADD comp7_4 (
    .a(net_a7_4),
    .b(net_sum6_4),
    .c(net_cout7_3),
    .cout(net_cout7_4),
    .sum(net_sum7_4));
  AL_FADD comp7_5 (
    .a(net_a7_5),
    .b(net_sum6_5),
    .c(net_cout7_4),
    .cout(net_cout7_5),
    .sum(net_sum7_5));
  AL_FADD comp7_6 (
    .a(net_a7_6),
    .b(net_sum6_6),
    .c(net_cout7_5),
    .cout(net_cout7_6),
    .sum(net_sum7_6));
  AL_FADD comp7_7 (
    .a(net_a7_7),
    .b(net_sum6_7),
    .c(net_cout7_6),
    .cout(net_cout7_7),
    .sum(net_sum7_7));
  AL_FADD comp7_8 (
    .a(net_a7_8),
    .b(net_sum6_8),
    .c(net_cout7_7),
    .cout(net_cout7_8),
    .sum(net_sum7_8));
  AL_FADD comp7_9 (
    .a(net_a7_9),
    .b(net_sum6_9),
    .c(net_cout7_8),
    .cout(net_cout7_9),
    .sum(net_sum7_9));
  AL_FADD comp8_0 (
    .a(net_a8_0),
    .b(net_sum7_0),
    .c(1'b0),
    .cout(net_cout8_0),
    .sum(net_sum8_0));
  AL_FADD comp8_1 (
    .a(net_a8_1),
    .b(net_sum7_1),
    .c(net_cout8_0),
    .cout(net_cout8_1),
    .sum(net_sum8_1));
  AL_FADD comp8_10 (
    .a(net_a8_10),
    .b(net_sum7_10),
    .c(net_cout8_9),
    .cout(net_cout8_10),
    .sum(net_sum8_10));
  AL_FADD comp8_11 (
    .a(net_a8_11),
    .b(net_sum7_11),
    .c(net_cout8_10),
    .cout(net_cout8_11),
    .sum(net_sum8_11));
  AL_FADD comp8_12 (
    .a(net_a8_12),
    .b(net_sum7_12),
    .c(net_cout8_11),
    .cout(net_cout8_12),
    .sum(net_sum8_12));
  AL_FADD comp8_13 (
    .a(net_a8_13),
    .b(net_sum7_13),
    .c(net_cout8_12),
    .cout(net_cout8_13),
    .sum(net_sum8_13));
  AL_FADD comp8_14 (
    .a(net_a8_14),
    .b(net_sum7_14),
    .c(net_cout8_13),
    .cout(net_cout8_14),
    .sum(net_sum8_14));
  AL_FADD comp8_15 (
    .a(1'b0),
    .b(net_sum7_15),
    .c(net_cout8_14),
    .cout(net_cout8_15),
    .sum(net_sum8_15));
  AL_FADD comp8_16 (
    .a(1'b0),
    .b(net_sum7_16),
    .c(net_cout8_15),
    .cout(net_cout8_16),
    .sum(net_sum8_16));
  AL_FADD comp8_17 (
    .a(1'b0),
    .b(net_sum7_17),
    .c(net_cout8_16),
    .cout(net_cout8_17),
    .sum(net_sum8_17));
  AL_FADD comp8_18 (
    .a(1'b0),
    .b(net_sum7_18),
    .c(net_cout8_17),
    .cout(net_cout8_18),
    .sum(net_sum8_18));
  AL_FADD comp8_19 (
    .a(1'b0),
    .b(net_sum7_19),
    .c(net_cout8_18),
    .cout(net_cout8_19),
    .sum(net_sum8_19));
  AL_FADD comp8_2 (
    .a(net_a8_2),
    .b(net_sum7_2),
    .c(net_cout8_1),
    .cout(net_cout8_2),
    .sum(net_sum8_2));
  AL_FADD comp8_20 (
    .a(1'b0),
    .b(net_sum7_20),
    .c(net_cout8_19),
    .cout(net_cout8_20),
    .sum(net_sum8_20));
  AL_FADD comp8_21 (
    .a(1'b0),
    .b(net_sum7_21),
    .c(net_cout8_20),
    .cout(net_cout8_21),
    .sum(net_sum8_21));
  AL_FADD comp8_22 (
    .a(1'b0),
    .b(net_sum7_22),
    .c(net_cout8_21),
    .cout(net_cout8_22),
    .sum(net_sum8_22));
  AL_FADD comp8_23 (
    .a(1'b0),
    .b(net_sum7_23),
    .c(net_cout8_22),
    .cout(net_cout8_23),
    .sum(net_sum8_23));
  AL_FADD comp8_3 (
    .a(net_a8_3),
    .b(net_sum7_3),
    .c(net_cout8_2),
    .cout(net_cout8_3),
    .sum(net_sum8_3));
  AL_FADD comp8_4 (
    .a(net_a8_4),
    .b(net_sum7_4),
    .c(net_cout8_3),
    .cout(net_cout8_4),
    .sum(net_sum8_4));
  AL_FADD comp8_5 (
    .a(net_a8_5),
    .b(net_sum7_5),
    .c(net_cout8_4),
    .cout(net_cout8_5),
    .sum(net_sum8_5));
  AL_FADD comp8_6 (
    .a(net_a8_6),
    .b(net_sum7_6),
    .c(net_cout8_5),
    .cout(net_cout8_6),
    .sum(net_sum8_6));
  AL_FADD comp8_7 (
    .a(net_a8_7),
    .b(net_sum7_7),
    .c(net_cout8_6),
    .cout(net_cout8_7),
    .sum(net_sum8_7));
  AL_FADD comp8_8 (
    .a(net_a8_8),
    .b(net_sum7_8),
    .c(net_cout8_7),
    .cout(net_cout8_8),
    .sum(net_sum8_8));
  AL_FADD comp8_9 (
    .a(net_a8_9),
    .b(net_sum7_9),
    .c(net_cout8_8),
    .cout(net_cout8_9),
    .sum(net_sum8_9));
  AL_FADD comp9_0 (
    .a(net_a9_0),
    .b(net_sum8_0),
    .c(1'b0),
    .cout(net_cout9_0),
    .sum(net_sum9_0));
  AL_FADD comp9_1 (
    .a(net_a9_1),
    .b(net_sum8_1),
    .c(net_cout9_0),
    .cout(net_cout9_1),
    .sum(net_sum9_1));
  AL_FADD comp9_10 (
    .a(net_a9_10),
    .b(net_sum8_10),
    .c(net_cout9_9),
    .cout(net_cout9_10),
    .sum(net_sum9_10));
  AL_FADD comp9_11 (
    .a(net_a9_11),
    .b(net_sum8_11),
    .c(net_cout9_10),
    .cout(net_cout9_11),
    .sum(net_sum9_11));
  AL_FADD comp9_12 (
    .a(net_a9_12),
    .b(net_sum8_12),
    .c(net_cout9_11),
    .cout(net_cout9_12),
    .sum(net_sum9_12));
  AL_FADD comp9_13 (
    .a(net_a9_13),
    .b(net_sum8_13),
    .c(net_cout9_12),
    .cout(net_cout9_13),
    .sum(net_sum9_13));
  AL_FADD comp9_14 (
    .a(1'b0),
    .b(net_sum8_14),
    .c(net_cout9_13),
    .cout(net_cout9_14),
    .sum(net_sum9_14));
  AL_FADD comp9_15 (
    .a(1'b0),
    .b(net_sum8_15),
    .c(net_cout9_14),
    .cout(net_cout9_15),
    .sum(net_sum9_15));
  AL_FADD comp9_16 (
    .a(1'b0),
    .b(net_sum8_16),
    .c(net_cout9_15),
    .cout(net_cout9_16),
    .sum(net_sum9_16));
  AL_FADD comp9_17 (
    .a(1'b0),
    .b(net_sum8_17),
    .c(net_cout9_16),
    .cout(net_cout9_17),
    .sum(net_sum9_17));
  AL_FADD comp9_18 (
    .a(1'b0),
    .b(net_sum8_18),
    .c(net_cout9_17),
    .cout(net_cout9_18),
    .sum(net_sum9_18));
  AL_FADD comp9_19 (
    .a(1'b0),
    .b(net_sum8_19),
    .c(net_cout9_18),
    .cout(net_cout9_19),
    .sum(net_sum9_19));
  AL_FADD comp9_2 (
    .a(net_a9_2),
    .b(net_sum8_2),
    .c(net_cout9_1),
    .cout(net_cout9_2),
    .sum(net_sum9_2));
  AL_FADD comp9_20 (
    .a(1'b0),
    .b(net_sum8_20),
    .c(net_cout9_19),
    .cout(net_cout9_20),
    .sum(net_sum9_20));
  AL_FADD comp9_21 (
    .a(1'b0),
    .b(net_sum8_21),
    .c(net_cout9_20),
    .cout(net_cout9_21),
    .sum(net_sum9_21));
  AL_FADD comp9_22 (
    .a(1'b0),
    .b(net_sum8_22),
    .c(net_cout9_21),
    .cout(net_cout9_22),
    .sum(net_sum9_22));
  AL_FADD comp9_23 (
    .a(1'b0),
    .b(net_sum8_23),
    .c(net_cout9_22),
    .cout(net_cout9_23),
    .sum(net_sum9_23));
  AL_FADD comp9_3 (
    .a(net_a9_3),
    .b(net_sum8_3),
    .c(net_cout9_2),
    .cout(net_cout9_3),
    .sum(net_sum9_3));
  AL_FADD comp9_4 (
    .a(net_a9_4),
    .b(net_sum8_4),
    .c(net_cout9_3),
    .cout(net_cout9_4),
    .sum(net_sum9_4));
  AL_FADD comp9_5 (
    .a(net_a9_5),
    .b(net_sum8_5),
    .c(net_cout9_4),
    .cout(net_cout9_5),
    .sum(net_sum9_5));
  AL_FADD comp9_6 (
    .a(net_a9_6),
    .b(net_sum8_6),
    .c(net_cout9_5),
    .cout(net_cout9_6),
    .sum(net_sum9_6));
  AL_FADD comp9_7 (
    .a(net_a9_7),
    .b(net_sum8_7),
    .c(net_cout9_6),
    .cout(net_cout9_7),
    .sum(net_sum9_7));
  AL_FADD comp9_8 (
    .a(net_a9_8),
    .b(net_sum8_8),
    .c(net_cout9_7),
    .cout(net_cout9_8),
    .sum(net_sum9_8));
  AL_FADD comp9_9 (
    .a(net_a9_9),
    .b(net_sum8_9),
    .c(net_cout9_8),
    .cout(net_cout9_9),
    .sum(net_sum9_9));

endmodule 

module AL_MUX
  (
  input i0,
  input i1,
  input sel,
  output o
  );

  wire not_sel, sel_i0, sel_i1;
  not u0 (not_sel, sel);
  and u1 (sel_i1, sel, i1);
  and u2 (sel_i0, not_sel, i0);
  or u3 (o, sel_i1, sel_i0);

endmodule

module AL_DFF
  (
  input reset,
  input set,
  input clk,
  input d,
  output reg q
  );

  parameter INI = 1'b0;

  tri0 gsrn = glbl.gsrn;

  always @(gsrn)
  begin
    if(!gsrn)
      assign q = INI;
    else
      deassign q;
  end

  always @(posedge reset or posedge set or posedge clk)
  begin
    if (reset)
      q <= 1'b0;
    else if (set)
      q <= 1'b1;
    else
      q <= d;
  end

endmodule

module AL_FADD
  (
  input a,
  input b,
  input c,
  output sum,
  output cout
  );

  wire prop;
  wire not_prop;
  wire sel_i0;
  wire sel_i1;

  xor u0 (prop, a, b);
  xor u1 (sum, prop, c);
  not u2 (not_prop, prop);
  and u3 (sel_i1, prop, c);
  and u4 (sel_i0, not_prop, a);
  or  u5 (cout, sel_i0, sel_i1);

endmodule

