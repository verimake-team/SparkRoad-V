// Verilog netlist created by TD v4.5.12562
// Mon Sep 30 17:08:18 2019

`timescale 1ns / 1ps
module M0demo  // ../RTL/M0demo.v(4)
  (
  NRST,
  SWCLKTCK,
  TDI,
  XTAL1,
  nTRST,
  uart0_rxd,
  P0,
  TDO,
  XTAL2,
  uart0_txd,
  uart0_txen,
  SWDIOTMS,
  b_pad_gpio_porta
  );

  input NRST;  // ../RTL/M0demo.v(7)
  input SWCLKTCK;  // ../RTL/M0demo.v(15)
  input TDI;  // ../RTL/M0demo.v(12)
  input XTAL1;  // ../RTL/M0demo.v(5)
  input nTRST;  // ../RTL/M0demo.v(11)
  input uart0_rxd;  // ../RTL/M0demo.v(19)
  output [15:0] P0;  // ../RTL/M0demo.v(8)
  output TDO;  // ../RTL/M0demo.v(13)
  output XTAL2;  // ../RTL/M0demo.v(6)
  output uart0_txd;  // ../RTL/M0demo.v(20)
  output uart0_txen;  // ../RTL/M0demo.v(21)
  inout SWDIOTMS;  // ../RTL/M0demo.v(14)
  inout [7:0] b_pad_gpio_porta;  // ../RTL/M0demo.v(17)

  parameter BE = 0;
  parameter BKPT = 4;
  parameter DBG = 1;
  parameter NUMIRQ = 32;
  parameter SMUL = 0;
  parameter SYST = 1;
  parameter WIC = 1;
  parameter WICLINES = 34;
  parameter WPT = 2;
  wire XTAL1_wire;  // ../RTL/M0demo.v(25)

  M0clkpll u_M0clkpll (
    .refclk(XTAL1),
    .clk0_out(XTAL1_wire));  // ../RTL/M0demo.v(74)
  \cmsdk_mcu(WIC=1)  u_cmsdk_mcu (
    .NRST(NRST),
    .TCK(SWCLKTCK),
    .TDI(TDI),
    .XTAL1(XTAL1_wire),
    .nTRST(nTRST),
    .uart0_rxd(uart0_rxd),
    .TDO(TDO),
    .XTAL2(XTAL2),
    .uart0_txd(uart0_txd),
    .uart0_txen(uart0_txen),
    .P0(P0),
    .TMS(SWDIOTMS),
    .b_pad_gpio_porta(b_pad_gpio_porta));  // ../RTL/M0demo.v(53)

endmodule 

module M0clkpll  // al_ip/M0clkpll.v(22)
  (
  refclk,
  reset,
  stdby,
  clk0_out,
  extlock
  );

  input refclk;  // al_ip/M0clkpll.v(28)
  input reset;  // al_ip/M0clkpll.v(29)
  input stdby;  // al_ip/M0clkpll.v(30)
  output clk0_out;  // al_ip/M0clkpll.v(32)
  output extlock;  // al_ip/M0clkpll.v(31)

  wire clk0_buf;  // al_ip/M0clkpll.v(34)

  EG_LOGIC_BUFG bufg_feedback (
    .i(clk0_buf),
    .o(clk0_out));  // al_ip/M0clkpll.v(36)
  EG_PHY_PLL #(
    .CLKC0_CPHASE(124),
    .CLKC0_DIV(125),
    .CLKC0_DIV2_ENABLE("DISABLE"),
    .CLKC0_ENABLE("ENABLE"),
    .CLKC0_FPHASE(0),
    .CLKC1_CPHASE(1),
    .CLKC1_DIV(1),
    .CLKC1_DIV2_ENABLE("DISABLE"),
    .CLKC1_ENABLE("DISABLE"),
    .CLKC1_FPHASE(0),
    .CLKC2_CPHASE(1),
    .CLKC2_DIV(1),
    .CLKC2_DIV2_ENABLE("DISABLE"),
    .CLKC2_ENABLE("DISABLE"),
    .CLKC2_FPHASE(0),
    .CLKC3_CPHASE(1),
    .CLKC3_DIV(1),
    .CLKC3_DIV2_ENABLE("DISABLE"),
    .CLKC3_ENABLE("DISABLE"),
    .CLKC3_FPHASE(0),
    .CLKC4_CPHASE(1),
    .CLKC4_DIV(1),
    .CLKC4_DIV2_ENABLE("DISABLE"),
    .CLKC4_ENABLE("DISABLE"),
    .CLKC4_FPHASE(0),
    .DERIVE_PLL_CLOCKS("DISABLE"),
    .DPHASE_SOURCE("DISABLE"),
    .DYNCFG("DISABLE"),
    .FBCLK_DIV(1),
    .FEEDBK_MODE("NORMAL"),
    .FEEDBK_PATH("CLKC0_EXT"),
    .FIN("24.000"),
    .FREQ_LOCK_ACCURACY(2),
    .GEN_BASIC_CLOCK("DISABLE"),
    .GMC_GAIN(6),
    .GMC_TEST(14),
    .ICP_CURRENT(3),
    .IF_ESCLKSTSW("DISABLE"),
    .INTFB_WAKE("DISABLE"),
    .KVCO(6),
    .LPF_CAPACITOR(3),
    .LPF_RESISTOR(2),
    .NORESET("DISABLE"),
    .ODIV_MUXC0("DIV"),
    .ODIV_MUXC1("DIV"),
    .ODIV_MUXC2("DIV"),
    .ODIV_MUXC3("DIV"),
    .ODIV_MUXC4("DIV"),
    .PLLC2RST_ENA("DISABLE"),
    .PLLC34RST_ENA("DISABLE"),
    .PLLMRST_ENA("DISABLE"),
    .PLLRST_ENA("ENABLE"),
    .PLL_LOCK_MODE(0),
    .PREDIV_MUXC0("VCO"),
    .PREDIV_MUXC1("VCO"),
    .PREDIV_MUXC2("VCO"),
    .PREDIV_MUXC3("VCO"),
    .PREDIV_MUXC4("VCO"),
    .REFCLK_DIV(3),
    .REFCLK_SEL("INTERNAL"),
    .STDBY_ENABLE("ENABLE"),
    .STDBY_VCO_ENA("DISABLE"),
    .SYNC_ENABLE("DISABLE"),
    .VCO_NORESET("DISABLE"))
    pll_inst (
    .daddr(6'b000000),
    .dclk(1'b0),
    .dcs(1'b0),
    .di(8'b00000000),
    .dwe(1'b0),
    .fbclk(clk0_out),
    .psclk(1'b0),
    .psclksel(3'b000),
    .psdown(1'b0),
    .psstep(1'b0),
    .refclk(refclk),
    .reset(reset),
    .stdby(stdby),
    .clkc({open_n0,open_n1,open_n2,open_n3,clk0_buf}),
    .extlock(extlock));  // al_ip/M0clkpll.v(59)

endmodule 

module \cmsdk_mcu(WIC=1)   // ../RTL/cmsdk_mcu.v(32)
  (
  NRST,
  SWCLKTCK,
  TCK,
  TDI,
  XTAL1,
  nTRST,
  uart0_rxd,
  TDO,
  XTAL2,
  uart0_txd,
  uart0_txen,
  P0,
  P1,
  SWDIOTMS,
  TMS,
  b_pad_gpio_porta
  );

  input NRST;  // ../RTL/cmsdk_mcu.v(50)
  input SWCLKTCK;  // ../RTL/cmsdk_mcu.v(60)
  input TCK;  // ../RTL/cmsdk_mcu.v(58)
  input TDI;  // ../RTL/cmsdk_mcu.v(55)
  input XTAL1;  // ../RTL/cmsdk_mcu.v(48)
  input nTRST;  // ../RTL/cmsdk_mcu.v(54)
  input uart0_rxd;  // ../RTL/cmsdk_mcu.v(66)
  output TDO;  // ../RTL/cmsdk_mcu.v(56)
  output XTAL2;  // ../RTL/cmsdk_mcu.v(49)
  output uart0_txd;  // ../RTL/cmsdk_mcu.v(67)
  output uart0_txen;  // ../RTL/cmsdk_mcu.v(68)
  inout [15:0] P0;  // ../RTL/cmsdk_mcu.v(51)
  inout [15:0] P1;  // ../RTL/cmsdk_mcu.v(52)
  inout SWDIOTMS;  // ../RTL/cmsdk_mcu.v(59)
  inout TMS;  // ../RTL/cmsdk_mcu.v(57)
  inout [7:0] b_pad_gpio_porta;  // ../RTL/cmsdk_mcu.v(64)

  parameter BE = 0;
  parameter BKPT = 4;
  parameter DBG = 1;
  parameter NUMIRQ = 32;
  parameter SMUL = 0;
  parameter SYST = 1;
  parameter WIC = 1;
  parameter WICLINES = 34;
  parameter WPT = 2;
  // localparam BASEADDR_GPIO0 = 32'b01000000000000010000000000000000;
  // localparam BASEADDR_GPIO1 = 32'b01000000000000010001000000000000;
  // localparam BASEADDR_SYSROMTABLE = 32'b11110000000000000000000000000000;
  wire [31:0] HADDR;  // ../RTL/cmsdk_mcu.v(103)
  wire [2:0] HSIZE;  // ../RTL/cmsdk_mcu.v(105)
  wire [1:0] HTRANS;  // ../RTL/cmsdk_mcu.v(104)
  wire [31:0] HWDATA;  // ../RTL/cmsdk_mcu.v(107)
  wire [31:0] flash_hrdata;  // ../RTL/cmsdk_mcu.v(113)
  wire [15:0] p0_altfunc;  // ../RTL/cmsdk_mcu.v(140)
  wire [15:0] p0_in;  // ../RTL/cmsdk_mcu.v(137)
  wire [15:0] p0_out;  // ../RTL/cmsdk_mcu.v(138)
  wire [15:0] p0_outen;  // ../RTL/cmsdk_mcu.v(139)
  wire [15:0] p1_altfunc;  // ../RTL/cmsdk_mcu.v(145)
  wire [15:0] p1_in;  // ../RTL/cmsdk_mcu.v(142)
  wire [15:0] p1_out;  // ../RTL/cmsdk_mcu.v(143)
  wire [15:0] p1_outen;  // ../RTL/cmsdk_mcu.v(144)
  wire [31:0] sram_hrdata;  // ../RTL/cmsdk_mcu.v(119)
  wire APBACTIVE;  // ../RTL/cmsdk_mcu.v(77)
  wire DBGRESETn;  // ../RTL/cmsdk_mcu.v(93)
  wire DCLK;  // ../RTL/cmsdk_mcu.v(96)
  wire FCLK;  // ../RTL/cmsdk_mcu.v(94)
  wire HCLK;  // ../RTL/cmsdk_mcu.v(95)
  wire HCLKSYS;  // ../RTL/cmsdk_mcu.v(100)
  wire HREADY;  // ../RTL/cmsdk_mcu.v(108)
  wire HRESETn;  // ../RTL/cmsdk_mcu.v(91)
  wire HWRITE;  // ../RTL/cmsdk_mcu.v(106)
  wire LOCKUP;  // ../RTL/cmsdk_mcu.v(85)
  wire LOCKUPRESET;  // ../RTL/cmsdk_mcu.v(86)
  wire PCLK;  // ../RTL/cmsdk_mcu.v(98)
  wire PCLKEN;  // ../RTL/cmsdk_mcu.v(101)
  wire PCLKG;  // ../RTL/cmsdk_mcu.v(99)
  wire PMUDBGRESETREQ;  // ../RTL/cmsdk_mcu.v(84)
  wire PMUHRESETREQ;  // ../RTL/cmsdk_mcu.v(83)
  wire PORESETn;  // ../RTL/cmsdk_mcu.v(90)
  wire PRESETn;  // ../RTL/cmsdk_mcu.v(92)
  wire SCLK;  // ../RTL/cmsdk_mcu.v(97)
  wire SLEEPDEEP;  // ../RTL/cmsdk_mcu.v(88)
  wire SLEEPING;  // ../RTL/cmsdk_mcu.v(76)
  wire SYSRESETREQ;  // ../RTL/cmsdk_mcu.v(78)
  wire TESTMODE;  // ../RTL/cmsdk_mcu.v(161)
  wire WDOGRESETREQ;  // ../RTL/cmsdk_mcu.v(79)
  wire clk_ctrl_sys_reset_req;  // ../RTL/cmsdk_mcu.v(82)
  wire cmsdk_SYSRESETREQ;  // ../RTL/cmsdk_mcu.v(81)
  wire dbg_swdo;  // ../RTL/cmsdk_mcu.v(166)
  wire dbg_swdo_en;  // ../RTL/cmsdk_mcu.v(165)
  wire flash_hreadyout;  // ../RTL/cmsdk_mcu.v(112)
  wire flash_hresp;  // ../RTL/cmsdk_mcu.v(114)
  wire flash_hsel;  // ../RTL/cmsdk_mcu.v(111)
  wire i_tdi;  // ../RTL/cmsdk_mcu.v(155)
  wire i_tdo;  // ../RTL/cmsdk_mcu.v(156)
  wire i_tdoen_n;  // ../RTL/cmsdk_mcu.v(157)
  wire i_trst_n;  // ../RTL/cmsdk_mcu.v(152)
  wire n0;
  wire n1;
  wire sram_hreadyout;  // ../RTL/cmsdk_mcu.v(118)
  wire sram_hresp;  // ../RTL/cmsdk_mcu.v(120)
  wire sram_hsel;  // ../RTL/cmsdk_mcu.v(117)
  wire timer1_extin;  // ../RTL/cmsdk_mcu.v(135)

  buf u1 (TESTMODE, 1'b0);  // ../RTL/cmsdk_mcu.v(163)
  buf u10 (PMUDBGRESETREQ, 1'b0);  // ../RTL/cmsdk_mcu.v(224)
  buf u11 (PMUHRESETREQ, 1'b0);  // ../RTL/cmsdk_mcu.v(225)
  buf u12 (HCLKSYS, HCLK);  // ../RTL/cmsdk_mcu.v(333)
  bufif1 u2 (TMS, dbg_swdo, dbg_swdo_en);  // ../RTL/cmsdk_mcu.v(167)
  or u3 (clk_ctrl_sys_reset_req, PMUHRESETREQ, cmsdk_SYSRESETREQ);  // ../RTL/cmsdk_mcu.v(177)
  or u4 (n0, SYSRESETREQ, WDOGRESETREQ);  // ../RTL/cmsdk_mcu.v(215)
  and u5 (n1, LOCKUP, LOCKUPRESET);  // ../RTL/cmsdk_mcu.v(216)
  or u6 (cmsdk_SYSRESETREQ, n0, n1);  // ../RTL/cmsdk_mcu.v(216)
  buf u7 (HCLK, FCLK);  // ../RTL/cmsdk_mcu.v(219)
  buf u8 (DCLK, FCLK);  // ../RTL/cmsdk_mcu.v(220)
  buf u9 (SCLK, FCLK);  // ../RTL/cmsdk_mcu.v(221)
  AHB2MEM u_ahb_ram (
    .HADDR({16'b0000000000000000,HADDR[15:0]}),
    .HCLK(HCLKSYS),
    .HREADY(HREADY),
    .HRESETn(HRESETn),
    .HSEL(sram_hsel),
    .HSIZE(HSIZE),
    .HTRANS(HTRANS),
    .HWDATA(HWDATA),
    .HWRITE(HWRITE),
    .HRDATA(sram_hrdata),
    .HREADYOUT(sram_hreadyout),
    .HRESP(sram_hresp));  // ../RTL/cmsdk_mcu.v(361)
  AHB2MEM u_ahb_rom (
    .HADDR({16'b0000000000000000,HADDR[15:0]}),
    .HCLK(HCLKSYS),
    .HREADY(HREADY),
    .HRESETn(HRESETn),
    .HSEL(flash_hsel),
    .HSIZE(HSIZE),
    .HTRANS(HTRANS),
    .HWDATA(HWDATA),
    .HWRITE(HWRITE),
    .HRDATA(flash_hrdata),
    .HREADYOUT(flash_hreadyout),
    .HRESP(flash_hresp));  // ../RTL/cmsdk_mcu.v(340)
  cmsdk_mcu_clkctrl u_cmsdk_mcu_clkctrl (
    .APBACTIVE(APBACTIVE),
    .CGBYPASS(TESTMODE),
    .DBGRESETREQ(PMUDBGRESETREQ),
    .LOCKUP(LOCKUP),
    .LOCKUPRESET(LOCKUPRESET),
    .NRST(NRST),
    .RSTBYPASS(TESTMODE),
    .SLEEPDEEP(SLEEPDEEP),
    .SLEEPING(SLEEPING),
    .SYSRESETREQ(clk_ctrl_sys_reset_req),
    .XTAL1(XTAL1),
    .DBGRESETn(DBGRESETn),
    .FCLK(FCLK),
    .HRESETn(HRESETn),
    .PCLK(PCLK),
    .PCLKEN(PCLKEN),
    .PCLKG(PCLKG),
    .PORESETn(PORESETn),
    .PRESETn(PRESETn),
    .XTAL2(XTAL2));  // ../RTL/cmsdk_mcu.v(182)
  \cmsdk_mcu_system(WIC=1)  u_cmsdk_mcu_system (
    .DBGRESETn(DBGRESETn),
    .DCLK(DCLK),
    .DFTSE(1'b0),
    .FCLK(FCLK),
    .HCLK(HCLK),
    .HRESETn(HRESETn),
    .PCLK(PCLK),
    .PCLKEN(PCLKEN),
    .PCLKG(PCLKG),
    .PORESETn(PORESETn),
    .PRESETn(PRESETn),
    .SCLK(SCLK),
    .SWCLKTCK(TCK),
    .SWDITMS(TMS),
    .TDI(i_tdi),
    .boot_hrdata(32'b00000000000000000000000000000000),
    .boot_hreadyout(1'b0),
    .boot_hresp(1'b0),
    .flash_hrdata(flash_hrdata),
    .flash_hreadyout(flash_hreadyout),
    .flash_hresp(flash_hresp),
    .nTRST(i_trst_n),
    .p0_in(p0_in),
    .p1_in(p1_in),
    .sram_hrdata(sram_hrdata),
    .sram_hreadyout(sram_hreadyout),
    .sram_hresp(sram_hresp),
    .timer1_extin(timer1_extin),
    .uart0_rxd(uart0_rxd),
    .APBACTIVE(APBACTIVE),
    .HADDR({open_n18,open_n19,open_n20,open_n21,open_n22,open_n23,open_n24,open_n25,open_n26,open_n27,open_n28,open_n29,open_n30,open_n31,open_n32,open_n33,HADDR[15:0]}),
    .HREADY(HREADY),
    .HSIZE(HSIZE),
    .HTRANS(HTRANS),
    .HWDATA(HWDATA),
    .HWRITE(HWRITE),
    .LOCKUP(LOCKUP),
    .LOCKUPRESET(LOCKUPRESET),
    .SLEEPDEEP(SLEEPDEEP),
    .SLEEPING(SLEEPING),
    .SWDO(dbg_swdo),
    .SWDOEN(dbg_swdo_en),
    .SYSRESETREQ(SYSRESETREQ),
    .TDO(i_tdo),
    .WDOGRESETREQ(WDOGRESETREQ),
    .flash_hsel(flash_hsel),
    .nTDOEN(i_tdoen_n),
    .p0_altfunc(p0_altfunc),
    .p0_out(p0_out),
    .p0_outen(p0_outen),
    .p1_altfunc(p1_altfunc),
    .p1_out(p1_out),
    .p1_outen(p1_outen),
    .sram_hsel(sram_hsel),
    .uart0_txd(uart0_txd),
    .uart0_txen(uart0_txen),
    .b_pad_gpio_porta(b_pad_gpio_porta));  // ../RTL/cmsdk_mcu.v(244)
  cmsdk_mcu_pin_mux u_pin_mux (
    .SWCLKTCK(SWCLKTCK),
    .TDI(TDI),
    .i_swdo(1'bx),
    .i_swdoen(1'bx),
    .i_tdo(i_tdo),
    .i_tdoen_n(i_tdoen_n),
    .nTRST(nTRST),
    .p0_altfunc(p0_altfunc),
    .p0_out(p0_out),
    .p0_outen(p0_outen),
    .p1_altfunc(p1_altfunc),
    .p1_out(p1_out),
    .p1_outen(p1_outen),
    .P0(P0),
    .TDO(TDO),
    .i_tdi(i_tdi),
    .i_trst_n(i_trst_n),
    .p0_in(p0_in),
    .p1_in(p1_in),
    .timer1_extin(timer1_extin),
    .P1(P1),
    .SWDIOTMS(SWDIOTMS));  // ../RTL/cmsdk_mcu.v(382)

endmodule 

module AHB2MEM  // ../RTL/AHB2MEM.v(5)
  (
  HADDR,
  HCLK,
  HREADY,
  HRESETn,
  HSEL,
  HSIZE,
  HTRANS,
  HWDATA,
  HWRITE,
  HRDATA,
  HREADYOUT,
  HRESP
  );

  input [31:0] HADDR;  // ../RTL/AHB2MEM.v(12)
  input HCLK;  // ../RTL/AHB2MEM.v(9)
  input HREADY;  // ../RTL/AHB2MEM.v(11)
  input HRESETn;  // ../RTL/AHB2MEM.v(10)
  input HSEL;  // ../RTL/AHB2MEM.v(8)
  input [2:0] HSIZE;  // ../RTL/AHB2MEM.v(15)
  input [1:0] HTRANS;  // ../RTL/AHB2MEM.v(13)
  input [31:0] HWDATA;  // ../RTL/AHB2MEM.v(16)
  input HWRITE;  // ../RTL/AHB2MEM.v(14)
  output [31:0] HRDATA;  // ../RTL/AHB2MEM.v(18)
  output HREADYOUT;  // ../RTL/AHB2MEM.v(17)
  output HRESP;  // ../RTL/AHB2MEM.v(19)

  parameter MEMWIDTH = 12;
  wire [31:0] buf_hwaddr;  // ../RTL/AHB2MEM.v(30)
  wire [31:0] hwdata_mask;  // ../RTL/AHB2MEM.v(28)
  wire [31:0] n10;
  wire [31:0] n11;
  wire [31:0] n12;
  wire [31:0] n13;
  wire [31:0] n17;
  wire [31:0] n3;
  wire [31:0] n4;
  wire [31:0] n5;
  wire [31:0] n7;
  wire [31:0] n8;
  wire [31:0] n9;
  wire n0;
  wire n1;
  wire n14;
  wire n15;
  wire n16;
  wire n18;
  wire n19;
  wire n2;
  wire n20;
  wire n21;
  wire n22;
  wire n23;
  wire n24;
  wire n25;
  wire n6;
  wire we;  // ../RTL/AHB2MEM.v(29)

  binary_mux_s2_w32 mux0 (
    .i0(n4),
    .i1({HADDR[1],HADDR[1],HADDR[1],HADDR[1],HADDR[1],HADDR[1],HADDR[1],HADDR[1],HADDR[1],HADDR[1],HADDR[1],HADDR[1],HADDR[1],HADDR[1],HADDR[1],HADDR[1],n3[15:0]}),
    .i2(32'b11111111111111111111111111111111),
    .i3(32'b11111111111111111111111111111111),
    .sel(HSIZE[1:0]),
    .o(n5));  // ../RTL/AHB2MEM.v(50)
  binary_mux_s1_w32 mux1 (
    .i0(buf_hwaddr),
    .i1(HADDR),
    .sel(HREADY),
    .o(n7));  // ../RTL/AHB2MEM.v(51)
  binary_mux_s1_w32 mux2 (
    .i0(hwdata_mask),
    .i1(n5),
    .sel(HREADY),
    .o(n8));  // ../RTL/AHB2MEM.v(51)
  binary_mux_s1_w32 mux3 (
    .i0(n8),
    .i1(hwdata_mask),
    .sel(n0),
    .o(n9));  // ../RTL/AHB2MEM.v(51)
  ram_w10x32_r10x32 #(
    .DATA_DEPTH_LEFT("0"),
    .DATA_DEPTH_RIGHT("1023"),
    .DATA_WIDTH_LEFT("31"),
    .DATA_WIDTH_RIGHT("0"))
    ram_memory (
    .clk1(HCLK),
    .ra1(HADDR[11:2]),
    .re1(1'b1),
    .wa1(buf_hwaddr[11:2]),
    .wd1(n13),
    .we1(n16),
    .rd1(n17));  // ../RTL/AHB2MEM.v(25)
  reg_ar_as_w32 reg0 (
    .clk(HCLK),
    .d(n7),
    .reset({n0,n0,n0,n0,n0,n0,n0,n0,n0,n0,n0,n0,n0,n0,n0,n0,n0,n0,n0,n0,n0,n0,n0,n0,n0,n0,n0,n0,n0,n0,n0,n0}),
    .set(32'b00000000000000000000000000000000),
    .q(buf_hwaddr));  // ../RTL/AHB2MEM.v(51)
  reg_ar_as_w32 reg1 (
    .clk(HCLK),
    .d(n9),
    .reset(32'b00000000000000000000000000000000),
    .set(32'b00000000000000000000000000000000),
    .q(hwdata_mask));  // ../RTL/AHB2MEM.v(51)
  reg_ar_as_w32 reg2 (
    .clk(HCLK),
    .d(n17),
    .reset(32'b00000000000000000000000000000000),
    .set(32'b00000000000000000000000000000000),
    .q(HRDATA));  // ../RTL/AHB2MEM.v(61)
  AL_MUX u10 (
    .i0(we),
    .i1(n2),
    .sel(HREADY),
    .o(n6));  // ../RTL/AHB2MEM.v(51)
  not u100 (n11[24], hwdata_mask[24]);  // ../RTL/AHB2MEM.v(58)
  not u101 (n11[25], hwdata_mask[25]);  // ../RTL/AHB2MEM.v(58)
  not u102 (n11[26], hwdata_mask[26]);  // ../RTL/AHB2MEM.v(58)
  not u103 (n11[27], hwdata_mask[27]);  // ../RTL/AHB2MEM.v(58)
  not u104 (n11[28], hwdata_mask[28]);  // ../RTL/AHB2MEM.v(58)
  not u105 (n11[29], hwdata_mask[29]);  // ../RTL/AHB2MEM.v(58)
  not u106 (n11[30], hwdata_mask[30]);  // ../RTL/AHB2MEM.v(58)
  not u107 (n11[31], hwdata_mask[31]);  // ../RTL/AHB2MEM.v(58)
  and u108 (n10[1], HWDATA[1], hwdata_mask[1]);  // ../RTL/AHB2MEM.v(58)
  and u109 (n10[2], HWDATA[2], hwdata_mask[2]);  // ../RTL/AHB2MEM.v(58)
  and u11 (n10[0], HWDATA[0], hwdata_mask[0]);  // ../RTL/AHB2MEM.v(58)
  and u110 (n10[3], HWDATA[3], hwdata_mask[3]);  // ../RTL/AHB2MEM.v(58)
  and u111 (n10[4], HWDATA[4], hwdata_mask[4]);  // ../RTL/AHB2MEM.v(58)
  and u112 (n10[5], HWDATA[5], hwdata_mask[5]);  // ../RTL/AHB2MEM.v(58)
  and u113 (n10[6], HWDATA[6], hwdata_mask[6]);  // ../RTL/AHB2MEM.v(58)
  and u114 (n10[7], HWDATA[7], hwdata_mask[7]);  // ../RTL/AHB2MEM.v(58)
  and u115 (n10[8], HWDATA[8], hwdata_mask[8]);  // ../RTL/AHB2MEM.v(58)
  and u116 (n10[9], HWDATA[9], hwdata_mask[9]);  // ../RTL/AHB2MEM.v(58)
  and u117 (n10[10], HWDATA[10], hwdata_mask[10]);  // ../RTL/AHB2MEM.v(58)
  and u118 (n10[11], HWDATA[11], hwdata_mask[11]);  // ../RTL/AHB2MEM.v(58)
  and u119 (n10[12], HWDATA[12], hwdata_mask[12]);  // ../RTL/AHB2MEM.v(58)
  not u12 (n11[0], hwdata_mask[0]);  // ../RTL/AHB2MEM.v(58)
  and u120 (n10[13], HWDATA[13], hwdata_mask[13]);  // ../RTL/AHB2MEM.v(58)
  and u121 (n10[14], HWDATA[14], hwdata_mask[14]);  // ../RTL/AHB2MEM.v(58)
  and u122 (n10[15], HWDATA[15], hwdata_mask[15]);  // ../RTL/AHB2MEM.v(58)
  and u123 (n10[16], HWDATA[16], hwdata_mask[16]);  // ../RTL/AHB2MEM.v(58)
  and u124 (n10[17], HWDATA[17], hwdata_mask[17]);  // ../RTL/AHB2MEM.v(58)
  and u125 (n10[18], HWDATA[18], hwdata_mask[18]);  // ../RTL/AHB2MEM.v(58)
  and u126 (n10[19], HWDATA[19], hwdata_mask[19]);  // ../RTL/AHB2MEM.v(58)
  and u127 (n10[20], HWDATA[20], hwdata_mask[20]);  // ../RTL/AHB2MEM.v(58)
  and u128 (n10[21], HWDATA[21], hwdata_mask[21]);  // ../RTL/AHB2MEM.v(58)
  and u129 (n10[22], HWDATA[22], hwdata_mask[22]);  // ../RTL/AHB2MEM.v(58)
  and u13 (n12[0], HRDATA[0], n11[0]);  // ../RTL/AHB2MEM.v(58)
  and u130 (n10[23], HWDATA[23], hwdata_mask[23]);  // ../RTL/AHB2MEM.v(58)
  and u131 (n10[24], HWDATA[24], hwdata_mask[24]);  // ../RTL/AHB2MEM.v(58)
  and u132 (n10[25], HWDATA[25], hwdata_mask[25]);  // ../RTL/AHB2MEM.v(58)
  and u133 (n10[26], HWDATA[26], hwdata_mask[26]);  // ../RTL/AHB2MEM.v(58)
  and u134 (n10[27], HWDATA[27], hwdata_mask[27]);  // ../RTL/AHB2MEM.v(58)
  and u135 (n10[28], HWDATA[28], hwdata_mask[28]);  // ../RTL/AHB2MEM.v(58)
  and u136 (n10[29], HWDATA[29], hwdata_mask[29]);  // ../RTL/AHB2MEM.v(58)
  and u137 (n10[30], HWDATA[30], hwdata_mask[30]);  // ../RTL/AHB2MEM.v(58)
  and u138 (n10[31], HWDATA[31], hwdata_mask[31]);  // ../RTL/AHB2MEM.v(58)
  not u139 (n18, HADDR[0]);  // ../RTL/AHB2MEM.v(49)
  or u14 (n13[0], n10[0], n12[0]);  // ../RTL/AHB2MEM.v(58)
  not u140 (n19, HADDR[0]);  // ../RTL/AHB2MEM.v(49)
  not u141 (n20, HADDR[0]);  // ../RTL/AHB2MEM.v(49)
  not u142 (n21, HADDR[0]);  // ../RTL/AHB2MEM.v(49)
  not u143 (n22, HADDR[0]);  // ../RTL/AHB2MEM.v(49)
  not u144 (n23, HADDR[0]);  // ../RTL/AHB2MEM.v(49)
  not u145 (n24, HADDR[0]);  // ../RTL/AHB2MEM.v(49)
  not u146 (n25, HADDR[0]);  // ../RTL/AHB2MEM.v(49)
  AL_MUX u147 (
    .i0(1'b0),
    .i1(HADDR[0]),
    .sel(HADDR[1]),
    .o(n4[31]));  // ../RTL/AHB2MEM.v(49)
  AL_MUX u148 (
    .i0(1'b0),
    .i1(HADDR[0]),
    .sel(HADDR[1]),
    .o(n4[30]));  // ../RTL/AHB2MEM.v(49)
  AL_MUX u149 (
    .i0(1'b0),
    .i1(HADDR[0]),
    .sel(HADDR[1]),
    .o(n4[29]));  // ../RTL/AHB2MEM.v(49)
  and u15 (n16, n14, n15);  // ../RTL/AHB2MEM.v(58)
  AL_MUX u150 (
    .i0(1'b0),
    .i1(HADDR[0]),
    .sel(HADDR[1]),
    .o(n4[28]));  // ../RTL/AHB2MEM.v(49)
  AL_MUX u151 (
    .i0(1'b0),
    .i1(HADDR[0]),
    .sel(HADDR[1]),
    .o(n4[27]));  // ../RTL/AHB2MEM.v(49)
  AL_MUX u152 (
    .i0(1'b0),
    .i1(HADDR[0]),
    .sel(HADDR[1]),
    .o(n4[26]));  // ../RTL/AHB2MEM.v(49)
  AL_MUX u153 (
    .i0(1'b0),
    .i1(HADDR[0]),
    .sel(HADDR[1]),
    .o(n4[25]));  // ../RTL/AHB2MEM.v(49)
  AL_MUX u154 (
    .i0(1'b0),
    .i1(HADDR[0]),
    .sel(HADDR[1]),
    .o(n4[24]));  // ../RTL/AHB2MEM.v(49)
  AL_MUX u155 (
    .i0(1'b0),
    .i1(n18),
    .sel(HADDR[1]),
    .o(n4[23]));  // ../RTL/AHB2MEM.v(49)
  AL_MUX u156 (
    .i0(1'b0),
    .i1(n19),
    .sel(HADDR[1]),
    .o(n4[22]));  // ../RTL/AHB2MEM.v(49)
  AL_MUX u157 (
    .i0(1'b0),
    .i1(n20),
    .sel(HADDR[1]),
    .o(n4[21]));  // ../RTL/AHB2MEM.v(49)
  AL_MUX u158 (
    .i0(1'b0),
    .i1(n21),
    .sel(HADDR[1]),
    .o(n4[20]));  // ../RTL/AHB2MEM.v(49)
  AL_MUX u159 (
    .i0(1'b0),
    .i1(n22),
    .sel(HADDR[1]),
    .o(n4[19]));  // ../RTL/AHB2MEM.v(49)
  buf u16 (n15, we);  // ../RTL/AHB2MEM.v(61)
  AL_MUX u160 (
    .i0(1'b0),
    .i1(n23),
    .sel(HADDR[1]),
    .o(n4[18]));  // ../RTL/AHB2MEM.v(49)
  AL_MUX u161 (
    .i0(1'b0),
    .i1(n24),
    .sel(HADDR[1]),
    .o(n4[17]));  // ../RTL/AHB2MEM.v(49)
  AL_MUX u162 (
    .i0(1'b0),
    .i1(n25),
    .sel(HADDR[1]),
    .o(n4[16]));  // ../RTL/AHB2MEM.v(49)
  AL_MUX u163 (
    .i0(HADDR[0]),
    .i1(1'b0),
    .sel(HADDR[1]),
    .o(n4[15]));  // ../RTL/AHB2MEM.v(49)
  AL_MUX u164 (
    .i0(HADDR[0]),
    .i1(1'b0),
    .sel(HADDR[1]),
    .o(n4[14]));  // ../RTL/AHB2MEM.v(49)
  AL_MUX u165 (
    .i0(HADDR[0]),
    .i1(1'b0),
    .sel(HADDR[1]),
    .o(n4[13]));  // ../RTL/AHB2MEM.v(49)
  AL_MUX u166 (
    .i0(HADDR[0]),
    .i1(1'b0),
    .sel(HADDR[1]),
    .o(n4[12]));  // ../RTL/AHB2MEM.v(49)
  AL_MUX u167 (
    .i0(HADDR[0]),
    .i1(1'b0),
    .sel(HADDR[1]),
    .o(n4[11]));  // ../RTL/AHB2MEM.v(49)
  AL_MUX u168 (
    .i0(HADDR[0]),
    .i1(1'b0),
    .sel(HADDR[1]),
    .o(n4[10]));  // ../RTL/AHB2MEM.v(49)
  AL_MUX u169 (
    .i0(HADDR[0]),
    .i1(1'b0),
    .sel(HADDR[1]),
    .o(n4[9]));  // ../RTL/AHB2MEM.v(49)
  or u17 (n13[3], n10[3], n12[3]);  // ../RTL/AHB2MEM.v(58)
  AL_MUX u170 (
    .i0(HADDR[0]),
    .i1(1'b0),
    .sel(HADDR[1]),
    .o(n4[8]));  // ../RTL/AHB2MEM.v(49)
  AL_MUX u171 (
    .i0(n18),
    .i1(1'b0),
    .sel(HADDR[1]),
    .o(n4[7]));  // ../RTL/AHB2MEM.v(49)
  AL_MUX u172 (
    .i0(n19),
    .i1(1'b0),
    .sel(HADDR[1]),
    .o(n4[6]));  // ../RTL/AHB2MEM.v(49)
  AL_MUX u173 (
    .i0(n20),
    .i1(1'b0),
    .sel(HADDR[1]),
    .o(n4[5]));  // ../RTL/AHB2MEM.v(49)
  AL_MUX u174 (
    .i0(n21),
    .i1(1'b0),
    .sel(HADDR[1]),
    .o(n4[4]));  // ../RTL/AHB2MEM.v(49)
  AL_MUX u175 (
    .i0(n22),
    .i1(1'b0),
    .sel(HADDR[1]),
    .o(n4[3]));  // ../RTL/AHB2MEM.v(49)
  AL_MUX u176 (
    .i0(n23),
    .i1(1'b0),
    .sel(HADDR[1]),
    .o(n4[2]));  // ../RTL/AHB2MEM.v(49)
  AL_MUX u177 (
    .i0(n24),
    .i1(1'b0),
    .sel(HADDR[1]),
    .o(n4[1]));  // ../RTL/AHB2MEM.v(49)
  AL_MUX u178 (
    .i0(n25),
    .i1(1'b0),
    .sel(HADDR[1]),
    .o(n4[0]));  // ../RTL/AHB2MEM.v(49)
  not u179 (n3[15], HADDR[1]);  // ../RTL/AHB2MEM.v(48)
  or u18 (n13[4], n10[4], n12[4]);  // ../RTL/AHB2MEM.v(58)
  not u180 (n3[14], HADDR[1]);  // ../RTL/AHB2MEM.v(48)
  not u181 (n3[13], HADDR[1]);  // ../RTL/AHB2MEM.v(48)
  not u182 (n3[12], HADDR[1]);  // ../RTL/AHB2MEM.v(48)
  not u183 (n3[11], HADDR[1]);  // ../RTL/AHB2MEM.v(48)
  not u184 (n3[10], HADDR[1]);  // ../RTL/AHB2MEM.v(48)
  not u185 (n3[9], HADDR[1]);  // ../RTL/AHB2MEM.v(48)
  not u186 (n3[8], HADDR[1]);  // ../RTL/AHB2MEM.v(48)
  not u187 (n3[7], HADDR[1]);  // ../RTL/AHB2MEM.v(48)
  not u188 (n3[6], HADDR[1]);  // ../RTL/AHB2MEM.v(48)
  not u189 (n3[5], HADDR[1]);  // ../RTL/AHB2MEM.v(48)
  or u19 (n13[5], n10[5], n12[5]);  // ../RTL/AHB2MEM.v(58)
  not u190 (n3[4], HADDR[1]);  // ../RTL/AHB2MEM.v(48)
  not u191 (n3[3], HADDR[1]);  // ../RTL/AHB2MEM.v(48)
  not u192 (n3[2], HADDR[1]);  // ../RTL/AHB2MEM.v(48)
  not u193 (n3[1], HADDR[1]);  // ../RTL/AHB2MEM.v(48)
  not u194 (n3[0], HADDR[1]);  // ../RTL/AHB2MEM.v(48)
  or u2 (n13[2], n10[2], n12[2]);  // ../RTL/AHB2MEM.v(58)
  or u20 (n13[6], n10[6], n12[6]);  // ../RTL/AHB2MEM.v(58)
  or u21 (n13[7], n10[7], n12[7]);  // ../RTL/AHB2MEM.v(58)
  or u22 (n13[8], n10[8], n12[8]);  // ../RTL/AHB2MEM.v(58)
  or u23 (n13[9], n10[9], n12[9]);  // ../RTL/AHB2MEM.v(58)
  or u24 (n13[10], n10[10], n12[10]);  // ../RTL/AHB2MEM.v(58)
  or u25 (n13[11], n10[11], n12[11]);  // ../RTL/AHB2MEM.v(58)
  or u26 (n13[12], n10[12], n12[12]);  // ../RTL/AHB2MEM.v(58)
  or u27 (n13[13], n10[13], n12[13]);  // ../RTL/AHB2MEM.v(58)
  or u28 (n13[14], n10[14], n12[14]);  // ../RTL/AHB2MEM.v(58)
  or u29 (n13[15], n10[15], n12[15]);  // ../RTL/AHB2MEM.v(58)
  or u3 (n13[1], n10[1], n12[1]);  // ../RTL/AHB2MEM.v(58)
  or u30 (n13[16], n10[16], n12[16]);  // ../RTL/AHB2MEM.v(58)
  or u31 (n13[17], n10[17], n12[17]);  // ../RTL/AHB2MEM.v(58)
  or u32 (n13[18], n10[18], n12[18]);  // ../RTL/AHB2MEM.v(58)
  or u33 (n13[19], n10[19], n12[19]);  // ../RTL/AHB2MEM.v(58)
  or u34 (n13[20], n10[20], n12[20]);  // ../RTL/AHB2MEM.v(58)
  or u35 (n13[21], n10[21], n12[21]);  // ../RTL/AHB2MEM.v(58)
  or u36 (n13[22], n10[22], n12[22]);  // ../RTL/AHB2MEM.v(58)
  or u37 (n13[23], n10[23], n12[23]);  // ../RTL/AHB2MEM.v(58)
  or u38 (n13[24], n10[24], n12[24]);  // ../RTL/AHB2MEM.v(58)
  or u39 (n13[25], n10[25], n12[25]);  // ../RTL/AHB2MEM.v(58)
  buf u4 (HREADYOUT, 1'b1);  // ../RTL/AHB2MEM.v(22)
  or u40 (n13[26], n10[26], n12[26]);  // ../RTL/AHB2MEM.v(58)
  or u41 (n13[27], n10[27], n12[27]);  // ../RTL/AHB2MEM.v(58)
  or u42 (n13[28], n10[28], n12[28]);  // ../RTL/AHB2MEM.v(58)
  or u43 (n13[29], n10[29], n12[29]);  // ../RTL/AHB2MEM.v(58)
  or u44 (n13[30], n10[30], n12[30]);  // ../RTL/AHB2MEM.v(58)
  or u45 (n13[31], n10[31], n12[31]);  // ../RTL/AHB2MEM.v(58)
  and u46 (n12[1], HRDATA[1], n11[1]);  // ../RTL/AHB2MEM.v(58)
  and u47 (n12[2], HRDATA[2], n11[2]);  // ../RTL/AHB2MEM.v(58)
  and u48 (n12[3], HRDATA[3], n11[3]);  // ../RTL/AHB2MEM.v(58)
  and u49 (n12[4], HRDATA[4], n11[4]);  // ../RTL/AHB2MEM.v(58)
  buf u5 (HRESP, 1'b0);  // ../RTL/AHB2MEM.v(23)
  and u50 (n12[5], HRDATA[5], n11[5]);  // ../RTL/AHB2MEM.v(58)
  and u51 (n12[6], HRDATA[6], n11[6]);  // ../RTL/AHB2MEM.v(58)
  and u52 (n12[7], HRDATA[7], n11[7]);  // ../RTL/AHB2MEM.v(58)
  and u53 (n12[8], HRDATA[8], n11[8]);  // ../RTL/AHB2MEM.v(58)
  and u54 (n12[9], HRDATA[9], n11[9]);  // ../RTL/AHB2MEM.v(58)
  and u55 (n12[10], HRDATA[10], n11[10]);  // ../RTL/AHB2MEM.v(58)
  and u56 (n12[11], HRDATA[11], n11[11]);  // ../RTL/AHB2MEM.v(58)
  and u57 (n12[12], HRDATA[12], n11[12]);  // ../RTL/AHB2MEM.v(58)
  and u58 (n12[13], HRDATA[13], n11[13]);  // ../RTL/AHB2MEM.v(58)
  and u59 (n12[14], HRDATA[14], n11[14]);  // ../RTL/AHB2MEM.v(58)
  not u6 (n14, buf_hwaddr[12]);  // ../RTL/AHB2MEM.v(58)
  and u60 (n12[15], HRDATA[15], n11[15]);  // ../RTL/AHB2MEM.v(58)
  and u61 (n12[16], HRDATA[16], n11[16]);  // ../RTL/AHB2MEM.v(58)
  and u62 (n12[17], HRDATA[17], n11[17]);  // ../RTL/AHB2MEM.v(58)
  and u63 (n12[18], HRDATA[18], n11[18]);  // ../RTL/AHB2MEM.v(58)
  and u64 (n12[19], HRDATA[19], n11[19]);  // ../RTL/AHB2MEM.v(58)
  and u65 (n12[20], HRDATA[20], n11[20]);  // ../RTL/AHB2MEM.v(58)
  and u66 (n12[21], HRDATA[21], n11[21]);  // ../RTL/AHB2MEM.v(58)
  and u67 (n12[22], HRDATA[22], n11[22]);  // ../RTL/AHB2MEM.v(58)
  and u68 (n12[23], HRDATA[23], n11[23]);  // ../RTL/AHB2MEM.v(58)
  and u69 (n12[24], HRDATA[24], n11[24]);  // ../RTL/AHB2MEM.v(58)
  not u7 (n0, HRESETn);  // ../RTL/AHB2MEM.v(35)
  and u70 (n12[25], HRDATA[25], n11[25]);  // ../RTL/AHB2MEM.v(58)
  and u71 (n12[26], HRDATA[26], n11[26]);  // ../RTL/AHB2MEM.v(58)
  and u72 (n12[27], HRDATA[27], n11[27]);  // ../RTL/AHB2MEM.v(58)
  and u73 (n12[28], HRDATA[28], n11[28]);  // ../RTL/AHB2MEM.v(58)
  and u74 (n12[29], HRDATA[29], n11[29]);  // ../RTL/AHB2MEM.v(58)
  and u75 (n12[30], HRDATA[30], n11[30]);  // ../RTL/AHB2MEM.v(58)
  and u76 (n12[31], HRDATA[31], n11[31]);  // ../RTL/AHB2MEM.v(58)
  not u77 (n11[1], hwdata_mask[1]);  // ../RTL/AHB2MEM.v(58)
  not u78 (n11[2], hwdata_mask[2]);  // ../RTL/AHB2MEM.v(58)
  not u79 (n11[3], hwdata_mask[3]);  // ../RTL/AHB2MEM.v(58)
  and u8 (n1, HSEL, HWRITE);  // ../RTL/AHB2MEM.v(43)
  not u80 (n11[4], hwdata_mask[4]);  // ../RTL/AHB2MEM.v(58)
  not u81 (n11[5], hwdata_mask[5]);  // ../RTL/AHB2MEM.v(58)
  not u82 (n11[6], hwdata_mask[6]);  // ../RTL/AHB2MEM.v(58)
  not u83 (n11[7], hwdata_mask[7]);  // ../RTL/AHB2MEM.v(58)
  not u84 (n11[8], hwdata_mask[8]);  // ../RTL/AHB2MEM.v(58)
  not u85 (n11[9], hwdata_mask[9]);  // ../RTL/AHB2MEM.v(58)
  not u86 (n11[10], hwdata_mask[10]);  // ../RTL/AHB2MEM.v(58)
  not u87 (n11[11], hwdata_mask[11]);  // ../RTL/AHB2MEM.v(58)
  not u88 (n11[12], hwdata_mask[12]);  // ../RTL/AHB2MEM.v(58)
  not u89 (n11[13], hwdata_mask[13]);  // ../RTL/AHB2MEM.v(58)
  and u9 (n2, n1, HTRANS[1]);  // ../RTL/AHB2MEM.v(43)
  not u90 (n11[14], hwdata_mask[14]);  // ../RTL/AHB2MEM.v(58)
  not u91 (n11[15], hwdata_mask[15]);  // ../RTL/AHB2MEM.v(58)
  not u92 (n11[16], hwdata_mask[16]);  // ../RTL/AHB2MEM.v(58)
  not u93 (n11[17], hwdata_mask[17]);  // ../RTL/AHB2MEM.v(58)
  not u94 (n11[18], hwdata_mask[18]);  // ../RTL/AHB2MEM.v(58)
  not u95 (n11[19], hwdata_mask[19]);  // ../RTL/AHB2MEM.v(58)
  not u96 (n11[20], hwdata_mask[20]);  // ../RTL/AHB2MEM.v(58)
  not u97 (n11[21], hwdata_mask[21]);  // ../RTL/AHB2MEM.v(58)
  not u98 (n11[22], hwdata_mask[22]);  // ../RTL/AHB2MEM.v(58)
  not u99 (n11[23], hwdata_mask[23]);  // ../RTL/AHB2MEM.v(58)
  AL_DFF we_reg (
    .clk(HCLK),
    .d(n6),
    .reset(n0),
    .set(1'b0),
    .q(we));  // ../RTL/AHB2MEM.v(51)

endmodule 

module cmsdk_mcu_clkctrl  // ../RTL/cmsdk_mcu_clkctrl.v(33)
  (
  APBACTIVE,
  CGBYPASS,
  DBGRESETREQ,
  LOCKUP,
  LOCKUPRESET,
  NRST,
  RSTBYPASS,
  SLEEPDEEP,
  SLEEPING,
  SYSRESETREQ,
  XTAL1,
  DBGRESETn,
  FCLK,
  HRESETn,
  PCLK,
  PCLKEN,
  PCLKG,
  PORESETn,
  PRESETn,
  XTAL2
  );

  input APBACTIVE;  // ../RTL/cmsdk_mcu_clkctrl.v(39)
  input CGBYPASS;  // ../RTL/cmsdk_mcu_clkctrl.v(47)
  input DBGRESETREQ;  // ../RTL/cmsdk_mcu_clkctrl.v(43)
  input LOCKUP;  // ../RTL/cmsdk_mcu_clkctrl.v(44)
  input LOCKUPRESET;  // ../RTL/cmsdk_mcu_clkctrl.v(45)
  input NRST;  // ../RTL/cmsdk_mcu_clkctrl.v(37)
  input RSTBYPASS;  // ../RTL/cmsdk_mcu_clkctrl.v(48)
  input SLEEPDEEP;  // ../RTL/cmsdk_mcu_clkctrl.v(41)
  input SLEEPING;  // ../RTL/cmsdk_mcu_clkctrl.v(40)
  input SYSRESETREQ;  // ../RTL/cmsdk_mcu_clkctrl.v(42)
  input XTAL1;  // ../RTL/cmsdk_mcu_clkctrl.v(36)
  output DBGRESETn;  // ../RTL/cmsdk_mcu_clkctrl.v(56)
  output FCLK;  // ../RTL/cmsdk_mcu_clkctrl.v(51)
  output HRESETn;  // ../RTL/cmsdk_mcu_clkctrl.v(57)
  output PCLK;  // ../RTL/cmsdk_mcu_clkctrl.v(52)
  output PCLKEN;  // ../RTL/cmsdk_mcu_clkctrl.v(54)
  output PCLKG;  // ../RTL/cmsdk_mcu_clkctrl.v(53)
  output PORESETn;  // ../RTL/cmsdk_mcu_clkctrl.v(55)
  output PRESETn;  // ../RTL/cmsdk_mcu_clkctrl.v(58)
  output XTAL2;  // ../RTL/cmsdk_mcu_clkctrl.v(50)

  parameter CLKGATE_PRESENT = 0;
  wire [2:0] nxt_reset_sync;  // ../RTL/cmsdk_mcu_clkctrl.v(63)
  wire [2:0] reset_sync_reg;  // ../RTL/cmsdk_mcu_clkctrl.v(62)
  wire clk;  // ../RTL/cmsdk_mcu_clkctrl.v(60)
  wire dbgrst_reg;  // ../RTL/cmsdk_mcu_clkctrl.v(66)
  wire i_pclken;  // ../RTL/cmsdk_mcu_clkctrl.v(69)
  wire n0;
  wire n1;
  wire n2;
  wire n3;
  wire n4;
  wire n5;
  wire nxt_hrst;  // ../RTL/cmsdk_mcu_clkctrl.v(65)
  wire prst_reg;  // ../RTL/cmsdk_mcu_clkctrl.v(67)
  wire reset_n;  // ../RTL/cmsdk_mcu_clkctrl.v(61)

  assign PRESETn = HRESETn;
  AL_DFF dbgrst_reg_reg (
    .clk(clk),
    .d(n5),
    .reset(n4),
    .set(1'b0),
    .q(dbgrst_reg));  // ../RTL/cmsdk_mcu_clkctrl.v(108)
  AL_DFF prst_reg_reg (
    .clk(clk),
    .d(nxt_hrst),
    .reset(n4),
    .set(1'b0),
    .q(prst_reg));  // ../RTL/cmsdk_mcu_clkctrl.v(119)
  reg_ar_as_w3 reg0 (
    .clk(clk),
    .d(nxt_reset_sync),
    .reset({n1,n1,n1}),
    .set(3'b000),
    .q(reset_sync_reg));  // ../RTL/cmsdk_mcu_clkctrl.v(86)
  not u10 (nxt_hrst, n3);  // ../RTL/cmsdk_mcu_clkctrl.v(92)
  not u11 (n4, reset_n);  // ../RTL/cmsdk_mcu_clkctrl.v(96)
  not u12 (n5, DBGRESETREQ);  // ../RTL/cmsdk_mcu_clkctrl.v(108)
  buf u13 (nxt_reset_sync[2], reset_sync_reg[1]);  // ../RTL/cmsdk_mcu_clkctrl.v(79)
  buf u14 (i_pclken, 1'b1);  // ../RTL/cmsdk_mcu_clkctrl.v(125)
  buf u15 (PCLK, clk);  // ../RTL/cmsdk_mcu_clkctrl.v(127)
  buf u16 (PCLKG, clk);  // ../RTL/cmsdk_mcu_clkctrl.v(128)
  AL_MUX u17 (
    .i0(reset_n),
    .i1(NRST),
    .sel(RSTBYPASS),
    .o(PORESETn));  // ../RTL/cmsdk_mcu_clkctrl.v(158)
  AL_MUX u18 (
    .i0(prst_reg),
    .i1(NRST),
    .sel(RSTBYPASS),
    .o(HRESETn));  // ../RTL/cmsdk_mcu_clkctrl.v(159)
  AL_MUX u19 (
    .i0(dbgrst_reg),
    .i1(NRST),
    .sel(RSTBYPASS),
    .o(DBGRESETn));  // ../RTL/cmsdk_mcu_clkctrl.v(160)
  or u2 (n0, XTAL1, SLEEPDEEP);  // ../RTL/cmsdk_mcu_clkctrl.v(73)
  buf u20 (nxt_reset_sync[0], 1'b1);  // ../RTL/cmsdk_mcu_clkctrl.v(79)
  buf u21 (FCLK, clk);  // ../RTL/cmsdk_mcu_clkctrl.v(162)
  buf u22 (PCLKEN, i_pclken);  // ../RTL/cmsdk_mcu_clkctrl.v(163)
  not u3 (XTAL2, n0);  // ../RTL/cmsdk_mcu_clkctrl.v(73)
  buf u4 (clk, XTAL1);  // ../RTL/cmsdk_mcu_clkctrl.v(76)
  not u5 (n1, NRST);  // ../RTL/cmsdk_mcu_clkctrl.v(83)
  buf u6 (nxt_reset_sync[1], reset_sync_reg[0]);  // ../RTL/cmsdk_mcu_clkctrl.v(79)
  buf u7 (reset_n, reset_sync_reg[2]);  // ../RTL/cmsdk_mcu_clkctrl.v(89)
  and u8 (n2, LOCKUP, LOCKUPRESET);  // ../RTL/cmsdk_mcu_clkctrl.v(92)
  or u9 (n3, SYSRESETREQ, n2);  // ../RTL/cmsdk_mcu_clkctrl.v(92)

endmodule 

module \cmsdk_mcu_system(WIC=1)   // ../RTL/cmsdk_mcu_system.v(29)
  (
  CDBGPWRUPACK,
  DBGRESETn,
  DBGRESTART,
  DCLK,
  DFTSE,
  EDBGRQ,
  FCLK,
  HCLK,
  HRESETn,
  PCLK,
  PCLKEN,
  PCLKG,
  PORESETn,
  PRESETn,
  RSTBYPASS,
  SCLK,
  SLEEPHOLDREQn,
  SLOWCLK,
  SLOWCLKG,
  SWCLKTCK,
  SWDITMS,
  TDI,
  WICENREQ,
  boot_hrdata,
  boot_hreadyout,
  boot_hresp,
  eth_interrupt,
  flash_hrdata,
  flash_hreadyout,
  flash_hresp,
  gpio2_interrupt,
  gpio3_interrupt,
  i2s_interrupt,
  nTRST,
  p0_in,
  p1_in,
  spi_interrupt,
  sram_hrdata,
  sram_hreadyout,
  sram_hresp,
  timer1_extin,
  ts_interrupt,
  uart0_rxd,
  zbt_boot_ctrl,
  APBACTIVE,
  CDBGPWRUPREQ,
  DBGRESTARTED,
  GATEHCLK,
  HADDR,
  HREADY,
  HSIZE,
  HTRANS,
  HWDATA,
  HWRITE,
  LOCKUP,
  LOCKUPRESET,
  PMUENABLE,
  SLEEPDEEP,
  SLEEPHOLDACKn,
  SLEEPING,
  SWDO,
  SWDOEN,
  SYSRESETREQ,
  TDO,
  WAKEUP,
  WDOGRESETREQ,
  WICENACK,
  boot_hsel,
  flash_hsel,
  nTDOEN,
  p0_altfunc,
  p0_out,
  p0_outen,
  p1_altfunc,
  p1_out,
  p1_outen,
  sram_hsel,
  uart0_txd,
  uart0_txen,
  b_pad_gpio_porta
  );

  input CDBGPWRUPACK;  // ../RTL/cmsdk_mcu_system.v(119)
  input DBGRESETn;  // ../RTL/cmsdk_mcu_system.v(69)
  input DBGRESTART;  // ../RTL/cmsdk_mcu_system.v(170)
  input DCLK;  // ../RTL/cmsdk_mcu_system.v(65)
  input DFTSE;  // ../RTL/cmsdk_mcu_system.v(174)
  input EDBGRQ;  // ../RTL/cmsdk_mcu_system.v(172)
  input FCLK;  // ../RTL/cmsdk_mcu_system.v(63)
  input HCLK;  // ../RTL/cmsdk_mcu_system.v(64)
  input HRESETn;  // ../RTL/cmsdk_mcu_system.v(67)
  input PCLK;  // ../RTL/cmsdk_mcu_system.v(71)
  input PCLKEN;  // ../RTL/cmsdk_mcu_system.v(76)
  input PCLKG;  // ../RTL/cmsdk_mcu_system.v(72)
  input PORESETn;  // ../RTL/cmsdk_mcu_system.v(68)
  input PRESETn;  // ../RTL/cmsdk_mcu_system.v(75)
  input RSTBYPASS;  // ../RTL/cmsdk_mcu_system.v(70)
  input SCLK;  // ../RTL/cmsdk_mcu_system.v(66)
  input SLEEPHOLDREQn;  // ../RTL/cmsdk_mcu_system.v(120)
  input SLOWCLK;  // ../RTL/cmsdk_mcu_system.v(73)
  input SLOWCLKG;  // ../RTL/cmsdk_mcu_system.v(74)
  input SWCLKTCK;  // ../RTL/cmsdk_mcu_system.v(162)
  input SWDITMS;  // ../RTL/cmsdk_mcu_system.v(163)
  input TDI;  // ../RTL/cmsdk_mcu_system.v(164)
  input WICENREQ;  // ../RTL/cmsdk_mcu_system.v(116)
  input [31:0] boot_hrdata;  // ../RTL/cmsdk_mcu_system.v(100)
  input boot_hreadyout;  // ../RTL/cmsdk_mcu_system.v(99)
  input boot_hresp;  // ../RTL/cmsdk_mcu_system.v(101)
  input eth_interrupt;  // ../RTL/cmsdk_mcu_system.v(155)
  input [31:0] flash_hrdata;  // ../RTL/cmsdk_mcu_system.v(89)
  input flash_hreadyout;  // ../RTL/cmsdk_mcu_system.v(88)
  input flash_hresp;  // ../RTL/cmsdk_mcu_system.v(90)
  input gpio2_interrupt;  // ../RTL/cmsdk_mcu_system.v(157)
  input gpio3_interrupt;  // ../RTL/cmsdk_mcu_system.v(158)
  input i2s_interrupt;  // ../RTL/cmsdk_mcu_system.v(154)
  input nTRST;  // ../RTL/cmsdk_mcu_system.v(161)
  input [15:0] p0_in;  // ../RTL/cmsdk_mcu_system.v(144)
  input [15:0] p1_in;  // ../RTL/cmsdk_mcu_system.v(148)
  input spi_interrupt;  // ../RTL/cmsdk_mcu_system.v(153)
  input [31:0] sram_hrdata;  // ../RTL/cmsdk_mcu_system.v(94)
  input sram_hreadyout;  // ../RTL/cmsdk_mcu_system.v(93)
  input sram_hresp;  // ../RTL/cmsdk_mcu_system.v(95)
  input timer1_extin;  // ../RTL/cmsdk_mcu_system.v(142)
  input ts_interrupt;  // ../RTL/cmsdk_mcu_system.v(156)
  input uart0_rxd;  // ../RTL/cmsdk_mcu_system.v(123)
  input zbt_boot_ctrl;  // ../RTL/cmsdk_mcu_system.v(78)
  output APBACTIVE;  // ../RTL/cmsdk_mcu_system.v(104)
  output CDBGPWRUPREQ;  // ../RTL/cmsdk_mcu_system.v(118)
  output DBGRESTARTED;  // ../RTL/cmsdk_mcu_system.v(171)
  output GATEHCLK;  // ../RTL/cmsdk_mcu_system.v(114)
  output [31:0] HADDR;  // ../RTL/cmsdk_mcu_system.v(80)
  output HREADY;  // ../RTL/cmsdk_mcu_system.v(85)
  output [2:0] HSIZE;  // ../RTL/cmsdk_mcu_system.v(82)
  output [1:0] HTRANS;  // ../RTL/cmsdk_mcu_system.v(81)
  output [31:0] HWDATA;  // ../RTL/cmsdk_mcu_system.v(84)
  output HWRITE;  // ../RTL/cmsdk_mcu_system.v(83)
  output LOCKUP;  // ../RTL/cmsdk_mcu_system.v(109)
  output LOCKUPRESET;  // ../RTL/cmsdk_mcu_system.v(110)
  output PMUENABLE;  // ../RTL/cmsdk_mcu_system.v(111)
  output SLEEPDEEP;  // ../RTL/cmsdk_mcu_system.v(106)
  output SLEEPHOLDACKn;  // ../RTL/cmsdk_mcu_system.v(121)
  output SLEEPING;  // ../RTL/cmsdk_mcu_system.v(105)
  output SWDO;  // ../RTL/cmsdk_mcu_system.v(165)
  output SWDOEN;  // ../RTL/cmsdk_mcu_system.v(166)
  output SYSRESETREQ;  // ../RTL/cmsdk_mcu_system.v(107)
  output TDO;  // ../RTL/cmsdk_mcu_system.v(167)
  output WAKEUP;  // ../RTL/cmsdk_mcu_system.v(115)
  output WDOGRESETREQ;  // ../RTL/cmsdk_mcu_system.v(108)
  output WICENACK;  // ../RTL/cmsdk_mcu_system.v(117)
  output boot_hsel;  // ../RTL/cmsdk_mcu_system.v(98)
  output flash_hsel;  // ../RTL/cmsdk_mcu_system.v(87)
  output nTDOEN;  // ../RTL/cmsdk_mcu_system.v(168)
  output [15:0] p0_altfunc;  // ../RTL/cmsdk_mcu_system.v(147)
  output [15:0] p0_out;  // ../RTL/cmsdk_mcu_system.v(145)
  output [15:0] p0_outen;  // ../RTL/cmsdk_mcu_system.v(146)
  output [15:0] p1_altfunc;  // ../RTL/cmsdk_mcu_system.v(151)
  output [15:0] p1_out;  // ../RTL/cmsdk_mcu_system.v(149)
  output [15:0] p1_outen;  // ../RTL/cmsdk_mcu_system.v(150)
  output sram_hsel;  // ../RTL/cmsdk_mcu_system.v(92)
  output uart0_txd;  // ../RTL/cmsdk_mcu_system.v(124)
  output uart0_txen;  // ../RTL/cmsdk_mcu_system.v(125)
  inout [7:0] b_pad_gpio_porta;  // ../RTL/cmsdk_mcu_system.v(139)

  parameter BASEADDR_GPIO0 = 32'b01000000000000010000000000000000;
  parameter BASEADDR_GPIO1 = 32'b01000000000000010001000000000000;
  parameter BASEADDR_SYSROMTABLE = 32'b11110000000000000000000000000000;
  parameter BE = 0;
  parameter BKPT = 4;
  parameter BOOT_LOADER_PRESENT = 0;
  parameter BOOT_MEM_TYPE = 0;
  parameter CLKGATE_PRESENT = 0;
  parameter DBG = 1;
  parameter DMA_CHANNEL_NUM = 0;
  parameter INCLUDE_BITBAND = 0;
  parameter INCLUDE_DMA = 0;
  parameter INCLUDE_JTAG = 0;
  parameter NUMIRQ = 32;
  parameter SMUL = 0;
  parameter SYST = 1;
  parameter WIC = 1;
  parameter WICLINES = 34;
  parameter WPT = 2;
  wire [31:0] HRDATAMTB;  // ../RTL/cmsdk_mcu_system.v(276)
  wire [31:0] apbsubsys_interrupt;  // ../RTL/cmsdk_mcu_system.v(307)
  wire [31:0] apbsys_hrdata;  // ../RTL/cmsdk_mcu_system.v(252)
  wire [31:0] cm0_haddr;  // ../RTL/cmsdk_mcu_system.v(197)
  wire [2:0] cm0_hburst;  // ../RTL/cmsdk_mcu_system.v(198)
  wire [3:0] cm0_hprot;  // ../RTL/cmsdk_mcu_system.v(200)
  wire [31:0] cm0_hrdata;  // ../RTL/cmsdk_mcu_system.v(205)
  wire [2:0] cm0_hsize;  // ../RTL/cmsdk_mcu_system.v(201)
  wire [1:0] cm0_htrans;  // ../RTL/cmsdk_mcu_system.v(202)
  wire [31:0] cm0_hwdata;  // ../RTL/cmsdk_mcu_system.v(203)
  wire [31:0] cm_haddr;  // ../RTL/cmsdk_mcu_system.v(183)
  wire [2:0] cm_hburst;  // ../RTL/cmsdk_mcu_system.v(186)
  wire [3:0] cm_hprot;  // ../RTL/cmsdk_mcu_system.v(187)
  wire [31:0] cm_hrdata;  // ../RTL/cmsdk_mcu_system.v(192)
  wire [2:0] cm_hsize;  // ../RTL/cmsdk_mcu_system.v(185)
  wire [1:0] cm_htrans;  // ../RTL/cmsdk_mcu_system.v(184)
  wire [31:0] cm_hwdata;  // ../RTL/cmsdk_mcu_system.v(191)
  wire [31:0] defslv_hrdata;  // ../RTL/cmsdk_mcu_system.v(247)
  wire [31:0] dmac_prdata;  // ../RTL/cmsdk_mcu_system.v(227)
  wire [31:0] gpio0_hrdata;  // ../RTL/cmsdk_mcu_system.v(257)
  wire [15:0] gpio0_intr;  // ../RTL/cmsdk_mcu_system.v(304)
  wire [31:0] gpio1_hrdata;  // ../RTL/cmsdk_mcu_system.v(262)
  wire [31:0] intisr_cm0;  // ../RTL/cmsdk_mcu_system.v(270)
  wire [31:0] sys_haddr;  // ../RTL/cmsdk_mcu_system.v(231)
  wire [2:0] sys_hburst;  // ../RTL/cmsdk_mcu_system.v(234)
  wire [3:0] sys_hprot;  // ../RTL/cmsdk_mcu_system.v(235)
  wire [31:0] sys_hrdata;  // ../RTL/cmsdk_mcu_system.v(240)
  wire [2:0] sys_hsize;  // ../RTL/cmsdk_mcu_system.v(233)
  wire [1:0] sys_htrans;  // ../RTL/cmsdk_mcu_system.v(232)
  wire [31:0] sys_hwdata;  // ../RTL/cmsdk_mcu_system.v(239)
  wire [31:0] sysctrl_hrdata;  // ../RTL/cmsdk_mcu_system.v(267)
  wire [31:0] sysrom_hrdata;  // ../RTL/cmsdk_mcu_system.v(288)
  wire DMA_DONE;  // ../RTL/cmsdk_mcu_system.v(324)
  wire HCLKSYS;  // ../RTL/cmsdk_mcu_system.v(180)
  wire HREADYOUTMTB;  // ../RTL/cmsdk_mcu_system.v(275)
  wire HRESPMTB;  // ../RTL/cmsdk_mcu_system.v(277)
  wire HSELMTB;  // ../RTL/cmsdk_mcu_system.v(274)
  wire RXEV;  // ../RTL/cmsdk_mcu_system.v(326)
  wire STCLKEN;  // ../RTL/cmsdk_mcu_system.v(282)
  wire apbsys_hreadyout;  // ../RTL/cmsdk_mcu_system.v(251)
  wire apbsys_hresp;  // ../RTL/cmsdk_mcu_system.v(253)
  wire apbsys_hsel;  // ../RTL/cmsdk_mcu_system.v(250)
  wire cm0_hmastlock;  // ../RTL/cmsdk_mcu_system.v(199)
  wire cm0_hready;  // ../RTL/cmsdk_mcu_system.v(206)
  wire cm0_hresp;  // ../RTL/cmsdk_mcu_system.v(207)
  wire cm0_hwrite;  // ../RTL/cmsdk_mcu_system.v(204)
  wire cm_hmastlock;  // ../RTL/cmsdk_mcu_system.v(188)
  wire cm_hready;  // ../RTL/cmsdk_mcu_system.v(193)
  wire cm_hreadyout;  // ../RTL/cmsdk_mcu_system.v(194)
  wire cm_hresp;  // ../RTL/cmsdk_mcu_system.v(195)
  wire cm_hwrite;  // ../RTL/cmsdk_mcu_system.v(190)
  wire cpu0cdbgpwrupack;  // ../RTL/cmsdk_mcu_system.v(343)
  wire cpu0cdbgpwrupreq;  // ../RTL/cmsdk_mcu_system.v(342)
  wire defslv_hreadyout;  // ../RTL/cmsdk_mcu_system.v(246)
  wire defslv_hresp;  // ../RTL/cmsdk_mcu_system.v(248)
  wire defslv_hsel;  // ../RTL/cmsdk_mcu_system.v(245)
  wire dma_err;  // ../RTL/cmsdk_mcu_system.v(308)
  wire dmac_pready;  // ../RTL/cmsdk_mcu_system.v(225)
  wire dmac_pslverr;  // ../RTL/cmsdk_mcu_system.v(226)
  wire gpio0_combintr;  // ../RTL/cmsdk_mcu_system.v(305)
  wire gpio0_hreadyout;  // ../RTL/cmsdk_mcu_system.v(256)
  wire gpio0_hresp;  // ../RTL/cmsdk_mcu_system.v(258)
  wire gpio0_hsel;  // ../RTL/cmsdk_mcu_system.v(255)
  wire gpio1_combintr;  // ../RTL/cmsdk_mcu_system.v(306)
  wire gpio1_hreadyout;  // ../RTL/cmsdk_mcu_system.v(261)
  wire gpio1_hresp;  // ../RTL/cmsdk_mcu_system.v(263)
  wire gpio1_hsel;  // ../RTL/cmsdk_mcu_system.v(260)
  wire intnmi_cm0;  // ../RTL/cmsdk_mcu_system.v(271)
  wire n0;
  wire n1;
  wire n2;
  wire n3;
  wire n4;
  wire n5;
  wire remap_ctrl;  // ../RTL/cmsdk_mcu_system.v(301)
  wire sys_hmastlock;  // ../RTL/cmsdk_mcu_system.v(237)
  wire sys_hready;  // ../RTL/cmsdk_mcu_system.v(241)
  wire sys_hreadyout;  // ../RTL/cmsdk_mcu_system.v(242)
  wire sys_hresp;  // ../RTL/cmsdk_mcu_system.v(243)
  wire sys_hwrite;  // ../RTL/cmsdk_mcu_system.v(238)
  wire sysctrl_hreadyout;  // ../RTL/cmsdk_mcu_system.v(266)
  wire sysctrl_hresp;  // ../RTL/cmsdk_mcu_system.v(268)
  wire sysctrl_hsel;  // ../RTL/cmsdk_mcu_system.v(265)
  wire sysrom_hreadyout;  // ../RTL/cmsdk_mcu_system.v(287)
  wire sysrom_hresp;  // ../RTL/cmsdk_mcu_system.v(289)
  wire sysrom_hsel;  // ../RTL/cmsdk_mcu_system.v(286)
  wire watchdog_interrupt;  // ../RTL/cmsdk_mcu_system.v(309)

  buf u10 (cm_haddr[0], cm0_haddr[0]);  // ../RTL/cmsdk_mcu_system.v(515)
  buf u100 (dmac_prdata[18], 1'b0);  // ../RTL/cmsdk_mcu_system.v(1067)
  buf u101 (dmac_prdata[19], 1'b0);  // ../RTL/cmsdk_mcu_system.v(1067)
  buf u102 (dmac_prdata[20], 1'b0);  // ../RTL/cmsdk_mcu_system.v(1067)
  buf u103 (dmac_prdata[21], 1'b0);  // ../RTL/cmsdk_mcu_system.v(1067)
  buf u104 (dmac_prdata[22], 1'b0);  // ../RTL/cmsdk_mcu_system.v(1067)
  buf u105 (dmac_prdata[23], 1'b0);  // ../RTL/cmsdk_mcu_system.v(1067)
  buf u106 (dmac_prdata[24], 1'b0);  // ../RTL/cmsdk_mcu_system.v(1067)
  buf u107 (dmac_prdata[25], 1'b0);  // ../RTL/cmsdk_mcu_system.v(1067)
  buf u108 (dmac_prdata[26], 1'b0);  // ../RTL/cmsdk_mcu_system.v(1067)
  buf u109 (dmac_prdata[27], 1'b0);  // ../RTL/cmsdk_mcu_system.v(1067)
  buf u11 (cm_htrans[0], cm0_htrans[0]);  // ../RTL/cmsdk_mcu_system.v(516)
  buf u110 (dmac_prdata[28], 1'b0);  // ../RTL/cmsdk_mcu_system.v(1067)
  buf u111 (dmac_prdata[29], 1'b0);  // ../RTL/cmsdk_mcu_system.v(1067)
  buf u112 (dmac_prdata[30], 1'b0);  // ../RTL/cmsdk_mcu_system.v(1067)
  buf u113 (dmac_prdata[31], 1'b0);  // ../RTL/cmsdk_mcu_system.v(1067)
  buf u114 (HWDATA[1], sys_hwdata[1]);  // ../RTL/cmsdk_mcu_system.v(997)
  buf u115 (HWDATA[2], sys_hwdata[2]);  // ../RTL/cmsdk_mcu_system.v(997)
  buf u116 (HWDATA[3], sys_hwdata[3]);  // ../RTL/cmsdk_mcu_system.v(997)
  buf u117 (HWDATA[4], sys_hwdata[4]);  // ../RTL/cmsdk_mcu_system.v(997)
  buf u118 (HWDATA[5], sys_hwdata[5]);  // ../RTL/cmsdk_mcu_system.v(997)
  buf u119 (HWDATA[6], sys_hwdata[6]);  // ../RTL/cmsdk_mcu_system.v(997)
  buf u12 (cm_hsize[0], cm0_hsize[0]);  // ../RTL/cmsdk_mcu_system.v(517)
  buf u120 (HWDATA[7], sys_hwdata[7]);  // ../RTL/cmsdk_mcu_system.v(997)
  buf u121 (HWDATA[8], sys_hwdata[8]);  // ../RTL/cmsdk_mcu_system.v(997)
  buf u122 (HWDATA[9], sys_hwdata[9]);  // ../RTL/cmsdk_mcu_system.v(997)
  buf u123 (HWDATA[10], sys_hwdata[10]);  // ../RTL/cmsdk_mcu_system.v(997)
  buf u124 (HWDATA[11], sys_hwdata[11]);  // ../RTL/cmsdk_mcu_system.v(997)
  buf u125 (HWDATA[12], sys_hwdata[12]);  // ../RTL/cmsdk_mcu_system.v(997)
  buf u126 (HWDATA[13], sys_hwdata[13]);  // ../RTL/cmsdk_mcu_system.v(997)
  buf u127 (HWDATA[14], sys_hwdata[14]);  // ../RTL/cmsdk_mcu_system.v(997)
  buf u128 (HWDATA[15], sys_hwdata[15]);  // ../RTL/cmsdk_mcu_system.v(997)
  buf u129 (HWDATA[16], sys_hwdata[16]);  // ../RTL/cmsdk_mcu_system.v(997)
  buf u13 (cm_hburst[0], cm0_hburst[0]);  // ../RTL/cmsdk_mcu_system.v(518)
  buf u130 (HWDATA[17], sys_hwdata[17]);  // ../RTL/cmsdk_mcu_system.v(997)
  buf u131 (HWDATA[18], sys_hwdata[18]);  // ../RTL/cmsdk_mcu_system.v(997)
  buf u132 (HWDATA[19], sys_hwdata[19]);  // ../RTL/cmsdk_mcu_system.v(997)
  buf u133 (HWDATA[20], sys_hwdata[20]);  // ../RTL/cmsdk_mcu_system.v(997)
  buf u134 (HWDATA[21], sys_hwdata[21]);  // ../RTL/cmsdk_mcu_system.v(997)
  buf u135 (HWDATA[22], sys_hwdata[22]);  // ../RTL/cmsdk_mcu_system.v(997)
  buf u136 (HWDATA[23], sys_hwdata[23]);  // ../RTL/cmsdk_mcu_system.v(997)
  buf u137 (HWDATA[24], sys_hwdata[24]);  // ../RTL/cmsdk_mcu_system.v(997)
  buf u138 (HWDATA[25], sys_hwdata[25]);  // ../RTL/cmsdk_mcu_system.v(997)
  buf u139 (HWDATA[26], sys_hwdata[26]);  // ../RTL/cmsdk_mcu_system.v(997)
  buf u14 (intisr_cm0[4], apbsubsys_interrupt[4]);  // ../RTL/cmsdk_mcu_system.v(1088)
  buf u140 (HWDATA[27], sys_hwdata[27]);  // ../RTL/cmsdk_mcu_system.v(997)
  buf u141 (HWDATA[28], sys_hwdata[28]);  // ../RTL/cmsdk_mcu_system.v(997)
  buf u142 (HWDATA[29], sys_hwdata[29]);  // ../RTL/cmsdk_mcu_system.v(997)
  buf u143 (HWDATA[30], sys_hwdata[30]);  // ../RTL/cmsdk_mcu_system.v(997)
  buf u144 (HWDATA[31], sys_hwdata[31]);  // ../RTL/cmsdk_mcu_system.v(997)
  buf u145 (HSIZE[1], sys_hsize[1]);  // ../RTL/cmsdk_mcu_system.v(995)
  buf u146 (HSIZE[2], sys_hsize[2]);  // ../RTL/cmsdk_mcu_system.v(995)
  buf u147 (HTRANS[1], sys_htrans[1]);  // ../RTL/cmsdk_mcu_system.v(994)
  buf u148 (HADDR[1], sys_haddr[1]);  // ../RTL/cmsdk_mcu_system.v(993)
  buf u149 (HADDR[2], sys_haddr[2]);  // ../RTL/cmsdk_mcu_system.v(993)
  buf u15 (cm_hmastlock, cm0_hmastlock);  // ../RTL/cmsdk_mcu_system.v(521)
  buf u150 (HADDR[3], sys_haddr[3]);  // ../RTL/cmsdk_mcu_system.v(993)
  buf u151 (HADDR[4], sys_haddr[4]);  // ../RTL/cmsdk_mcu_system.v(993)
  buf u152 (HADDR[5], sys_haddr[5]);  // ../RTL/cmsdk_mcu_system.v(993)
  buf u153 (HADDR[6], sys_haddr[6]);  // ../RTL/cmsdk_mcu_system.v(993)
  buf u154 (HADDR[7], sys_haddr[7]);  // ../RTL/cmsdk_mcu_system.v(993)
  buf u155 (HADDR[8], sys_haddr[8]);  // ../RTL/cmsdk_mcu_system.v(993)
  buf u156 (HADDR[9], sys_haddr[9]);  // ../RTL/cmsdk_mcu_system.v(993)
  buf u157 (HADDR[10], sys_haddr[10]);  // ../RTL/cmsdk_mcu_system.v(993)
  buf u158 (HADDR[11], sys_haddr[11]);  // ../RTL/cmsdk_mcu_system.v(993)
  buf u159 (HADDR[12], sys_haddr[12]);  // ../RTL/cmsdk_mcu_system.v(993)
  buf u16 (cm_hwrite, cm0_hwrite);  // ../RTL/cmsdk_mcu_system.v(522)
  buf u160 (HADDR[13], sys_haddr[13]);  // ../RTL/cmsdk_mcu_system.v(993)
  buf u161 (HADDR[14], sys_haddr[14]);  // ../RTL/cmsdk_mcu_system.v(993)
  buf u162 (HADDR[15], sys_haddr[15]);  // ../RTL/cmsdk_mcu_system.v(993)
  buf u163 (HADDR[16], sys_haddr[16]);  // ../RTL/cmsdk_mcu_system.v(993)
  buf u164 (HADDR[17], sys_haddr[17]);  // ../RTL/cmsdk_mcu_system.v(993)
  buf u165 (HADDR[18], sys_haddr[18]);  // ../RTL/cmsdk_mcu_system.v(993)
  buf u166 (HADDR[19], sys_haddr[19]);  // ../RTL/cmsdk_mcu_system.v(993)
  buf u167 (HADDR[20], sys_haddr[20]);  // ../RTL/cmsdk_mcu_system.v(993)
  buf u168 (HADDR[21], sys_haddr[21]);  // ../RTL/cmsdk_mcu_system.v(993)
  buf u169 (HADDR[22], sys_haddr[22]);  // ../RTL/cmsdk_mcu_system.v(993)
  buf u17 (cm_hprot[0], cm0_hprot[0]);  // ../RTL/cmsdk_mcu_system.v(519)
  buf u170 (HADDR[23], sys_haddr[23]);  // ../RTL/cmsdk_mcu_system.v(993)
  buf u171 (HADDR[24], sys_haddr[24]);  // ../RTL/cmsdk_mcu_system.v(993)
  buf u172 (HADDR[25], sys_haddr[25]);  // ../RTL/cmsdk_mcu_system.v(993)
  buf u173 (HADDR[26], sys_haddr[26]);  // ../RTL/cmsdk_mcu_system.v(993)
  buf u174 (HADDR[27], sys_haddr[27]);  // ../RTL/cmsdk_mcu_system.v(993)
  buf u175 (HADDR[28], sys_haddr[28]);  // ../RTL/cmsdk_mcu_system.v(993)
  buf u176 (HADDR[29], sys_haddr[29]);  // ../RTL/cmsdk_mcu_system.v(993)
  buf u177 (HADDR[30], sys_haddr[30]);  // ../RTL/cmsdk_mcu_system.v(993)
  buf u178 (HADDR[31], sys_haddr[31]);  // ../RTL/cmsdk_mcu_system.v(993)
  buf u179 (defslv_hrdata[1], 1'b0);  // ../RTL/cmsdk_mcu_system.v(734)
  buf u18 (cm_hready, cm0_hready);  // ../RTL/cmsdk_mcu_system.v(524)
  buf u180 (defslv_hrdata[2], 1'b0);  // ../RTL/cmsdk_mcu_system.v(734)
  buf u181 (defslv_hrdata[3], 1'b0);  // ../RTL/cmsdk_mcu_system.v(734)
  buf u182 (defslv_hrdata[4], 1'b0);  // ../RTL/cmsdk_mcu_system.v(734)
  buf u183 (defslv_hrdata[5], 1'b0);  // ../RTL/cmsdk_mcu_system.v(734)
  buf u184 (defslv_hrdata[6], 1'b0);  // ../RTL/cmsdk_mcu_system.v(734)
  buf u185 (defslv_hrdata[7], 1'b0);  // ../RTL/cmsdk_mcu_system.v(734)
  buf u186 (defslv_hrdata[8], 1'b0);  // ../RTL/cmsdk_mcu_system.v(734)
  buf u187 (defslv_hrdata[9], 1'b0);  // ../RTL/cmsdk_mcu_system.v(734)
  buf u188 (defslv_hrdata[10], 1'b0);  // ../RTL/cmsdk_mcu_system.v(734)
  buf u189 (defslv_hrdata[11], 1'b0);  // ../RTL/cmsdk_mcu_system.v(734)
  buf u19 (cm_hwdata[0], cm0_hwdata[0]);  // ../RTL/cmsdk_mcu_system.v(523)
  buf u190 (defslv_hrdata[12], 1'b0);  // ../RTL/cmsdk_mcu_system.v(734)
  buf u191 (defslv_hrdata[13], 1'b0);  // ../RTL/cmsdk_mcu_system.v(734)
  buf u192 (defslv_hrdata[14], 1'b0);  // ../RTL/cmsdk_mcu_system.v(734)
  buf u193 (defslv_hrdata[15], 1'b0);  // ../RTL/cmsdk_mcu_system.v(734)
  buf u194 (defslv_hrdata[16], 1'b0);  // ../RTL/cmsdk_mcu_system.v(734)
  buf u195 (defslv_hrdata[17], 1'b0);  // ../RTL/cmsdk_mcu_system.v(734)
  buf u196 (defslv_hrdata[18], 1'b0);  // ../RTL/cmsdk_mcu_system.v(734)
  buf u197 (defslv_hrdata[19], 1'b0);  // ../RTL/cmsdk_mcu_system.v(734)
  buf u198 (defslv_hrdata[20], 1'b0);  // ../RTL/cmsdk_mcu_system.v(734)
  buf u199 (defslv_hrdata[21], 1'b0);  // ../RTL/cmsdk_mcu_system.v(734)
  buf u2 (intisr_cm0[8], apbsubsys_interrupt[8]);  // ../RTL/cmsdk_mcu_system.v(1088)
  buf u20 (cm0_hready, cm_hreadyout);  // ../RTL/cmsdk_mcu_system.v(526)
  buf u200 (defslv_hrdata[22], 1'b0);  // ../RTL/cmsdk_mcu_system.v(734)
  buf u201 (defslv_hrdata[23], 1'b0);  // ../RTL/cmsdk_mcu_system.v(734)
  buf u202 (defslv_hrdata[24], 1'b0);  // ../RTL/cmsdk_mcu_system.v(734)
  buf u203 (defslv_hrdata[25], 1'b0);  // ../RTL/cmsdk_mcu_system.v(734)
  buf u204 (defslv_hrdata[26], 1'b0);  // ../RTL/cmsdk_mcu_system.v(734)
  buf u205 (defslv_hrdata[27], 1'b0);  // ../RTL/cmsdk_mcu_system.v(734)
  buf u206 (defslv_hrdata[28], 1'b0);  // ../RTL/cmsdk_mcu_system.v(734)
  buf u207 (defslv_hrdata[29], 1'b0);  // ../RTL/cmsdk_mcu_system.v(734)
  buf u208 (defslv_hrdata[30], 1'b0);  // ../RTL/cmsdk_mcu_system.v(734)
  buf u209 (defslv_hrdata[31], 1'b0);  // ../RTL/cmsdk_mcu_system.v(734)
  buf u21 (cm0_hresp, cm_hresp);  // ../RTL/cmsdk_mcu_system.v(527)
  buf u210 (cm_hrdata[1], sys_hrdata[1]);  // ../RTL/cmsdk_mcu_system.v(625)
  buf u211 (cm_hrdata[2], sys_hrdata[2]);  // ../RTL/cmsdk_mcu_system.v(625)
  buf u212 (cm_hrdata[3], sys_hrdata[3]);  // ../RTL/cmsdk_mcu_system.v(625)
  buf u213 (cm_hrdata[4], sys_hrdata[4]);  // ../RTL/cmsdk_mcu_system.v(625)
  buf u214 (cm_hrdata[5], sys_hrdata[5]);  // ../RTL/cmsdk_mcu_system.v(625)
  buf u215 (cm_hrdata[6], sys_hrdata[6]);  // ../RTL/cmsdk_mcu_system.v(625)
  buf u216 (cm_hrdata[7], sys_hrdata[7]);  // ../RTL/cmsdk_mcu_system.v(625)
  buf u217 (cm_hrdata[8], sys_hrdata[8]);  // ../RTL/cmsdk_mcu_system.v(625)
  buf u218 (cm_hrdata[9], sys_hrdata[9]);  // ../RTL/cmsdk_mcu_system.v(625)
  buf u219 (cm_hrdata[10], sys_hrdata[10]);  // ../RTL/cmsdk_mcu_system.v(625)
  buf u22 (cm0_hrdata[0], cm_hrdata[0]);  // ../RTL/cmsdk_mcu_system.v(525)
  buf u220 (cm_hrdata[11], sys_hrdata[11]);  // ../RTL/cmsdk_mcu_system.v(625)
  buf u221 (cm_hrdata[12], sys_hrdata[12]);  // ../RTL/cmsdk_mcu_system.v(625)
  buf u222 (cm_hrdata[13], sys_hrdata[13]);  // ../RTL/cmsdk_mcu_system.v(625)
  buf u223 (cm_hrdata[14], sys_hrdata[14]);  // ../RTL/cmsdk_mcu_system.v(625)
  buf u224 (cm_hrdata[15], sys_hrdata[15]);  // ../RTL/cmsdk_mcu_system.v(625)
  buf u225 (cm_hrdata[16], sys_hrdata[16]);  // ../RTL/cmsdk_mcu_system.v(625)
  buf u226 (cm_hrdata[17], sys_hrdata[17]);  // ../RTL/cmsdk_mcu_system.v(625)
  buf u227 (cm_hrdata[18], sys_hrdata[18]);  // ../RTL/cmsdk_mcu_system.v(625)
  buf u228 (cm_hrdata[19], sys_hrdata[19]);  // ../RTL/cmsdk_mcu_system.v(625)
  buf u229 (cm_hrdata[20], sys_hrdata[20]);  // ../RTL/cmsdk_mcu_system.v(625)
  buf u23 (sys_haddr[0], cm_haddr[0]);  // ../RTL/cmsdk_mcu_system.v(615)
  buf u230 (cm_hrdata[21], sys_hrdata[21]);  // ../RTL/cmsdk_mcu_system.v(625)
  buf u231 (cm_hrdata[22], sys_hrdata[22]);  // ../RTL/cmsdk_mcu_system.v(625)
  buf u232 (cm_hrdata[23], sys_hrdata[23]);  // ../RTL/cmsdk_mcu_system.v(625)
  buf u233 (cm_hrdata[24], sys_hrdata[24]);  // ../RTL/cmsdk_mcu_system.v(625)
  buf u234 (cm_hrdata[25], sys_hrdata[25]);  // ../RTL/cmsdk_mcu_system.v(625)
  buf u235 (cm_hrdata[26], sys_hrdata[26]);  // ../RTL/cmsdk_mcu_system.v(625)
  buf u236 (cm_hrdata[27], sys_hrdata[27]);  // ../RTL/cmsdk_mcu_system.v(625)
  buf u237 (cm_hrdata[28], sys_hrdata[28]);  // ../RTL/cmsdk_mcu_system.v(625)
  buf u238 (cm_hrdata[29], sys_hrdata[29]);  // ../RTL/cmsdk_mcu_system.v(625)
  buf u239 (cm_hrdata[30], sys_hrdata[30]);  // ../RTL/cmsdk_mcu_system.v(625)
  buf u24 (sys_htrans[0], cm_htrans[0]);  // ../RTL/cmsdk_mcu_system.v(616)
  buf u240 (cm_hrdata[31], sys_hrdata[31]);  // ../RTL/cmsdk_mcu_system.v(625)
  buf u241 (sys_hwdata[1], cm_hwdata[1]);  // ../RTL/cmsdk_mcu_system.v(623)
  buf u242 (sys_hwdata[2], cm_hwdata[2]);  // ../RTL/cmsdk_mcu_system.v(623)
  buf u243 (sys_hwdata[3], cm_hwdata[3]);  // ../RTL/cmsdk_mcu_system.v(623)
  buf u244 (sys_hwdata[4], cm_hwdata[4]);  // ../RTL/cmsdk_mcu_system.v(623)
  buf u245 (sys_hwdata[5], cm_hwdata[5]);  // ../RTL/cmsdk_mcu_system.v(623)
  buf u246 (sys_hwdata[6], cm_hwdata[6]);  // ../RTL/cmsdk_mcu_system.v(623)
  buf u247 (sys_hwdata[7], cm_hwdata[7]);  // ../RTL/cmsdk_mcu_system.v(623)
  buf u248 (sys_hwdata[8], cm_hwdata[8]);  // ../RTL/cmsdk_mcu_system.v(623)
  buf u249 (sys_hwdata[9], cm_hwdata[9]);  // ../RTL/cmsdk_mcu_system.v(623)
  buf u25 (sys_hsize[0], cm_hsize[0]);  // ../RTL/cmsdk_mcu_system.v(617)
  buf u250 (sys_hwdata[10], cm_hwdata[10]);  // ../RTL/cmsdk_mcu_system.v(623)
  buf u251 (sys_hwdata[11], cm_hwdata[11]);  // ../RTL/cmsdk_mcu_system.v(623)
  buf u252 (sys_hwdata[12], cm_hwdata[12]);  // ../RTL/cmsdk_mcu_system.v(623)
  buf u253 (sys_hwdata[13], cm_hwdata[13]);  // ../RTL/cmsdk_mcu_system.v(623)
  buf u254 (sys_hwdata[14], cm_hwdata[14]);  // ../RTL/cmsdk_mcu_system.v(623)
  buf u255 (sys_hwdata[15], cm_hwdata[15]);  // ../RTL/cmsdk_mcu_system.v(623)
  buf u256 (sys_hwdata[16], cm_hwdata[16]);  // ../RTL/cmsdk_mcu_system.v(623)
  buf u257 (sys_hwdata[17], cm_hwdata[17]);  // ../RTL/cmsdk_mcu_system.v(623)
  buf u258 (sys_hwdata[18], cm_hwdata[18]);  // ../RTL/cmsdk_mcu_system.v(623)
  buf u259 (sys_hwdata[19], cm_hwdata[19]);  // ../RTL/cmsdk_mcu_system.v(623)
  buf u26 (sys_hburst[0], cm_hburst[0]);  // ../RTL/cmsdk_mcu_system.v(618)
  buf u260 (sys_hwdata[20], cm_hwdata[20]);  // ../RTL/cmsdk_mcu_system.v(623)
  buf u261 (sys_hwdata[21], cm_hwdata[21]);  // ../RTL/cmsdk_mcu_system.v(623)
  buf u262 (sys_hwdata[22], cm_hwdata[22]);  // ../RTL/cmsdk_mcu_system.v(623)
  buf u263 (sys_hwdata[23], cm_hwdata[23]);  // ../RTL/cmsdk_mcu_system.v(623)
  buf u264 (sys_hwdata[24], cm_hwdata[24]);  // ../RTL/cmsdk_mcu_system.v(623)
  buf u265 (sys_hwdata[25], cm_hwdata[25]);  // ../RTL/cmsdk_mcu_system.v(623)
  buf u266 (sys_hwdata[26], cm_hwdata[26]);  // ../RTL/cmsdk_mcu_system.v(623)
  buf u267 (sys_hwdata[27], cm_hwdata[27]);  // ../RTL/cmsdk_mcu_system.v(623)
  buf u268 (sys_hwdata[28], cm_hwdata[28]);  // ../RTL/cmsdk_mcu_system.v(623)
  buf u269 (sys_hwdata[29], cm_hwdata[29]);  // ../RTL/cmsdk_mcu_system.v(623)
  buf u27 (intisr_cm0[3], apbsubsys_interrupt[3]);  // ../RTL/cmsdk_mcu_system.v(1088)
  buf u270 (sys_hwdata[30], cm_hwdata[30]);  // ../RTL/cmsdk_mcu_system.v(623)
  buf u271 (sys_hwdata[31], cm_hwdata[31]);  // ../RTL/cmsdk_mcu_system.v(623)
  buf u272 (sys_hprot[1], cm_hprot[1]);  // ../RTL/cmsdk_mcu_system.v(619)
  buf u273 (sys_hprot[2], cm_hprot[2]);  // ../RTL/cmsdk_mcu_system.v(619)
  buf u274 (sys_hprot[3], cm_hprot[3]);  // ../RTL/cmsdk_mcu_system.v(619)
  buf u275 (sys_hburst[1], cm_hburst[1]);  // ../RTL/cmsdk_mcu_system.v(618)
  buf u276 (sys_hburst[2], cm_hburst[2]);  // ../RTL/cmsdk_mcu_system.v(618)
  buf u277 (sys_hsize[1], cm_hsize[1]);  // ../RTL/cmsdk_mcu_system.v(617)
  buf u278 (sys_hsize[2], cm_hsize[2]);  // ../RTL/cmsdk_mcu_system.v(617)
  buf u279 (sys_htrans[1], cm_htrans[1]);  // ../RTL/cmsdk_mcu_system.v(616)
  buf u28 (sys_hmastlock, cm_hmastlock);  // ../RTL/cmsdk_mcu_system.v(621)
  buf u280 (sys_haddr[1], cm_haddr[1]);  // ../RTL/cmsdk_mcu_system.v(615)
  buf u281 (sys_haddr[2], cm_haddr[2]);  // ../RTL/cmsdk_mcu_system.v(615)
  buf u282 (sys_haddr[3], cm_haddr[3]);  // ../RTL/cmsdk_mcu_system.v(615)
  buf u283 (sys_haddr[4], cm_haddr[4]);  // ../RTL/cmsdk_mcu_system.v(615)
  buf u284 (sys_haddr[5], cm_haddr[5]);  // ../RTL/cmsdk_mcu_system.v(615)
  buf u285 (sys_haddr[6], cm_haddr[6]);  // ../RTL/cmsdk_mcu_system.v(615)
  buf u286 (sys_haddr[7], cm_haddr[7]);  // ../RTL/cmsdk_mcu_system.v(615)
  buf u287 (sys_haddr[8], cm_haddr[8]);  // ../RTL/cmsdk_mcu_system.v(615)
  buf u288 (sys_haddr[9], cm_haddr[9]);  // ../RTL/cmsdk_mcu_system.v(615)
  buf u289 (sys_haddr[10], cm_haddr[10]);  // ../RTL/cmsdk_mcu_system.v(615)
  buf u29 (sys_hwrite, cm_hwrite);  // ../RTL/cmsdk_mcu_system.v(622)
  buf u290 (sys_haddr[11], cm_haddr[11]);  // ../RTL/cmsdk_mcu_system.v(615)
  buf u291 (sys_haddr[12], cm_haddr[12]);  // ../RTL/cmsdk_mcu_system.v(615)
  buf u292 (sys_haddr[13], cm_haddr[13]);  // ../RTL/cmsdk_mcu_system.v(615)
  buf u293 (sys_haddr[14], cm_haddr[14]);  // ../RTL/cmsdk_mcu_system.v(615)
  buf u294 (sys_haddr[15], cm_haddr[15]);  // ../RTL/cmsdk_mcu_system.v(615)
  buf u295 (sys_haddr[16], cm_haddr[16]);  // ../RTL/cmsdk_mcu_system.v(615)
  buf u296 (sys_haddr[17], cm_haddr[17]);  // ../RTL/cmsdk_mcu_system.v(615)
  buf u297 (sys_haddr[18], cm_haddr[18]);  // ../RTL/cmsdk_mcu_system.v(615)
  buf u298 (sys_haddr[19], cm_haddr[19]);  // ../RTL/cmsdk_mcu_system.v(615)
  buf u299 (sys_haddr[20], cm_haddr[20]);  // ../RTL/cmsdk_mcu_system.v(615)
  buf u3 (intisr_cm0[5], apbsubsys_interrupt[5]);  // ../RTL/cmsdk_mcu_system.v(1088)
  buf u30 (sys_hprot[0], cm_hprot[0]);  // ../RTL/cmsdk_mcu_system.v(619)
  buf u300 (sys_haddr[21], cm_haddr[21]);  // ../RTL/cmsdk_mcu_system.v(615)
  buf u301 (sys_haddr[22], cm_haddr[22]);  // ../RTL/cmsdk_mcu_system.v(615)
  buf u302 (sys_haddr[23], cm_haddr[23]);  // ../RTL/cmsdk_mcu_system.v(615)
  buf u303 (sys_haddr[24], cm_haddr[24]);  // ../RTL/cmsdk_mcu_system.v(615)
  buf u304 (sys_haddr[25], cm_haddr[25]);  // ../RTL/cmsdk_mcu_system.v(615)
  buf u305 (sys_haddr[26], cm_haddr[26]);  // ../RTL/cmsdk_mcu_system.v(615)
  buf u306 (sys_haddr[27], cm_haddr[27]);  // ../RTL/cmsdk_mcu_system.v(615)
  buf u307 (sys_haddr[28], cm_haddr[28]);  // ../RTL/cmsdk_mcu_system.v(615)
  buf u308 (sys_haddr[29], cm_haddr[29]);  // ../RTL/cmsdk_mcu_system.v(615)
  buf u309 (sys_haddr[30], cm_haddr[30]);  // ../RTL/cmsdk_mcu_system.v(615)
  buf u31 (sys_hready, cm_hready);  // ../RTL/cmsdk_mcu_system.v(624)
  buf u310 (sys_haddr[31], cm_haddr[31]);  // ../RTL/cmsdk_mcu_system.v(615)
  buf u311 (cm0_hrdata[1], cm_hrdata[1]);  // ../RTL/cmsdk_mcu_system.v(525)
  buf u312 (cm0_hrdata[2], cm_hrdata[2]);  // ../RTL/cmsdk_mcu_system.v(525)
  buf u313 (cm0_hrdata[3], cm_hrdata[3]);  // ../RTL/cmsdk_mcu_system.v(525)
  buf u314 (cm0_hrdata[4], cm_hrdata[4]);  // ../RTL/cmsdk_mcu_system.v(525)
  buf u315 (cm0_hrdata[5], cm_hrdata[5]);  // ../RTL/cmsdk_mcu_system.v(525)
  buf u316 (cm0_hrdata[6], cm_hrdata[6]);  // ../RTL/cmsdk_mcu_system.v(525)
  buf u317 (cm0_hrdata[7], cm_hrdata[7]);  // ../RTL/cmsdk_mcu_system.v(525)
  buf u318 (cm0_hrdata[8], cm_hrdata[8]);  // ../RTL/cmsdk_mcu_system.v(525)
  buf u319 (cm0_hrdata[9], cm_hrdata[9]);  // ../RTL/cmsdk_mcu_system.v(525)
  buf u32 (sys_hwdata[0], cm_hwdata[0]);  // ../RTL/cmsdk_mcu_system.v(623)
  buf u320 (cm0_hrdata[10], cm_hrdata[10]);  // ../RTL/cmsdk_mcu_system.v(525)
  buf u321 (cm0_hrdata[11], cm_hrdata[11]);  // ../RTL/cmsdk_mcu_system.v(525)
  buf u322 (cm0_hrdata[12], cm_hrdata[12]);  // ../RTL/cmsdk_mcu_system.v(525)
  buf u323 (cm0_hrdata[13], cm_hrdata[13]);  // ../RTL/cmsdk_mcu_system.v(525)
  buf u324 (cm0_hrdata[14], cm_hrdata[14]);  // ../RTL/cmsdk_mcu_system.v(525)
  buf u325 (cm0_hrdata[15], cm_hrdata[15]);  // ../RTL/cmsdk_mcu_system.v(525)
  buf u326 (cm0_hrdata[16], cm_hrdata[16]);  // ../RTL/cmsdk_mcu_system.v(525)
  buf u327 (cm0_hrdata[17], cm_hrdata[17]);  // ../RTL/cmsdk_mcu_system.v(525)
  buf u328 (cm0_hrdata[18], cm_hrdata[18]);  // ../RTL/cmsdk_mcu_system.v(525)
  buf u329 (cm0_hrdata[19], cm_hrdata[19]);  // ../RTL/cmsdk_mcu_system.v(525)
  buf u33 (cm_hreadyout, sys_hreadyout);  // ../RTL/cmsdk_mcu_system.v(626)
  buf u330 (cm0_hrdata[20], cm_hrdata[20]);  // ../RTL/cmsdk_mcu_system.v(525)
  buf u331 (cm0_hrdata[21], cm_hrdata[21]);  // ../RTL/cmsdk_mcu_system.v(525)
  buf u332 (cm0_hrdata[22], cm_hrdata[22]);  // ../RTL/cmsdk_mcu_system.v(525)
  buf u333 (cm0_hrdata[23], cm_hrdata[23]);  // ../RTL/cmsdk_mcu_system.v(525)
  buf u334 (cm0_hrdata[24], cm_hrdata[24]);  // ../RTL/cmsdk_mcu_system.v(525)
  buf u335 (cm0_hrdata[25], cm_hrdata[25]);  // ../RTL/cmsdk_mcu_system.v(525)
  buf u336 (cm0_hrdata[26], cm_hrdata[26]);  // ../RTL/cmsdk_mcu_system.v(525)
  buf u337 (cm0_hrdata[27], cm_hrdata[27]);  // ../RTL/cmsdk_mcu_system.v(525)
  buf u338 (cm0_hrdata[28], cm_hrdata[28]);  // ../RTL/cmsdk_mcu_system.v(525)
  buf u339 (cm0_hrdata[29], cm_hrdata[29]);  // ../RTL/cmsdk_mcu_system.v(525)
  buf u34 (cm_hresp, sys_hresp);  // ../RTL/cmsdk_mcu_system.v(627)
  buf u340 (cm0_hrdata[30], cm_hrdata[30]);  // ../RTL/cmsdk_mcu_system.v(525)
  buf u341 (cm0_hrdata[31], cm_hrdata[31]);  // ../RTL/cmsdk_mcu_system.v(525)
  buf u342 (cm_hwdata[1], cm0_hwdata[1]);  // ../RTL/cmsdk_mcu_system.v(523)
  buf u343 (cm_hwdata[2], cm0_hwdata[2]);  // ../RTL/cmsdk_mcu_system.v(523)
  buf u344 (cm_hwdata[3], cm0_hwdata[3]);  // ../RTL/cmsdk_mcu_system.v(523)
  buf u345 (cm_hwdata[4], cm0_hwdata[4]);  // ../RTL/cmsdk_mcu_system.v(523)
  buf u346 (cm_hwdata[5], cm0_hwdata[5]);  // ../RTL/cmsdk_mcu_system.v(523)
  buf u347 (cm_hwdata[6], cm0_hwdata[6]);  // ../RTL/cmsdk_mcu_system.v(523)
  buf u348 (cm_hwdata[7], cm0_hwdata[7]);  // ../RTL/cmsdk_mcu_system.v(523)
  buf u349 (cm_hwdata[8], cm0_hwdata[8]);  // ../RTL/cmsdk_mcu_system.v(523)
  buf u35 (intisr_cm0[2], apbsubsys_interrupt[2]);  // ../RTL/cmsdk_mcu_system.v(1088)
  buf u350 (cm_hwdata[9], cm0_hwdata[9]);  // ../RTL/cmsdk_mcu_system.v(523)
  buf u351 (cm_hwdata[10], cm0_hwdata[10]);  // ../RTL/cmsdk_mcu_system.v(523)
  buf u352 (cm_hwdata[11], cm0_hwdata[11]);  // ../RTL/cmsdk_mcu_system.v(523)
  buf u353 (cm_hwdata[12], cm0_hwdata[12]);  // ../RTL/cmsdk_mcu_system.v(523)
  buf u354 (cm_hwdata[13], cm0_hwdata[13]);  // ../RTL/cmsdk_mcu_system.v(523)
  buf u355 (cm_hwdata[14], cm0_hwdata[14]);  // ../RTL/cmsdk_mcu_system.v(523)
  buf u356 (cm_hwdata[15], cm0_hwdata[15]);  // ../RTL/cmsdk_mcu_system.v(523)
  buf u357 (cm_hwdata[16], cm0_hwdata[16]);  // ../RTL/cmsdk_mcu_system.v(523)
  buf u358 (cm_hwdata[17], cm0_hwdata[17]);  // ../RTL/cmsdk_mcu_system.v(523)
  buf u359 (cm_hwdata[18], cm0_hwdata[18]);  // ../RTL/cmsdk_mcu_system.v(523)
  buf u36 (cm_hrdata[0], sys_hrdata[0]);  // ../RTL/cmsdk_mcu_system.v(625)
  buf u360 (cm_hwdata[19], cm0_hwdata[19]);  // ../RTL/cmsdk_mcu_system.v(523)
  buf u361 (cm_hwdata[20], cm0_hwdata[20]);  // ../RTL/cmsdk_mcu_system.v(523)
  buf u362 (cm_hwdata[21], cm0_hwdata[21]);  // ../RTL/cmsdk_mcu_system.v(523)
  buf u363 (cm_hwdata[22], cm0_hwdata[22]);  // ../RTL/cmsdk_mcu_system.v(523)
  buf u364 (cm_hwdata[23], cm0_hwdata[23]);  // ../RTL/cmsdk_mcu_system.v(523)
  buf u365 (cm_hwdata[24], cm0_hwdata[24]);  // ../RTL/cmsdk_mcu_system.v(523)
  buf u366 (cm_hwdata[25], cm0_hwdata[25]);  // ../RTL/cmsdk_mcu_system.v(523)
  buf u367 (cm_hwdata[26], cm0_hwdata[26]);  // ../RTL/cmsdk_mcu_system.v(523)
  buf u368 (cm_hwdata[27], cm0_hwdata[27]);  // ../RTL/cmsdk_mcu_system.v(523)
  buf u369 (cm_hwdata[28], cm0_hwdata[28]);  // ../RTL/cmsdk_mcu_system.v(523)
  buf u37 (intisr_cm0[1], apbsubsys_interrupt[1]);  // ../RTL/cmsdk_mcu_system.v(1088)
  buf u370 (cm_hwdata[29], cm0_hwdata[29]);  // ../RTL/cmsdk_mcu_system.v(523)
  buf u371 (cm_hwdata[30], cm0_hwdata[30]);  // ../RTL/cmsdk_mcu_system.v(523)
  buf u372 (cm_hwdata[31], cm0_hwdata[31]);  // ../RTL/cmsdk_mcu_system.v(523)
  buf u373 (cm_hprot[1], cm0_hprot[1]);  // ../RTL/cmsdk_mcu_system.v(519)
  buf u374 (cm_hprot[2], cm0_hprot[2]);  // ../RTL/cmsdk_mcu_system.v(519)
  buf u375 (cm_hprot[3], cm0_hprot[3]);  // ../RTL/cmsdk_mcu_system.v(519)
  buf u376 (cm_hburst[1], cm0_hburst[1]);  // ../RTL/cmsdk_mcu_system.v(518)
  buf u377 (cm_hburst[2], cm0_hburst[2]);  // ../RTL/cmsdk_mcu_system.v(518)
  buf u378 (cm_hsize[1], cm0_hsize[1]);  // ../RTL/cmsdk_mcu_system.v(517)
  buf u379 (cm_hsize[2], cm0_hsize[2]);  // ../RTL/cmsdk_mcu_system.v(517)
  or u38 (intisr_cm0[31], apbsubsys_interrupt[31], gpio0_intr[15]);  // ../RTL/cmsdk_mcu_system.v(1089)
  buf u380 (cm_htrans[1], cm0_htrans[1]);  // ../RTL/cmsdk_mcu_system.v(516)
  buf u381 (cm_haddr[1], cm0_haddr[1]);  // ../RTL/cmsdk_mcu_system.v(515)
  buf u382 (cm_haddr[2], cm0_haddr[2]);  // ../RTL/cmsdk_mcu_system.v(515)
  buf u383 (cm_haddr[3], cm0_haddr[3]);  // ../RTL/cmsdk_mcu_system.v(515)
  buf u384 (cm_haddr[4], cm0_haddr[4]);  // ../RTL/cmsdk_mcu_system.v(515)
  buf u385 (cm_haddr[5], cm0_haddr[5]);  // ../RTL/cmsdk_mcu_system.v(515)
  buf u386 (cm_haddr[6], cm0_haddr[6]);  // ../RTL/cmsdk_mcu_system.v(515)
  buf u387 (cm_haddr[7], cm0_haddr[7]);  // ../RTL/cmsdk_mcu_system.v(515)
  buf u388 (cm_haddr[8], cm0_haddr[8]);  // ../RTL/cmsdk_mcu_system.v(515)
  buf u389 (cm_haddr[9], cm0_haddr[9]);  // ../RTL/cmsdk_mcu_system.v(515)
  buf u39 (defslv_hrdata[0], 1'b0);  // ../RTL/cmsdk_mcu_system.v(734)
  buf u390 (cm_haddr[10], cm0_haddr[10]);  // ../RTL/cmsdk_mcu_system.v(515)
  buf u391 (cm_haddr[11], cm0_haddr[11]);  // ../RTL/cmsdk_mcu_system.v(515)
  buf u392 (cm_haddr[12], cm0_haddr[12]);  // ../RTL/cmsdk_mcu_system.v(515)
  buf u393 (cm_haddr[13], cm0_haddr[13]);  // ../RTL/cmsdk_mcu_system.v(515)
  buf u394 (cm_haddr[14], cm0_haddr[14]);  // ../RTL/cmsdk_mcu_system.v(515)
  buf u395 (cm_haddr[15], cm0_haddr[15]);  // ../RTL/cmsdk_mcu_system.v(515)
  buf u396 (cm_haddr[16], cm0_haddr[16]);  // ../RTL/cmsdk_mcu_system.v(515)
  buf u397 (cm_haddr[17], cm0_haddr[17]);  // ../RTL/cmsdk_mcu_system.v(515)
  buf u398 (cm_haddr[18], cm0_haddr[18]);  // ../RTL/cmsdk_mcu_system.v(515)
  buf u399 (cm_haddr[19], cm0_haddr[19]);  // ../RTL/cmsdk_mcu_system.v(515)
  buf u4 (cpu0cdbgpwrupack, cpu0cdbgpwrupreq);  // ../RTL/cmsdk_mcu_system.v(344)
  buf u40 (HADDR[0], sys_haddr[0]);  // ../RTL/cmsdk_mcu_system.v(993)
  buf u400 (cm_haddr[20], cm0_haddr[20]);  // ../RTL/cmsdk_mcu_system.v(515)
  buf u401 (cm_haddr[21], cm0_haddr[21]);  // ../RTL/cmsdk_mcu_system.v(515)
  buf u402 (cm_haddr[22], cm0_haddr[22]);  // ../RTL/cmsdk_mcu_system.v(515)
  buf u403 (cm_haddr[23], cm0_haddr[23]);  // ../RTL/cmsdk_mcu_system.v(515)
  buf u404 (cm_haddr[24], cm0_haddr[24]);  // ../RTL/cmsdk_mcu_system.v(515)
  buf u405 (cm_haddr[25], cm0_haddr[25]);  // ../RTL/cmsdk_mcu_system.v(515)
  buf u406 (cm_haddr[26], cm0_haddr[26]);  // ../RTL/cmsdk_mcu_system.v(515)
  buf u407 (cm_haddr[27], cm0_haddr[27]);  // ../RTL/cmsdk_mcu_system.v(515)
  buf u408 (cm_haddr[28], cm0_haddr[28]);  // ../RTL/cmsdk_mcu_system.v(515)
  buf u409 (cm_haddr[29], cm0_haddr[29]);  // ../RTL/cmsdk_mcu_system.v(515)
  buf u41 (HTRANS[0], sys_htrans[0]);  // ../RTL/cmsdk_mcu_system.v(994)
  buf u410 (cm_haddr[30], cm0_haddr[30]);  // ../RTL/cmsdk_mcu_system.v(515)
  buf u411 (cm_haddr[31], cm0_haddr[31]);  // ../RTL/cmsdk_mcu_system.v(515)
  buf u412 (HRDATAMTB[1], 1'b0);  // ../RTL/cmsdk_mcu_system.v(466)
  buf u413 (HRDATAMTB[2], 1'b0);  // ../RTL/cmsdk_mcu_system.v(466)
  buf u414 (HRDATAMTB[3], 1'b0);  // ../RTL/cmsdk_mcu_system.v(466)
  buf u415 (HRDATAMTB[4], 1'b0);  // ../RTL/cmsdk_mcu_system.v(466)
  buf u416 (HRDATAMTB[5], 1'b0);  // ../RTL/cmsdk_mcu_system.v(466)
  buf u417 (HRDATAMTB[6], 1'b0);  // ../RTL/cmsdk_mcu_system.v(466)
  buf u418 (HRDATAMTB[7], 1'b0);  // ../RTL/cmsdk_mcu_system.v(466)
  buf u419 (HRDATAMTB[8], 1'b0);  // ../RTL/cmsdk_mcu_system.v(466)
  buf u42 (HWRITE, sys_hwrite);  // ../RTL/cmsdk_mcu_system.v(996)
  buf u420 (HRDATAMTB[9], 1'b0);  // ../RTL/cmsdk_mcu_system.v(466)
  buf u421 (HRDATAMTB[10], 1'b0);  // ../RTL/cmsdk_mcu_system.v(466)
  buf u422 (HRDATAMTB[11], 1'b0);  // ../RTL/cmsdk_mcu_system.v(466)
  buf u423 (HRDATAMTB[12], 1'b0);  // ../RTL/cmsdk_mcu_system.v(466)
  buf u424 (HRDATAMTB[13], 1'b0);  // ../RTL/cmsdk_mcu_system.v(466)
  buf u425 (HRDATAMTB[14], 1'b0);  // ../RTL/cmsdk_mcu_system.v(466)
  buf u426 (HRDATAMTB[15], 1'b0);  // ../RTL/cmsdk_mcu_system.v(466)
  buf u427 (HRDATAMTB[16], 1'b0);  // ../RTL/cmsdk_mcu_system.v(466)
  buf u428 (HRDATAMTB[17], 1'b0);  // ../RTL/cmsdk_mcu_system.v(466)
  buf u429 (HRDATAMTB[18], 1'b0);  // ../RTL/cmsdk_mcu_system.v(466)
  buf u43 (HSIZE[0], sys_hsize[0]);  // ../RTL/cmsdk_mcu_system.v(995)
  buf u430 (HRDATAMTB[19], 1'b0);  // ../RTL/cmsdk_mcu_system.v(466)
  buf u431 (HRDATAMTB[20], 1'b0);  // ../RTL/cmsdk_mcu_system.v(466)
  buf u432 (HRDATAMTB[21], 1'b0);  // ../RTL/cmsdk_mcu_system.v(466)
  buf u433 (HRDATAMTB[22], 1'b0);  // ../RTL/cmsdk_mcu_system.v(466)
  buf u434 (HRDATAMTB[23], 1'b0);  // ../RTL/cmsdk_mcu_system.v(466)
  buf u435 (HRDATAMTB[24], 1'b0);  // ../RTL/cmsdk_mcu_system.v(466)
  buf u436 (HRDATAMTB[25], 1'b0);  // ../RTL/cmsdk_mcu_system.v(466)
  buf u437 (HRDATAMTB[26], 1'b0);  // ../RTL/cmsdk_mcu_system.v(466)
  buf u438 (HRDATAMTB[27], 1'b0);  // ../RTL/cmsdk_mcu_system.v(466)
  buf u439 (HRDATAMTB[28], 1'b0);  // ../RTL/cmsdk_mcu_system.v(466)
  buf u44 (HREADY, sys_hready);  // ../RTL/cmsdk_mcu_system.v(998)
  buf u440 (HRDATAMTB[29], 1'b0);  // ../RTL/cmsdk_mcu_system.v(466)
  buf u441 (HRDATAMTB[30], 1'b0);  // ../RTL/cmsdk_mcu_system.v(466)
  buf u442 (HRDATAMTB[31], 1'b0);  // ../RTL/cmsdk_mcu_system.v(466)
  or u45 (intisr_cm0[30], apbsubsys_interrupt[30], gpio0_intr[14]);  // ../RTL/cmsdk_mcu_system.v(1089)
  or u46 (intisr_cm0[29], apbsubsys_interrupt[29], gpio0_intr[13]);  // ../RTL/cmsdk_mcu_system.v(1089)
  or u47 (intisr_cm0[28], apbsubsys_interrupt[28], gpio0_intr[12]);  // ../RTL/cmsdk_mcu_system.v(1089)
  or u48 (intisr_cm0[27], apbsubsys_interrupt[27], gpio0_intr[11]);  // ../RTL/cmsdk_mcu_system.v(1089)
  or u49 (intisr_cm0[26], apbsubsys_interrupt[26], gpio0_intr[10]);  // ../RTL/cmsdk_mcu_system.v(1089)
  buf u5 (HCLKSYS, HCLK);  // ../RTL/cmsdk_mcu_system.v(355)
  or u50 (intisr_cm0[25], apbsubsys_interrupt[25], gpio0_intr[9]);  // ../RTL/cmsdk_mcu_system.v(1089)
  or u51 (intisr_cm0[24], apbsubsys_interrupt[24], gpio0_intr[8]);  // ../RTL/cmsdk_mcu_system.v(1089)
  or u52 (intisr_cm0[23], apbsubsys_interrupt[23], gpio0_intr[7]);  // ../RTL/cmsdk_mcu_system.v(1089)
  or u53 (intisr_cm0[22], apbsubsys_interrupt[22], gpio0_intr[6]);  // ../RTL/cmsdk_mcu_system.v(1089)
  buf u54 (DMA_DONE, 1'b0);  // ../RTL/cmsdk_mcu_system.v(1063)
  buf u55 (dma_err, 1'b0);  // ../RTL/cmsdk_mcu_system.v(1064)
  buf u56 (dmac_pready, 1'b1);  // ../RTL/cmsdk_mcu_system.v(1065)
  buf u57 (dmac_pslverr, 1'b0);  // ../RTL/cmsdk_mcu_system.v(1066)
  buf u58 (HWDATA[0], sys_hwdata[0]);  // ../RTL/cmsdk_mcu_system.v(997)
  or u59 (intisr_cm0[21], apbsubsys_interrupt[21], gpio0_intr[5]);  // ../RTL/cmsdk_mcu_system.v(1089)
  buf u6 (RXEV, DMA_DONE);  // ../RTL/cmsdk_mcu_system.v(358)
  buf u60 (intnmi_cm0, watchdog_interrupt);  // ../RTL/cmsdk_mcu_system.v(1076)
  buf u61 (intisr_cm0[18], gpio0_intr[2]);  // ../RTL/cmsdk_mcu_system.v(1088)
  or u62 (n0, apbsubsys_interrupt[6], gpio0_combintr);  // ../RTL/cmsdk_mcu_system.v(1078)
  buf u63 (dmac_prdata[4], 1'b0);  // ../RTL/cmsdk_mcu_system.v(1067)
  or u64 (n1, apbsubsys_interrupt[7], gpio1_combintr);  // ../RTL/cmsdk_mcu_system.v(1079)
  buf u65 (dmac_prdata[3], 1'b0);  // ../RTL/cmsdk_mcu_system.v(1067)
  buf u66 (intisr_cm0[14], i2s_interrupt);  // ../RTL/cmsdk_mcu_system.v(1088)
  buf u67 (intisr_cm0[13], eth_interrupt);  // ../RTL/cmsdk_mcu_system.v(1088)
  buf u68 (dmac_prdata[0], 1'b0);  // ../RTL/cmsdk_mcu_system.v(1067)
  buf u69 (dmac_prdata[2], 1'b0);  // ../RTL/cmsdk_mcu_system.v(1067)
  buf u7 (HREADYOUTMTB, 1'b0);  // ../RTL/cmsdk_mcu_system.v(467)
  buf u70 (intisr_cm0[11], spi_interrupt);  // ../RTL/cmsdk_mcu_system.v(1088)
  buf u71 (intisr_cm0[10], apbsubsys_interrupt[10]);  // ../RTL/cmsdk_mcu_system.v(1088)
  or u72 (n3, DMA_DONE, dma_err);  // ../RTL/cmsdk_mcu_system.v(1085)
  buf u73 (dmac_prdata[1], 1'b0);  // ../RTL/cmsdk_mcu_system.v(1067)
  or u74 (n2, n5, n4);  // ../RTL/cmsdk_mcu_system.v(1082)
  or u75 (n4, apbsubsys_interrupt[14], apbsubsys_interrupt[15]);  // ../RTL/cmsdk_mcu_system.v(1082)
  buf u76 (intisr_cm0[9], apbsubsys_interrupt[9]);  // ../RTL/cmsdk_mcu_system.v(1088)
  or u77 (n5, apbsubsys_interrupt[12], apbsubsys_interrupt[13]);  // ../RTL/cmsdk_mcu_system.v(1082)
  or u78 (intisr_cm0[20], apbsubsys_interrupt[20], gpio0_intr[4]);  // ../RTL/cmsdk_mcu_system.v(1089)
  or u79 (intisr_cm0[19], apbsubsys_interrupt[19], gpio0_intr[3]);  // ../RTL/cmsdk_mcu_system.v(1089)
  buf u8 (HRESPMTB, 1'b0);  // ../RTL/cmsdk_mcu_system.v(468)
  or u80 (intisr_cm0[17], apbsubsys_interrupt[17], gpio0_intr[1]);  // ../RTL/cmsdk_mcu_system.v(1089)
  or u81 (intisr_cm0[16], apbsubsys_interrupt[16], gpio0_intr[0]);  // ../RTL/cmsdk_mcu_system.v(1089)
  or u82 (intisr_cm0[15], n3, ts_interrupt);  // ../RTL/cmsdk_mcu_system.v(1089)
  or u83 (intisr_cm0[12], n2, apbsubsys_interrupt[18]);  // ../RTL/cmsdk_mcu_system.v(1089)
  or u84 (intisr_cm0[7], n1, gpio3_interrupt);  // ../RTL/cmsdk_mcu_system.v(1089)
  or u85 (intisr_cm0[6], n0, gpio2_interrupt);  // ../RTL/cmsdk_mcu_system.v(1089)
  buf u86 (intisr_cm0[0], apbsubsys_interrupt[0]);  // ../RTL/cmsdk_mcu_system.v(1088)
  buf u87 (dmac_prdata[5], 1'b0);  // ../RTL/cmsdk_mcu_system.v(1067)
  buf u88 (dmac_prdata[6], 1'b0);  // ../RTL/cmsdk_mcu_system.v(1067)
  buf u89 (dmac_prdata[7], 1'b0);  // ../RTL/cmsdk_mcu_system.v(1067)
  buf u9 (HRDATAMTB[0], 1'b0);  // ../RTL/cmsdk_mcu_system.v(466)
  buf u90 (dmac_prdata[8], 1'b0);  // ../RTL/cmsdk_mcu_system.v(1067)
  buf u91 (dmac_prdata[9], 1'b0);  // ../RTL/cmsdk_mcu_system.v(1067)
  buf u92 (dmac_prdata[10], 1'b0);  // ../RTL/cmsdk_mcu_system.v(1067)
  buf u93 (dmac_prdata[11], 1'b0);  // ../RTL/cmsdk_mcu_system.v(1067)
  buf u94 (dmac_prdata[12], 1'b0);  // ../RTL/cmsdk_mcu_system.v(1067)
  buf u95 (dmac_prdata[13], 1'b0);  // ../RTL/cmsdk_mcu_system.v(1067)
  buf u96 (dmac_prdata[14], 1'b0);  // ../RTL/cmsdk_mcu_system.v(1067)
  buf u97 (dmac_prdata[15], 1'b0);  // ../RTL/cmsdk_mcu_system.v(1067)
  buf u98 (dmac_prdata[16], 1'b0);  // ../RTL/cmsdk_mcu_system.v(1067)
  buf u99 (dmac_prdata[17], 1'b0);  // ../RTL/cmsdk_mcu_system.v(1067)
  cmsdk_mcu_addr_decode u_addr_decode (
    .haddr(sys_haddr),
    .remap_ctrl(remap_ctrl),
    .zbt_boot_ctrl(zbt_boot_ctrl),
    .apbsys_hsel(apbsys_hsel),
    .boot_hsel(boot_hsel),
    .defslv_hsel(defslv_hsel),
    .flash_hsel(flash_hsel),
    .gpio0_hsel(gpio0_hsel),
    .gpio1_hsel(gpio1_hsel),
    .hselmtb(HSELMTB),
    .sram_hsel(sram_hsel),
    .sysctrl_hsel(sysctrl_hsel),
    .sysrom_hsel(sysrom_hsel));  // ../RTL/cmsdk_mcu_system.v(639)
  cmsdk_ahb_default_slave u_ahb_default_slave_1 (
    .HCLK(HCLKSYS),
    .HREADY(sys_hready),
    .HRESETn(HRESETn),
    .HSEL(defslv_hsel),
    .HTRANS(sys_htrans),
    .HREADYOUT(defslv_hreadyout),
    .HRESP(defslv_hresp));  // ../RTL/cmsdk_mcu_system.v(724)
  cmsdk_ahb_gpio u_ahb_gpio_0 (
    .ECOREVNUM(4'b0000),
    .FCLK(FCLK),
    .HADDR(sys_haddr[11:0]),
    .HCLK(HCLKSYS),
    .HREADY(sys_hready),
    .HRESETn(HRESETn),
    .HSEL(gpio0_hsel),
    .HSIZE(sys_hsize),
    .HTRANS(sys_htrans),
    .HWDATA(sys_hwdata),
    .HWRITE(sys_hwrite),
    .PORTIN(p0_in),
    .COMBINT(gpio0_combintr),
    .GPIOINT(gpio0_intr),
    .HRDATA(gpio0_hrdata),
    .HREADYOUT(gpio0_hreadyout),
    .HRESP(gpio0_hresp),
    .PORTEN(p0_outen),
    .PORTFUNC(p0_altfunc),
    .PORTOUT(p0_out));  // ../RTL/cmsdk_mcu_system.v(815)
  cmsdk_ahb_gpio u_ahb_gpio_1 (
    .ECOREVNUM(4'b0000),
    .FCLK(FCLK),
    .HADDR(sys_haddr[11:0]),
    .HCLK(HCLKSYS),
    .HREADY(sys_hready),
    .HRESETn(HRESETn),
    .HSEL(gpio1_hsel),
    .HSIZE(sys_hsize),
    .HTRANS(sys_htrans),
    .HWDATA(sys_hwdata),
    .HWRITE(sys_hwrite),
    .PORTIN(p1_in),
    .COMBINT(gpio1_combintr),
    .HRDATA(gpio1_hrdata),
    .HREADYOUT(gpio1_hreadyout),
    .HRESP(gpio1_hresp),
    .PORTEN(p1_outen),
    .PORTFUNC(p1_altfunc),
    .PORTOUT(p1_out));  // ../RTL/cmsdk_mcu_system.v(848)
  \cmsdk_ahb_slave_mux(PORT2_ENABLE=0,PORT9_ENABLE=0)  u_ahb_slave_mux_sys_bus (
    .HCLK(HCLKSYS),
    .HRDATA0(flash_hrdata),
    .HRDATA1(sram_hrdata),
    .HRDATA2(boot_hrdata),
    .HRDATA3(defslv_hrdata),
    .HRDATA4(apbsys_hrdata),
    .HRDATA5(gpio0_hrdata),
    .HRDATA6(gpio1_hrdata),
    .HRDATA7(sysctrl_hrdata),
    .HRDATA8(sysrom_hrdata),
    .HRDATA9(HRDATAMTB),
    .HREADY(sys_hready),
    .HREADYOUT0(flash_hreadyout),
    .HREADYOUT1(sram_hreadyout),
    .HREADYOUT2(boot_hreadyout),
    .HREADYOUT3(defslv_hreadyout),
    .HREADYOUT4(apbsys_hreadyout),
    .HREADYOUT5(gpio0_hreadyout),
    .HREADYOUT6(gpio1_hreadyout),
    .HREADYOUT7(sysctrl_hreadyout),
    .HREADYOUT8(sysrom_hreadyout),
    .HREADYOUT9(HREADYOUTMTB),
    .HRESETn(HRESETn),
    .HRESP0(flash_hresp),
    .HRESP1(sram_hresp),
    .HRESP2(boot_hresp),
    .HRESP3(defslv_hresp),
    .HRESP4(apbsys_hresp),
    .HRESP5(gpio0_hresp),
    .HRESP6(gpio1_hresp),
    .HRESP7(sysctrl_hresp),
    .HRESP8(sysrom_hresp),
    .HRESP9(HRESPMTB),
    .HSEL0(flash_hsel),
    .HSEL1(sram_hsel),
    .HSEL2(boot_hsel),
    .HSEL3(defslv_hsel),
    .HSEL4(apbsys_hsel),
    .HSEL5(gpio0_hsel),
    .HSEL6(gpio1_hsel),
    .HSEL7(sysctrl_hsel),
    .HSEL8(sysrom_hsel),
    .HSEL9(HSELMTB),
    .HRDATA(sys_hrdata),
    .HREADYOUT(sys_hreadyout),
    .HRESP(sys_hresp));  // ../RTL/cmsdk_mcu_system.v(673)
  \cmsdk_apb_subsystem_m0ds(INCLUDE_APB_TEST_SLAVE=0,INCLUDE_APB_TIMER1=0,INCLUDE_APB_DUALTIMER0=0,INCLUDE_APB_UART1=0,INCLUDE_APB_UART2=0,INCLUDE_APB_UART3=0,INCLUDE_APB_UART4=0,INCLUDE_APB_WATCHDOG=0)  u_apb_subsystem (
    .HADDR(sys_haddr[15:0]),
    .HCLK(HCLKSYS),
    .HPROT(sys_hprot),
    .HREADY(sys_hready),
    .HRESETn(HRESETn),
    .HSEL(apbsys_hsel),
    .HSIZE(sys_hsize),
    .HTRANS(sys_htrans),
    .HWDATA(sys_hwdata),
    .HWRITE(sys_hwrite),
    .PCLK(PCLK),
    .PCLKEN(PCLKEN),
    .PCLKG(PCLKG),
    .PRESETn(PRESETn),
    .ext12_prdata(32'b00000000000000000000000000000000),
    .ext12_pready(1'b1),
    .ext12_pslverr(1'b0),
    .ext13_prdata(32'b00000000000000000000000000000000),
    .ext13_pready(1'b1),
    .ext13_pslverr(1'b0),
    .ext14_prdata(32'b00000000000000000000000000000000),
    .ext14_pready(1'b1),
    .ext14_pslverr(1'b0),
    .ext15_prdata(dmac_prdata),
    .ext15_pready(dmac_pready),
    .ext15_pslverr(dmac_pslverr),
    .timer0_extin(1'bx),
    .timer1_extin(timer1_extin),
    .uart0_rxd(uart0_rxd),
    .APBACTIVE(APBACTIVE),
    .HRDATA(apbsys_hrdata),
    .HREADYOUT(apbsys_hreadyout),
    .HRESP(apbsys_hresp),
    .apbsubsys_interrupt({apbsubsys_interrupt[31:12],open_n64,apbsubsys_interrupt[10:0]}),
    .uart0_txd(uart0_txd),
    .uart0_txen(uart0_txen),
    .watchdog_interrupt(watchdog_interrupt),
    .watchdog_reset(WDOGRESETREQ),
    .b_pad_gpio_porta(b_pad_gpio_porta));  // ../RTL/cmsdk_mcu_system.v(901)
  cmsdk_mcu_stclkctrl u_cmsdk_mcu_stclkctrl (
    .FCLK(FCLK),
    .SYSRESETn(HRESETn),
    .STCLKEN(STCLKEN));  // ../RTL/cmsdk_mcu_system.v(1097)
  cmsdk_mcu_sysctrl u_cmsdk_mcu_sysctrl (
    .ECOREVNUM(4'b0000),
    .FCLK(FCLK),
    .HADDR(sys_haddr[11:0]),
    .HCLK(HCLKSYS),
    .HREADY(sys_hready),
    .HRESETn(HRESETn),
    .HSEL(sysctrl_hsel),
    .HSIZE(sys_hsize),
    .HTRANS(sys_htrans),
    .HWDATA(sys_hwdata),
    .HWRITE(sys_hwrite),
    .LOCKUP(LOCKUP),
    .PORESETn(PORESETn),
    .SYSRESETREQ(SYSRESETREQ),
    .WDOGRESETREQ(WDOGRESETREQ),
    .HRDATA(sysctrl_hrdata),
    .HREADYOUT(sysctrl_hreadyout),
    .HRESP(sysctrl_hresp),
    .LOCKUPRESET(LOCKUPRESET),
    .PMUENABLE(PMUENABLE),
    .REMAP(remap_ctrl));  // ../RTL/cmsdk_mcu_system.v(776)
  CORTEXM0INTEGRATION u_cortex_m0_integration (
    .CDBGPWRUPACK(cpu0cdbgpwrupack),
    .DBGRESETn(DBGRESETn),
    .DBGRESTART(DBGRESTART),
    .DCLK(DCLK),
    .ECOREVNUM(28'b0000000000000000000000000000),
    .EDBGRQ(EDBGRQ),
    .FCLK(FCLK),
    .HCLK(HCLK),
    .HRDATA(cm0_hrdata),
    .HREADY(cm0_hready),
    .HRESETn(HRESETn),
    .HRESP(cm0_hresp),
    .IRQ(intisr_cm0),
    .IRQLATENCY(8'b00000000),
    .NMI(intnmi_cm0),
    .PORESETn(PORESETn),
    .RSTBYPASS(RSTBYPASS),
    .RXEV(RXEV),
    .SCLK(SCLK),
    .SE(DFTSE),
    .SLEEPHOLDREQn(SLEEPHOLDREQn),
    .STCALIB(26'b10000000111101000010001111),
    .STCLKEN(STCLKEN),
    .SWCLKTCK(SWCLKTCK),
    .SWDITMS(SWDITMS),
    .TDI(TDI),
    .WICENREQ(WICENREQ),
    .nTRST(nTRST),
    .CDBGPWRUPREQ(cpu0cdbgpwrupreq),
    .DBGRESTARTED(DBGRESTARTED),
    .GATEHCLK(GATEHCLK),
    .HADDR(cm0_haddr),
    .HBURST(cm0_hburst),
    .HMASTLOCK(cm0_hmastlock),
    .HPROT(cm0_hprot),
    .HSIZE(cm0_hsize),
    .HTRANS(cm0_htrans),
    .HWDATA(cm0_hwdata),
    .HWRITE(cm0_hwrite),
    .LOCKUP(LOCKUP),
    .SLEEPDEEP(SLEEPDEEP),
    .SLEEPHOLDACKn(SLEEPHOLDACKn),
    .SLEEPING(SLEEPING),
    .SWDO(SWDO),
    .SWDOEN(SWDOEN),
    .SYSRESETREQ(SYSRESETREQ),
    .TDO(TDO),
    .WAKEUP(WAKEUP),
    .WICENACK(WICENACK),
    .nTDOEN(nTDOEN));  // ../RTL/cmsdk_mcu_system.v(384)
  \cmsdk_ahb_cs_rom_table(BASE=32'b11110000000000000000000000000000,ENTRY0BASEADDR=32'b11100000000011111111000000000000,ENTRY0PRESENT=1'b1,ENTRY1BASEADDR=32'b11110000001000000000000000000000,ENTRY1PRESENT=0)  u_system_rom_table (
    .ECOREVNUM(4'b0000),
    .HADDR(sys_haddr),
    .HBURST(sys_hburst),
    .HCLK(HCLKSYS),
    .HMASTLOCK(sys_hmastlock),
    .HPROT(sys_hprot),
    .HREADY(sys_hready),
    .HSEL(sysrom_hsel),
    .HSIZE(sys_hsize),
    .HTRANS(sys_htrans),
    .HWDATA(sys_hwdata),
    .HWRITE(sys_hwrite),
    .HRDATA(sysrom_hrdata),
    .HREADYOUT(sysrom_hreadyout),
    .HRESP(sysrom_hresp));  // ../RTL/cmsdk_mcu_system.v(752)

endmodule 

module cmsdk_mcu_pin_mux  // ../RTL/cmsdk_mcu_pin_mux.v(30)
  (
  SWCLKTCK,
  TDI,
  i_swdo,
  i_swdoen,
  i_tdo,
  i_tdoen_n,
  nTRST,
  p0_altfunc,
  p0_out,
  p0_outen,
  p1_altfunc,
  p1_out,
  p1_outen,
  uart0_txd,
  uart0_txen,
  uart1_txd,
  uart1_txen,
  uart2_txd,
  uart2_txen,
  P0,
  TDO,
  i_swclktck,
  i_swditms,
  i_tdi,
  i_trst_n,
  p0_in,
  p1_in,
  timer0_extin,
  timer1_extin,
  uart0_rxd,
  uart1_rxd,
  uart2_rxd,
  P1,
  SWDIOTMS
  );

  input SWCLKTCK;  // ../RTL/cmsdk_mcu_pin_mux.v(78)
  input TDI;  // ../RTL/cmsdk_mcu_pin_mux.v(76)
  input i_swdo;  // ../RTL/cmsdk_mcu_pin_mux.v(68)
  input i_swdoen;  // ../RTL/cmsdk_mcu_pin_mux.v(69)
  input i_tdo;  // ../RTL/cmsdk_mcu_pin_mux.v(66)
  input i_tdoen_n;  // ../RTL/cmsdk_mcu_pin_mux.v(67)
  input nTRST;  // ../RTL/cmsdk_mcu_pin_mux.v(75)
  input [15:0] p0_altfunc;  // ../RTL/cmsdk_mcu_pin_mux.v(54)
  input [15:0] p0_out;  // ../RTL/cmsdk_mcu_pin_mux.v(52)
  input [15:0] p0_outen;  // ../RTL/cmsdk_mcu_pin_mux.v(53)
  input [15:0] p1_altfunc;  // ../RTL/cmsdk_mcu_pin_mux.v(59)
  input [15:0] p1_out;  // ../RTL/cmsdk_mcu_pin_mux.v(57)
  input [15:0] p1_outen;  // ../RTL/cmsdk_mcu_pin_mux.v(58)
  input uart0_txd;  // ../RTL/cmsdk_mcu_pin_mux.v(37)
  input uart0_txen;  // ../RTL/cmsdk_mcu_pin_mux.v(38)
  input uart1_txd;  // ../RTL/cmsdk_mcu_pin_mux.v(40)
  input uart1_txen;  // ../RTL/cmsdk_mcu_pin_mux.v(41)
  input uart2_txd;  // ../RTL/cmsdk_mcu_pin_mux.v(43)
  input uart2_txen;  // ../RTL/cmsdk_mcu_pin_mux.v(44)
  output [15:0] P0;  // ../RTL/cmsdk_mcu_pin_mux.v(72)
  output TDO;  // ../RTL/cmsdk_mcu_pin_mux.v(79)
  output i_swclktck;  // ../RTL/cmsdk_mcu_pin_mux.v(64)
  output i_swditms;  // ../RTL/cmsdk_mcu_pin_mux.v(63)
  output i_tdi;  // ../RTL/cmsdk_mcu_pin_mux.v(65)
  output i_trst_n;  // ../RTL/cmsdk_mcu_pin_mux.v(62)
  output [15:0] p0_in;  // ../RTL/cmsdk_mcu_pin_mux.v(51)
  output [15:0] p1_in;  // ../RTL/cmsdk_mcu_pin_mux.v(56)
  output timer0_extin;  // ../RTL/cmsdk_mcu_pin_mux.v(47)
  output timer1_extin;  // ../RTL/cmsdk_mcu_pin_mux.v(48)
  output uart0_rxd;  // ../RTL/cmsdk_mcu_pin_mux.v(36)
  output uart1_rxd;  // ../RTL/cmsdk_mcu_pin_mux.v(39)
  output uart2_rxd;  // ../RTL/cmsdk_mcu_pin_mux.v(42)
  inout [15:0] P1;  // ../RTL/cmsdk_mcu_pin_mux.v(73)
  inout SWDIOTMS;  // ../RTL/cmsdk_mcu_pin_mux.v(77)

  wire [15:0] p0_out_en_mux;  // ../RTL/cmsdk_mcu_pin_mux.v(87)
  wire [15:0] p0_out_mux;  // ../RTL/cmsdk_mcu_pin_mux.v(84)
  wire [15:0] p1_out_en_mux;  // ../RTL/cmsdk_mcu_pin_mux.v(88)
  wire [15:0] p1_out_mux;  // ../RTL/cmsdk_mcu_pin_mux.v(85)
  wire n0;

  buf u0 (uart0_rxd, p1_in[0]);  // ../RTL/cmsdk_mcu_pin_mux.v(94)
  buf u1 (uart1_rxd, p1_in[2]);  // ../RTL/cmsdk_mcu_pin_mux.v(95)
  buf u10 (p1_out_en_mux[0], p1_outen[0]);  // ../RTL/cmsdk_mcu_pin_mux.v(123)
  buf u100 (p1_out_mux[14], p1_out[14]);  // ../RTL/cmsdk_mcu_pin_mux.v(112)
  buf u101 (p1_out_mux[13], p1_out[13]);  // ../RTL/cmsdk_mcu_pin_mux.v(112)
  buf u102 (p1_out_mux[12], p1_out[12]);  // ../RTL/cmsdk_mcu_pin_mux.v(112)
  bufif1 u103 (P1[12], p1_out_mux[12], p1_out_en_mux[12]);  // ../RTL/cmsdk_mcu_pin_mux.v(155)
  buf u104 (p1_out_mux[11], p1_out[11]);  // ../RTL/cmsdk_mcu_pin_mux.v(112)
  buf u105 (p1_out_mux[10], p1_out[10]);  // ../RTL/cmsdk_mcu_pin_mux.v(112)
  buf u106 (p1_out_mux[9], p1_out[9]);  // ../RTL/cmsdk_mcu_pin_mux.v(112)
  bufif1 u107 (P1[13], p1_out_mux[13], p1_out_en_mux[13]);  // ../RTL/cmsdk_mcu_pin_mux.v(156)
  buf u108 (p1_out_mux[8], p1_out[8]);  // ../RTL/cmsdk_mcu_pin_mux.v(112)
  buf u109 (p1_out_mux[7], p1_out[7]);  // ../RTL/cmsdk_mcu_pin_mux.v(112)
  AL_MUX u11 (
    .i0(p1_outen[1]),
    .i1(uart0_txen),
    .sel(p1_altfunc[1]),
    .o(p1_out_en_mux[1]));  // ../RTL/cmsdk_mcu_pin_mux.v(118)
  buf u110 (p1_out_mux[6], p1_out[6]);  // ../RTL/cmsdk_mcu_pin_mux.v(112)
  bufif1 u111 (P1[14], p1_out_mux[14], p1_out_en_mux[14]);  // ../RTL/cmsdk_mcu_pin_mux.v(157)
  buf u112 (p1_out_mux[4], p1_out[4]);  // ../RTL/cmsdk_mcu_pin_mux.v(112)
  buf u113 (p1_out_mux[2], p1_out[2]);  // ../RTL/cmsdk_mcu_pin_mux.v(112)
  buf u114 (p1_out_mux[0], p1_out[0]);  // ../RTL/cmsdk_mcu_pin_mux.v(112)
  bufif1 u115 (P1[15], p1_out_mux[15], p1_out_en_mux[15]);  // ../RTL/cmsdk_mcu_pin_mux.v(158)
  buf u116 (i_trst_n, nTRST);  // ../RTL/cmsdk_mcu_pin_mux.v(204)
  buf u117 (i_tdi, TDI);  // ../RTL/cmsdk_mcu_pin_mux.v(205)
  buf u118 (i_swclktck, SWCLKTCK);  // ../RTL/cmsdk_mcu_pin_mux.v(206)
  buf u119 (i_swditms, SWDIOTMS);  // ../RTL/cmsdk_mcu_pin_mux.v(207)
  AL_MUX u12 (
    .i0(p1_outen[3]),
    .i1(uart1_txen),
    .sel(p1_altfunc[3]),
    .o(p1_out_en_mux[3]));  // ../RTL/cmsdk_mcu_pin_mux.v(120)
  bufif1 u120 (SWDIOTMS, i_swdo, i_swdoen);  // ../RTL/cmsdk_mcu_pin_mux.v(210)
  not u121 (n0, i_tdoen_n);  // ../RTL/cmsdk_mcu_pin_mux.v(211)
  bufif1 u122 (TDO, i_tdo, n0);  // ../RTL/cmsdk_mcu_pin_mux.v(211)
  buf u123 (p0_out_en_mux[0], p0_outen[0]);  // ../RTL/cmsdk_mcu_pin_mux.v(115)
  AL_MUX u13 (
    .i0(p1_outen[5]),
    .i1(uart2_txen),
    .sel(p1_altfunc[5]),
    .o(p1_out_en_mux[5]));  // ../RTL/cmsdk_mcu_pin_mux.v(122)
  bufif1 u14 (P0[0], p0_out_mux[0], p0_out_en_mux[0]);  // ../RTL/cmsdk_mcu_pin_mux.v(126)
  bufif1 u15 (P0[1], p0_out_mux[1], p0_out_en_mux[1]);  // ../RTL/cmsdk_mcu_pin_mux.v(127)
  bufif1 u16 (P0[2], p0_out_mux[2], p0_out_en_mux[2]);  // ../RTL/cmsdk_mcu_pin_mux.v(128)
  bufif1 u17 (P0[3], p0_out_mux[3], p0_out_en_mux[3]);  // ../RTL/cmsdk_mcu_pin_mux.v(129)
  bufif1 u18 (P0[4], p0_out_mux[4], p0_out_en_mux[4]);  // ../RTL/cmsdk_mcu_pin_mux.v(130)
  bufif1 u19 (P0[5], p0_out_mux[5], p0_out_en_mux[5]);  // ../RTL/cmsdk_mcu_pin_mux.v(131)
  buf u2 (uart2_rxd, p1_in[4]);  // ../RTL/cmsdk_mcu_pin_mux.v(96)
  bufif1 u20 (P0[6], p0_out_mux[6], p0_out_en_mux[6]);  // ../RTL/cmsdk_mcu_pin_mux.v(132)
  bufif1 u21 (P0[7], p0_out_mux[7], p0_out_en_mux[7]);  // ../RTL/cmsdk_mcu_pin_mux.v(133)
  buf u22 (p1_in[15], P1[15]);  // ../RTL/cmsdk_mcu_pin_mux.v(101)
  bufif1 u23 (P0[8], p0_out_mux[8], p0_out_en_mux[8]);  // ../RTL/cmsdk_mcu_pin_mux.v(134)
  buf u24 (p1_in[14], P1[14]);  // ../RTL/cmsdk_mcu_pin_mux.v(101)
  buf u25 (p1_in[13], P1[13]);  // ../RTL/cmsdk_mcu_pin_mux.v(101)
  buf u26 (p1_in[12], P1[12]);  // ../RTL/cmsdk_mcu_pin_mux.v(101)
  bufif1 u27 (P0[9], p0_out_mux[9], p0_out_en_mux[9]);  // ../RTL/cmsdk_mcu_pin_mux.v(135)
  buf u28 (p1_in[11], P1[11]);  // ../RTL/cmsdk_mcu_pin_mux.v(101)
  buf u29 (p1_in[10], P1[10]);  // ../RTL/cmsdk_mcu_pin_mux.v(101)
  buf u3 (timer0_extin, p1_in[8]);  // ../RTL/cmsdk_mcu_pin_mux.v(97)
  buf u30 (p1_in[9], P1[9]);  // ../RTL/cmsdk_mcu_pin_mux.v(101)
  bufif1 u31 (P0[10], p0_out_mux[10], p0_out_en_mux[10]);  // ../RTL/cmsdk_mcu_pin_mux.v(136)
  buf u32 (p1_in[8], P1[8]);  // ../RTL/cmsdk_mcu_pin_mux.v(101)
  buf u33 (p1_in[7], P1[7]);  // ../RTL/cmsdk_mcu_pin_mux.v(101)
  buf u34 (p1_in[6], P1[6]);  // ../RTL/cmsdk_mcu_pin_mux.v(101)
  bufif1 u35 (P0[11], p0_out_mux[11], p0_out_en_mux[11]);  // ../RTL/cmsdk_mcu_pin_mux.v(137)
  buf u36 (p1_in[5], P1[5]);  // ../RTL/cmsdk_mcu_pin_mux.v(101)
  buf u37 (p1_in[4], P1[4]);  // ../RTL/cmsdk_mcu_pin_mux.v(101)
  buf u38 (p1_in[3], P1[3]);  // ../RTL/cmsdk_mcu_pin_mux.v(101)
  bufif1 u39 (P0[12], p0_out_mux[12], p0_out_en_mux[12]);  // ../RTL/cmsdk_mcu_pin_mux.v(138)
  buf u4 (timer1_extin, p1_in[9]);  // ../RTL/cmsdk_mcu_pin_mux.v(98)
  buf u40 (p1_in[2], P1[2]);  // ../RTL/cmsdk_mcu_pin_mux.v(101)
  buf u41 (p1_in[1], P1[1]);  // ../RTL/cmsdk_mcu_pin_mux.v(101)
  buf u42 (p0_out_mux[15], p0_out[15]);  // ../RTL/cmsdk_mcu_pin_mux.v(104)
  bufif1 u43 (P0[13], p0_out_mux[13], p0_out_en_mux[13]);  // ../RTL/cmsdk_mcu_pin_mux.v(139)
  buf u44 (p0_out_mux[14], p0_out[14]);  // ../RTL/cmsdk_mcu_pin_mux.v(104)
  buf u45 (p0_out_mux[13], p0_out[13]);  // ../RTL/cmsdk_mcu_pin_mux.v(104)
  buf u46 (p0_out_mux[12], p0_out[12]);  // ../RTL/cmsdk_mcu_pin_mux.v(104)
  bufif1 u47 (P0[14], p0_out_mux[14], p0_out_en_mux[14]);  // ../RTL/cmsdk_mcu_pin_mux.v(140)
  buf u48 (p0_out_mux[11], p0_out[11]);  // ../RTL/cmsdk_mcu_pin_mux.v(104)
  buf u49 (p0_out_mux[10], p0_out[10]);  // ../RTL/cmsdk_mcu_pin_mux.v(104)
  buf u5 (p1_in[0], P1[0]);  // ../RTL/cmsdk_mcu_pin_mux.v(101)
  buf u50 (p0_out_mux[9], p0_out[9]);  // ../RTL/cmsdk_mcu_pin_mux.v(104)
  bufif1 u51 (P0[15], p0_out_mux[15], p0_out_en_mux[15]);  // ../RTL/cmsdk_mcu_pin_mux.v(141)
  buf u52 (p0_out_mux[8], p0_out[8]);  // ../RTL/cmsdk_mcu_pin_mux.v(104)
  buf u53 (p0_out_mux[7], p0_out[7]);  // ../RTL/cmsdk_mcu_pin_mux.v(104)
  buf u54 (p0_out_mux[6], p0_out[6]);  // ../RTL/cmsdk_mcu_pin_mux.v(104)
  bufif1 u55 (P1[0], p1_out_mux[0], p1_out_en_mux[0]);  // ../RTL/cmsdk_mcu_pin_mux.v(143)
  buf u56 (p0_out_mux[5], p0_out[5]);  // ../RTL/cmsdk_mcu_pin_mux.v(104)
  buf u57 (p0_out_mux[4], p0_out[4]);  // ../RTL/cmsdk_mcu_pin_mux.v(104)
  buf u58 (p0_out_mux[3], p0_out[3]);  // ../RTL/cmsdk_mcu_pin_mux.v(104)
  bufif1 u59 (P1[1], p1_out_mux[1], p1_out_en_mux[1]);  // ../RTL/cmsdk_mcu_pin_mux.v(144)
  AL_MUX u6 (
    .i0(p1_out[1]),
    .i1(uart0_txd),
    .sel(p1_altfunc[1]),
    .o(p1_out_mux[1]));  // ../RTL/cmsdk_mcu_pin_mux.v(107)
  buf u60 (p0_out_mux[2], p0_out[2]);  // ../RTL/cmsdk_mcu_pin_mux.v(104)
  buf u61 (p0_out_mux[1], p0_out[1]);  // ../RTL/cmsdk_mcu_pin_mux.v(104)
  buf u62 (p1_out_en_mux[15], p1_outen[15]);  // ../RTL/cmsdk_mcu_pin_mux.v(123)
  bufif1 u63 (P1[2], p1_out_mux[2], p1_out_en_mux[2]);  // ../RTL/cmsdk_mcu_pin_mux.v(145)
  buf u64 (p1_out_en_mux[14], p1_outen[14]);  // ../RTL/cmsdk_mcu_pin_mux.v(123)
  buf u65 (p1_out_en_mux[13], p1_outen[13]);  // ../RTL/cmsdk_mcu_pin_mux.v(123)
  buf u66 (p1_out_en_mux[12], p1_outen[12]);  // ../RTL/cmsdk_mcu_pin_mux.v(123)
  bufif1 u67 (P1[3], p1_out_mux[3], p1_out_en_mux[3]);  // ../RTL/cmsdk_mcu_pin_mux.v(146)
  buf u68 (p1_out_en_mux[11], p1_outen[11]);  // ../RTL/cmsdk_mcu_pin_mux.v(123)
  buf u69 (p1_out_en_mux[10], p1_outen[10]);  // ../RTL/cmsdk_mcu_pin_mux.v(123)
  AL_MUX u7 (
    .i0(p1_out[3]),
    .i1(uart1_txd),
    .sel(p1_altfunc[3]),
    .o(p1_out_mux[3]));  // ../RTL/cmsdk_mcu_pin_mux.v(109)
  buf u70 (p1_out_en_mux[9], p1_outen[9]);  // ../RTL/cmsdk_mcu_pin_mux.v(123)
  bufif1 u71 (P1[4], p1_out_mux[4], p1_out_en_mux[4]);  // ../RTL/cmsdk_mcu_pin_mux.v(147)
  buf u72 (p1_out_en_mux[8], p1_outen[8]);  // ../RTL/cmsdk_mcu_pin_mux.v(123)
  buf u73 (p1_out_en_mux[7], p1_outen[7]);  // ../RTL/cmsdk_mcu_pin_mux.v(123)
  buf u74 (p1_out_en_mux[6], p1_outen[6]);  // ../RTL/cmsdk_mcu_pin_mux.v(123)
  bufif1 u75 (P1[5], p1_out_mux[5], p1_out_en_mux[5]);  // ../RTL/cmsdk_mcu_pin_mux.v(148)
  buf u76 (p1_out_en_mux[4], p1_outen[4]);  // ../RTL/cmsdk_mcu_pin_mux.v(123)
  buf u77 (p1_out_en_mux[2], p1_outen[2]);  // ../RTL/cmsdk_mcu_pin_mux.v(123)
  buf u78 (p0_out_en_mux[15], p0_outen[15]);  // ../RTL/cmsdk_mcu_pin_mux.v(115)
  bufif1 u79 (P1[6], p1_out_mux[6], p1_out_en_mux[6]);  // ../RTL/cmsdk_mcu_pin_mux.v(149)
  AL_MUX u8 (
    .i0(p1_out[5]),
    .i1(uart2_txd),
    .sel(p1_altfunc[5]),
    .o(p1_out_mux[5]));  // ../RTL/cmsdk_mcu_pin_mux.v(111)
  buf u80 (p0_out_en_mux[14], p0_outen[14]);  // ../RTL/cmsdk_mcu_pin_mux.v(115)
  buf u81 (p0_out_en_mux[13], p0_outen[13]);  // ../RTL/cmsdk_mcu_pin_mux.v(115)
  buf u82 (p0_out_en_mux[12], p0_outen[12]);  // ../RTL/cmsdk_mcu_pin_mux.v(115)
  bufif1 u83 (P1[7], p1_out_mux[7], p1_out_en_mux[7]);  // ../RTL/cmsdk_mcu_pin_mux.v(150)
  buf u84 (p0_out_en_mux[11], p0_outen[11]);  // ../RTL/cmsdk_mcu_pin_mux.v(115)
  buf u85 (p0_out_en_mux[10], p0_outen[10]);  // ../RTL/cmsdk_mcu_pin_mux.v(115)
  buf u86 (p0_out_en_mux[9], p0_outen[9]);  // ../RTL/cmsdk_mcu_pin_mux.v(115)
  bufif1 u87 (P1[8], p1_out_mux[8], p1_out_en_mux[8]);  // ../RTL/cmsdk_mcu_pin_mux.v(151)
  buf u88 (p0_out_en_mux[8], p0_outen[8]);  // ../RTL/cmsdk_mcu_pin_mux.v(115)
  buf u89 (p0_out_en_mux[7], p0_outen[7]);  // ../RTL/cmsdk_mcu_pin_mux.v(115)
  buf u9 (p0_out_mux[0], p0_out[0]);  // ../RTL/cmsdk_mcu_pin_mux.v(104)
  buf u90 (p0_out_en_mux[6], p0_outen[6]);  // ../RTL/cmsdk_mcu_pin_mux.v(115)
  bufif1 u91 (P1[9], p1_out_mux[9], p1_out_en_mux[9]);  // ../RTL/cmsdk_mcu_pin_mux.v(152)
  buf u92 (p0_out_en_mux[5], p0_outen[5]);  // ../RTL/cmsdk_mcu_pin_mux.v(115)
  buf u93 (p0_out_en_mux[4], p0_outen[4]);  // ../RTL/cmsdk_mcu_pin_mux.v(115)
  buf u94 (p0_out_en_mux[3], p0_outen[3]);  // ../RTL/cmsdk_mcu_pin_mux.v(115)
  bufif1 u95 (P1[10], p1_out_mux[10], p1_out_en_mux[10]);  // ../RTL/cmsdk_mcu_pin_mux.v(153)
  buf u96 (p0_out_en_mux[2], p0_outen[2]);  // ../RTL/cmsdk_mcu_pin_mux.v(115)
  buf u97 (p0_out_en_mux[1], p0_outen[1]);  // ../RTL/cmsdk_mcu_pin_mux.v(115)
  buf u98 (p1_out_mux[15], p1_out[15]);  // ../RTL/cmsdk_mcu_pin_mux.v(112)
  bufif1 u99 (P1[11], p1_out_mux[11], p1_out_en_mux[11]);  // ../RTL/cmsdk_mcu_pin_mux.v(154)

endmodule 

module binary_mux_s2_w32
  (
  i0,
  i1,
  i2,
  i3,
  sel,
  o
  );

  input [31:0] i0;
  input [31:0] i1;
  input [31:0] i2;
  input [31:0] i3;
  input [1:0] sel;
  output [31:0] o;



endmodule 

module binary_mux_s1_w32
  (
  i0,
  i1,
  sel,
  o
  );

  input [31:0] i0;
  input [31:0] i1;
  input sel;
  output [31:0] o;



endmodule 

module ram_w10x32_r10x32
  (
  clk1,
  ra1,
  re1,
  wa1,
  wd1,
  we1,
  rd1
  );

  input clk1;
  input [9:0] ra1;
  input re1;
  input [9:0] wa1;
  input [31:0] wd1;
  input we1;
  output [31:0] rd1;



endmodule 

module reg_ar_as_w32
  (
  clk,
  d,
  en,
  reset,
  set,
  q
  );

  input clk;
  input [31:0] d;
  input en;
  input [31:0] reset;
  input [31:0] set;
  output [31:0] q;



endmodule 

module reg_ar_as_w3
  (
  clk,
  d,
  en,
  reset,
  set,
  q
  );

  input clk;
  input [2:0] d;
  input en;
  input [2:0] reset;
  input [2:0] set;
  output [2:0] q;



endmodule 

module cmsdk_mcu_addr_decode  // ../RTL/cmsdk_mcu_addr_decode.v(32)
  (
  haddr,
  remap_ctrl,
  zbt_boot_ctrl,
  apbsys_hsel,
  boot_hsel,
  defslv_hsel,
  flash_hsel,
  gpio0_hsel,
  gpio1_hsel,
  hselmtb,
  hselram,
  hselsfr,
  sram_hsel,
  sysctrl_hsel,
  sysrom_hsel
  );

  input [31:0] haddr;  // ../RTL/cmsdk_mcu_addr_decode.v(47)
  input remap_ctrl;  // ../RTL/cmsdk_mcu_addr_decode.v(49)
  input zbt_boot_ctrl;  // ../RTL/cmsdk_mcu_addr_decode.v(50)
  output apbsys_hsel;  // ../RTL/cmsdk_mcu_addr_decode.v(58)
  output boot_hsel;  // ../RTL/cmsdk_mcu_addr_decode.v(53)
  output defslv_hsel;  // ../RTL/cmsdk_mcu_addr_decode.v(65)
  output flash_hsel;  // ../RTL/cmsdk_mcu_addr_decode.v(54)
  output gpio0_hsel;  // ../RTL/cmsdk_mcu_addr_decode.v(59)
  output gpio1_hsel;  // ../RTL/cmsdk_mcu_addr_decode.v(60)
  output hselmtb;  // ../RTL/cmsdk_mcu_addr_decode.v(68)
  output hselram;  // ../RTL/cmsdk_mcu_addr_decode.v(69)
  output hselsfr;  // ../RTL/cmsdk_mcu_addr_decode.v(70)
  output sram_hsel;  // ../RTL/cmsdk_mcu_addr_decode.v(55)
  output sysctrl_hsel;  // ../RTL/cmsdk_mcu_addr_decode.v(61)
  output sysrom_hsel;  // ../RTL/cmsdk_mcu_addr_decode.v(62)

  parameter BASEADDR_GPIO0 = 32'b01000000000000010000000000000000;
  parameter BASEADDR_GPIO1 = 32'b01000000000000010001000000000000;
  parameter BASEADDR_SYSROMTABLE = 32'b11110000000000000000000000000000;
  parameter BOOT_LOADER_PRESENT = 0;
  wire n0;
  wire n1;
  wire n2;
  wire n3;
  wire n4;
  wire n5;
  wire n6;

  eq_w9 eq0 (
    .i0(haddr[31:23]),
    .i1(9'b000000000),
    .o(flash_hsel));  // ../RTL/cmsdk_mcu_addr_decode.v(96)
  eq_w16 eq1 (
    .i0(haddr[31:16]),
    .i1(16'b0100000000000000),
    .o(apbsys_hsel));  // ../RTL/cmsdk_mcu_addr_decode.v(105)
  eq_w20 eq2 (
    .i0(haddr[31:12]),
    .i1(20'b01000000000000010000),
    .o(gpio0_hsel));  // ../RTL/cmsdk_mcu_addr_decode.v(107)
  eq_w20 eq3 (
    .i0(haddr[31:12]),
    .i1(20'b01000000000000010001),
    .o(gpio1_hsel));  // ../RTL/cmsdk_mcu_addr_decode.v(109)
  eq_w20 eq4 (
    .i0(haddr[31:12]),
    .i1(20'b01000000000000011111),
    .o(sysctrl_hsel));  // ../RTL/cmsdk_mcu_addr_decode.v(110)
  eq_w20 eq5 (
    .i0(haddr[31:12]),
    .i1(20'b11110000000000000000),
    .o(sysrom_hsel));  // ../RTL/cmsdk_mcu_addr_decode.v(112)
  or u10 (n6, n5, sysrom_hsel);  // ../RTL/cmsdk_mcu_addr_decode.v(128)
  not u11 (sram_hsel, n6);  // ../RTL/cmsdk_mcu_addr_decode.v(128)
  buf u12 (hselmtb, 1'b0);  // ../RTL/cmsdk_mcu_addr_decode.v(155)
  buf u13 (hselram, 1'b0);  // ../RTL/cmsdk_mcu_addr_decode.v(156)
  buf u14 (hselsfr, 1'b0);  // ../RTL/cmsdk_mcu_addr_decode.v(157)
  buf u2 (boot_hsel, 1'b0);  // ../RTL/cmsdk_mcu_addr_decode.v(92)
  buf u3 (defslv_hsel, 1'b0);  // ../RTL/cmsdk_mcu_addr_decode.v(120)
  or u4 (n0, flash_hsel, hselmtb);  // ../RTL/cmsdk_mcu_addr_decode.v(125)
  or u5 (n1, n0, boot_hsel);  // ../RTL/cmsdk_mcu_addr_decode.v(126)
  or u6 (n2, n1, apbsys_hsel);  // ../RTL/cmsdk_mcu_addr_decode.v(126)
  or u7 (n3, n2, gpio0_hsel);  // ../RTL/cmsdk_mcu_addr_decode.v(127)
  or u8 (n4, n3, gpio1_hsel);  // ../RTL/cmsdk_mcu_addr_decode.v(127)
  or u9 (n5, n4, sysctrl_hsel);  // ../RTL/cmsdk_mcu_addr_decode.v(128)

endmodule 

module cmsdk_ahb_default_slave  // ../RTL/cmsdk_ahb_default_slave.v(30)
  (
  HCLK,
  HREADY,
  HRESETn,
  HSEL,
  HTRANS,
  HREADYOUT,
  HRESP
  );

  input HCLK;  // ../RTL/cmsdk_ahb_default_slave.v(32)
  input HREADY;  // ../RTL/cmsdk_ahb_default_slave.v(36)
  input HRESETn;  // ../RTL/cmsdk_ahb_default_slave.v(33)
  input HSEL;  // ../RTL/cmsdk_ahb_default_slave.v(34)
  input [1:0] HTRANS;  // ../RTL/cmsdk_ahb_default_slave.v(35)
  output HREADYOUT;  // ../RTL/cmsdk_ahb_default_slave.v(39)
  output HRESP;  // ../RTL/cmsdk_ahb_default_slave.v(40)

  wire [1:0] next_state;  // ../RTL/cmsdk_ahb_default_slave.v(49)
  wire [1:0] resp_state;  // ../RTL/cmsdk_ahb_default_slave.v(48)
  wire n0;
  wire n1;
  wire n2;
  wire trans_req;  // ../RTL/cmsdk_ahb_default_slave.v(47)

  reg_ar_as_w2 reg0 (
    .clk(HCLK),
    .d(next_state),
    .reset({n2,1'b0}),
    .set({1'b0,n2}),
    .q(resp_state));  // ../RTL/cmsdk_ahb_default_slave.v(68)
  and u1 (n0, HSEL, HTRANS[1]);  // ../RTL/cmsdk_ahb_default_slave.v(52)
  and u2 (trans_req, n0, HREADY);  // ../RTL/cmsdk_ahb_default_slave.v(52)
  not u3 (n1, resp_state[0]);  // ../RTL/cmsdk_ahb_default_slave.v(60)
  or u4 (next_state[1], trans_req, n1);  // ../RTL/cmsdk_ahb_default_slave.v(60)
  not u5 (next_state[0], trans_req);  // ../RTL/cmsdk_ahb_default_slave.v(61)
  not u6 (n2, HRESETn);  // ../RTL/cmsdk_ahb_default_slave.v(65)
  buf u7 (HREADYOUT, resp_state[0]);  // ../RTL/cmsdk_ahb_default_slave.v(71)
  buf u8 (HRESP, resp_state[1]);  // ../RTL/cmsdk_ahb_default_slave.v(72)

endmodule 

module cmsdk_ahb_gpio  // ../RTL/cmsdk_ahb_gpio.v(24)
  (
  ECOREVNUM,
  FCLK,
  HADDR,
  HCLK,
  HREADY,
  HRESETn,
  HSEL,
  HSIZE,
  HTRANS,
  HWDATA,
  HWRITE,
  PORTIN,
  COMBINT,
  GPIOINT,
  HRDATA,
  HREADYOUT,
  HRESP,
  PORTEN,
  PORTFUNC,
  PORTOUT
  );

  input [3:0] ECOREVNUM;  // ../RTL/cmsdk_ahb_gpio.v(54)
  input FCLK;  // ../RTL/cmsdk_ahb_gpio.v(45)
  input [11:0] HADDR;  // ../RTL/cmsdk_ahb_gpio.v(51)
  input HCLK;  // ../RTL/cmsdk_ahb_gpio.v(43)
  input HREADY;  // ../RTL/cmsdk_ahb_gpio.v(47)
  input HRESETn;  // ../RTL/cmsdk_ahb_gpio.v(44)
  input HSEL;  // ../RTL/cmsdk_ahb_gpio.v(46)
  input [2:0] HSIZE;  // ../RTL/cmsdk_ahb_gpio.v(49)
  input [1:0] HTRANS;  // ../RTL/cmsdk_ahb_gpio.v(48)
  input [31:0] HWDATA;  // ../RTL/cmsdk_ahb_gpio.v(52)
  input HWRITE;  // ../RTL/cmsdk_ahb_gpio.v(50)
  input [15:0] PORTIN;  // ../RTL/cmsdk_ahb_gpio.v(56)
  output COMBINT;  // ../RTL/cmsdk_ahb_gpio.v(68)
  output [15:0] GPIOINT;  // ../RTL/cmsdk_ahb_gpio.v(67)
  output [31:0] HRDATA;  // ../RTL/cmsdk_ahb_gpio.v(61)
  output HREADYOUT;  // ../RTL/cmsdk_ahb_gpio.v(59)
  output HRESP;  // ../RTL/cmsdk_ahb_gpio.v(60)
  output [15:0] PORTEN;  // ../RTL/cmsdk_ahb_gpio.v(64)
  output [15:0] PORTFUNC;  // ../RTL/cmsdk_ahb_gpio.v(65)
  output [15:0] PORTOUT;  // ../RTL/cmsdk_ahb_gpio.v(63)

  parameter ALTERNATE_FUNC_DEFAULT = 16'b0000000000000000;
  parameter ALTERNATE_FUNC_MASK = 16'b1111111111111111;
  parameter BE = 0;
  wire [11:0] IOADDR;  // ../RTL/cmsdk_ahb_gpio.v(76)
  wire [31:0] IORDATA;  // ../RTL/cmsdk_ahb_gpio.v(74)
  wire [1:0] IOSIZE;  // ../RTL/cmsdk_ahb_gpio.v(78)
  wire [31:0] IOWDATA;  // ../RTL/cmsdk_ahb_gpio.v(80)
  wire IOSEL;  // ../RTL/cmsdk_ahb_gpio.v(75)
  wire IOTRANS;  // ../RTL/cmsdk_ahb_gpio.v(79)
  wire IOWRITE;  // ../RTL/cmsdk_ahb_gpio.v(77)

  cmsdk_ahb_to_iop u_ahb_to_gpio (
    .HADDR(HADDR),
    .HCLK(HCLK),
    .HREADY(HREADY),
    .HRESETn(HRESETn),
    .HSEL(HSEL),
    .HSIZE(HSIZE),
    .HTRANS(HTRANS),
    .HWDATA(HWDATA),
    .HWRITE(HWRITE),
    .IORDATA(IORDATA),
    .HRDATA(HRDATA),
    .HREADYOUT(HREADYOUT),
    .HRESP(HRESP),
    .IOADDR(IOADDR),
    .IOSEL(IOSEL),
    .IOSIZE(IOSIZE),
    .IOTRANS(IOTRANS),
    .IOWDATA(IOWDATA),
    .IOWRITE(IOWRITE));  // ../RTL/cmsdk_ahb_gpio.v(87)
  cmsdk_iop_gpio u_iop_gpio (
    .ECOREVNUM(ECOREVNUM),
    .FCLK(FCLK),
    .HCLK(HCLK),
    .HRESETn(HRESETn),
    .IOADDR(IOADDR),
    .IOSEL(IOSEL),
    .IOSIZE(IOSIZE),
    .IOTRANS(IOTRANS),
    .IOWDATA(IOWDATA),
    .IOWRITE(IOWRITE),
    .PORTIN(PORTIN),
    .COMBINT(COMBINT),
    .GPIOINT(GPIOINT),
    .IORDATA(IORDATA),
    .PORTEN(PORTEN),
    .PORTFUNC(PORTFUNC),
    .PORTOUT(PORTOUT));  // ../RTL/cmsdk_ahb_gpio.v(118)

endmodule 

module \cmsdk_ahb_slave_mux(PORT2_ENABLE=0,PORT9_ENABLE=0)   // ../RTL/cmsdk_ahb_slave_mux.v(28)
  (
  HCLK,
  HRDATA0,
  HRDATA1,
  HRDATA2,
  HRDATA3,
  HRDATA4,
  HRDATA5,
  HRDATA6,
  HRDATA7,
  HRDATA8,
  HRDATA9,
  HREADY,
  HREADYOUT0,
  HREADYOUT1,
  HREADYOUT2,
  HREADYOUT3,
  HREADYOUT4,
  HREADYOUT5,
  HREADYOUT6,
  HREADYOUT7,
  HREADYOUT8,
  HREADYOUT9,
  HRESETn,
  HRESP0,
  HRESP1,
  HRESP2,
  HRESP3,
  HRESP4,
  HRESP5,
  HRESP6,
  HRESP7,
  HRESP8,
  HRESP9,
  HSEL0,
  HSEL1,
  HSEL2,
  HSEL3,
  HSEL4,
  HSEL5,
  HSEL6,
  HSEL7,
  HSEL8,
  HSEL9,
  HRDATA,
  HREADYOUT,
  HRESP
  );

  input HCLK;  // ../RTL/cmsdk_ahb_slave_mux.v(46)
  input [31:0] HRDATA0;  // ../RTL/cmsdk_ahb_slave_mux.v(52)
  input [31:0] HRDATA1;  // ../RTL/cmsdk_ahb_slave_mux.v(56)
  input [31:0] HRDATA2;  // ../RTL/cmsdk_ahb_slave_mux.v(60)
  input [31:0] HRDATA3;  // ../RTL/cmsdk_ahb_slave_mux.v(64)
  input [31:0] HRDATA4;  // ../RTL/cmsdk_ahb_slave_mux.v(68)
  input [31:0] HRDATA5;  // ../RTL/cmsdk_ahb_slave_mux.v(72)
  input [31:0] HRDATA6;  // ../RTL/cmsdk_ahb_slave_mux.v(76)
  input [31:0] HRDATA7;  // ../RTL/cmsdk_ahb_slave_mux.v(80)
  input [31:0] HRDATA8;  // ../RTL/cmsdk_ahb_slave_mux.v(84)
  input [31:0] HRDATA9;  // ../RTL/cmsdk_ahb_slave_mux.v(88)
  input HREADY;  // ../RTL/cmsdk_ahb_slave_mux.v(48)
  input HREADYOUT0;  // ../RTL/cmsdk_ahb_slave_mux.v(50)
  input HREADYOUT1;  // ../RTL/cmsdk_ahb_slave_mux.v(54)
  input HREADYOUT2;  // ../RTL/cmsdk_ahb_slave_mux.v(58)
  input HREADYOUT3;  // ../RTL/cmsdk_ahb_slave_mux.v(62)
  input HREADYOUT4;  // ../RTL/cmsdk_ahb_slave_mux.v(66)
  input HREADYOUT5;  // ../RTL/cmsdk_ahb_slave_mux.v(70)
  input HREADYOUT6;  // ../RTL/cmsdk_ahb_slave_mux.v(74)
  input HREADYOUT7;  // ../RTL/cmsdk_ahb_slave_mux.v(78)
  input HREADYOUT8;  // ../RTL/cmsdk_ahb_slave_mux.v(82)
  input HREADYOUT9;  // ../RTL/cmsdk_ahb_slave_mux.v(86)
  input HRESETn;  // ../RTL/cmsdk_ahb_slave_mux.v(47)
  input HRESP0;  // ../RTL/cmsdk_ahb_slave_mux.v(51)
  input HRESP1;  // ../RTL/cmsdk_ahb_slave_mux.v(55)
  input HRESP2;  // ../RTL/cmsdk_ahb_slave_mux.v(59)
  input HRESP3;  // ../RTL/cmsdk_ahb_slave_mux.v(63)
  input HRESP4;  // ../RTL/cmsdk_ahb_slave_mux.v(67)
  input HRESP5;  // ../RTL/cmsdk_ahb_slave_mux.v(71)
  input HRESP6;  // ../RTL/cmsdk_ahb_slave_mux.v(75)
  input HRESP7;  // ../RTL/cmsdk_ahb_slave_mux.v(79)
  input HRESP8;  // ../RTL/cmsdk_ahb_slave_mux.v(83)
  input HRESP9;  // ../RTL/cmsdk_ahb_slave_mux.v(87)
  input HSEL0;  // ../RTL/cmsdk_ahb_slave_mux.v(49)
  input HSEL1;  // ../RTL/cmsdk_ahb_slave_mux.v(53)
  input HSEL2;  // ../RTL/cmsdk_ahb_slave_mux.v(57)
  input HSEL3;  // ../RTL/cmsdk_ahb_slave_mux.v(61)
  input HSEL4;  // ../RTL/cmsdk_ahb_slave_mux.v(65)
  input HSEL5;  // ../RTL/cmsdk_ahb_slave_mux.v(69)
  input HSEL6;  // ../RTL/cmsdk_ahb_slave_mux.v(73)
  input HSEL7;  // ../RTL/cmsdk_ahb_slave_mux.v(77)
  input HSEL8;  // ../RTL/cmsdk_ahb_slave_mux.v(81)
  input HSEL9;  // ../RTL/cmsdk_ahb_slave_mux.v(85)
  output [31:0] HRDATA;  // ../RTL/cmsdk_ahb_slave_mux.v(91)
  output HREADYOUT;  // ../RTL/cmsdk_ahb_slave_mux.v(89)
  output HRESP;  // ../RTL/cmsdk_ahb_slave_mux.v(90)

  parameter DW = 32;
  parameter PORT0_ENABLE = 1;
  parameter PORT1_ENABLE = 1;
  parameter PORT2_ENABLE = 0;
  parameter PORT3_ENABLE = 1;
  parameter PORT4_ENABLE = 1;
  parameter PORT5_ENABLE = 1;
  parameter PORT6_ENABLE = 1;
  parameter PORT7_ENABLE = 1;
  parameter PORT8_ENABLE = 1;
  parameter PORT9_ENABLE = 0;
  wire [9:0] n1;
  wire [31:0] n24;
  wire [31:0] n25;
  wire [31:0] n26;
  wire [31:0] n27;
  wire [31:0] n28;
  wire [31:0] n29;
  wire [31:0] n30;
  wire [31:0] n31;
  wire [31:0] n32;
  wire [31:0] n33;
  wire [31:0] n34;
  wire [31:0] n35;
  wire [31:0] n36;
  wire [31:0] n37;
  wire [9:0] nxt_hsel_reg;  // ../RTL/cmsdk_ahb_slave_mux.v(96)
  wire [9:0] reg_hsel;  // ../RTL/cmsdk_ahb_slave_mux.v(95)
  wire mux_hready;  // ../RTL/cmsdk_ahb_slave_mux.v(94)
  wire n0;
  wire n10;
  wire n11;
  wire n12;
  wire n13;
  wire n14;
  wire n15;
  wire n16;
  wire n17;
  wire n18;
  wire n19;
  wire n2;
  wire n20;
  wire n21;
  wire n22;
  wire n23;
  wire n3;
  wire n38;
  wire n39;
  wire n4;
  wire n40;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n5;
  wire n50;
  wire n51;
  wire n6;
  wire n7;
  wire n8;
  wire n9;

  binary_mux_s1_w10 mux0 (
    .i0(reg_hsel),
    .i1(nxt_hsel_reg),
    .sel(HREADY),
    .o(n1));  // ../RTL/cmsdk_ahb_slave_mux.v(115)
  reg_ar_as_w10 reg0 (
    .clk(HCLK),
    .d(n1),
    .reset({n0,n0,n0,n0,n0,n0,n0,n0,n0,n0}),
    .set(10'b0000000000),
    .q(reg_hsel));  // ../RTL/cmsdk_ahb_slave_mux.v(115)
  or u1 (HRDATA[9], n36[9], n37[9]);  // ../RTL/cmsdk_ahb_slave_mux.v(141)
  or u10 (HRDATA[13], n36[13], n37[13]);  // ../RTL/cmsdk_ahb_slave_mux.v(141)
  and u100 (n37[14], reg_hsel[8], HRDATA8[14]);  // ../RTL/cmsdk_ahb_slave_mux.v(141)
  and u101 (n37[15], reg_hsel[8], HRDATA8[15]);  // ../RTL/cmsdk_ahb_slave_mux.v(141)
  and u102 (n37[16], reg_hsel[8], HRDATA8[16]);  // ../RTL/cmsdk_ahb_slave_mux.v(141)
  and u103 (n37[17], reg_hsel[8], HRDATA8[17]);  // ../RTL/cmsdk_ahb_slave_mux.v(141)
  and u104 (n37[18], reg_hsel[8], HRDATA8[18]);  // ../RTL/cmsdk_ahb_slave_mux.v(141)
  and u105 (n37[19], reg_hsel[8], HRDATA8[19]);  // ../RTL/cmsdk_ahb_slave_mux.v(141)
  and u106 (n37[20], reg_hsel[8], HRDATA8[20]);  // ../RTL/cmsdk_ahb_slave_mux.v(141)
  and u107 (n37[21], reg_hsel[8], HRDATA8[21]);  // ../RTL/cmsdk_ahb_slave_mux.v(141)
  and u108 (n37[22], reg_hsel[8], HRDATA8[22]);  // ../RTL/cmsdk_ahb_slave_mux.v(141)
  and u109 (n37[23], reg_hsel[8], HRDATA8[23]);  // ../RTL/cmsdk_ahb_slave_mux.v(141)
  or u11 (HRDATA[12], n36[12], n37[12]);  // ../RTL/cmsdk_ahb_slave_mux.v(141)
  and u110 (n37[24], reg_hsel[8], HRDATA8[24]);  // ../RTL/cmsdk_ahb_slave_mux.v(141)
  and u111 (n37[25], reg_hsel[8], HRDATA8[25]);  // ../RTL/cmsdk_ahb_slave_mux.v(141)
  and u112 (n37[26], reg_hsel[8], HRDATA8[26]);  // ../RTL/cmsdk_ahb_slave_mux.v(141)
  and u113 (n37[27], reg_hsel[8], HRDATA8[27]);  // ../RTL/cmsdk_ahb_slave_mux.v(141)
  and u114 (n37[28], reg_hsel[8], HRDATA8[28]);  // ../RTL/cmsdk_ahb_slave_mux.v(141)
  and u115 (n37[29], reg_hsel[8], HRDATA8[29]);  // ../RTL/cmsdk_ahb_slave_mux.v(141)
  and u116 (n37[30], reg_hsel[8], HRDATA8[30]);  // ../RTL/cmsdk_ahb_slave_mux.v(141)
  and u117 (n37[31], reg_hsel[8], HRDATA8[31]);  // ../RTL/cmsdk_ahb_slave_mux.v(141)
  or u118 (n36[1], n34[1], n35[1]);  // ../RTL/cmsdk_ahb_slave_mux.v(140)
  or u119 (n36[2], n34[2], n35[2]);  // ../RTL/cmsdk_ahb_slave_mux.v(140)
  or u12 (HRDATA[11], n36[11], n37[11]);  // ../RTL/cmsdk_ahb_slave_mux.v(141)
  or u120 (n36[3], n34[3], n35[3]);  // ../RTL/cmsdk_ahb_slave_mux.v(140)
  or u121 (n36[4], n34[4], n35[4]);  // ../RTL/cmsdk_ahb_slave_mux.v(140)
  or u122 (n36[5], n34[5], n35[5]);  // ../RTL/cmsdk_ahb_slave_mux.v(140)
  or u123 (n36[6], n34[6], n35[6]);  // ../RTL/cmsdk_ahb_slave_mux.v(140)
  or u124 (n36[7], n34[7], n35[7]);  // ../RTL/cmsdk_ahb_slave_mux.v(140)
  or u125 (n36[8], n34[8], n35[8]);  // ../RTL/cmsdk_ahb_slave_mux.v(140)
  or u126 (n36[9], n34[9], n35[9]);  // ../RTL/cmsdk_ahb_slave_mux.v(140)
  or u127 (n36[10], n34[10], n35[10]);  // ../RTL/cmsdk_ahb_slave_mux.v(140)
  or u128 (n36[11], n34[11], n35[11]);  // ../RTL/cmsdk_ahb_slave_mux.v(140)
  or u129 (n36[12], n34[12], n35[12]);  // ../RTL/cmsdk_ahb_slave_mux.v(140)
  or u13 (HRDATA[10], n36[10], n37[10]);  // ../RTL/cmsdk_ahb_slave_mux.v(141)
  or u130 (n36[13], n34[13], n35[13]);  // ../RTL/cmsdk_ahb_slave_mux.v(140)
  or u131 (n36[14], n34[14], n35[14]);  // ../RTL/cmsdk_ahb_slave_mux.v(140)
  or u132 (n36[15], n34[15], n35[15]);  // ../RTL/cmsdk_ahb_slave_mux.v(140)
  or u133 (n36[16], n34[16], n35[16]);  // ../RTL/cmsdk_ahb_slave_mux.v(140)
  or u134 (n36[17], n34[17], n35[17]);  // ../RTL/cmsdk_ahb_slave_mux.v(140)
  or u135 (n36[18], n34[18], n35[18]);  // ../RTL/cmsdk_ahb_slave_mux.v(140)
  or u136 (n36[19], n34[19], n35[19]);  // ../RTL/cmsdk_ahb_slave_mux.v(140)
  or u137 (n36[20], n34[20], n35[20]);  // ../RTL/cmsdk_ahb_slave_mux.v(140)
  or u138 (n36[21], n34[21], n35[21]);  // ../RTL/cmsdk_ahb_slave_mux.v(140)
  or u139 (n36[22], n34[22], n35[22]);  // ../RTL/cmsdk_ahb_slave_mux.v(140)
  or u14 (HRDATA[6], n36[6], n37[6]);  // ../RTL/cmsdk_ahb_slave_mux.v(141)
  or u140 (n36[23], n34[23], n35[23]);  // ../RTL/cmsdk_ahb_slave_mux.v(140)
  or u141 (n36[24], n34[24], n35[24]);  // ../RTL/cmsdk_ahb_slave_mux.v(140)
  or u142 (n36[25], n34[25], n35[25]);  // ../RTL/cmsdk_ahb_slave_mux.v(140)
  or u143 (n36[26], n34[26], n35[26]);  // ../RTL/cmsdk_ahb_slave_mux.v(140)
  or u144 (n36[27], n34[27], n35[27]);  // ../RTL/cmsdk_ahb_slave_mux.v(140)
  or u145 (n36[28], n34[28], n35[28]);  // ../RTL/cmsdk_ahb_slave_mux.v(140)
  or u146 (n36[29], n34[29], n35[29]);  // ../RTL/cmsdk_ahb_slave_mux.v(140)
  or u147 (n36[30], n34[30], n35[30]);  // ../RTL/cmsdk_ahb_slave_mux.v(140)
  or u148 (n36[31], n34[31], n35[31]);  // ../RTL/cmsdk_ahb_slave_mux.v(140)
  and u149 (n35[1], reg_hsel[7], HRDATA7[1]);  // ../RTL/cmsdk_ahb_slave_mux.v(140)
  not u15 (n0, HRESETn);  // ../RTL/cmsdk_ahb_slave_mux.v(112)
  and u150 (n35[2], reg_hsel[7], HRDATA7[2]);  // ../RTL/cmsdk_ahb_slave_mux.v(140)
  and u151 (n35[3], reg_hsel[7], HRDATA7[3]);  // ../RTL/cmsdk_ahb_slave_mux.v(140)
  and u152 (n35[4], reg_hsel[7], HRDATA7[4]);  // ../RTL/cmsdk_ahb_slave_mux.v(140)
  and u153 (n35[5], reg_hsel[7], HRDATA7[5]);  // ../RTL/cmsdk_ahb_slave_mux.v(140)
  and u154 (n35[6], reg_hsel[7], HRDATA7[6]);  // ../RTL/cmsdk_ahb_slave_mux.v(140)
  and u155 (n35[7], reg_hsel[7], HRDATA7[7]);  // ../RTL/cmsdk_ahb_slave_mux.v(140)
  and u156 (n35[8], reg_hsel[7], HRDATA7[8]);  // ../RTL/cmsdk_ahb_slave_mux.v(140)
  and u157 (n35[9], reg_hsel[7], HRDATA7[9]);  // ../RTL/cmsdk_ahb_slave_mux.v(140)
  and u158 (n35[10], reg_hsel[7], HRDATA7[10]);  // ../RTL/cmsdk_ahb_slave_mux.v(140)
  and u159 (n35[11], reg_hsel[7], HRDATA7[11]);  // ../RTL/cmsdk_ahb_slave_mux.v(140)
  not u16 (n2, reg_hsel[0]);  // ../RTL/cmsdk_ahb_slave_mux.v(119)
  and u160 (n35[12], reg_hsel[7], HRDATA7[12]);  // ../RTL/cmsdk_ahb_slave_mux.v(140)
  and u161 (n35[13], reg_hsel[7], HRDATA7[13]);  // ../RTL/cmsdk_ahb_slave_mux.v(140)
  and u162 (n35[14], reg_hsel[7], HRDATA7[14]);  // ../RTL/cmsdk_ahb_slave_mux.v(140)
  and u163 (n35[15], reg_hsel[7], HRDATA7[15]);  // ../RTL/cmsdk_ahb_slave_mux.v(140)
  and u164 (n35[16], reg_hsel[7], HRDATA7[16]);  // ../RTL/cmsdk_ahb_slave_mux.v(140)
  and u165 (n35[17], reg_hsel[7], HRDATA7[17]);  // ../RTL/cmsdk_ahb_slave_mux.v(140)
  and u166 (n35[18], reg_hsel[7], HRDATA7[18]);  // ../RTL/cmsdk_ahb_slave_mux.v(140)
  and u167 (n35[19], reg_hsel[7], HRDATA7[19]);  // ../RTL/cmsdk_ahb_slave_mux.v(140)
  and u168 (n35[20], reg_hsel[7], HRDATA7[20]);  // ../RTL/cmsdk_ahb_slave_mux.v(140)
  and u169 (n35[21], reg_hsel[7], HRDATA7[21]);  // ../RTL/cmsdk_ahb_slave_mux.v(140)
  or u17 (n3, n2, HREADYOUT0);  // ../RTL/cmsdk_ahb_slave_mux.v(119)
  and u170 (n35[22], reg_hsel[7], HRDATA7[22]);  // ../RTL/cmsdk_ahb_slave_mux.v(140)
  and u171 (n35[23], reg_hsel[7], HRDATA7[23]);  // ../RTL/cmsdk_ahb_slave_mux.v(140)
  and u172 (n35[24], reg_hsel[7], HRDATA7[24]);  // ../RTL/cmsdk_ahb_slave_mux.v(140)
  and u173 (n35[25], reg_hsel[7], HRDATA7[25]);  // ../RTL/cmsdk_ahb_slave_mux.v(140)
  and u174 (n35[26], reg_hsel[7], HRDATA7[26]);  // ../RTL/cmsdk_ahb_slave_mux.v(140)
  and u175 (n35[27], reg_hsel[7], HRDATA7[27]);  // ../RTL/cmsdk_ahb_slave_mux.v(140)
  and u176 (n35[28], reg_hsel[7], HRDATA7[28]);  // ../RTL/cmsdk_ahb_slave_mux.v(140)
  and u177 (n35[29], reg_hsel[7], HRDATA7[29]);  // ../RTL/cmsdk_ahb_slave_mux.v(140)
  and u178 (n35[30], reg_hsel[7], HRDATA7[30]);  // ../RTL/cmsdk_ahb_slave_mux.v(140)
  and u179 (n35[31], reg_hsel[7], HRDATA7[31]);  // ../RTL/cmsdk_ahb_slave_mux.v(140)
  not u18 (n4, reg_hsel[1]);  // ../RTL/cmsdk_ahb_slave_mux.v(120)
  or u180 (n34[1], n32[1], n33[1]);  // ../RTL/cmsdk_ahb_slave_mux.v(139)
  or u181 (n34[2], n32[2], n33[2]);  // ../RTL/cmsdk_ahb_slave_mux.v(139)
  or u182 (n34[3], n32[3], n33[3]);  // ../RTL/cmsdk_ahb_slave_mux.v(139)
  or u183 (n34[4], n32[4], n33[4]);  // ../RTL/cmsdk_ahb_slave_mux.v(139)
  or u184 (n34[5], n32[5], n33[5]);  // ../RTL/cmsdk_ahb_slave_mux.v(139)
  or u185 (n34[6], n32[6], n33[6]);  // ../RTL/cmsdk_ahb_slave_mux.v(139)
  or u186 (n34[7], n32[7], n33[7]);  // ../RTL/cmsdk_ahb_slave_mux.v(139)
  or u187 (n34[8], n32[8], n33[8]);  // ../RTL/cmsdk_ahb_slave_mux.v(139)
  or u188 (n34[9], n32[9], n33[9]);  // ../RTL/cmsdk_ahb_slave_mux.v(139)
  or u189 (n34[10], n32[10], n33[10]);  // ../RTL/cmsdk_ahb_slave_mux.v(139)
  or u19 (n5, n4, HREADYOUT1);  // ../RTL/cmsdk_ahb_slave_mux.v(120)
  or u190 (n34[11], n32[11], n33[11]);  // ../RTL/cmsdk_ahb_slave_mux.v(139)
  or u191 (n34[12], n32[12], n33[12]);  // ../RTL/cmsdk_ahb_slave_mux.v(139)
  or u192 (n34[13], n32[13], n33[13]);  // ../RTL/cmsdk_ahb_slave_mux.v(139)
  or u193 (n34[14], n32[14], n33[14]);  // ../RTL/cmsdk_ahb_slave_mux.v(139)
  or u194 (n34[15], n32[15], n33[15]);  // ../RTL/cmsdk_ahb_slave_mux.v(139)
  or u195 (n34[16], n32[16], n33[16]);  // ../RTL/cmsdk_ahb_slave_mux.v(139)
  or u196 (n34[17], n32[17], n33[17]);  // ../RTL/cmsdk_ahb_slave_mux.v(139)
  or u197 (n34[18], n32[18], n33[18]);  // ../RTL/cmsdk_ahb_slave_mux.v(139)
  or u198 (n34[19], n32[19], n33[19]);  // ../RTL/cmsdk_ahb_slave_mux.v(139)
  or u199 (n34[20], n32[20], n33[20]);  // ../RTL/cmsdk_ahb_slave_mux.v(139)
  or u2 (HRDATA[8], n36[8], n37[8]);  // ../RTL/cmsdk_ahb_slave_mux.v(141)
  and u20 (n6, n3, n5);  // ../RTL/cmsdk_ahb_slave_mux.v(120)
  or u200 (n34[21], n32[21], n33[21]);  // ../RTL/cmsdk_ahb_slave_mux.v(139)
  or u201 (n34[22], n32[22], n33[22]);  // ../RTL/cmsdk_ahb_slave_mux.v(139)
  or u202 (n34[23], n32[23], n33[23]);  // ../RTL/cmsdk_ahb_slave_mux.v(139)
  or u203 (n34[24], n32[24], n33[24]);  // ../RTL/cmsdk_ahb_slave_mux.v(139)
  or u204 (n34[25], n32[25], n33[25]);  // ../RTL/cmsdk_ahb_slave_mux.v(139)
  or u205 (n34[26], n32[26], n33[26]);  // ../RTL/cmsdk_ahb_slave_mux.v(139)
  or u206 (n34[27], n32[27], n33[27]);  // ../RTL/cmsdk_ahb_slave_mux.v(139)
  or u207 (n34[28], n32[28], n33[28]);  // ../RTL/cmsdk_ahb_slave_mux.v(139)
  or u208 (n34[29], n32[29], n33[29]);  // ../RTL/cmsdk_ahb_slave_mux.v(139)
  or u209 (n34[30], n32[30], n33[30]);  // ../RTL/cmsdk_ahb_slave_mux.v(139)
  or u21 (HRDATA[5], n36[5], n37[5]);  // ../RTL/cmsdk_ahb_slave_mux.v(141)
  or u210 (n34[31], n32[31], n33[31]);  // ../RTL/cmsdk_ahb_slave_mux.v(139)
  and u211 (n33[1], reg_hsel[6], HRDATA6[1]);  // ../RTL/cmsdk_ahb_slave_mux.v(139)
  and u212 (n33[2], reg_hsel[6], HRDATA6[2]);  // ../RTL/cmsdk_ahb_slave_mux.v(139)
  and u213 (n33[3], reg_hsel[6], HRDATA6[3]);  // ../RTL/cmsdk_ahb_slave_mux.v(139)
  and u214 (n33[4], reg_hsel[6], HRDATA6[4]);  // ../RTL/cmsdk_ahb_slave_mux.v(139)
  and u215 (n33[5], reg_hsel[6], HRDATA6[5]);  // ../RTL/cmsdk_ahb_slave_mux.v(139)
  and u216 (n33[6], reg_hsel[6], HRDATA6[6]);  // ../RTL/cmsdk_ahb_slave_mux.v(139)
  and u217 (n33[7], reg_hsel[6], HRDATA6[7]);  // ../RTL/cmsdk_ahb_slave_mux.v(139)
  and u218 (n33[8], reg_hsel[6], HRDATA6[8]);  // ../RTL/cmsdk_ahb_slave_mux.v(139)
  and u219 (n33[9], reg_hsel[6], HRDATA6[9]);  // ../RTL/cmsdk_ahb_slave_mux.v(139)
  or u22 (HRDATA[4], n36[4], n37[4]);  // ../RTL/cmsdk_ahb_slave_mux.v(141)
  and u220 (n33[10], reg_hsel[6], HRDATA6[10]);  // ../RTL/cmsdk_ahb_slave_mux.v(139)
  and u221 (n33[11], reg_hsel[6], HRDATA6[11]);  // ../RTL/cmsdk_ahb_slave_mux.v(139)
  and u222 (n33[12], reg_hsel[6], HRDATA6[12]);  // ../RTL/cmsdk_ahb_slave_mux.v(139)
  and u223 (n33[13], reg_hsel[6], HRDATA6[13]);  // ../RTL/cmsdk_ahb_slave_mux.v(139)
  and u224 (n33[14], reg_hsel[6], HRDATA6[14]);  // ../RTL/cmsdk_ahb_slave_mux.v(139)
  and u225 (n33[15], reg_hsel[6], HRDATA6[15]);  // ../RTL/cmsdk_ahb_slave_mux.v(139)
  and u226 (n33[16], reg_hsel[6], HRDATA6[16]);  // ../RTL/cmsdk_ahb_slave_mux.v(139)
  and u227 (n33[17], reg_hsel[6], HRDATA6[17]);  // ../RTL/cmsdk_ahb_slave_mux.v(139)
  and u228 (n33[18], reg_hsel[6], HRDATA6[18]);  // ../RTL/cmsdk_ahb_slave_mux.v(139)
  and u229 (n33[19], reg_hsel[6], HRDATA6[19]);  // ../RTL/cmsdk_ahb_slave_mux.v(139)
  not u23 (n7, reg_hsel[3]);  // ../RTL/cmsdk_ahb_slave_mux.v(122)
  and u230 (n33[20], reg_hsel[6], HRDATA6[20]);  // ../RTL/cmsdk_ahb_slave_mux.v(139)
  and u231 (n33[21], reg_hsel[6], HRDATA6[21]);  // ../RTL/cmsdk_ahb_slave_mux.v(139)
  and u232 (n33[22], reg_hsel[6], HRDATA6[22]);  // ../RTL/cmsdk_ahb_slave_mux.v(139)
  and u233 (n33[23], reg_hsel[6], HRDATA6[23]);  // ../RTL/cmsdk_ahb_slave_mux.v(139)
  and u234 (n33[24], reg_hsel[6], HRDATA6[24]);  // ../RTL/cmsdk_ahb_slave_mux.v(139)
  and u235 (n33[25], reg_hsel[6], HRDATA6[25]);  // ../RTL/cmsdk_ahb_slave_mux.v(139)
  and u236 (n33[26], reg_hsel[6], HRDATA6[26]);  // ../RTL/cmsdk_ahb_slave_mux.v(139)
  and u237 (n33[27], reg_hsel[6], HRDATA6[27]);  // ../RTL/cmsdk_ahb_slave_mux.v(139)
  and u238 (n33[28], reg_hsel[6], HRDATA6[28]);  // ../RTL/cmsdk_ahb_slave_mux.v(139)
  and u239 (n33[29], reg_hsel[6], HRDATA6[29]);  // ../RTL/cmsdk_ahb_slave_mux.v(139)
  or u24 (n8, n7, HREADYOUT3);  // ../RTL/cmsdk_ahb_slave_mux.v(122)
  and u240 (n33[30], reg_hsel[6], HRDATA6[30]);  // ../RTL/cmsdk_ahb_slave_mux.v(139)
  and u241 (n33[31], reg_hsel[6], HRDATA6[31]);  // ../RTL/cmsdk_ahb_slave_mux.v(139)
  or u242 (n32[1], n30[1], n31[1]);  // ../RTL/cmsdk_ahb_slave_mux.v(138)
  or u243 (n32[2], n30[2], n31[2]);  // ../RTL/cmsdk_ahb_slave_mux.v(138)
  or u244 (n32[3], n30[3], n31[3]);  // ../RTL/cmsdk_ahb_slave_mux.v(138)
  or u245 (n32[4], n30[4], n31[4]);  // ../RTL/cmsdk_ahb_slave_mux.v(138)
  or u246 (n32[5], n30[5], n31[5]);  // ../RTL/cmsdk_ahb_slave_mux.v(138)
  or u247 (n32[6], n30[6], n31[6]);  // ../RTL/cmsdk_ahb_slave_mux.v(138)
  or u248 (n32[7], n30[7], n31[7]);  // ../RTL/cmsdk_ahb_slave_mux.v(138)
  or u249 (n32[8], n30[8], n31[8]);  // ../RTL/cmsdk_ahb_slave_mux.v(138)
  and u25 (n9, n6, n8);  // ../RTL/cmsdk_ahb_slave_mux.v(122)
  or u250 (n32[9], n30[9], n31[9]);  // ../RTL/cmsdk_ahb_slave_mux.v(138)
  or u251 (n32[10], n30[10], n31[10]);  // ../RTL/cmsdk_ahb_slave_mux.v(138)
  or u252 (n32[11], n30[11], n31[11]);  // ../RTL/cmsdk_ahb_slave_mux.v(138)
  or u253 (n32[12], n30[12], n31[12]);  // ../RTL/cmsdk_ahb_slave_mux.v(138)
  or u254 (n32[13], n30[13], n31[13]);  // ../RTL/cmsdk_ahb_slave_mux.v(138)
  or u255 (n32[14], n30[14], n31[14]);  // ../RTL/cmsdk_ahb_slave_mux.v(138)
  or u256 (n32[15], n30[15], n31[15]);  // ../RTL/cmsdk_ahb_slave_mux.v(138)
  or u257 (n32[16], n30[16], n31[16]);  // ../RTL/cmsdk_ahb_slave_mux.v(138)
  or u258 (n32[17], n30[17], n31[17]);  // ../RTL/cmsdk_ahb_slave_mux.v(138)
  or u259 (n32[18], n30[18], n31[18]);  // ../RTL/cmsdk_ahb_slave_mux.v(138)
  not u26 (n10, reg_hsel[4]);  // ../RTL/cmsdk_ahb_slave_mux.v(123)
  or u260 (n32[19], n30[19], n31[19]);  // ../RTL/cmsdk_ahb_slave_mux.v(138)
  or u261 (n32[20], n30[20], n31[20]);  // ../RTL/cmsdk_ahb_slave_mux.v(138)
  or u262 (n32[21], n30[21], n31[21]);  // ../RTL/cmsdk_ahb_slave_mux.v(138)
  or u263 (n32[22], n30[22], n31[22]);  // ../RTL/cmsdk_ahb_slave_mux.v(138)
  or u264 (n32[23], n30[23], n31[23]);  // ../RTL/cmsdk_ahb_slave_mux.v(138)
  or u265 (n32[24], n30[24], n31[24]);  // ../RTL/cmsdk_ahb_slave_mux.v(138)
  or u266 (n32[25], n30[25], n31[25]);  // ../RTL/cmsdk_ahb_slave_mux.v(138)
  or u267 (n32[26], n30[26], n31[26]);  // ../RTL/cmsdk_ahb_slave_mux.v(138)
  or u268 (n32[27], n30[27], n31[27]);  // ../RTL/cmsdk_ahb_slave_mux.v(138)
  or u269 (n32[28], n30[28], n31[28]);  // ../RTL/cmsdk_ahb_slave_mux.v(138)
  or u27 (n11, n10, HREADYOUT4);  // ../RTL/cmsdk_ahb_slave_mux.v(123)
  or u270 (n32[29], n30[29], n31[29]);  // ../RTL/cmsdk_ahb_slave_mux.v(138)
  or u271 (n32[30], n30[30], n31[30]);  // ../RTL/cmsdk_ahb_slave_mux.v(138)
  or u272 (n32[31], n30[31], n31[31]);  // ../RTL/cmsdk_ahb_slave_mux.v(138)
  and u273 (n31[1], reg_hsel[5], HRDATA5[1]);  // ../RTL/cmsdk_ahb_slave_mux.v(138)
  and u274 (n31[2], reg_hsel[5], HRDATA5[2]);  // ../RTL/cmsdk_ahb_slave_mux.v(138)
  and u275 (n31[3], reg_hsel[5], HRDATA5[3]);  // ../RTL/cmsdk_ahb_slave_mux.v(138)
  and u276 (n31[4], reg_hsel[5], HRDATA5[4]);  // ../RTL/cmsdk_ahb_slave_mux.v(138)
  and u277 (n31[5], reg_hsel[5], HRDATA5[5]);  // ../RTL/cmsdk_ahb_slave_mux.v(138)
  and u278 (n31[6], reg_hsel[5], HRDATA5[6]);  // ../RTL/cmsdk_ahb_slave_mux.v(138)
  and u279 (n31[7], reg_hsel[5], HRDATA5[7]);  // ../RTL/cmsdk_ahb_slave_mux.v(138)
  and u28 (n12, n9, n11);  // ../RTL/cmsdk_ahb_slave_mux.v(123)
  and u280 (n31[8], reg_hsel[5], HRDATA5[8]);  // ../RTL/cmsdk_ahb_slave_mux.v(138)
  and u281 (n31[9], reg_hsel[5], HRDATA5[9]);  // ../RTL/cmsdk_ahb_slave_mux.v(138)
  and u282 (n31[10], reg_hsel[5], HRDATA5[10]);  // ../RTL/cmsdk_ahb_slave_mux.v(138)
  and u283 (n31[11], reg_hsel[5], HRDATA5[11]);  // ../RTL/cmsdk_ahb_slave_mux.v(138)
  and u284 (n31[12], reg_hsel[5], HRDATA5[12]);  // ../RTL/cmsdk_ahb_slave_mux.v(138)
  and u285 (n31[13], reg_hsel[5], HRDATA5[13]);  // ../RTL/cmsdk_ahb_slave_mux.v(138)
  and u286 (n31[14], reg_hsel[5], HRDATA5[14]);  // ../RTL/cmsdk_ahb_slave_mux.v(138)
  and u287 (n31[15], reg_hsel[5], HRDATA5[15]);  // ../RTL/cmsdk_ahb_slave_mux.v(138)
  and u288 (n31[16], reg_hsel[5], HRDATA5[16]);  // ../RTL/cmsdk_ahb_slave_mux.v(138)
  and u289 (n31[17], reg_hsel[5], HRDATA5[17]);  // ../RTL/cmsdk_ahb_slave_mux.v(138)
  not u29 (n13, reg_hsel[5]);  // ../RTL/cmsdk_ahb_slave_mux.v(124)
  and u290 (n31[18], reg_hsel[5], HRDATA5[18]);  // ../RTL/cmsdk_ahb_slave_mux.v(138)
  and u291 (n31[19], reg_hsel[5], HRDATA5[19]);  // ../RTL/cmsdk_ahb_slave_mux.v(138)
  and u292 (n31[20], reg_hsel[5], HRDATA5[20]);  // ../RTL/cmsdk_ahb_slave_mux.v(138)
  and u293 (n31[21], reg_hsel[5], HRDATA5[21]);  // ../RTL/cmsdk_ahb_slave_mux.v(138)
  and u294 (n31[22], reg_hsel[5], HRDATA5[22]);  // ../RTL/cmsdk_ahb_slave_mux.v(138)
  and u295 (n31[23], reg_hsel[5], HRDATA5[23]);  // ../RTL/cmsdk_ahb_slave_mux.v(138)
  and u296 (n31[24], reg_hsel[5], HRDATA5[24]);  // ../RTL/cmsdk_ahb_slave_mux.v(138)
  and u297 (n31[25], reg_hsel[5], HRDATA5[25]);  // ../RTL/cmsdk_ahb_slave_mux.v(138)
  and u298 (n31[26], reg_hsel[5], HRDATA5[26]);  // ../RTL/cmsdk_ahb_slave_mux.v(138)
  and u299 (n31[27], reg_hsel[5], HRDATA5[27]);  // ../RTL/cmsdk_ahb_slave_mux.v(138)
  or u3 (HRDATA[7], n36[7], n37[7]);  // ../RTL/cmsdk_ahb_slave_mux.v(141)
  or u30 (n14, n13, HREADYOUT5);  // ../RTL/cmsdk_ahb_slave_mux.v(124)
  and u300 (n31[28], reg_hsel[5], HRDATA5[28]);  // ../RTL/cmsdk_ahb_slave_mux.v(138)
  and u301 (n31[29], reg_hsel[5], HRDATA5[29]);  // ../RTL/cmsdk_ahb_slave_mux.v(138)
  and u302 (n31[30], reg_hsel[5], HRDATA5[30]);  // ../RTL/cmsdk_ahb_slave_mux.v(138)
  and u303 (n31[31], reg_hsel[5], HRDATA5[31]);  // ../RTL/cmsdk_ahb_slave_mux.v(138)
  or u304 (n30[1], n28[1], n29[1]);  // ../RTL/cmsdk_ahb_slave_mux.v(137)
  or u305 (n30[2], n28[2], n29[2]);  // ../RTL/cmsdk_ahb_slave_mux.v(137)
  or u306 (n30[3], n28[3], n29[3]);  // ../RTL/cmsdk_ahb_slave_mux.v(137)
  or u307 (n30[4], n28[4], n29[4]);  // ../RTL/cmsdk_ahb_slave_mux.v(137)
  or u308 (n30[5], n28[5], n29[5]);  // ../RTL/cmsdk_ahb_slave_mux.v(137)
  or u309 (n30[6], n28[6], n29[6]);  // ../RTL/cmsdk_ahb_slave_mux.v(137)
  and u31 (n15, n12, n14);  // ../RTL/cmsdk_ahb_slave_mux.v(124)
  or u310 (n30[7], n28[7], n29[7]);  // ../RTL/cmsdk_ahb_slave_mux.v(137)
  or u311 (n30[8], n28[8], n29[8]);  // ../RTL/cmsdk_ahb_slave_mux.v(137)
  or u312 (n30[9], n28[9], n29[9]);  // ../RTL/cmsdk_ahb_slave_mux.v(137)
  or u313 (n30[10], n28[10], n29[10]);  // ../RTL/cmsdk_ahb_slave_mux.v(137)
  or u314 (n30[11], n28[11], n29[11]);  // ../RTL/cmsdk_ahb_slave_mux.v(137)
  or u315 (n30[12], n28[12], n29[12]);  // ../RTL/cmsdk_ahb_slave_mux.v(137)
  or u316 (n30[13], n28[13], n29[13]);  // ../RTL/cmsdk_ahb_slave_mux.v(137)
  or u317 (n30[14], n28[14], n29[14]);  // ../RTL/cmsdk_ahb_slave_mux.v(137)
  or u318 (n30[15], n28[15], n29[15]);  // ../RTL/cmsdk_ahb_slave_mux.v(137)
  or u319 (n30[16], n28[16], n29[16]);  // ../RTL/cmsdk_ahb_slave_mux.v(137)
  not u32 (n16, reg_hsel[6]);  // ../RTL/cmsdk_ahb_slave_mux.v(125)
  or u320 (n30[17], n28[17], n29[17]);  // ../RTL/cmsdk_ahb_slave_mux.v(137)
  or u321 (n30[18], n28[18], n29[18]);  // ../RTL/cmsdk_ahb_slave_mux.v(137)
  or u322 (n30[19], n28[19], n29[19]);  // ../RTL/cmsdk_ahb_slave_mux.v(137)
  or u323 (n30[20], n28[20], n29[20]);  // ../RTL/cmsdk_ahb_slave_mux.v(137)
  or u324 (n30[21], n28[21], n29[21]);  // ../RTL/cmsdk_ahb_slave_mux.v(137)
  or u325 (n30[22], n28[22], n29[22]);  // ../RTL/cmsdk_ahb_slave_mux.v(137)
  or u326 (n30[23], n28[23], n29[23]);  // ../RTL/cmsdk_ahb_slave_mux.v(137)
  or u327 (n30[24], n28[24], n29[24]);  // ../RTL/cmsdk_ahb_slave_mux.v(137)
  or u328 (n30[25], n28[25], n29[25]);  // ../RTL/cmsdk_ahb_slave_mux.v(137)
  or u329 (n30[26], n28[26], n29[26]);  // ../RTL/cmsdk_ahb_slave_mux.v(137)
  or u33 (n17, n16, HREADYOUT6);  // ../RTL/cmsdk_ahb_slave_mux.v(125)
  or u330 (n30[27], n28[27], n29[27]);  // ../RTL/cmsdk_ahb_slave_mux.v(137)
  or u331 (n30[28], n28[28], n29[28]);  // ../RTL/cmsdk_ahb_slave_mux.v(137)
  or u332 (n30[29], n28[29], n29[29]);  // ../RTL/cmsdk_ahb_slave_mux.v(137)
  or u333 (n30[30], n28[30], n29[30]);  // ../RTL/cmsdk_ahb_slave_mux.v(137)
  or u334 (n30[31], n28[31], n29[31]);  // ../RTL/cmsdk_ahb_slave_mux.v(137)
  and u335 (n29[1], reg_hsel[4], HRDATA4[1]);  // ../RTL/cmsdk_ahb_slave_mux.v(137)
  and u336 (n29[2], reg_hsel[4], HRDATA4[2]);  // ../RTL/cmsdk_ahb_slave_mux.v(137)
  and u337 (n29[3], reg_hsel[4], HRDATA4[3]);  // ../RTL/cmsdk_ahb_slave_mux.v(137)
  and u338 (n29[4], reg_hsel[4], HRDATA4[4]);  // ../RTL/cmsdk_ahb_slave_mux.v(137)
  and u339 (n29[5], reg_hsel[4], HRDATA4[5]);  // ../RTL/cmsdk_ahb_slave_mux.v(137)
  and u34 (n18, n15, n17);  // ../RTL/cmsdk_ahb_slave_mux.v(125)
  and u340 (n29[6], reg_hsel[4], HRDATA4[6]);  // ../RTL/cmsdk_ahb_slave_mux.v(137)
  and u341 (n29[7], reg_hsel[4], HRDATA4[7]);  // ../RTL/cmsdk_ahb_slave_mux.v(137)
  and u342 (n29[8], reg_hsel[4], HRDATA4[8]);  // ../RTL/cmsdk_ahb_slave_mux.v(137)
  and u343 (n29[9], reg_hsel[4], HRDATA4[9]);  // ../RTL/cmsdk_ahb_slave_mux.v(137)
  and u344 (n29[10], reg_hsel[4], HRDATA4[10]);  // ../RTL/cmsdk_ahb_slave_mux.v(137)
  and u345 (n29[11], reg_hsel[4], HRDATA4[11]);  // ../RTL/cmsdk_ahb_slave_mux.v(137)
  and u346 (n29[12], reg_hsel[4], HRDATA4[12]);  // ../RTL/cmsdk_ahb_slave_mux.v(137)
  and u347 (n29[13], reg_hsel[4], HRDATA4[13]);  // ../RTL/cmsdk_ahb_slave_mux.v(137)
  and u348 (n29[14], reg_hsel[4], HRDATA4[14]);  // ../RTL/cmsdk_ahb_slave_mux.v(137)
  and u349 (n29[15], reg_hsel[4], HRDATA4[15]);  // ../RTL/cmsdk_ahb_slave_mux.v(137)
  not u35 (n19, reg_hsel[7]);  // ../RTL/cmsdk_ahb_slave_mux.v(126)
  and u350 (n29[16], reg_hsel[4], HRDATA4[16]);  // ../RTL/cmsdk_ahb_slave_mux.v(137)
  and u351 (n29[17], reg_hsel[4], HRDATA4[17]);  // ../RTL/cmsdk_ahb_slave_mux.v(137)
  and u352 (n29[18], reg_hsel[4], HRDATA4[18]);  // ../RTL/cmsdk_ahb_slave_mux.v(137)
  and u353 (n29[19], reg_hsel[4], HRDATA4[19]);  // ../RTL/cmsdk_ahb_slave_mux.v(137)
  and u354 (n29[20], reg_hsel[4], HRDATA4[20]);  // ../RTL/cmsdk_ahb_slave_mux.v(137)
  and u355 (n29[21], reg_hsel[4], HRDATA4[21]);  // ../RTL/cmsdk_ahb_slave_mux.v(137)
  and u356 (n29[22], reg_hsel[4], HRDATA4[22]);  // ../RTL/cmsdk_ahb_slave_mux.v(137)
  and u357 (n29[23], reg_hsel[4], HRDATA4[23]);  // ../RTL/cmsdk_ahb_slave_mux.v(137)
  and u358 (n29[24], reg_hsel[4], HRDATA4[24]);  // ../RTL/cmsdk_ahb_slave_mux.v(137)
  and u359 (n29[25], reg_hsel[4], HRDATA4[25]);  // ../RTL/cmsdk_ahb_slave_mux.v(137)
  or u36 (n20, n19, HREADYOUT7);  // ../RTL/cmsdk_ahb_slave_mux.v(126)
  and u360 (n29[26], reg_hsel[4], HRDATA4[26]);  // ../RTL/cmsdk_ahb_slave_mux.v(137)
  and u361 (n29[27], reg_hsel[4], HRDATA4[27]);  // ../RTL/cmsdk_ahb_slave_mux.v(137)
  and u362 (n29[28], reg_hsel[4], HRDATA4[28]);  // ../RTL/cmsdk_ahb_slave_mux.v(137)
  and u363 (n29[29], reg_hsel[4], HRDATA4[29]);  // ../RTL/cmsdk_ahb_slave_mux.v(137)
  and u364 (n29[30], reg_hsel[4], HRDATA4[30]);  // ../RTL/cmsdk_ahb_slave_mux.v(137)
  and u365 (n29[31], reg_hsel[4], HRDATA4[31]);  // ../RTL/cmsdk_ahb_slave_mux.v(137)
  or u366 (n28[1], n26[1], n27[1]);  // ../RTL/cmsdk_ahb_slave_mux.v(136)
  or u367 (n28[2], n26[2], n27[2]);  // ../RTL/cmsdk_ahb_slave_mux.v(136)
  or u368 (n28[3], n26[3], n27[3]);  // ../RTL/cmsdk_ahb_slave_mux.v(136)
  or u369 (n28[4], n26[4], n27[4]);  // ../RTL/cmsdk_ahb_slave_mux.v(136)
  and u37 (n21, n18, n20);  // ../RTL/cmsdk_ahb_slave_mux.v(126)
  or u370 (n28[5], n26[5], n27[5]);  // ../RTL/cmsdk_ahb_slave_mux.v(136)
  or u371 (n28[6], n26[6], n27[6]);  // ../RTL/cmsdk_ahb_slave_mux.v(136)
  or u372 (n28[7], n26[7], n27[7]);  // ../RTL/cmsdk_ahb_slave_mux.v(136)
  or u373 (n28[8], n26[8], n27[8]);  // ../RTL/cmsdk_ahb_slave_mux.v(136)
  or u374 (n28[9], n26[9], n27[9]);  // ../RTL/cmsdk_ahb_slave_mux.v(136)
  or u375 (n28[10], n26[10], n27[10]);  // ../RTL/cmsdk_ahb_slave_mux.v(136)
  or u376 (n28[11], n26[11], n27[11]);  // ../RTL/cmsdk_ahb_slave_mux.v(136)
  or u377 (n28[12], n26[12], n27[12]);  // ../RTL/cmsdk_ahb_slave_mux.v(136)
  or u378 (n28[13], n26[13], n27[13]);  // ../RTL/cmsdk_ahb_slave_mux.v(136)
  or u379 (n28[14], n26[14], n27[14]);  // ../RTL/cmsdk_ahb_slave_mux.v(136)
  not u38 (n22, reg_hsel[8]);  // ../RTL/cmsdk_ahb_slave_mux.v(127)
  or u380 (n28[15], n26[15], n27[15]);  // ../RTL/cmsdk_ahb_slave_mux.v(136)
  or u381 (n28[16], n26[16], n27[16]);  // ../RTL/cmsdk_ahb_slave_mux.v(136)
  or u382 (n28[17], n26[17], n27[17]);  // ../RTL/cmsdk_ahb_slave_mux.v(136)
  or u383 (n28[18], n26[18], n27[18]);  // ../RTL/cmsdk_ahb_slave_mux.v(136)
  or u384 (n28[19], n26[19], n27[19]);  // ../RTL/cmsdk_ahb_slave_mux.v(136)
  or u385 (n28[20], n26[20], n27[20]);  // ../RTL/cmsdk_ahb_slave_mux.v(136)
  or u386 (n28[21], n26[21], n27[21]);  // ../RTL/cmsdk_ahb_slave_mux.v(136)
  or u387 (n28[22], n26[22], n27[22]);  // ../RTL/cmsdk_ahb_slave_mux.v(136)
  or u388 (n28[23], n26[23], n27[23]);  // ../RTL/cmsdk_ahb_slave_mux.v(136)
  or u389 (n28[24], n26[24], n27[24]);  // ../RTL/cmsdk_ahb_slave_mux.v(136)
  or u39 (n23, n22, HREADYOUT8);  // ../RTL/cmsdk_ahb_slave_mux.v(127)
  or u390 (n28[25], n26[25], n27[25]);  // ../RTL/cmsdk_ahb_slave_mux.v(136)
  or u391 (n28[26], n26[26], n27[26]);  // ../RTL/cmsdk_ahb_slave_mux.v(136)
  or u392 (n28[27], n26[27], n27[27]);  // ../RTL/cmsdk_ahb_slave_mux.v(136)
  or u393 (n28[28], n26[28], n27[28]);  // ../RTL/cmsdk_ahb_slave_mux.v(136)
  or u394 (n28[29], n26[29], n27[29]);  // ../RTL/cmsdk_ahb_slave_mux.v(136)
  or u395 (n28[30], n26[30], n27[30]);  // ../RTL/cmsdk_ahb_slave_mux.v(136)
  or u396 (n28[31], n26[31], n27[31]);  // ../RTL/cmsdk_ahb_slave_mux.v(136)
  and u397 (n27[1], reg_hsel[3], HRDATA3[1]);  // ../RTL/cmsdk_ahb_slave_mux.v(136)
  and u398 (n27[2], reg_hsel[3], HRDATA3[2]);  // ../RTL/cmsdk_ahb_slave_mux.v(136)
  and u399 (n27[3], reg_hsel[3], HRDATA3[3]);  // ../RTL/cmsdk_ahb_slave_mux.v(136)
  or u4 (HRDATA[19], n36[19], n37[19]);  // ../RTL/cmsdk_ahb_slave_mux.v(141)
  and u40 (mux_hready, n21, n23);  // ../RTL/cmsdk_ahb_slave_mux.v(127)
  and u400 (n27[4], reg_hsel[3], HRDATA3[4]);  // ../RTL/cmsdk_ahb_slave_mux.v(136)
  and u401 (n27[5], reg_hsel[3], HRDATA3[5]);  // ../RTL/cmsdk_ahb_slave_mux.v(136)
  and u402 (n27[6], reg_hsel[3], HRDATA3[6]);  // ../RTL/cmsdk_ahb_slave_mux.v(136)
  and u403 (n27[7], reg_hsel[3], HRDATA3[7]);  // ../RTL/cmsdk_ahb_slave_mux.v(136)
  and u404 (n27[8], reg_hsel[3], HRDATA3[8]);  // ../RTL/cmsdk_ahb_slave_mux.v(136)
  and u405 (n27[9], reg_hsel[3], HRDATA3[9]);  // ../RTL/cmsdk_ahb_slave_mux.v(136)
  and u406 (n27[10], reg_hsel[3], HRDATA3[10]);  // ../RTL/cmsdk_ahb_slave_mux.v(136)
  and u407 (n27[11], reg_hsel[3], HRDATA3[11]);  // ../RTL/cmsdk_ahb_slave_mux.v(136)
  and u408 (n27[12], reg_hsel[3], HRDATA3[12]);  // ../RTL/cmsdk_ahb_slave_mux.v(136)
  and u409 (n27[13], reg_hsel[3], HRDATA3[13]);  // ../RTL/cmsdk_ahb_slave_mux.v(136)
  or u41 (HRDATA[3], n36[3], n37[3]);  // ../RTL/cmsdk_ahb_slave_mux.v(141)
  and u410 (n27[14], reg_hsel[3], HRDATA3[14]);  // ../RTL/cmsdk_ahb_slave_mux.v(136)
  and u411 (n27[15], reg_hsel[3], HRDATA3[15]);  // ../RTL/cmsdk_ahb_slave_mux.v(136)
  and u412 (n27[16], reg_hsel[3], HRDATA3[16]);  // ../RTL/cmsdk_ahb_slave_mux.v(136)
  and u413 (n27[17], reg_hsel[3], HRDATA3[17]);  // ../RTL/cmsdk_ahb_slave_mux.v(136)
  and u414 (n27[18], reg_hsel[3], HRDATA3[18]);  // ../RTL/cmsdk_ahb_slave_mux.v(136)
  and u415 (n27[19], reg_hsel[3], HRDATA3[19]);  // ../RTL/cmsdk_ahb_slave_mux.v(136)
  and u416 (n27[20], reg_hsel[3], HRDATA3[20]);  // ../RTL/cmsdk_ahb_slave_mux.v(136)
  and u417 (n27[21], reg_hsel[3], HRDATA3[21]);  // ../RTL/cmsdk_ahb_slave_mux.v(136)
  and u418 (n27[22], reg_hsel[3], HRDATA3[22]);  // ../RTL/cmsdk_ahb_slave_mux.v(136)
  and u419 (n27[23], reg_hsel[3], HRDATA3[23]);  // ../RTL/cmsdk_ahb_slave_mux.v(136)
  or u42 (HRDATA[2], n36[2], n37[2]);  // ../RTL/cmsdk_ahb_slave_mux.v(141)
  and u420 (n27[24], reg_hsel[3], HRDATA3[24]);  // ../RTL/cmsdk_ahb_slave_mux.v(136)
  and u421 (n27[25], reg_hsel[3], HRDATA3[25]);  // ../RTL/cmsdk_ahb_slave_mux.v(136)
  and u422 (n27[26], reg_hsel[3], HRDATA3[26]);  // ../RTL/cmsdk_ahb_slave_mux.v(136)
  and u423 (n27[27], reg_hsel[3], HRDATA3[27]);  // ../RTL/cmsdk_ahb_slave_mux.v(136)
  and u424 (n27[28], reg_hsel[3], HRDATA3[28]);  // ../RTL/cmsdk_ahb_slave_mux.v(136)
  and u425 (n27[29], reg_hsel[3], HRDATA3[29]);  // ../RTL/cmsdk_ahb_slave_mux.v(136)
  and u426 (n27[30], reg_hsel[3], HRDATA3[30]);  // ../RTL/cmsdk_ahb_slave_mux.v(136)
  and u427 (n27[31], reg_hsel[3], HRDATA3[31]);  // ../RTL/cmsdk_ahb_slave_mux.v(136)
  or u428 (n26[1], n24[1], n25[1]);  // ../RTL/cmsdk_ahb_slave_mux.v(134)
  or u429 (n26[2], n24[2], n25[2]);  // ../RTL/cmsdk_ahb_slave_mux.v(134)
  buf u43 (HREADYOUT, mux_hready);  // ../RTL/cmsdk_ahb_slave_mux.v(130)
  or u430 (n26[3], n24[3], n25[3]);  // ../RTL/cmsdk_ahb_slave_mux.v(134)
  or u431 (n26[4], n24[4], n25[4]);  // ../RTL/cmsdk_ahb_slave_mux.v(134)
  or u432 (n26[5], n24[5], n25[5]);  // ../RTL/cmsdk_ahb_slave_mux.v(134)
  or u433 (n26[6], n24[6], n25[6]);  // ../RTL/cmsdk_ahb_slave_mux.v(134)
  or u434 (n26[7], n24[7], n25[7]);  // ../RTL/cmsdk_ahb_slave_mux.v(134)
  or u435 (n26[8], n24[8], n25[8]);  // ../RTL/cmsdk_ahb_slave_mux.v(134)
  or u436 (n26[9], n24[9], n25[9]);  // ../RTL/cmsdk_ahb_slave_mux.v(134)
  or u437 (n26[10], n24[10], n25[10]);  // ../RTL/cmsdk_ahb_slave_mux.v(134)
  or u438 (n26[11], n24[11], n25[11]);  // ../RTL/cmsdk_ahb_slave_mux.v(134)
  or u439 (n26[12], n24[12], n25[12]);  // ../RTL/cmsdk_ahb_slave_mux.v(134)
  and u44 (n25[0], reg_hsel[1], HRDATA1[0]);  // ../RTL/cmsdk_ahb_slave_mux.v(133)
  or u440 (n26[13], n24[13], n25[13]);  // ../RTL/cmsdk_ahb_slave_mux.v(134)
  or u441 (n26[14], n24[14], n25[14]);  // ../RTL/cmsdk_ahb_slave_mux.v(134)
  or u442 (n26[15], n24[15], n25[15]);  // ../RTL/cmsdk_ahb_slave_mux.v(134)
  or u443 (n26[16], n24[16], n25[16]);  // ../RTL/cmsdk_ahb_slave_mux.v(134)
  or u444 (n26[17], n24[17], n25[17]);  // ../RTL/cmsdk_ahb_slave_mux.v(134)
  or u445 (n26[18], n24[18], n25[18]);  // ../RTL/cmsdk_ahb_slave_mux.v(134)
  or u446 (n26[19], n24[19], n25[19]);  // ../RTL/cmsdk_ahb_slave_mux.v(134)
  or u447 (n26[20], n24[20], n25[20]);  // ../RTL/cmsdk_ahb_slave_mux.v(134)
  or u448 (n26[21], n24[21], n25[21]);  // ../RTL/cmsdk_ahb_slave_mux.v(134)
  or u449 (n26[22], n24[22], n25[22]);  // ../RTL/cmsdk_ahb_slave_mux.v(134)
  or u45 (HRDATA[20], n36[20], n37[20]);  // ../RTL/cmsdk_ahb_slave_mux.v(141)
  or u450 (n26[23], n24[23], n25[23]);  // ../RTL/cmsdk_ahb_slave_mux.v(134)
  or u451 (n26[24], n24[24], n25[24]);  // ../RTL/cmsdk_ahb_slave_mux.v(134)
  or u452 (n26[25], n24[25], n25[25]);  // ../RTL/cmsdk_ahb_slave_mux.v(134)
  or u453 (n26[26], n24[26], n25[26]);  // ../RTL/cmsdk_ahb_slave_mux.v(134)
  or u454 (n26[27], n24[27], n25[27]);  // ../RTL/cmsdk_ahb_slave_mux.v(134)
  or u455 (n26[28], n24[28], n25[28]);  // ../RTL/cmsdk_ahb_slave_mux.v(134)
  or u456 (n26[29], n24[29], n25[29]);  // ../RTL/cmsdk_ahb_slave_mux.v(134)
  or u457 (n26[30], n24[30], n25[30]);  // ../RTL/cmsdk_ahb_slave_mux.v(134)
  or u458 (n26[31], n24[31], n25[31]);  // ../RTL/cmsdk_ahb_slave_mux.v(134)
  buf u459 (nxt_hsel_reg[1], HSEL1);  // ../RTL/cmsdk_ahb_slave_mux.v(107)
  buf u46 (nxt_hsel_reg[0], HSEL0);  // ../RTL/cmsdk_ahb_slave_mux.v(107)
  buf u460 (nxt_hsel_reg[2], 1'b0);  // ../RTL/cmsdk_ahb_slave_mux.v(107)
  buf u461 (nxt_hsel_reg[3], HSEL3);  // ../RTL/cmsdk_ahb_slave_mux.v(107)
  buf u462 (nxt_hsel_reg[4], HSEL4);  // ../RTL/cmsdk_ahb_slave_mux.v(107)
  buf u463 (nxt_hsel_reg[5], HSEL5);  // ../RTL/cmsdk_ahb_slave_mux.v(107)
  buf u464 (nxt_hsel_reg[6], HSEL6);  // ../RTL/cmsdk_ahb_slave_mux.v(107)
  buf u465 (nxt_hsel_reg[7], HSEL7);  // ../RTL/cmsdk_ahb_slave_mux.v(107)
  buf u466 (nxt_hsel_reg[8], HSEL8);  // ../RTL/cmsdk_ahb_slave_mux.v(107)
  buf u467 (nxt_hsel_reg[9], 1'b0);  // ../RTL/cmsdk_ahb_slave_mux.v(107)
  and u468 (n25[1], reg_hsel[1], HRDATA1[1]);  // ../RTL/cmsdk_ahb_slave_mux.v(133)
  and u469 (n25[2], reg_hsel[1], HRDATA1[2]);  // ../RTL/cmsdk_ahb_slave_mux.v(133)
  or u47 (n26[0], n24[0], n25[0]);  // ../RTL/cmsdk_ahb_slave_mux.v(134)
  and u470 (n25[3], reg_hsel[1], HRDATA1[3]);  // ../RTL/cmsdk_ahb_slave_mux.v(133)
  and u471 (n25[4], reg_hsel[1], HRDATA1[4]);  // ../RTL/cmsdk_ahb_slave_mux.v(133)
  and u472 (n25[5], reg_hsel[1], HRDATA1[5]);  // ../RTL/cmsdk_ahb_slave_mux.v(133)
  and u473 (n25[6], reg_hsel[1], HRDATA1[6]);  // ../RTL/cmsdk_ahb_slave_mux.v(133)
  and u474 (n25[7], reg_hsel[1], HRDATA1[7]);  // ../RTL/cmsdk_ahb_slave_mux.v(133)
  and u475 (n25[8], reg_hsel[1], HRDATA1[8]);  // ../RTL/cmsdk_ahb_slave_mux.v(133)
  and u476 (n25[9], reg_hsel[1], HRDATA1[9]);  // ../RTL/cmsdk_ahb_slave_mux.v(133)
  and u477 (n25[10], reg_hsel[1], HRDATA1[10]);  // ../RTL/cmsdk_ahb_slave_mux.v(133)
  and u478 (n25[11], reg_hsel[1], HRDATA1[11]);  // ../RTL/cmsdk_ahb_slave_mux.v(133)
  and u479 (n25[12], reg_hsel[1], HRDATA1[12]);  // ../RTL/cmsdk_ahb_slave_mux.v(133)
  and u48 (n27[0], reg_hsel[3], HRDATA3[0]);  // ../RTL/cmsdk_ahb_slave_mux.v(136)
  and u480 (n25[13], reg_hsel[1], HRDATA1[13]);  // ../RTL/cmsdk_ahb_slave_mux.v(133)
  and u481 (n25[14], reg_hsel[1], HRDATA1[14]);  // ../RTL/cmsdk_ahb_slave_mux.v(133)
  and u482 (n25[15], reg_hsel[1], HRDATA1[15]);  // ../RTL/cmsdk_ahb_slave_mux.v(133)
  and u483 (n25[16], reg_hsel[1], HRDATA1[16]);  // ../RTL/cmsdk_ahb_slave_mux.v(133)
  and u484 (n25[17], reg_hsel[1], HRDATA1[17]);  // ../RTL/cmsdk_ahb_slave_mux.v(133)
  and u485 (n25[18], reg_hsel[1], HRDATA1[18]);  // ../RTL/cmsdk_ahb_slave_mux.v(133)
  and u486 (n25[19], reg_hsel[1], HRDATA1[19]);  // ../RTL/cmsdk_ahb_slave_mux.v(133)
  and u487 (n25[20], reg_hsel[1], HRDATA1[20]);  // ../RTL/cmsdk_ahb_slave_mux.v(133)
  and u488 (n25[21], reg_hsel[1], HRDATA1[21]);  // ../RTL/cmsdk_ahb_slave_mux.v(133)
  and u489 (n25[22], reg_hsel[1], HRDATA1[22]);  // ../RTL/cmsdk_ahb_slave_mux.v(133)
  or u49 (n28[0], n26[0], n27[0]);  // ../RTL/cmsdk_ahb_slave_mux.v(136)
  and u490 (n25[23], reg_hsel[1], HRDATA1[23]);  // ../RTL/cmsdk_ahb_slave_mux.v(133)
  and u491 (n25[24], reg_hsel[1], HRDATA1[24]);  // ../RTL/cmsdk_ahb_slave_mux.v(133)
  and u492 (n25[25], reg_hsel[1], HRDATA1[25]);  // ../RTL/cmsdk_ahb_slave_mux.v(133)
  and u493 (n25[26], reg_hsel[1], HRDATA1[26]);  // ../RTL/cmsdk_ahb_slave_mux.v(133)
  and u494 (n25[27], reg_hsel[1], HRDATA1[27]);  // ../RTL/cmsdk_ahb_slave_mux.v(133)
  and u495 (n25[28], reg_hsel[1], HRDATA1[28]);  // ../RTL/cmsdk_ahb_slave_mux.v(133)
  and u496 (n25[29], reg_hsel[1], HRDATA1[29]);  // ../RTL/cmsdk_ahb_slave_mux.v(133)
  and u497 (n25[30], reg_hsel[1], HRDATA1[30]);  // ../RTL/cmsdk_ahb_slave_mux.v(133)
  and u498 (n25[31], reg_hsel[1], HRDATA1[31]);  // ../RTL/cmsdk_ahb_slave_mux.v(133)
  and u499 (n24[0], reg_hsel[0], HRDATA0[0]);  // ../RTL/cmsdk_ahb_slave_mux.v(133)
  or u5 (HRDATA[18], n36[18], n37[18]);  // ../RTL/cmsdk_ahb_slave_mux.v(141)
  and u50 (n29[0], reg_hsel[4], HRDATA4[0]);  // ../RTL/cmsdk_ahb_slave_mux.v(137)
  and u500 (n24[1], reg_hsel[0], HRDATA0[1]);  // ../RTL/cmsdk_ahb_slave_mux.v(133)
  and u501 (n24[2], reg_hsel[0], HRDATA0[2]);  // ../RTL/cmsdk_ahb_slave_mux.v(133)
  and u502 (n24[3], reg_hsel[0], HRDATA0[3]);  // ../RTL/cmsdk_ahb_slave_mux.v(133)
  and u503 (n24[4], reg_hsel[0], HRDATA0[4]);  // ../RTL/cmsdk_ahb_slave_mux.v(133)
  and u504 (n24[5], reg_hsel[0], HRDATA0[5]);  // ../RTL/cmsdk_ahb_slave_mux.v(133)
  and u505 (n24[6], reg_hsel[0], HRDATA0[6]);  // ../RTL/cmsdk_ahb_slave_mux.v(133)
  and u506 (n24[7], reg_hsel[0], HRDATA0[7]);  // ../RTL/cmsdk_ahb_slave_mux.v(133)
  and u507 (n24[8], reg_hsel[0], HRDATA0[8]);  // ../RTL/cmsdk_ahb_slave_mux.v(133)
  and u508 (n24[9], reg_hsel[0], HRDATA0[9]);  // ../RTL/cmsdk_ahb_slave_mux.v(133)
  and u509 (n24[10], reg_hsel[0], HRDATA0[10]);  // ../RTL/cmsdk_ahb_slave_mux.v(133)
  or u51 (n30[0], n28[0], n29[0]);  // ../RTL/cmsdk_ahb_slave_mux.v(137)
  and u510 (n24[11], reg_hsel[0], HRDATA0[11]);  // ../RTL/cmsdk_ahb_slave_mux.v(133)
  and u511 (n24[12], reg_hsel[0], HRDATA0[12]);  // ../RTL/cmsdk_ahb_slave_mux.v(133)
  and u512 (n24[13], reg_hsel[0], HRDATA0[13]);  // ../RTL/cmsdk_ahb_slave_mux.v(133)
  and u513 (n24[14], reg_hsel[0], HRDATA0[14]);  // ../RTL/cmsdk_ahb_slave_mux.v(133)
  and u514 (n24[15], reg_hsel[0], HRDATA0[15]);  // ../RTL/cmsdk_ahb_slave_mux.v(133)
  and u515 (n24[16], reg_hsel[0], HRDATA0[16]);  // ../RTL/cmsdk_ahb_slave_mux.v(133)
  and u516 (n24[17], reg_hsel[0], HRDATA0[17]);  // ../RTL/cmsdk_ahb_slave_mux.v(133)
  and u517 (n24[18], reg_hsel[0], HRDATA0[18]);  // ../RTL/cmsdk_ahb_slave_mux.v(133)
  and u518 (n24[19], reg_hsel[0], HRDATA0[19]);  // ../RTL/cmsdk_ahb_slave_mux.v(133)
  and u519 (n24[20], reg_hsel[0], HRDATA0[20]);  // ../RTL/cmsdk_ahb_slave_mux.v(133)
  and u52 (n31[0], reg_hsel[5], HRDATA5[0]);  // ../RTL/cmsdk_ahb_slave_mux.v(138)
  and u520 (n24[21], reg_hsel[0], HRDATA0[21]);  // ../RTL/cmsdk_ahb_slave_mux.v(133)
  and u521 (n24[22], reg_hsel[0], HRDATA0[22]);  // ../RTL/cmsdk_ahb_slave_mux.v(133)
  and u522 (n24[23], reg_hsel[0], HRDATA0[23]);  // ../RTL/cmsdk_ahb_slave_mux.v(133)
  and u523 (n24[24], reg_hsel[0], HRDATA0[24]);  // ../RTL/cmsdk_ahb_slave_mux.v(133)
  and u524 (n24[25], reg_hsel[0], HRDATA0[25]);  // ../RTL/cmsdk_ahb_slave_mux.v(133)
  and u525 (n24[26], reg_hsel[0], HRDATA0[26]);  // ../RTL/cmsdk_ahb_slave_mux.v(133)
  and u526 (n24[27], reg_hsel[0], HRDATA0[27]);  // ../RTL/cmsdk_ahb_slave_mux.v(133)
  and u527 (n24[28], reg_hsel[0], HRDATA0[28]);  // ../RTL/cmsdk_ahb_slave_mux.v(133)
  and u528 (n24[29], reg_hsel[0], HRDATA0[29]);  // ../RTL/cmsdk_ahb_slave_mux.v(133)
  and u529 (n24[30], reg_hsel[0], HRDATA0[30]);  // ../RTL/cmsdk_ahb_slave_mux.v(133)
  or u53 (n32[0], n30[0], n31[0]);  // ../RTL/cmsdk_ahb_slave_mux.v(138)
  and u530 (n24[31], reg_hsel[0], HRDATA0[31]);  // ../RTL/cmsdk_ahb_slave_mux.v(133)
  and u54 (n33[0], reg_hsel[6], HRDATA6[0]);  // ../RTL/cmsdk_ahb_slave_mux.v(139)
  or u55 (n34[0], n32[0], n33[0]);  // ../RTL/cmsdk_ahb_slave_mux.v(139)
  and u56 (n35[0], reg_hsel[7], HRDATA7[0]);  // ../RTL/cmsdk_ahb_slave_mux.v(140)
  or u57 (n36[0], n34[0], n35[0]);  // ../RTL/cmsdk_ahb_slave_mux.v(140)
  and u58 (n37[0], reg_hsel[8], HRDATA8[0]);  // ../RTL/cmsdk_ahb_slave_mux.v(141)
  and u59 (n38, reg_hsel[0], HRESP0);  // ../RTL/cmsdk_ahb_slave_mux.v(145)
  or u6 (HRDATA[17], n36[17], n37[17]);  // ../RTL/cmsdk_ahb_slave_mux.v(141)
  and u60 (n39, reg_hsel[1], HRESP1);  // ../RTL/cmsdk_ahb_slave_mux.v(146)
  or u61 (n40, n38, n39);  // ../RTL/cmsdk_ahb_slave_mux.v(146)
  or u62 (HRDATA[1], n36[1], n37[1]);  // ../RTL/cmsdk_ahb_slave_mux.v(141)
  and u63 (n41, reg_hsel[3], HRESP3);  // ../RTL/cmsdk_ahb_slave_mux.v(148)
  or u64 (n42, n40, n41);  // ../RTL/cmsdk_ahb_slave_mux.v(148)
  and u65 (n43, reg_hsel[4], HRESP4);  // ../RTL/cmsdk_ahb_slave_mux.v(149)
  or u66 (n44, n42, n43);  // ../RTL/cmsdk_ahb_slave_mux.v(149)
  and u67 (n45, reg_hsel[5], HRESP5);  // ../RTL/cmsdk_ahb_slave_mux.v(150)
  or u68 (n46, n44, n45);  // ../RTL/cmsdk_ahb_slave_mux.v(150)
  and u69 (n47, reg_hsel[6], HRESP6);  // ../RTL/cmsdk_ahb_slave_mux.v(151)
  or u7 (HRDATA[16], n36[16], n37[16]);  // ../RTL/cmsdk_ahb_slave_mux.v(141)
  or u70 (n48, n46, n47);  // ../RTL/cmsdk_ahb_slave_mux.v(151)
  and u71 (n49, reg_hsel[7], HRESP7);  // ../RTL/cmsdk_ahb_slave_mux.v(152)
  or u72 (n50, n48, n49);  // ../RTL/cmsdk_ahb_slave_mux.v(152)
  and u73 (n51, reg_hsel[8], HRESP8);  // ../RTL/cmsdk_ahb_slave_mux.v(153)
  or u74 (HRESP, n50, n51);  // ../RTL/cmsdk_ahb_slave_mux.v(153)
  or u75 (HRDATA[0], n36[0], n37[0]);  // ../RTL/cmsdk_ahb_slave_mux.v(141)
  or u76 (HRDATA[21], n36[21], n37[21]);  // ../RTL/cmsdk_ahb_slave_mux.v(141)
  or u77 (HRDATA[22], n36[22], n37[22]);  // ../RTL/cmsdk_ahb_slave_mux.v(141)
  or u78 (HRDATA[23], n36[23], n37[23]);  // ../RTL/cmsdk_ahb_slave_mux.v(141)
  or u79 (HRDATA[24], n36[24], n37[24]);  // ../RTL/cmsdk_ahb_slave_mux.v(141)
  or u8 (HRDATA[15], n36[15], n37[15]);  // ../RTL/cmsdk_ahb_slave_mux.v(141)
  or u80 (HRDATA[25], n36[25], n37[25]);  // ../RTL/cmsdk_ahb_slave_mux.v(141)
  or u81 (HRDATA[26], n36[26], n37[26]);  // ../RTL/cmsdk_ahb_slave_mux.v(141)
  or u82 (HRDATA[27], n36[27], n37[27]);  // ../RTL/cmsdk_ahb_slave_mux.v(141)
  or u83 (HRDATA[28], n36[28], n37[28]);  // ../RTL/cmsdk_ahb_slave_mux.v(141)
  or u84 (HRDATA[29], n36[29], n37[29]);  // ../RTL/cmsdk_ahb_slave_mux.v(141)
  or u85 (HRDATA[30], n36[30], n37[30]);  // ../RTL/cmsdk_ahb_slave_mux.v(141)
  or u86 (HRDATA[31], n36[31], n37[31]);  // ../RTL/cmsdk_ahb_slave_mux.v(141)
  and u87 (n37[1], reg_hsel[8], HRDATA8[1]);  // ../RTL/cmsdk_ahb_slave_mux.v(141)
  and u88 (n37[2], reg_hsel[8], HRDATA8[2]);  // ../RTL/cmsdk_ahb_slave_mux.v(141)
  and u89 (n37[3], reg_hsel[8], HRDATA8[3]);  // ../RTL/cmsdk_ahb_slave_mux.v(141)
  or u9 (HRDATA[14], n36[14], n37[14]);  // ../RTL/cmsdk_ahb_slave_mux.v(141)
  and u90 (n37[4], reg_hsel[8], HRDATA8[4]);  // ../RTL/cmsdk_ahb_slave_mux.v(141)
  and u91 (n37[5], reg_hsel[8], HRDATA8[5]);  // ../RTL/cmsdk_ahb_slave_mux.v(141)
  and u92 (n37[6], reg_hsel[8], HRDATA8[6]);  // ../RTL/cmsdk_ahb_slave_mux.v(141)
  and u93 (n37[7], reg_hsel[8], HRDATA8[7]);  // ../RTL/cmsdk_ahb_slave_mux.v(141)
  and u94 (n37[8], reg_hsel[8], HRDATA8[8]);  // ../RTL/cmsdk_ahb_slave_mux.v(141)
  and u95 (n37[9], reg_hsel[8], HRDATA8[9]);  // ../RTL/cmsdk_ahb_slave_mux.v(141)
  and u96 (n37[10], reg_hsel[8], HRDATA8[10]);  // ../RTL/cmsdk_ahb_slave_mux.v(141)
  and u97 (n37[11], reg_hsel[8], HRDATA8[11]);  // ../RTL/cmsdk_ahb_slave_mux.v(141)
  and u98 (n37[12], reg_hsel[8], HRDATA8[12]);  // ../RTL/cmsdk_ahb_slave_mux.v(141)
  and u99 (n37[13], reg_hsel[8], HRDATA8[13]);  // ../RTL/cmsdk_ahb_slave_mux.v(141)

endmodule 

module \cmsdk_apb_subsystem_m0ds(INCLUDE_APB_TEST_SLAVE=0,INCLUDE_APB_TIMER1=0,INCLUDE_APB_DUALTIMER0=0,INCLUDE_APB_UART1=0,INCLUDE_APB_UART2=0,INCLUDE_APB_UART3=0,INCLUDE_APB_UART4=0,INCLUDE_APB_WATCHDOG=0)   // ../RTL/cmsdk_apb_subsystem_m0ds.v(26)
  (
  HADDR,
  HCLK,
  HPROT,
  HREADY,
  HRESETn,
  HSEL,
  HSIZE,
  HTRANS,
  HWDATA,
  HWRITE,
  PCLK,
  PCLKEN,
  PCLKG,
  PRESETn,
  ext12_prdata,
  ext12_pready,
  ext12_pslverr,
  ext13_prdata,
  ext13_pready,
  ext13_pslverr,
  ext14_prdata,
  ext14_pready,
  ext14_pslverr,
  ext15_prdata,
  ext15_pready,
  ext15_pslverr,
  timer0_extin,
  timer1_extin,
  uart0_rxd,
  APBACTIVE,
  HRDATA,
  HREADYOUT,
  HRESP,
  PADDR,
  PENABLE,
  PWDATA,
  PWRITE,
  apbsubsys_interrupt,
  ext12_psel,
  ext13_psel,
  ext14_psel,
  ext15_psel,
  uart0_txd,
  uart0_txen,
  watchdog_interrupt,
  watchdog_reset,
  b_pad_gpio_porta
  );

  input [15:0] HADDR;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(88)
  input HCLK;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(84)
  input [3:0] HPROT;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(92)
  input HREADY;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(93)
  input HRESETn;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(85)
  input HSEL;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(87)
  input [2:0] HSIZE;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(91)
  input [1:0] HTRANS;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(89)
  input [31:0] HWDATA;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(94)
  input HWRITE;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(90)
  input PCLK;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(99)
  input PCLKEN;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(101)
  input PCLKG;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(100)
  input PRESETn;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(102)
  input [31:0] ext12_prdata;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(114)
  input ext12_pready;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(115)
  input ext12_pslverr;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(116)
  input [31:0] ext13_prdata;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(118)
  input ext13_pready;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(119)
  input ext13_pslverr;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(120)
  input [31:0] ext14_prdata;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(122)
  input ext14_pready;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(123)
  input ext14_pslverr;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(124)
  input [31:0] ext15_prdata;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(126)
  input ext15_pready;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(127)
  input ext15_pslverr;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(128)
  input timer0_extin;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(159)
  input timer1_extin;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(160)
  input uart0_rxd;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(134)
  output APBACTIVE;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(130)
  output [31:0] HRDATA;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(96)
  output HREADYOUT;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(95)
  output HRESP;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(97)
  output [11:0] PADDR;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(104)
  output PENABLE;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(107)
  output [31:0] PWDATA;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(106)
  output PWRITE;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(105)
  output [31:0] apbsubsys_interrupt;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(163)
  output ext12_psel;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(109)
  output ext13_psel;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(110)
  output ext14_psel;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(111)
  output ext15_psel;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(112)
  output uart0_txd;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(135)
  output uart0_txen;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(136)
  output watchdog_interrupt;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(164)
  output watchdog_reset;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(165)
  inout [7:0] b_pad_gpio_porta;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(156)

  parameter APB_EXT_PORT12_ENABLE = 0;
  parameter APB_EXT_PORT13_ENABLE = 0;
  parameter APB_EXT_PORT14_ENABLE = 0;
  parameter APB_EXT_PORT15_ENABLE = 0;
  parameter BE = 0;
  parameter INCLUDE_APB_DUALTIMER0 = 0;
  parameter INCLUDE_APB_GPIO0 = 1;
  parameter INCLUDE_APB_TEST_SLAVE = 0;
  parameter INCLUDE_APB_TIMER1 = 0;
  parameter INCLUDE_APB_UART0 = 1;
  parameter INCLUDE_APB_UART1 = 0;
  parameter INCLUDE_APB_UART2 = 0;
  parameter INCLUDE_APB_UART3 = 0;
  parameter INCLUDE_APB_UART4 = 0;
  parameter INCLUDE_APB_WATCHDOG = 0;
  parameter INCLUDE_IRQ_SYNCHRONIZER = 0;
  wire [31:0] dualtimer2_prdata;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(195)
  wire [7:0] gpio0_intr;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(240)
  wire [31:0] gpio0_prdata;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(185)
  wire [31:0] hrdata_le;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(317)
  wire [31:0] hrdata_mux_1;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(343)
  wire [31:0] hwdata_le;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(316)
  wire [31:0] hwdata_mux_1;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(335)
  wire [7:0] i_gpio0_intr;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(306)
  wire [15:0] i_paddr;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(170)
  wire [31:0] i_prdata_mux;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(180)
  wire [31:0] i_pwdata;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(176)
  wire [1:0] n5;
  wire [1:0] nxt_be_swap_ctrl;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(320)
  wire [1:0] reg_be_swap_ctrl;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(319)
  wire [31:0] test_slave_prdata;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(230)
  wire [31:0] timer1_prdata;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(190)
  wire [31:0] uart0_prdata;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(205)
  wire bigendian;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(313)
  wire dualtimer2_comb_int;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(244)
  wire dualtimer2_pready;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(196)
  wire dualtimer2_pslverr;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(197)
  wire gpio0_pready;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(186)
  wire gpio0_psel;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(184)
  wire gpio0_pslverr;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(187)
  wire i_dualtimer2_int;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(308)
  wire i_penable;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(172)
  wire i_pready_mux;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(179)
  wire i_psel;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(171)
  wire i_pslverr_mux;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(181)
  wire i_pwrite;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(173)
  wire i_timer1_int;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(307)
  wire i_uart0_overflow_int;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(291)
  wire i_uart0_rxint;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(290)
  wire i_uart0_txint;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(289)
  wire i_watchdog_int;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(309)
  wire i_watchdog_rst;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(310)
  wire n0;
  wire n1;
  wire n2;
  wire n3;
  wire n4;
  wire n6;
  wire n7;
  wire reg_be_swap_ctrl_en;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(318)
  wire test_slave_pready;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(231)
  wire test_slave_pslverr;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(232)
  wire timer1_int;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(241)
  wire timer1_pready;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(191)
  wire timer1_pslverr;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(192)
  wire uart0_overflow_int;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(278)
  wire uart0_pready;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(206)
  wire uart0_psel;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(204)
  wire uart0_pslverr;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(207)
  wire uart0_rxint;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(247)
  wire uart0_rxovrint;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(249)
  wire uart0_txint;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(246)
  wire uart0_txovrint;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(248)
  wire watchdog_int;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(285)
  wire watchdog_rst;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(286)

  eq_w2 eq0 (
    .i0(HSIZE[1:0]),
    .i1(2'b10),
    .o(n2));  // ../RTL/cmsdk_apb_subsystem_m0ds.v(322)
  gpio gen_apb_gpio_0$u_gpio_0 (
    .paddr(i_paddr[6:2]),
    .pclk(PCLK),
    .pclk_intr(1'b1),
    .penable(i_penable),
    .presetn(PRESETn),
    .psel(gpio0_psel),
    .pwdata(i_pwdata),
    .pwrite(i_pwrite),
    .gpio_intr(gpio0_intr),
    .prdata(gpio0_prdata),
    .pready(gpio0_pready),
    .pslverr(gpio0_pslverr),
    .b_pad_gpio_porta(b_pad_gpio_porta));  // ../RTL/cmsdk_apb_subsystem_m0ds.v(503)
  cmsdk_apb_uart gen_apb_uart_0$u_apb_uart_0 (
    .ECOREVNUM(4'b0000),
    .PADDR(i_paddr[11:2]),
    .PCLK(PCLK),
    .PCLKG(PCLKG),
    .PENABLE(i_penable),
    .PRESETn(PRESETn),
    .PSEL(uart0_psel),
    .PWDATA(i_pwdata),
    .PWRITE(i_pwrite),
    .RXD(uart0_rxd),
    .PRDATA(uart0_prdata),
    .PREADY(uart0_pready),
    .PSLVERR(uart0_pslverr),
    .RXINT(uart0_rxint),
    .RXOVRINT(uart0_rxovrint),
    .TXD(uart0_txd),
    .TXEN(uart0_txen),
    .TXINT(uart0_txint),
    .TXOVRINT(uart0_txovrint));  // ../RTL/cmsdk_apb_subsystem_m0ds.v(643)
  binary_mux_s1_w2 mux0 (
    .i0(reg_be_swap_ctrl),
    .i1(nxt_be_swap_ctrl),
    .sel(reg_be_swap_ctrl_en),
    .o(n5));  // ../RTL/cmsdk_apb_subsystem_m0ds.v(331)
  binary_mux_s1_w32 mux1 (
    .i0(HWDATA),
    .i1({HWDATA[23:16],HWDATA[31:24],HWDATA[7:0],HWDATA[15:8]}),
    .sel(n6),
    .o(hwdata_mux_1));  // ../RTL/cmsdk_apb_subsystem_m0ds.v(337)
  binary_mux_s1_w32 mux2 (
    .i0(hwdata_mux_1),
    .i1({hwdata_mux_1[15:0],hwdata_mux_1[31:16]}),
    .sel(n7),
    .o(hwdata_le));  // ../RTL/cmsdk_apb_subsystem_m0ds.v(341)
  binary_mux_s1_w32 mux3 (
    .i0(hrdata_le),
    .i1({hrdata_le[23:16],hrdata_le[31:24],hrdata_le[7:0],hrdata_le[15:8]}),
    .sel(n6),
    .o(hrdata_mux_1));  // ../RTL/cmsdk_apb_subsystem_m0ds.v(345)
  binary_mux_s1_w32 mux4 (
    .i0(hrdata_mux_1),
    .i1({hrdata_mux_1[15:0],hrdata_mux_1[31:16]}),
    .sel(n7),
    .o(HRDATA));  // ../RTL/cmsdk_apb_subsystem_m0ds.v(349)
  ne_w2 neq0 (
    .i0(HSIZE[1:0]),
    .i1(2'b00),
    .o(n3));  // ../RTL/cmsdk_apb_subsystem_m0ds.v(323)
  reg_ar_as_w2 reg0 (
    .clk(HCLK),
    .d(n5),
    .reset({n4,n4}),
    .set(2'b00),
    .q(reg_be_swap_ctrl));  // ../RTL/cmsdk_apb_subsystem_m0ds.v(331)
  buf u10 (apbsubsys_interrupt[7], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(1064)
  buf u100 (PWDATA[24], i_pwdata[24]);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(903)
  buf u101 (PWDATA[25], i_pwdata[25]);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(903)
  buf u102 (PWDATA[26], i_pwdata[26]);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(903)
  buf u103 (PWDATA[27], i_pwdata[27]);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(903)
  buf u104 (PWDATA[28], i_pwdata[28]);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(903)
  buf u105 (PWDATA[29], i_pwdata[29]);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(903)
  buf u106 (PWDATA[30], i_pwdata[30]);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(903)
  buf u107 (PWDATA[31], i_pwdata[31]);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(903)
  buf u108 (PADDR[1], i_paddr[1]);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(900)
  buf u109 (PADDR[2], i_paddr[2]);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(900)
  not u11 (n4, HRESETn);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(328)
  buf u110 (PADDR[3], i_paddr[3]);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(900)
  buf u111 (PADDR[4], i_paddr[4]);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(900)
  buf u112 (PADDR[5], i_paddr[5]);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(900)
  buf u113 (PADDR[6], i_paddr[6]);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(900)
  buf u114 (PADDR[7], i_paddr[7]);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(900)
  buf u115 (PADDR[8], i_paddr[8]);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(900)
  buf u116 (PADDR[9], i_paddr[9]);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(900)
  buf u117 (PADDR[10], i_paddr[10]);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(900)
  buf u118 (PADDR[11], i_paddr[11]);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(900)
  buf u119 (test_slave_prdata[1], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(894)
  and u12 (n6, reg_be_swap_ctrl[0], bigendian);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(335)
  buf u120 (test_slave_prdata[2], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(894)
  buf u121 (test_slave_prdata[3], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(894)
  buf u122 (test_slave_prdata[4], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(894)
  buf u123 (test_slave_prdata[5], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(894)
  buf u124 (test_slave_prdata[6], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(894)
  buf u125 (test_slave_prdata[7], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(894)
  buf u126 (test_slave_prdata[8], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(894)
  buf u127 (test_slave_prdata[9], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(894)
  buf u128 (test_slave_prdata[10], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(894)
  buf u129 (test_slave_prdata[11], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(894)
  and u13 (n7, reg_be_swap_ctrl[1], bigendian);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(339)
  buf u130 (test_slave_prdata[12], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(894)
  buf u131 (test_slave_prdata[13], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(894)
  buf u132 (test_slave_prdata[14], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(894)
  buf u133 (test_slave_prdata[15], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(894)
  buf u134 (test_slave_prdata[16], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(894)
  buf u135 (test_slave_prdata[17], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(894)
  buf u136 (test_slave_prdata[18], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(894)
  buf u137 (test_slave_prdata[19], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(894)
  buf u138 (test_slave_prdata[20], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(894)
  buf u139 (test_slave_prdata[21], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(894)
  buf u14 (apbsubsys_interrupt[1], i_uart0_txint);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(1064)
  buf u140 (test_slave_prdata[22], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(894)
  buf u141 (test_slave_prdata[23], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(894)
  buf u142 (test_slave_prdata[24], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(894)
  buf u143 (test_slave_prdata[25], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(894)
  buf u144 (test_slave_prdata[26], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(894)
  buf u145 (test_slave_prdata[27], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(894)
  buf u146 (test_slave_prdata[28], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(894)
  buf u147 (test_slave_prdata[29], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(894)
  buf u148 (test_slave_prdata[30], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(894)
  buf u149 (test_slave_prdata[31], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(894)
  buf u15 (apbsubsys_interrupt[0], i_uart0_rxint);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(1064)
  buf u150 (dualtimer2_prdata[1], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(590)
  buf u151 (dualtimer2_prdata[2], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(590)
  buf u152 (dualtimer2_prdata[3], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(590)
  buf u153 (dualtimer2_prdata[4], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(590)
  buf u154 (dualtimer2_prdata[5], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(590)
  buf u155 (dualtimer2_prdata[6], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(590)
  buf u156 (dualtimer2_prdata[7], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(590)
  buf u157 (dualtimer2_prdata[8], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(590)
  buf u158 (dualtimer2_prdata[9], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(590)
  buf u159 (dualtimer2_prdata[10], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(590)
  and u16 (nxt_be_swap_ctrl[0], bigendian, n3);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(322)
  buf u160 (dualtimer2_prdata[11], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(590)
  buf u161 (dualtimer2_prdata[12], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(590)
  buf u162 (dualtimer2_prdata[13], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(590)
  buf u163 (dualtimer2_prdata[14], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(590)
  buf u164 (dualtimer2_prdata[15], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(590)
  buf u165 (dualtimer2_prdata[16], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(590)
  buf u166 (dualtimer2_prdata[17], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(590)
  buf u167 (dualtimer2_prdata[18], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(590)
  buf u168 (dualtimer2_prdata[19], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(590)
  buf u169 (dualtimer2_prdata[20], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(590)
  buf u17 (timer1_pready, 1'b1);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(556)
  buf u170 (dualtimer2_prdata[21], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(590)
  buf u171 (dualtimer2_prdata[22], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(590)
  buf u172 (dualtimer2_prdata[23], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(590)
  buf u173 (dualtimer2_prdata[24], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(590)
  buf u174 (dualtimer2_prdata[25], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(590)
  buf u175 (dualtimer2_prdata[26], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(590)
  buf u176 (dualtimer2_prdata[27], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(590)
  buf u177 (dualtimer2_prdata[28], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(590)
  buf u178 (dualtimer2_prdata[29], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(590)
  buf u179 (dualtimer2_prdata[30], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(590)
  buf u18 (timer1_pslverr, 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(557)
  buf u180 (dualtimer2_prdata[31], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(590)
  buf u181 (timer1_prdata[1], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(555)
  buf u182 (timer1_prdata[2], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(555)
  buf u183 (timer1_prdata[3], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(555)
  buf u184 (timer1_prdata[4], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(555)
  buf u185 (timer1_prdata[5], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(555)
  buf u186 (timer1_prdata[6], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(555)
  buf u187 (timer1_prdata[7], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(555)
  buf u188 (timer1_prdata[8], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(555)
  buf u189 (timer1_prdata[9], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(555)
  buf u19 (timer1_int, 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(558)
  buf u190 (timer1_prdata[10], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(555)
  buf u191 (timer1_prdata[11], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(555)
  buf u192 (timer1_prdata[12], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(555)
  buf u193 (timer1_prdata[13], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(555)
  buf u194 (timer1_prdata[14], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(555)
  buf u195 (timer1_prdata[15], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(555)
  buf u196 (timer1_prdata[16], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(555)
  buf u197 (timer1_prdata[17], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(555)
  buf u198 (timer1_prdata[18], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(555)
  buf u199 (timer1_prdata[19], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(555)
  buf u2 (apbsubsys_interrupt[9], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(1064)
  buf u20 (timer1_prdata[0], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(555)
  buf u200 (timer1_prdata[20], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(555)
  buf u201 (timer1_prdata[21], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(555)
  buf u202 (timer1_prdata[22], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(555)
  buf u203 (timer1_prdata[23], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(555)
  buf u204 (timer1_prdata[24], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(555)
  buf u205 (timer1_prdata[25], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(555)
  buf u206 (timer1_prdata[26], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(555)
  buf u207 (timer1_prdata[27], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(555)
  buf u208 (timer1_prdata[28], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(555)
  buf u209 (timer1_prdata[29], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(555)
  buf u21 (dualtimer2_comb_int, 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(591)
  buf u210 (timer1_prdata[30], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(555)
  buf u211 (timer1_prdata[31], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(555)
  and u212 (nxt_be_swap_ctrl[1], bigendian, n2);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(322)
  buf u22 (apbsubsys_interrupt[6], i_dualtimer2_int);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(1064)
  buf u23 (apbsubsys_interrupt[5], i_timer1_int);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(1064)
  buf u24 (dualtimer2_pslverr, 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(598)
  buf u25 (dualtimer2_pready, 1'b1);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(599)
  buf u26 (apbsubsys_interrupt[4], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(1064)
  buf u27 (watchdog_int, 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(631)
  buf u28 (watchdog_rst, 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(632)
  buf u29 (apbsubsys_interrupt[3], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(1064)
  buf u3 (apbsubsys_interrupt[8], i_uart0_overflow_int);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(1064)
  buf u30 (apbsubsys_interrupt[2], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(1064)
  buf u31 (dualtimer2_prdata[0], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(590)
  buf u32 (test_slave_pready, 1'b1);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(895)
  buf u33 (test_slave_pslverr, 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(896)
  buf u34 (test_slave_prdata[0], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(894)
  buf u35 (PENABLE, i_penable);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(901)
  buf u36 (PWRITE, i_pwrite);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(902)
  buf u37 (PADDR[0], i_paddr[0]);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(900)
  or u38 (uart0_overflow_int, uart0_txovrint, uart0_rxovrint);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(905)
  buf u39 (i_uart0_txint, uart0_txint);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(914)
  buf u4 (bigendian, 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(314)
  buf u40 (i_uart0_rxint, uart0_rxint);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(915)
  buf u41 (PWDATA[0], i_pwdata[0]);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(903)
  buf u42 (i_timer1_int, timer1_int);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(927)
  buf u43 (i_dualtimer2_int, dualtimer2_comb_int);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(928)
  buf u44 (i_uart0_overflow_int, uart0_overflow_int);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(929)
  buf u45 (i_watchdog_int, watchdog_int);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(936)
  buf u46 (i_watchdog_rst, watchdog_rst);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(937)
  buf u47 (i_gpio0_intr[0], gpio0_intr[0]);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(926)
  buf u48 (watchdog_interrupt, i_watchdog_int);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(1066)
  buf u49 (watchdog_reset, i_watchdog_rst);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(1067)
  and u5 (n0, HSEL, HTRANS[1]);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(318)
  buf u50 (apbsubsys_interrupt[12], i_gpio0_intr[2]);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(1064)
  buf u51 (apbsubsys_interrupt[13], i_gpio0_intr[3]);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(1064)
  buf u52 (apbsubsys_interrupt[14], i_gpio0_intr[4]);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(1064)
  buf u53 (apbsubsys_interrupt[15], i_gpio0_intr[5]);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(1064)
  buf u54 (apbsubsys_interrupt[16], i_gpio0_intr[6]);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(1064)
  buf u55 (apbsubsys_interrupt[17], i_gpio0_intr[7]);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(1064)
  buf u56 (apbsubsys_interrupt[18], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(1064)
  buf u57 (apbsubsys_interrupt[19], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(1064)
  buf u58 (apbsubsys_interrupt[20], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(1064)
  buf u59 (apbsubsys_interrupt[21], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(1064)
  and u6 (n1, n0, HREADY);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(318)
  buf u60 (apbsubsys_interrupt[22], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(1064)
  buf u61 (apbsubsys_interrupt[23], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(1064)
  buf u62 (apbsubsys_interrupt[24], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(1064)
  buf u63 (apbsubsys_interrupt[25], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(1064)
  buf u64 (apbsubsys_interrupt[26], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(1064)
  buf u65 (apbsubsys_interrupt[27], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(1064)
  buf u66 (apbsubsys_interrupt[28], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(1064)
  buf u67 (apbsubsys_interrupt[29], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(1064)
  buf u68 (apbsubsys_interrupt[30], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(1064)
  buf u69 (apbsubsys_interrupt[31], 1'b0);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(1064)
  and u7 (reg_be_swap_ctrl_en, n1, bigendian);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(318)
  buf u70 (i_gpio0_intr[1], gpio0_intr[1]);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(926)
  buf u71 (i_gpio0_intr[2], gpio0_intr[2]);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(926)
  buf u72 (i_gpio0_intr[3], gpio0_intr[3]);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(926)
  buf u73 (i_gpio0_intr[4], gpio0_intr[4]);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(926)
  buf u74 (i_gpio0_intr[5], gpio0_intr[5]);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(926)
  buf u75 (i_gpio0_intr[6], gpio0_intr[6]);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(926)
  buf u76 (i_gpio0_intr[7], gpio0_intr[7]);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(926)
  buf u77 (PWDATA[1], i_pwdata[1]);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(903)
  buf u78 (PWDATA[2], i_pwdata[2]);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(903)
  buf u79 (PWDATA[3], i_pwdata[3]);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(903)
  buf u8 (apbsubsys_interrupt[10], i_gpio0_intr[0]);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(1064)
  buf u80 (PWDATA[4], i_pwdata[4]);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(903)
  buf u81 (PWDATA[5], i_pwdata[5]);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(903)
  buf u82 (PWDATA[6], i_pwdata[6]);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(903)
  buf u83 (PWDATA[7], i_pwdata[7]);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(903)
  buf u84 (PWDATA[8], i_pwdata[8]);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(903)
  buf u85 (PWDATA[9], i_pwdata[9]);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(903)
  buf u86 (PWDATA[10], i_pwdata[10]);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(903)
  buf u87 (PWDATA[11], i_pwdata[11]);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(903)
  buf u88 (PWDATA[12], i_pwdata[12]);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(903)
  buf u89 (PWDATA[13], i_pwdata[13]);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(903)
  buf u9 (apbsubsys_interrupt[11], i_gpio0_intr[1]);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(1064)
  buf u90 (PWDATA[14], i_pwdata[14]);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(903)
  buf u91 (PWDATA[15], i_pwdata[15]);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(903)
  buf u92 (PWDATA[16], i_pwdata[16]);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(903)
  buf u93 (PWDATA[17], i_pwdata[17]);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(903)
  buf u94 (PWDATA[18], i_pwdata[18]);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(903)
  buf u95 (PWDATA[19], i_pwdata[19]);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(903)
  buf u96 (PWDATA[20], i_pwdata[20]);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(903)
  buf u97 (PWDATA[21], i_pwdata[21]);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(903)
  buf u98 (PWDATA[22], i_pwdata[22]);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(903)
  buf u99 (PWDATA[23], i_pwdata[23]);  // ../RTL/cmsdk_apb_subsystem_m0ds.v(903)
  cmsdk_ahb_to_apb u_ahb_to_apb (
    .HADDR(HADDR),
    .HCLK(HCLK),
    .HPROT(HPROT),
    .HREADY(HREADY),
    .HRESETn(HRESETn),
    .HSEL(HSEL),
    .HSIZE(HSIZE),
    .HTRANS(HTRANS),
    .HWDATA(hwdata_le),
    .HWRITE(HWRITE),
    .PCLKEN(PCLKEN),
    .PRDATA(i_prdata_mux),
    .PREADY(i_pready_mux),
    .PSLVERR(i_pslverr_mux),
    .APBACTIVE(APBACTIVE),
    .HRDATA(hrdata_le),
    .HREADYOUT(HREADYOUT),
    .HRESP(HRESP),
    .PADDR(i_paddr),
    .PENABLE(i_penable),
    .PSEL(i_psel),
    .PWDATA(i_pwdata),
    .PWRITE(i_pwrite));  // ../RTL/cmsdk_apb_subsystem_m0ds.v(356)
  \cmsdk_apb_slave_mux(PORT1_ENABLE=0,PORT2_ENABLE=0,PORT3_ENABLE=0,PORT5_ENABLE=0,PORT6_ENABLE=0,PORT7_ENABLE=0,PORT8_ENABLE=0,PORT9_ENABLE=0,PORT10_ENABLE=0,PORT11_ENABLE=0,PORT12_ENABLE=0,PORT13_ENABLE=0,PORT14_ENABLE=0,PORT15_ENABLE=0)  u_apb_slave_mux (
    .DECODE4BIT(i_paddr[15:12]),
    .PRDATA0(gpio0_prdata),
    .PRDATA1(timer1_prdata),
    .PRDATA10(32'b00000000000000000000000000000000),
    .PRDATA11(test_slave_prdata),
    .PRDATA12(ext12_prdata),
    .PRDATA13(ext13_prdata),
    .PRDATA14(ext14_prdata),
    .PRDATA15(ext15_prdata),
    .PRDATA2(dualtimer2_prdata),
    .PRDATA3(32'b00000000000000000000000000000000),
    .PRDATA4(uart0_prdata),
    .PREADY0(gpio0_pready),
    .PREADY1(timer1_pready),
    .PREADY10(1'b1),
    .PREADY11(test_slave_pready),
    .PREADY12(ext12_pready),
    .PREADY13(ext13_pready),
    .PREADY14(ext14_pready),
    .PREADY15(ext15_pready),
    .PREADY2(dualtimer2_pready),
    .PREADY3(1'b1),
    .PREADY4(uart0_pready),
    .PSEL(i_psel),
    .PSLVERR0(gpio0_pslverr),
    .PSLVERR1(timer1_pslverr),
    .PSLVERR10(1'b0),
    .PSLVERR11(test_slave_pslverr),
    .PSLVERR12(ext12_pslverr),
    .PSLVERR13(ext13_pslverr),
    .PSLVERR14(ext14_pslverr),
    .PSLVERR15(ext15_pslverr),
    .PSLVERR2(dualtimer2_pslverr),
    .PSLVERR3(1'b0),
    .PSLVERR4(uart0_pslverr),
    .PRDATA(i_prdata_mux),
    .PREADY(i_pready_mux),
    .PSEL0(gpio0_psel),
    .PSEL12(ext12_psel),
    .PSEL13(ext13_psel),
    .PSEL14(ext14_psel),
    .PSEL15(ext15_psel),
    .PSEL4(uart0_psel),
    .PSLVERR(i_pslverr_mux));  // ../RTL/cmsdk_apb_subsystem_m0ds.v(409)

endmodule 

module cmsdk_mcu_stclkctrl  // ../RTL/cmsdk_mcu_stclkctrl.v(26)
  (
  FCLK,
  SYSRESETn,
  STCALIB,
  STCLKEN
  );

  input FCLK;  // ../RTL/cmsdk_mcu_stclkctrl.v(34)
  input SYSRESETn;  // ../RTL/cmsdk_mcu_stclkctrl.v(35)
  output [25:0] STCALIB;  // ../RTL/cmsdk_mcu_stclkctrl.v(38)
  output STCLKEN;  // ../RTL/cmsdk_mcu_stclkctrl.v(37)

  parameter DIVIDER_RELOAD = 32'b00000000000000000000000111110011;
  parameter DIV_RATIO = 18'b000000001111101000;
  wire [17:0] n16;
  wire [17:0] reg_clk_div_min1;  // ../RTL/cmsdk_mcu_stclkctrl.v(49)
  wire [17:0] reg_clk_divider;  // ../RTL/cmsdk_mcu_stclkctrl.v(41)
  wire n0;
  wire n1;
  wire n10;
  wire n11;
  wire n12;
  wire n13;
  wire n14;
  wire n15;
  wire n17;
  wire n18;
  wire n19;
  wire n2;
  wire n20;
  wire n21;
  wire n3;
  wire n4;
  wire n5;
  wire n6;
  wire n7;
  wire n8;
  wire n9;
  wire reg_stclken;  // ../RTL/cmsdk_mcu_stclkctrl.v(42)

  eq_w18 eq0 (
    .i0(reg_clk_divider),
    .i1(18'b000000000000000000),
    .o(n19));  // ../RTL/cmsdk_mcu_stclkctrl.v(70)
  binary_mux_s1_w18 mux0 (
    .i0(18'b000000000111110011),
    .i1(reg_clk_div_min1),
    .sel(n15),
    .o(n16));  // ../RTL/cmsdk_mcu_stclkctrl.v(59)
  reg_ar_as_w18 reg0 (
    .clk(FCLK),
    .d(n16),
    .reset({n14,n14,n14,n14,n14,n14,n14,n14,n14,n14,n14,n14,n14,n14,n14,n14,n14,n14}),
    .set(18'b000000000000000000),
    .q(reg_clk_divider));  // ../RTL/cmsdk_mcu_stclkctrl.v(60)
  AL_DFF reg_stclken_reg (
    .clk(FCLK),
    .d(n21),
    .reset(n14),
    .set(1'b0),
    .q(reg_stclken));  // ../RTL/cmsdk_mcu_stclkctrl.v(72)
  add_pu18_mu18_o18 sub0 (
    .i0(reg_clk_divider),
    .i1(18'b000000000000000001),
    .o(reg_clk_div_min1));  // ../RTL/cmsdk_mcu_stclkctrl.v(49)
  buf u10 (STCALIB[0], 1'b0);  // ../RTL/cmsdk_mcu_stclkctrl.v(44)
  not u11 (n20, reg_stclken);  // ../RTL/cmsdk_mcu_stclkctrl.v(71)
  AL_MUX u12 (
    .i0(reg_stclken),
    .i1(n20),
    .sel(n19),
    .o(n21));  // ../RTL/cmsdk_mcu_stclkctrl.v(71)
  or u13 (n18, reg_clk_divider[0], reg_clk_divider[1]);  // ../RTL/cmsdk_mcu_stclkctrl.v(56)
  buf u14 (STCLKEN, reg_stclken);  // ../RTL/cmsdk_mcu_stclkctrl.v(76)
  buf u15 (STCALIB[8], 1'b0);  // ../RTL/cmsdk_mcu_stclkctrl.v(44)
  buf u16 (STCALIB[9], 1'b0);  // ../RTL/cmsdk_mcu_stclkctrl.v(44)
  buf u17 (STCALIB[10], 1'b0);  // ../RTL/cmsdk_mcu_stclkctrl.v(44)
  buf u18 (STCALIB[11], 1'b0);  // ../RTL/cmsdk_mcu_stclkctrl.v(44)
  buf u19 (STCALIB[12], 1'b0);  // ../RTL/cmsdk_mcu_stclkctrl.v(44)
  buf u2 (STCALIB[4], 1'b0);  // ../RTL/cmsdk_mcu_stclkctrl.v(44)
  buf u20 (STCALIB[13], 1'b0);  // ../RTL/cmsdk_mcu_stclkctrl.v(44)
  buf u21 (STCALIB[14], 1'b0);  // ../RTL/cmsdk_mcu_stclkctrl.v(44)
  buf u22 (STCALIB[15], 1'b0);  // ../RTL/cmsdk_mcu_stclkctrl.v(44)
  buf u23 (STCALIB[16], 1'b0);  // ../RTL/cmsdk_mcu_stclkctrl.v(44)
  buf u24 (STCALIB[17], 1'b0);  // ../RTL/cmsdk_mcu_stclkctrl.v(44)
  buf u25 (STCALIB[18], 1'b0);  // ../RTL/cmsdk_mcu_stclkctrl.v(44)
  buf u26 (STCALIB[19], 1'b0);  // ../RTL/cmsdk_mcu_stclkctrl.v(44)
  buf u27 (STCALIB[20], 1'b0);  // ../RTL/cmsdk_mcu_stclkctrl.v(44)
  buf u28 (STCALIB[21], 1'b0);  // ../RTL/cmsdk_mcu_stclkctrl.v(44)
  buf u29 (STCALIB[22], 1'b0);  // ../RTL/cmsdk_mcu_stclkctrl.v(44)
  buf u3 (STCALIB[3], 1'b0);  // ../RTL/cmsdk_mcu_stclkctrl.v(44)
  buf u30 (STCALIB[23], 1'b0);  // ../RTL/cmsdk_mcu_stclkctrl.v(44)
  buf u31 (STCALIB[24], 1'b1);  // ../RTL/cmsdk_mcu_stclkctrl.v(44)
  buf u32 (STCALIB[25], 1'b0);  // ../RTL/cmsdk_mcu_stclkctrl.v(44)
  or u33 (n17, reg_clk_divider[2], reg_clk_divider[3]);  // ../RTL/cmsdk_mcu_stclkctrl.v(56)
  or u34 (n13, n18, n17);  // ../RTL/cmsdk_mcu_stclkctrl.v(56)
  or u35 (n1, reg_clk_divider[4], reg_clk_divider[5]);  // ../RTL/cmsdk_mcu_stclkctrl.v(56)
  or u36 (n0, reg_clk_divider[7], reg_clk_divider[8]);  // ../RTL/cmsdk_mcu_stclkctrl.v(56)
  or u37 (n2, reg_clk_divider[6], n0);  // ../RTL/cmsdk_mcu_stclkctrl.v(56)
  or u38 (n3, n1, n2);  // ../RTL/cmsdk_mcu_stclkctrl.v(56)
  or u39 (n4, n13, n3);  // ../RTL/cmsdk_mcu_stclkctrl.v(56)
  buf u4 (STCALIB[5], 1'b0);  // ../RTL/cmsdk_mcu_stclkctrl.v(44)
  or u40 (n5, reg_clk_divider[9], reg_clk_divider[10]);  // ../RTL/cmsdk_mcu_stclkctrl.v(56)
  or u41 (n6, reg_clk_divider[11], reg_clk_divider[12]);  // ../RTL/cmsdk_mcu_stclkctrl.v(56)
  or u42 (n7, n5, n6);  // ../RTL/cmsdk_mcu_stclkctrl.v(56)
  or u43 (n8, reg_clk_divider[13], reg_clk_divider[14]);  // ../RTL/cmsdk_mcu_stclkctrl.v(56)
  or u44 (n9, reg_clk_divider[16], reg_clk_divider[17]);  // ../RTL/cmsdk_mcu_stclkctrl.v(56)
  or u45 (n10, reg_clk_divider[15], n9);  // ../RTL/cmsdk_mcu_stclkctrl.v(56)
  or u46 (n11, n8, n10);  // ../RTL/cmsdk_mcu_stclkctrl.v(56)
  or u47 (n12, n7, n11);  // ../RTL/cmsdk_mcu_stclkctrl.v(56)
  or u48 (n15, n4, n12);  // ../RTL/cmsdk_mcu_stclkctrl.v(56)
  buf u5 (STCALIB[6], 1'b0);  // ../RTL/cmsdk_mcu_stclkctrl.v(44)
  buf u6 (STCALIB[7], 1'b0);  // ../RTL/cmsdk_mcu_stclkctrl.v(44)
  buf u7 (STCALIB[2], 1'b0);  // ../RTL/cmsdk_mcu_stclkctrl.v(44)
  not u8 (n14, SYSRESETn);  // ../RTL/cmsdk_mcu_stclkctrl.v(52)
  buf u9 (STCALIB[1], 1'b0);  // ../RTL/cmsdk_mcu_stclkctrl.v(44)

endmodule 

module cmsdk_mcu_sysctrl  // ../RTL/cmsdk_mcu_sysctrl.v(44)
  (
  ECOREVNUM,
  FCLK,
  HADDR,
  HCLK,
  HREADY,
  HRESETn,
  HSEL,
  HSIZE,
  HTRANS,
  HWDATA,
  HWRITE,
  LOCKUP,
  PORESETn,
  SYSRESETREQ,
  WDOGRESETREQ,
  HRDATA,
  HREADYOUT,
  HRESP,
  LOCKUPRESET,
  PMUENABLE,
  REMAP
  );

  input [3:0] ECOREVNUM;  // ../RTL/cmsdk_mcu_sysctrl.v(70)
  input FCLK;  // ../RTL/cmsdk_mcu_sysctrl.v(53)
  input [11:0] HADDR;  // ../RTL/cmsdk_mcu_sysctrl.v(60)
  input HCLK;  // ../RTL/cmsdk_mcu_sysctrl.v(51)
  input HREADY;  // ../RTL/cmsdk_mcu_sysctrl.v(56)
  input HRESETn;  // ../RTL/cmsdk_mcu_sysctrl.v(52)
  input HSEL;  // ../RTL/cmsdk_mcu_sysctrl.v(55)
  input [2:0] HSIZE;  // ../RTL/cmsdk_mcu_sysctrl.v(58)
  input [1:0] HTRANS;  // ../RTL/cmsdk_mcu_sysctrl.v(57)
  input [31:0] HWDATA;  // ../RTL/cmsdk_mcu_sysctrl.v(61)
  input HWRITE;  // ../RTL/cmsdk_mcu_sysctrl.v(59)
  input LOCKUP;  // ../RTL/cmsdk_mcu_sysctrl.v(68)
  input PORESETn;  // ../RTL/cmsdk_mcu_sysctrl.v(54)
  input SYSRESETREQ;  // ../RTL/cmsdk_mcu_sysctrl.v(66)
  input WDOGRESETREQ;  // ../RTL/cmsdk_mcu_sysctrl.v(67)
  output [31:0] HRDATA;  // ../RTL/cmsdk_mcu_sysctrl.v(64)
  output HREADYOUT;  // ../RTL/cmsdk_mcu_sysctrl.v(62)
  output HRESP;  // ../RTL/cmsdk_mcu_sysctrl.v(63)
  output LOCKUPRESET;  // ../RTL/cmsdk_mcu_sysctrl.v(74)
  output PMUENABLE;  // ../RTL/cmsdk_mcu_sysctrl.v(73)
  output REMAP;  // ../RTL/cmsdk_mcu_sysctrl.v(72)

  parameter BE = 0;
  // localparam ARM_CMSDK_CM0_SYSCTRL_CID0 = 32'b00000000000000000000000000001101;
  // localparam ARM_CMSDK_CM0_SYSCTRL_CID1 = 32'b00000000000000000000000011110000;
  // localparam ARM_CMSDK_CM0_SYSCTRL_CID2 = 32'b00000000000000000000000000000101;
  // localparam ARM_CMSDK_CM0_SYSCTRL_CID3 = 32'b00000000000000000000000010110001;
  // localparam ARM_CMSDK_CM0_SYSCTRL_PID0 = 32'b00000000000000000000000000100110;
  // localparam ARM_CMSDK_CM0_SYSCTRL_PID1 = 32'b00000000000000000000000010111000;
  // localparam ARM_CMSDK_CM0_SYSCTRL_PID2 = 32'b00000000000000000000000000011011;
  // localparam ARM_CMSDK_CM0_SYSCTRL_PID3 = 32'b00000000000000000000000000000000;
  // localparam ARM_CMSDK_CM0_SYSCTRL_PID4 = 32'b00000000000000000000000000000100;
  // localparam ARM_CMSDK_CM0_SYSCTRL_PID5 = 32'b00000000000000000000000000000000;
  // localparam ARM_CMSDK_CM0_SYSCTRL_PID6 = 32'b00000000000000000000000000000000;
  // localparam ARM_CMSDK_CM0_SYSCTRL_PID7 = 32'b00000000000000000000000000000000;
  wire [31:0] HWDATALE;  // ../RTL/cmsdk_mcu_sysctrl.v(125)
  wire [3:0] n10;
  wire [9:0] n14;
  wire [1:0] n15;
  wire [31:0] n17;
  wire [31:0] n19;
  wire [31:0] n20;
  wire [31:0] n21;
  wire [31:0] n26;
  wire [31:0] n27;
  wire [2:0] n36;
  wire [2:0] n37;
  wire [2:0] n38;
  wire [3:0] n4;
  wire [2:0] n43;
  wire [3:0] n5;
  wire [3:0] n6;
  wire [3:0] nxt_byte_strobe;  // ../RTL/cmsdk_mcu_sysctrl.v(119)
  wire [2:0] nxt_resetinfo;  // ../RTL/cmsdk_mcu_sysctrl.v(302)
  wire [31:0] read_mux;  // ../RTL/cmsdk_mcu_sysctrl.v(100)
  wire [31:0] read_mux_le;  // ../RTL/cmsdk_mcu_sysctrl.v(101)
  wire [11:2] reg_addr;  // ../RTL/cmsdk_mcu_sysctrl.v(123)
  wire [3:0] reg_byte_strobe;  // ../RTL/cmsdk_mcu_sysctrl.v(120)
  wire [1:0] reg_hsize;  // ../RTL/cmsdk_mcu_sysctrl.v(124)
  wire [2:0] reg_resetinfo;  // ../RTL/cmsdk_mcu_sysctrl.v(109)
  wire ahb_access;  // ../RTL/cmsdk_mcu_sysctrl.v(116)
  wire ahb_read;  // ../RTL/cmsdk_mcu_sysctrl.v(118)
  wire ahb_write;  // ../RTL/cmsdk_mcu_sysctrl.v(117)
  wire bigendian;  // ../RTL/cmsdk_mcu_sysctrl.v(115)
  wire n0;
  wire n1;
  wire n11;
  wire n12;
  wire n13;
  wire n16;
  wire n18;
  wire n2;
  wire n22;
  wire n23;
  wire n24;
  wire n25;
  wire n28;
  wire n29;
  wire n3;
  wire n30;
  wire n31;
  wire n32;
  wire n33;
  wire n34;
  wire n35;
  wire n39;
  wire n40;
  wire n41;
  wire n42;
  wire n7;
  wire n8;
  wire n9;
  wire reg_lockupreset;  // ../RTL/cmsdk_mcu_sysctrl.v(108)
  wire reg_lockupreset_write;  // ../RTL/cmsdk_mcu_sysctrl.v(280)
  wire reg_pmuenable;  // ../RTL/cmsdk_mcu_sysctrl.v(104)
  wire reg_read_enable;  // ../RTL/cmsdk_mcu_sysctrl.v(121)
  wire reg_remap;  // ../RTL/cmsdk_mcu_sysctrl.v(102)
  wire reg_remap_write;  // ../RTL/cmsdk_mcu_sysctrl.v(240)
  wire reg_resetinfo_en;  // ../RTL/cmsdk_mcu_sysctrl.v(309)
  wire reg_resetinfo_write;  // ../RTL/cmsdk_mcu_sysctrl.v(297)
  wire reg_write_enable;  // ../RTL/cmsdk_mcu_sysctrl.v(122)

  eq_w2 eq0 (
    .i0(HADDR[1:0]),
    .i1(2'b00),
    .o(n3));  // ../RTL/cmsdk_mcu_sysctrl.v(128)
  eq_w2 eq1 (
    .i0(HADDR[1:0]),
    .i1(2'b01),
    .o(n7));  // ../RTL/cmsdk_mcu_sysctrl.v(129)
  eq_w10 eq10 (
    .i0(reg_addr),
    .i1(10'b0000000100),
    .o(n34));  // ../RTL/cmsdk_mcu_sysctrl.v(299)
  eq_w2 eq2 (
    .i0(HADDR[1:0]),
    .i1(2'b10),
    .o(n8));  // ../RTL/cmsdk_mcu_sysctrl.v(130)
  eq_w2 eq3 (
    .i0(HADDR[1:0]),
    .i1(2'b11),
    .o(n9));  // ../RTL/cmsdk_mcu_sysctrl.v(131)
  eq_w7 eq4 (
    .i0(reg_addr[11:5]),
    .i1(7'b0000000),
    .o(n16));  // ../RTL/cmsdk_mcu_sysctrl.v(175)
  eq_w6 eq5 (
    .i0(reg_addr[11:6]),
    .i1(6'b111111),
    .o(n18));  // ../RTL/cmsdk_mcu_sysctrl.v(185)
  eq_w2 eq6 (
    .i0(reg_hsize),
    .i1(2'b10),
    .o(n22));  // ../RTL/cmsdk_mcu_sysctrl.v(219)
  eq_w2 eq7 (
    .i0(reg_hsize),
    .i1(2'b01),
    .o(n24));  // ../RTL/cmsdk_mcu_sysctrl.v(225)
  eq_w10 eq8 (
    .i0(reg_addr),
    .i1(10'b0000000000),
    .o(n28));  // ../RTL/cmsdk_mcu_sysctrl.v(242)
  eq_w10 eq9 (
    .i0(reg_addr),
    .i1(10'b0000000010),
    .o(n31));  // ../RTL/cmsdk_mcu_sysctrl.v(282)
  binary_mux_s1_w4 mux0 (
    .i0(reg_byte_strobe),
    .i1(nxt_byte_strobe),
    .sel(HREADY),
    .o(n10));  // ../RTL/cmsdk_mcu_sysctrl.v(147)
  binary_mux_s1_w10 mux1 (
    .i0(reg_addr),
    .i1(HADDR[11:2]),
    .sel(ahb_access),
    .o(n14));  // ../RTL/cmsdk_mcu_sysctrl.v(156)
  binary_mux_s1_w32 mux10 (
    .i0(n26),
    .i1({read_mux_le[7:0],read_mux_le[15:8],read_mux_le[23:16],read_mux_le[31:24]}),
    .sel(n23),
    .o(read_mux));  // ../RTL/cmsdk_mcu_sysctrl.v(235)
  binary_mux_s1_w32 mux11 (
    .i0(n27),
    .i1({HWDATA[7:0],HWDATA[15:8],HWDATA[23:16],HWDATA[31:24]}),
    .sel(n23),
    .o({open_n0,open_n1,open_n2,open_n3,open_n4,open_n5,open_n6,open_n7,open_n8,open_n9,open_n10,open_n11,open_n12,open_n13,open_n14,open_n15,open_n16,open_n17,open_n18,open_n19,open_n20,open_n21,open_n22,open_n23,open_n24,open_n25,open_n26,open_n27,open_n28,HWDATALE[2:0]}));  // ../RTL/cmsdk_mcu_sysctrl.v(235)
  binary_mux_s1_w3 mux12 (
    .i0(reg_resetinfo),
    .i1(nxt_resetinfo),
    .sel(reg_resetinfo_en),
    .o(n43));  // ../RTL/cmsdk_mcu_sysctrl.v(318)
  binary_mux_s1_w2 mux2 (
    .i0(reg_hsize),
    .i1(HSIZE[1:0]),
    .sel(ahb_access),
    .o(n15));  // ../RTL/cmsdk_mcu_sysctrl.v(165)
  binary_mux_s3_w32 mux3 (
    .i0({31'b0000000000000000000000000000000,reg_remap}),
    .i1({31'b0000000000000000000000000000000,reg_pmuenable}),
    .i2({31'b0000000000000000000000000000000,reg_lockupreset}),
    .i3(32'b00000000000000000000000000000000),
    .i4({29'b00000000000000000000000000000,reg_resetinfo}),
    .i5(32'b00000000000000000000000000000000),
    .i6(32'b00000000000000000000000000000000),
    .i7(32'b00000000000000000000000000000000),
    .sel(reg_addr[4:2]),
    .o(n17));  // ../RTL/cmsdk_mcu_sysctrl.v(183)
  binary_mux_s4_w32 mux4 (
    .i0(32'b00000000000000000000000000000000),
    .i1(32'b00000000000000000000000000000000),
    .i10(32'b00000000000000000000000000011011),
    .i11({24'b000000000000000000000000,ECOREVNUM,4'b0000}),
    .i12(32'b00000000000000000000000000001101),
    .i13(32'b00000000000000000000000011110000),
    .i14(32'b00000000000000000000000000000101),
    .i15(32'b00000000000000000000000010110001),
    .i2(32'b00000000000000000000000000000000),
    .i3(32'b00000000000000000000000000000000),
    .i4(32'b00000000000000000000000000000100),
    .i5(32'b00000000000000000000000000000000),
    .i6(32'b00000000000000000000000000000000),
    .i7(32'b00000000000000000000000000000000),
    .i8(32'b00000000000000000000000000100110),
    .i9(32'b00000000000000000000000010111000),
    .sel(reg_addr[5:2]),
    .o(n19));  // ../RTL/cmsdk_mcu_sysctrl.v(201)
  binary_mux_s1_w32 mux5 (
    .i0(32'b00000000000000000000000000000000),
    .i1(n19),
    .sel(n18),
    .o(n20));  // ../RTL/cmsdk_mcu_sysctrl.v(205)
  binary_mux_s1_w32 mux6 (
    .i0(n20),
    .i1(n17),
    .sel(n16),
    .o(n21));  // ../RTL/cmsdk_mcu_sysctrl.v(205)
  binary_mux_s1_w32 mux7 (
    .i0(32'b00000000000000000000000000000000),
    .i1(n21),
    .sel(reg_read_enable),
    .o(read_mux_le));  // ../RTL/cmsdk_mcu_sysctrl.v(213)
  binary_mux_s1_w32 mux8 (
    .i0(read_mux_le),
    .i1({read_mux_le[23:16],read_mux_le[31:24],read_mux_le[7:0],read_mux_le[15:8]}),
    .sel(n25),
    .o(n26));  // ../RTL/cmsdk_mcu_sysctrl.v(235)
  binary_mux_s1_w32 mux9 (
    .i0(HWDATA),
    .i1({HWDATA[23:16],HWDATA[31:24],HWDATA[7:0],HWDATA[15:8]}),
    .sel(n25),
    .o(n27));  // ../RTL/cmsdk_mcu_sysctrl.v(235)
  reg_ar_as_w10 reg0 (
    .clk(HCLK),
    .d(n14),
    .reset({n13,n13,n13,n13,n13,n13,n13,n13,n13,n13}),
    .set(10'b0000000000),
    .q(reg_addr));  // ../RTL/cmsdk_mcu_sysctrl.v(156)
  reg_ar_as_w2 reg1 (
    .clk(HCLK),
    .d(n15),
    .reset({n13,n13}),
    .set(2'b00),
    .q(reg_hsize));  // ../RTL/cmsdk_mcu_sysctrl.v(165)
  reg_ar_as_w3 reg2 (
    .clk(FCLK),
    .d(n43),
    .reset({n42,n42,n42}),
    .set(3'b000),
    .q(reg_resetinfo));  // ../RTL/cmsdk_mcu_sysctrl.v(318)
  reg_ar_as_w4 reg3 (
    .clk(HCLK),
    .d(n10),
    .reset({n13,n13,n13,n13}),
    .set(4'b0000),
    .q(reg_byte_strobe));  // ../RTL/cmsdk_mcu_sysctrl.v(147)
  AL_DFF reg_lockupreset_reg (
    .clk(HCLK),
    .d(n33),
    .reset(n13),
    .set(1'b0),
    .q(reg_lockupreset));  // ../RTL/cmsdk_mcu_sysctrl.v(290)
  AL_DFF reg_read_enable_reg (
    .clk(HCLK),
    .d(n11),
    .reset(n13),
    .set(1'b0),
    .q(reg_read_enable));  // ../RTL/cmsdk_mcu_sysctrl.v(147)
  AL_DFF reg_remap_reg (
    .clk(HCLK),
    .d(n30),
    .reset(1'b0),
    .set(n13),
    .q(reg_remap));  // ../RTL/cmsdk_mcu_sysctrl.v(250)
  AL_DFF reg_write_enable_reg (
    .clk(HCLK),
    .d(n12),
    .reset(n13),
    .set(1'b0),
    .q(reg_write_enable));  // ../RTL/cmsdk_mcu_sysctrl.v(147)
  not u10 (n2, HADDR[1]);  // ../RTL/cmsdk_mcu_sysctrl.v(128)
  buf u11 (HRDATA[28], read_mux[28]);  // ../RTL/cmsdk_mcu_sysctrl.v(327)
  buf u12 (HRDATA[31], read_mux[31]);  // ../RTL/cmsdk_mcu_sysctrl.v(327)
  and u13 (nxt_byte_strobe[3], n4[3], ahb_access);  // ../RTL/cmsdk_mcu_sysctrl.v(131)
  and u14 (n38[1], n37[1], reg_resetinfo[1]);  // ../RTL/cmsdk_mcu_sysctrl.v(306)
  buf u15 (HRDATA[6], read_mux[6]);  // ../RTL/cmsdk_mcu_sysctrl.v(327)
  buf u16 (HRDATA[27], read_mux[27]);  // ../RTL/cmsdk_mcu_sysctrl.v(327)
  buf u17 (HRDATA[30], read_mux[30]);  // ../RTL/cmsdk_mcu_sysctrl.v(327)
  and u18 (nxt_byte_strobe[2], n4[2], ahb_access);  // ../RTL/cmsdk_mcu_sysctrl.v(131)
  and u19 (n5[3], HADDR[1], HSIZE[0]);  // ../RTL/cmsdk_mcu_sysctrl.v(131)
  buf u2 (HRDATA[16], read_mux[16]);  // ../RTL/cmsdk_mcu_sysctrl.v(327)
  buf u20 (HRDATA[14], read_mux[14]);  // ../RTL/cmsdk_mcu_sysctrl.v(327)
  buf u21 (HRDATA[26], read_mux[26]);  // ../RTL/cmsdk_mcu_sysctrl.v(327)
  buf u22 (HRDATA[29], read_mux[29]);  // ../RTL/cmsdk_mcu_sysctrl.v(327)
  and u23 (nxt_byte_strobe[1], n4[1], ahb_access);  // ../RTL/cmsdk_mcu_sysctrl.v(131)
  or u24 (n6[3], HSIZE[1], n5[3]);  // ../RTL/cmsdk_mcu_sysctrl.v(131)
  buf u25 (HRDATA[13], read_mux[13]);  // ../RTL/cmsdk_mcu_sysctrl.v(327)
  buf u26 (HRDATA[0], read_mux[0]);  // ../RTL/cmsdk_mcu_sysctrl.v(327)
  buf u27 (HRDATA[7], read_mux[7]);  // ../RTL/cmsdk_mcu_sysctrl.v(327)
  or u28 (nxt_resetinfo[0], n38[0], SYSRESETREQ);  // ../RTL/cmsdk_mcu_sysctrl.v(306)
  buf u29 (HRDATA[12], read_mux[12]);  // ../RTL/cmsdk_mcu_sysctrl.v(327)
  buf u3 (HRDATA[15], read_mux[15]);  // ../RTL/cmsdk_mcu_sysctrl.v(327)
  not u30 (n13, HRESETn);  // ../RTL/cmsdk_mcu_sysctrl.v(136)
  AL_MUX u31 (
    .i0(reg_read_enable),
    .i1(ahb_read),
    .sel(HREADY),
    .o(n11));  // ../RTL/cmsdk_mcu_sysctrl.v(147)
  AL_MUX u32 (
    .i0(reg_write_enable),
    .i1(ahb_write),
    .sel(HREADY),
    .o(n12));  // ../RTL/cmsdk_mcu_sysctrl.v(147)
  buf u33 (HRDATA[11], read_mux[11]);  // ../RTL/cmsdk_mcu_sysctrl.v(327)
  buf u34 (HRDATA[5], read_mux[5]);  // ../RTL/cmsdk_mcu_sysctrl.v(327)
  buf u35 (HRDATA[10], read_mux[10]);  // ../RTL/cmsdk_mcu_sysctrl.v(327)
  buf u36 (HRDATA[4], read_mux[4]);  // ../RTL/cmsdk_mcu_sysctrl.v(327)
  buf u37 (HRDATA[3], read_mux[3]);  // ../RTL/cmsdk_mcu_sysctrl.v(327)
  and u38 (n23, bigendian, n22);  // ../RTL/cmsdk_mcu_sysctrl.v(219)
  and u39 (n25, bigendian, n24);  // ../RTL/cmsdk_mcu_sysctrl.v(225)
  buf u4 (bigendian, 1'b0);  // ../RTL/cmsdk_mcu_sysctrl.v(115)
  and u40 (n29, reg_write_enable, n28);  // ../RTL/cmsdk_mcu_sysctrl.v(242)
  and u41 (reg_remap_write, n29, reg_byte_strobe[0]);  // ../RTL/cmsdk_mcu_sysctrl.v(242)
  buf u42 (HRDATA[9], read_mux[9]);  // ../RTL/cmsdk_mcu_sysctrl.v(327)
  buf u43 (HRDATA[2], read_mux[2]);  // ../RTL/cmsdk_mcu_sysctrl.v(327)
  AL_MUX u44 (
    .i0(reg_remap),
    .i1(HWDATALE[0]),
    .sel(reg_remap_write),
    .o(n30));  // ../RTL/cmsdk_mcu_sysctrl.v(250)
  buf u45 (reg_pmuenable, 1'b0);  // ../RTL/cmsdk_mcu_sysctrl.v(260)
  and u46 (n32, reg_write_enable, n31);  // ../RTL/cmsdk_mcu_sysctrl.v(282)
  and u47 (reg_lockupreset_write, n32, reg_byte_strobe[0]);  // ../RTL/cmsdk_mcu_sysctrl.v(282)
  buf u48 (HRDATA[8], read_mux[8]);  // ../RTL/cmsdk_mcu_sysctrl.v(327)
  buf u49 (HRDATA[1], read_mux[1]);  // ../RTL/cmsdk_mcu_sysctrl.v(327)
  and u5 (n0, HTRANS[1], HSEL);  // ../RTL/cmsdk_mcu_sysctrl.v(116)
  AL_MUX u50 (
    .i0(reg_lockupreset),
    .i1(HWDATALE[0]),
    .sel(reg_lockupreset_write),
    .o(n33));  // ../RTL/cmsdk_mcu_sysctrl.v(290)
  and u51 (n35, reg_write_enable, n34);  // ../RTL/cmsdk_mcu_sysctrl.v(299)
  and u52 (reg_resetinfo_write, n35, reg_byte_strobe[0]);  // ../RTL/cmsdk_mcu_sysctrl.v(299)
  buf u53 (HRDATA[19], read_mux[19]);  // ../RTL/cmsdk_mcu_sysctrl.v(327)
  buf u54 (HRDATA[21], read_mux[21]);  // ../RTL/cmsdk_mcu_sysctrl.v(327)
  buf u55 (HRDATA[23], read_mux[23]);  // ../RTL/cmsdk_mcu_sysctrl.v(327)
  buf u56 (HRDATA[25], read_mux[25]);  // ../RTL/cmsdk_mcu_sysctrl.v(327)
  buf u57 (HRDATA[18], read_mux[18]);  // ../RTL/cmsdk_mcu_sysctrl.v(327)
  buf u58 (HRDATA[20], read_mux[20]);  // ../RTL/cmsdk_mcu_sysctrl.v(327)
  buf u59 (HRDATA[22], read_mux[22]);  // ../RTL/cmsdk_mcu_sysctrl.v(327)
  and u6 (ahb_access, n0, HREADY);  // ../RTL/cmsdk_mcu_sysctrl.v(116)
  buf u60 (HRDATA[24], read_mux[24]);  // ../RTL/cmsdk_mcu_sysctrl.v(327)
  buf u61 (HRDATA[17], read_mux[17]);  // ../RTL/cmsdk_mcu_sysctrl.v(327)
  or u62 (n4[0], n6[1], n3);  // ../RTL/cmsdk_mcu_sysctrl.v(131)
  and u63 (n36[0], reg_resetinfo_write, HWDATALE[0]);  // ../RTL/cmsdk_mcu_sysctrl.v(306)
  and u64 (n39, reg_lockupreset, LOCKUP);  // ../RTL/cmsdk_mcu_sysctrl.v(306)
  not u65 (n37[0], n36[0]);  // ../RTL/cmsdk_mcu_sysctrl.v(306)
  or u66 (n40, reg_resetinfo_write, SYSRESETREQ);  // ../RTL/cmsdk_mcu_sysctrl.v(310)
  or u67 (n41, n40, WDOGRESETREQ);  // ../RTL/cmsdk_mcu_sysctrl.v(310)
  and u68 (n38[0], n37[0], reg_resetinfo[0]);  // ../RTL/cmsdk_mcu_sysctrl.v(306)
  or u69 (reg_resetinfo_en, n41, n39);  // ../RTL/cmsdk_mcu_sysctrl.v(310)
  and u7 (ahb_write, ahb_access, HWRITE);  // ../RTL/cmsdk_mcu_sysctrl.v(117)
  and u70 (n5[1], n2, HSIZE[0]);  // ../RTL/cmsdk_mcu_sysctrl.v(131)
  not u71 (n42, PORESETn);  // ../RTL/cmsdk_mcu_sysctrl.v(315)
  or u72 (n6[1], HSIZE[1], n5[1]);  // ../RTL/cmsdk_mcu_sysctrl.v(131)
  buf u73 (REMAP, reg_remap);  // ../RTL/cmsdk_mcu_sysctrl.v(322)
  buf u74 (PMUENABLE, reg_pmuenable);  // ../RTL/cmsdk_mcu_sysctrl.v(323)
  buf u75 (LOCKUPRESET, reg_lockupreset);  // ../RTL/cmsdk_mcu_sysctrl.v(324)
  buf u76 (HREADYOUT, 1'b1);  // ../RTL/cmsdk_mcu_sysctrl.v(326)
  and u77 (nxt_byte_strobe[0], n4[0], ahb_access);  // ../RTL/cmsdk_mcu_sysctrl.v(131)
  buf u78 (HRESP, 1'b0);  // ../RTL/cmsdk_mcu_sysctrl.v(328)
  and u79 (n38[2], n37[2], reg_resetinfo[2]);  // ../RTL/cmsdk_mcu_sysctrl.v(306)
  not u8 (n1, HWRITE);  // ../RTL/cmsdk_mcu_sysctrl.v(118)
  not u80 (n37[1], n36[1]);  // ../RTL/cmsdk_mcu_sysctrl.v(306)
  not u81 (n37[2], n36[2]);  // ../RTL/cmsdk_mcu_sysctrl.v(306)
  and u82 (n36[1], reg_resetinfo_write, HWDATALE[1]);  // ../RTL/cmsdk_mcu_sysctrl.v(306)
  and u83 (n36[2], reg_resetinfo_write, HWDATALE[2]);  // ../RTL/cmsdk_mcu_sysctrl.v(306)
  or u84 (n4[1], n6[1], n7);  // ../RTL/cmsdk_mcu_sysctrl.v(131)
  or u85 (n4[2], n6[3], n8);  // ../RTL/cmsdk_mcu_sysctrl.v(131)
  or u86 (n4[3], n6[3], n9);  // ../RTL/cmsdk_mcu_sysctrl.v(131)
  or u87 (nxt_resetinfo[1], n38[1], WDOGRESETREQ);  // ../RTL/cmsdk_mcu_sysctrl.v(306)
  or u88 (nxt_resetinfo[2], n38[2], n39);  // ../RTL/cmsdk_mcu_sysctrl.v(306)
  and u9 (ahb_read, ahb_access, n1);  // ../RTL/cmsdk_mcu_sysctrl.v(118)

endmodule 

module CORTEXM0INTEGRATION  // ../RTL/CORTEXM0INTEGRATION.v(29)
  (
  CDBGPWRUPACK,
  DBGRESETn,
  DBGRESTART,
  DCLK,
  ECOREVNUM,
  EDBGRQ,
  FCLK,
  HCLK,
  HRDATA,
  HREADY,
  HRESETn,
  HRESP,
  IRQ,
  IRQLATENCY,
  NMI,
  PORESETn,
  RSTBYPASS,
  RXEV,
  SCLK,
  SE,
  SLEEPHOLDREQn,
  STCALIB,
  STCLKEN,
  SWCLKTCK,
  SWDITMS,
  TDI,
  WICENREQ,
  nTRST,
  CDBGPWRUPREQ,
  CODEHINTDE,
  CODENSEQ,
  DBGRESTARTED,
  GATEHCLK,
  HADDR,
  HALTED,
  HBURST,
  HMASTER,
  HMASTLOCK,
  HPROT,
  HSIZE,
  HTRANS,
  HWDATA,
  HWRITE,
  LOCKUP,
  SLEEPDEEP,
  SLEEPHOLDACKn,
  SLEEPING,
  SPECHTRANS,
  SWDO,
  SWDOEN,
  SYSRESETREQ,
  TDO,
  TXEV,
  WAKEUP,
  WICENACK,
  WICSENSE,
  nTDOEN
  );

  input CDBGPWRUPACK;  // ../RTL/CORTEXM0INTEGRATION.v(95)
  input DBGRESETn;  // ../RTL/CORTEXM0INTEGRATION.v(36)
  input DBGRESTART;  // ../RTL/CORTEXM0INTEGRATION.v(67)
  input DCLK;  // ../RTL/CORTEXM0INTEGRATION.v(34)
  input [27:0] ECOREVNUM;  // ../RTL/CORTEXM0INTEGRATION.v(82)
  input EDBGRQ;  // ../RTL/CORTEXM0INTEGRATION.v(69)
  input FCLK;  // ../RTL/CORTEXM0INTEGRATION.v(31)
  input HCLK;  // ../RTL/CORTEXM0INTEGRATION.v(33)
  input [31:0] HRDATA;  // ../RTL/CORTEXM0INTEGRATION.v(50)
  input HREADY;  // ../RTL/CORTEXM0INTEGRATION.v(51)
  input HRESETn;  // ../RTL/CORTEXM0INTEGRATION.v(37)
  input HRESP;  // ../RTL/CORTEXM0INTEGRATION.v(52)
  input [31:0] IRQ;  // ../RTL/CORTEXM0INTEGRATION.v(74)
  input [7:0] IRQLATENCY;  // ../RTL/CORTEXM0INTEGRATION.v(81)
  input NMI;  // ../RTL/CORTEXM0INTEGRATION.v(73)
  input PORESETn;  // ../RTL/CORTEXM0INTEGRATION.v(35)
  input RSTBYPASS;  // ../RTL/CORTEXM0INTEGRATION.v(99)
  input RXEV;  // ../RTL/CORTEXM0INTEGRATION.v(76)
  input SCLK;  // ../RTL/CORTEXM0INTEGRATION.v(32)
  input SE;  // ../RTL/CORTEXM0INTEGRATION.v(98)
  input SLEEPHOLDREQn;  // ../RTL/CORTEXM0INTEGRATION.v(90)
  input [25:0] STCALIB;  // ../RTL/CORTEXM0INTEGRATION.v(79)
  input STCLKEN;  // ../RTL/CORTEXM0INTEGRATION.v(80)
  input SWCLKTCK;  // ../RTL/CORTEXM0INTEGRATION.v(38)
  input SWDITMS;  // ../RTL/CORTEXM0INTEGRATION.v(61)
  input TDI;  // ../RTL/CORTEXM0INTEGRATION.v(62)
  input WICENREQ;  // ../RTL/CORTEXM0INTEGRATION.v(92)
  input nTRST;  // ../RTL/CORTEXM0INTEGRATION.v(39)
  output CDBGPWRUPREQ;  // ../RTL/CORTEXM0INTEGRATION.v(94)
  output [2:0] CODEHINTDE;  // ../RTL/CORTEXM0INTEGRATION.v(57)
  output CODENSEQ;  // ../RTL/CORTEXM0INTEGRATION.v(56)
  output DBGRESTARTED;  // ../RTL/CORTEXM0INTEGRATION.v(68)
  output GATEHCLK;  // ../RTL/CORTEXM0INTEGRATION.v(85)
  output [31:0] HADDR;  // ../RTL/CORTEXM0INTEGRATION.v(42)
  output HALTED;  // ../RTL/CORTEXM0INTEGRATION.v(70)
  output [2:0] HBURST;  // ../RTL/CORTEXM0INTEGRATION.v(43)
  output HMASTER;  // ../RTL/CORTEXM0INTEGRATION.v(53)
  output HMASTLOCK;  // ../RTL/CORTEXM0INTEGRATION.v(44)
  output [3:0] HPROT;  // ../RTL/CORTEXM0INTEGRATION.v(45)
  output [2:0] HSIZE;  // ../RTL/CORTEXM0INTEGRATION.v(46)
  output [1:0] HTRANS;  // ../RTL/CORTEXM0INTEGRATION.v(47)
  output [31:0] HWDATA;  // ../RTL/CORTEXM0INTEGRATION.v(48)
  output HWRITE;  // ../RTL/CORTEXM0INTEGRATION.v(49)
  output LOCKUP;  // ../RTL/CORTEXM0INTEGRATION.v(77)
  output SLEEPDEEP;  // ../RTL/CORTEXM0INTEGRATION.v(87)
  output SLEEPHOLDACKn;  // ../RTL/CORTEXM0INTEGRATION.v(91)
  output SLEEPING;  // ../RTL/CORTEXM0INTEGRATION.v(86)
  output SPECHTRANS;  // ../RTL/CORTEXM0INTEGRATION.v(58)
  output SWDO;  // ../RTL/CORTEXM0INTEGRATION.v(63)
  output SWDOEN;  // ../RTL/CORTEXM0INTEGRATION.v(64)
  output SYSRESETREQ;  // ../RTL/CORTEXM0INTEGRATION.v(78)
  output TDO;  // ../RTL/CORTEXM0INTEGRATION.v(65)
  output TXEV;  // ../RTL/CORTEXM0INTEGRATION.v(75)
  output WAKEUP;  // ../RTL/CORTEXM0INTEGRATION.v(88)
  output WICENACK;  // ../RTL/CORTEXM0INTEGRATION.v(93)
  output [33:0] WICSENSE;  // ../RTL/CORTEXM0INTEGRATION.v(89)
  output nTDOEN;  // ../RTL/CORTEXM0INTEGRATION.v(66)


  cortexm0ds_logic u_logic (
    .CDBGPWRUPACK(CDBGPWRUPACK),
    .DBGRESETn(DBGRESETn),
    .DBGRESTART(DBGRESTART),
    .DCLK(DCLK),
    .ECOREVNUM(ECOREVNUM),
    .EDBGRQ(EDBGRQ),
    .FCLK(FCLK),
    .HCLK(HCLK),
    .HRDATA(HRDATA),
    .HREADY(HREADY),
    .HRESETn(HRESETn),
    .HRESP(HRESP),
    .IRQ(IRQ),
    .IRQLATENCY(IRQLATENCY),
    .NMI(NMI),
    .PORESETn(PORESETn),
    .RSTBYPASS(RSTBYPASS),
    .RXEV(RXEV),
    .SCLK(SCLK),
    .SE(SE),
    .SLEEPHOLDREQn(SLEEPHOLDREQn),
    .STCALIB(STCALIB),
    .STCLKEN(STCLKEN),
    .SWCLKTCK(SWCLKTCK),
    .SWDITMS(SWDITMS),
    .TDI(TDI),
    .WICENREQ(WICENREQ),
    .nTRST(nTRST),
    .CDBGPWRUPREQ(CDBGPWRUPREQ),
    .CODEHINTDE(CODEHINTDE),
    .CODENSEQ(CODENSEQ),
    .DBGRESTARTED(DBGRESTARTED),
    .GATEHCLK(GATEHCLK),
    .HADDR(HADDR),
    .HALTED(HALTED),
    .HBURST(HBURST),
    .HMASTER(HMASTER),
    .HMASTLOCK(HMASTLOCK),
    .HPROT(HPROT),
    .HSIZE(HSIZE),
    .HTRANS(HTRANS),
    .HWDATA(HWDATA),
    .HWRITE(HWRITE),
    .LOCKUP(LOCKUP),
    .SLEEPDEEP(SLEEPDEEP),
    .SLEEPHOLDACKn(SLEEPHOLDACKn),
    .SLEEPING(SLEEPING),
    .SPECHTRANS(SPECHTRANS),
    .SWDO(SWDO),
    .SWDOEN(SWDOEN),
    .SYSRESETREQ(SYSRESETREQ),
    .TDO(TDO),
    .TXEV(TXEV),
    .WAKEUP(WAKEUP),
    .WICENACK(WICENACK),
    .WICSENSE(WICSENSE),
    .nTDOEN(nTDOEN));  // ../RTL/CORTEXM0INTEGRATION.v(139)

endmodule 

module \cmsdk_ahb_cs_rom_table(BASE=32'b11110000000000000000000000000000,ENTRY0BASEADDR=32'b11100000000011111111000000000000,ENTRY0PRESENT=1'b1,ENTRY1BASEADDR=32'b11110000001000000000000000000000,ENTRY1PRESENT=0)   // ../RTL/cmsdk_ahb_cs_rom_table.v(67)
  (
  ECOREVNUM,
  HADDR,
  HBURST,
  HCLK,
  HMASTLOCK,
  HPROT,
  HREADY,
  HSEL,
  HSIZE,
  HTRANS,
  HWDATA,
  HWRITE,
  HRDATA,
  HREADYOUT,
  HRESP
  );

  input [3:0] ECOREVNUM;  // ../RTL/cmsdk_ahb_cs_rom_table.v(110)
  input [31:0] HADDR;  // ../RTL/cmsdk_ahb_cs_rom_table.v(101)
  input [2:0] HBURST;  // ../RTL/cmsdk_ahb_cs_rom_table.v(102)
  input HCLK;  // ../RTL/cmsdk_ahb_cs_rom_table.v(99)
  input HMASTLOCK;  // ../RTL/cmsdk_ahb_cs_rom_table.v(103)
  input [3:0] HPROT;  // ../RTL/cmsdk_ahb_cs_rom_table.v(104)
  input HREADY;  // ../RTL/cmsdk_ahb_cs_rom_table.v(109)
  input HSEL;  // ../RTL/cmsdk_ahb_cs_rom_table.v(100)
  input [2:0] HSIZE;  // ../RTL/cmsdk_ahb_cs_rom_table.v(105)
  input [1:0] HTRANS;  // ../RTL/cmsdk_ahb_cs_rom_table.v(106)
  input [31:0] HWDATA;  // ../RTL/cmsdk_ahb_cs_rom_table.v(107)
  input HWRITE;  // ../RTL/cmsdk_ahb_cs_rom_table.v(108)
  output [31:0] HRDATA;  // ../RTL/cmsdk_ahb_cs_rom_table.v(111)
  output HREADYOUT;  // ../RTL/cmsdk_ahb_cs_rom_table.v(113)
  output HRESP;  // ../RTL/cmsdk_ahb_cs_rom_table.v(112)

  parameter BASE = 32'b11110000000000000000000000000000;
  parameter ENTRY0BASEADDR = 32'b11100000000011111111000000000000;
  parameter ENTRY0PRESENT = 1'b1;
  parameter ENTRY1BASEADDR = 32'b11110000001000000000000000000000;
  parameter ENTRY1PRESENT = 0;
  parameter ENTRY2BASEADDR = 32'b00000000000000000000000000000000;
  parameter ENTRY2PRESENT = 1'b0;
  parameter ENTRY3BASEADDR = 32'b00000000000000000000000000000000;
  parameter ENTRY3PRESENT = 1'b0;
  parameter JEPCONTINUATION = 4'b0000;
  parameter JEPID = 7'b0000000;
  parameter PARTNUMBER = 12'b000000000000;
  parameter REVISION = 4'b0000;
  // localparam ENTRY0 = 32'b11110000000011111111000000000011;
  // localparam ENTRY0OFFSET = 20'b11110000000011111111;
  // localparam ENTRY1 = 32'b00000000001000000000000000000010;
  // localparam ENTRY1OFFSET = 20'b00000000001000000000;
  // localparam ENTRY2 = 32'b00010000000000000000000000000010;
  // localparam ENTRY2OFFSET = 20'b00010000000000000000;
  // localparam ENTRY3 = 32'b00010000000000000000000000000010;
  // localparam ENTRY3OFFSET = 20'b00010000000000000000;
  wire [9:0] haddr_reg;  // ../RTL/cmsdk_ahb_cs_rom_table.v(118)
  wire [7:0] ids;  // ../RTL/cmsdk_ahb_cs_rom_table.v(200)
  wire [9:0] n1;
  wire [7:0] n2;
  wire [7:0] n3;
  wire [7:0] n4;
  wire [31:0] n5;
  wire [31:0] n6;
  wire [31:0] n7;
  wire [31:0] rdata;  // ../RTL/cmsdk_ahb_cs_rom_table.v(119)
  wire [11:0] word_addr;  // ../RTL/cmsdk_ahb_cs_rom_table.v(167)
  wire cid0_en;  // ../RTL/cmsdk_ahb_cs_rom_table.v(182)
  wire cid1_en;  // ../RTL/cmsdk_ahb_cs_rom_table.v(181)
  wire cid2_en;  // ../RTL/cmsdk_ahb_cs_rom_table.v(180)
  wire cid3_en;  // ../RTL/cmsdk_ahb_cs_rom_table.v(179)
  wire entry1_en;  // ../RTL/cmsdk_ahb_cs_rom_table.v(196)
  wire entry2_en;  // ../RTL/cmsdk_ahb_cs_rom_table.v(197)
  wire entry3_en;  // ../RTL/cmsdk_ahb_cs_rom_table.v(198)
  wire n0;
  wire pid2_en;  // ../RTL/cmsdk_ahb_cs_rom_table.v(189)
  wire pid3_en;  // ../RTL/cmsdk_ahb_cs_rom_table.v(188)
  wire systemaccess_en;  // ../RTL/cmsdk_ahb_cs_rom_table.v(193)
  wire trans_valid;  // ../RTL/cmsdk_ahb_cs_rom_table.v(157)

  eq_w12 eq0 (
    .i0(word_addr),
    .i1(12'b111111111100),
    .o(cid3_en));  // ../RTL/cmsdk_ahb_cs_rom_table.v(179)
  eq_w12 eq1 (
    .i0(word_addr),
    .i1(12'b111111111000),
    .o(cid2_en));  // ../RTL/cmsdk_ahb_cs_rom_table.v(180)
  eq_w12 eq10 (
    .i0(word_addr),
    .i1(12'b000000001100),
    .o(entry3_en));  // ../RTL/cmsdk_ahb_cs_rom_table.v(198)
  eq_w12 eq2 (
    .i0(word_addr),
    .i1(12'b111111110100),
    .o(cid1_en));  // ../RTL/cmsdk_ahb_cs_rom_table.v(181)
  eq_w12 eq3 (
    .i0(word_addr),
    .i1(12'b111111110000),
    .o(cid0_en));  // ../RTL/cmsdk_ahb_cs_rom_table.v(182)
  eq_w12 eq4 (
    .i0(word_addr),
    .i1(12'b111111101100),
    .o(pid3_en));  // ../RTL/cmsdk_ahb_cs_rom_table.v(188)
  eq_w12 eq5 (
    .i0(word_addr),
    .i1(12'b111111101000),
    .o(pid2_en));  // ../RTL/cmsdk_ahb_cs_rom_table.v(189)
  eq_w12 eq6 (
    .i0(word_addr),
    .i1(12'b111111001100),
    .o(systemaccess_en));  // ../RTL/cmsdk_ahb_cs_rom_table.v(193)
  eq_w12 eq7 (
    .i0(word_addr),
    .i1(12'b000000000000),
    .o(rdata[31]));  // ../RTL/cmsdk_ahb_cs_rom_table.v(195)
  eq_w12 eq8 (
    .i0(word_addr),
    .i1(12'b000000000100),
    .o(entry1_en));  // ../RTL/cmsdk_ahb_cs_rom_table.v(196)
  eq_w12 eq9 (
    .i0(word_addr),
    .i1(12'b000000001000),
    .o(entry2_en));  // ../RTL/cmsdk_ahb_cs_rom_table.v(197)
  binary_mux_s1_w10 mux0 (
    .i0(haddr_reg),
    .i1(HADDR[11:2]),
    .sel(trans_valid),
    .o(n1));  // ../RTL/cmsdk_ahb_cs_rom_table.v(161)
  reg_ar_as_w10 reg0 (
    .clk(HCLK),
    .d(n1),
    .reset(10'b0000000000),
    .set(10'b0000000000),
    .q(haddr_reg));  // ../RTL/cmsdk_ahb_cs_rom_table.v(161)
  or u10 (ids[0], n2[0], cid0_en);  // ../RTL/cmsdk_ahb_cs_rom_table.v(204)
  or u11 (n5[0], ids[0], systemaccess_en);  // ../RTL/cmsdk_ahb_cs_rom_table.v(222)
  or u12 (rdata[0], n5[0], rdata[31]);  // ../RTL/cmsdk_ahb_cs_rom_table.v(224)
  or u13 (rdata[28], n7[28], entry3_en);  // ../RTL/cmsdk_ahb_cs_rom_table.v(228)
  or u14 (n7[1], n6[1], entry2_en);  // ../RTL/cmsdk_ahb_cs_rom_table.v(226)
  or u15 (n7[28], rdata[31], entry2_en);  // ../RTL/cmsdk_ahb_cs_rom_table.v(226)
  or u16 (n6[1], rdata[31], entry1_en);  // ../RTL/cmsdk_ahb_cs_rom_table.v(225)
  or u17 (ids[3], cid0_en, pid2_en);  // ../RTL/cmsdk_ahb_cs_rom_table.v(211)
  or u18 (ids[4], n3[4], n4[4]);  // ../RTL/cmsdk_ahb_cs_rom_table.v(210)
  or u19 (ids[5], cid3_en, n4[5]);  // ../RTL/cmsdk_ahb_cs_rom_table.v(210)
  and u2 (n0, HSEL, HTRANS[1]);  // ../RTL/cmsdk_ahb_cs_rom_table.v(157)
  or u20 (ids[7], cid3_en, n4[7]);  // ../RTL/cmsdk_ahb_cs_rom_table.v(210)
  and u21 (n4[4], pid3_en, ECOREVNUM[0]);  // ../RTL/cmsdk_ahb_cs_rom_table.v(210)
  and u22 (n4[5], pid3_en, ECOREVNUM[1]);  // ../RTL/cmsdk_ahb_cs_rom_table.v(210)
  and u23 (ids[6], pid3_en, ECOREVNUM[2]);  // ../RTL/cmsdk_ahb_cs_rom_table.v(210)
  and u24 (n4[7], pid3_en, ECOREVNUM[3]);  // ../RTL/cmsdk_ahb_cs_rom_table.v(210)
  or u25 (ids[2], cid2_en, cid0_en);  // ../RTL/cmsdk_ahb_cs_rom_table.v(204)
  or u26 (n3[4], cid3_en, cid1_en);  // ../RTL/cmsdk_ahb_cs_rom_table.v(203)
  buf u27 (word_addr[1], 1'b0);  // ../RTL/cmsdk_ahb_cs_rom_table.v(167)
  buf u28 (word_addr[2], haddr_reg[0]);  // ../RTL/cmsdk_ahb_cs_rom_table.v(167)
  buf u29 (word_addr[3], haddr_reg[1]);  // ../RTL/cmsdk_ahb_cs_rom_table.v(167)
  and u3 (trans_valid, n0, HREADY);  // ../RTL/cmsdk_ahb_cs_rom_table.v(157)
  buf u30 (word_addr[4], haddr_reg[2]);  // ../RTL/cmsdk_ahb_cs_rom_table.v(167)
  buf u31 (word_addr[5], haddr_reg[3]);  // ../RTL/cmsdk_ahb_cs_rom_table.v(167)
  buf u32 (word_addr[6], haddr_reg[4]);  // ../RTL/cmsdk_ahb_cs_rom_table.v(167)
  buf u33 (word_addr[7], haddr_reg[5]);  // ../RTL/cmsdk_ahb_cs_rom_table.v(167)
  buf u34 (word_addr[8], haddr_reg[6]);  // ../RTL/cmsdk_ahb_cs_rom_table.v(167)
  buf u35 (word_addr[9], haddr_reg[7]);  // ../RTL/cmsdk_ahb_cs_rom_table.v(167)
  buf u36 (word_addr[10], haddr_reg[8]);  // ../RTL/cmsdk_ahb_cs_rom_table.v(167)
  buf u37 (word_addr[11], haddr_reg[9]);  // ../RTL/cmsdk_ahb_cs_rom_table.v(167)
  buf u38 (HRDATA[1], rdata[1]);  // ../RTL/cmsdk_ahb_cs_rom_table.v(164)
  buf u39 (HRDATA[2], ids[2]);  // ../RTL/cmsdk_ahb_cs_rom_table.v(164)
  buf u4 (HREADYOUT, 1'b1);  // ../RTL/cmsdk_ahb_cs_rom_table.v(163)
  buf u40 (HRDATA[3], ids[3]);  // ../RTL/cmsdk_ahb_cs_rom_table.v(164)
  buf u41 (HRDATA[4], ids[4]);  // ../RTL/cmsdk_ahb_cs_rom_table.v(164)
  buf u42 (HRDATA[5], ids[5]);  // ../RTL/cmsdk_ahb_cs_rom_table.v(164)
  buf u43 (HRDATA[6], ids[6]);  // ../RTL/cmsdk_ahb_cs_rom_table.v(164)
  buf u44 (HRDATA[7], ids[7]);  // ../RTL/cmsdk_ahb_cs_rom_table.v(164)
  buf u45 (HRDATA[8], 1'b0);  // ../RTL/cmsdk_ahb_cs_rom_table.v(164)
  buf u46 (HRDATA[9], 1'b0);  // ../RTL/cmsdk_ahb_cs_rom_table.v(164)
  buf u47 (HRDATA[10], 1'b0);  // ../RTL/cmsdk_ahb_cs_rom_table.v(164)
  buf u48 (HRDATA[11], 1'b0);  // ../RTL/cmsdk_ahb_cs_rom_table.v(164)
  buf u49 (HRDATA[12], rdata[31]);  // ../RTL/cmsdk_ahb_cs_rom_table.v(164)
  buf u5 (HRESP, 1'b0);  // ../RTL/cmsdk_ahb_cs_rom_table.v(165)
  buf u50 (HRDATA[13], rdata[31]);  // ../RTL/cmsdk_ahb_cs_rom_table.v(164)
  buf u51 (HRDATA[14], rdata[31]);  // ../RTL/cmsdk_ahb_cs_rom_table.v(164)
  buf u52 (HRDATA[15], rdata[31]);  // ../RTL/cmsdk_ahb_cs_rom_table.v(164)
  buf u53 (HRDATA[16], rdata[31]);  // ../RTL/cmsdk_ahb_cs_rom_table.v(164)
  buf u54 (HRDATA[17], rdata[31]);  // ../RTL/cmsdk_ahb_cs_rom_table.v(164)
  buf u55 (HRDATA[18], rdata[31]);  // ../RTL/cmsdk_ahb_cs_rom_table.v(164)
  buf u56 (HRDATA[19], rdata[31]);  // ../RTL/cmsdk_ahb_cs_rom_table.v(164)
  buf u57 (HRDATA[20], 1'b0);  // ../RTL/cmsdk_ahb_cs_rom_table.v(164)
  buf u58 (HRDATA[21], entry1_en);  // ../RTL/cmsdk_ahb_cs_rom_table.v(164)
  buf u59 (HRDATA[22], 1'b0);  // ../RTL/cmsdk_ahb_cs_rom_table.v(164)
  buf u6 (HRDATA[0], rdata[0]);  // ../RTL/cmsdk_ahb_cs_rom_table.v(164)
  buf u60 (HRDATA[23], 1'b0);  // ../RTL/cmsdk_ahb_cs_rom_table.v(164)
  buf u61 (HRDATA[24], 1'b0);  // ../RTL/cmsdk_ahb_cs_rom_table.v(164)
  buf u62 (HRDATA[25], 1'b0);  // ../RTL/cmsdk_ahb_cs_rom_table.v(164)
  buf u63 (HRDATA[26], 1'b0);  // ../RTL/cmsdk_ahb_cs_rom_table.v(164)
  buf u64 (HRDATA[27], 1'b0);  // ../RTL/cmsdk_ahb_cs_rom_table.v(164)
  buf u65 (HRDATA[28], rdata[28]);  // ../RTL/cmsdk_ahb_cs_rom_table.v(164)
  buf u66 (HRDATA[29], rdata[31]);  // ../RTL/cmsdk_ahb_cs_rom_table.v(164)
  buf u67 (HRDATA[30], rdata[31]);  // ../RTL/cmsdk_ahb_cs_rom_table.v(164)
  buf u68 (HRDATA[31], rdata[31]);  // ../RTL/cmsdk_ahb_cs_rom_table.v(164)
  or u7 (rdata[1], n7[1], entry3_en);  // ../RTL/cmsdk_ahb_cs_rom_table.v(228)
  buf u8 (word_addr[0], 1'b0);  // ../RTL/cmsdk_ahb_cs_rom_table.v(167)
  or u9 (n2[0], cid3_en, cid2_en);  // ../RTL/cmsdk_ahb_cs_rom_table.v(202)

endmodule 

module eq_w9
  (
  i0,
  i1,
  o
  );

  input [8:0] i0;
  input [8:0] i1;
  output o;



endmodule 

module eq_w16
  (
  i0,
  i1,
  o
  );

  input [15:0] i0;
  input [15:0] i1;
  output o;



endmodule 

module eq_w20
  (
  i0,
  i1,
  o
  );

  input [19:0] i0;
  input [19:0] i1;
  output o;



endmodule 

module reg_ar_as_w2
  (
  clk,
  d,
  en,
  reset,
  set,
  q
  );

  input clk;
  input [1:0] d;
  input en;
  input [1:0] reset;
  input [1:0] set;
  output [1:0] q;



endmodule 

module cmsdk_ahb_to_iop  // ../RTL/cmsdk_ahb_to_iop.v(28)
  (
  HADDR,
  HCLK,
  HREADY,
  HRESETn,
  HSEL,
  HSIZE,
  HTRANS,
  HWDATA,
  HWRITE,
  IORDATA,
  HRDATA,
  HREADYOUT,
  HRESP,
  IOADDR,
  IOSEL,
  IOSIZE,
  IOTRANS,
  IOWDATA,
  IOWRITE
  );

  input [11:0] HADDR;  // ../RTL/cmsdk_ahb_to_iop.v(40)
  input HCLK;  // ../RTL/cmsdk_ahb_to_iop.v(33)
  input HREADY;  // ../RTL/cmsdk_ahb_to_iop.v(36)
  input HRESETn;  // ../RTL/cmsdk_ahb_to_iop.v(34)
  input HSEL;  // ../RTL/cmsdk_ahb_to_iop.v(35)
  input [2:0] HSIZE;  // ../RTL/cmsdk_ahb_to_iop.v(38)
  input [1:0] HTRANS;  // ../RTL/cmsdk_ahb_to_iop.v(37)
  input [31:0] HWDATA;  // ../RTL/cmsdk_ahb_to_iop.v(41)
  input HWRITE;  // ../RTL/cmsdk_ahb_to_iop.v(39)
  input [31:0] IORDATA;  // ../RTL/cmsdk_ahb_to_iop.v(44)
  output [31:0] HRDATA;  // ../RTL/cmsdk_ahb_to_iop.v(49)
  output HREADYOUT;  // ../RTL/cmsdk_ahb_to_iop.v(47)
  output HRESP;  // ../RTL/cmsdk_ahb_to_iop.v(48)
  output [11:0] IOADDR;  // ../RTL/cmsdk_ahb_to_iop.v(53)
  output IOSEL;  // ../RTL/cmsdk_ahb_to_iop.v(52)
  output [1:0] IOSIZE;  // ../RTL/cmsdk_ahb_to_iop.v(55)
  output IOTRANS;  // ../RTL/cmsdk_ahb_to_iop.v(56)
  output [31:0] IOWDATA;  // ../RTL/cmsdk_ahb_to_iop.v(57)
  output IOWRITE;  // ../RTL/cmsdk_ahb_to_iop.v(54)

  wire n0;
  wire n1;

  AL_DFF IOSEL_reg (
    .clk(HCLK),
    .d(n0),
    .reset(n1),
    .set(1'b0),
    .q(IOSEL));  // ../RTL/cmsdk_ahb_to_iop.v(69)
  AL_DFF IOTRANS_reg (
    .clk(HCLK),
    .d(HTRANS[1]),
    .reset(n1),
    .set(1'b0),
    .q(IOTRANS));  // ../RTL/cmsdk_ahb_to_iop.v(105)
  AL_DFF IOWRITE_reg (
    .clk(HCLK),
    .d(HWRITE),
    .reset(n1),
    .set(1'b0),
    .q(IOWRITE));  // ../RTL/cmsdk_ahb_to_iop.v(87)
  reg_ar_as_w12 reg0 (
    .clk(HCLK),
    .d(HADDR),
    .reset({n1,n1,n1,n1,n1,n1,n1,n1,n1,n1,n1,n1}),
    .set(12'b000000000000),
    .q(IOADDR));  // ../RTL/cmsdk_ahb_to_iop.v(78)
  reg_ar_as_w2 reg1 (
    .clk(HCLK),
    .d(HSIZE[1:0]),
    .reset({n1,n1}),
    .set(2'b00),
    .q(IOSIZE));  // ../RTL/cmsdk_ahb_to_iop.v(96)
  buf u10 (HRDATA[2], IORDATA[2]);  // ../RTL/cmsdk_ahb_to_iop.v(109)
  buf u11 (HRDATA[5], IORDATA[5]);  // ../RTL/cmsdk_ahb_to_iop.v(109)
  buf u12 (HRDATA[1], IORDATA[1]);  // ../RTL/cmsdk_ahb_to_iop.v(109)
  buf u13 (HRDATA[4], IORDATA[4]);  // ../RTL/cmsdk_ahb_to_iop.v(109)
  buf u14 (HRDATA[0], IORDATA[0]);  // ../RTL/cmsdk_ahb_to_iop.v(109)
  buf u15 (HRDATA[11], IORDATA[11]);  // ../RTL/cmsdk_ahb_to_iop.v(109)
  buf u16 (IOWDATA[0], HWDATA[0]);  // ../RTL/cmsdk_ahb_to_iop.v(108)
  buf u17 (HREADYOUT, 1'b1);  // ../RTL/cmsdk_ahb_to_iop.v(110)
  buf u18 (HRESP, 1'b0);  // ../RTL/cmsdk_ahb_to_iop.v(111)
  buf u19 (HRDATA[12], IORDATA[12]);  // ../RTL/cmsdk_ahb_to_iop.v(109)
  buf u2 (HRDATA[10], IORDATA[10]);  // ../RTL/cmsdk_ahb_to_iop.v(109)
  buf u20 (HRDATA[13], IORDATA[13]);  // ../RTL/cmsdk_ahb_to_iop.v(109)
  buf u21 (HRDATA[14], IORDATA[14]);  // ../RTL/cmsdk_ahb_to_iop.v(109)
  buf u22 (HRDATA[15], IORDATA[15]);  // ../RTL/cmsdk_ahb_to_iop.v(109)
  buf u23 (HRDATA[16], IORDATA[16]);  // ../RTL/cmsdk_ahb_to_iop.v(109)
  buf u24 (HRDATA[17], IORDATA[17]);  // ../RTL/cmsdk_ahb_to_iop.v(109)
  buf u25 (HRDATA[18], IORDATA[18]);  // ../RTL/cmsdk_ahb_to_iop.v(109)
  buf u26 (HRDATA[19], IORDATA[19]);  // ../RTL/cmsdk_ahb_to_iop.v(109)
  buf u27 (HRDATA[20], IORDATA[20]);  // ../RTL/cmsdk_ahb_to_iop.v(109)
  buf u28 (HRDATA[21], IORDATA[21]);  // ../RTL/cmsdk_ahb_to_iop.v(109)
  buf u29 (HRDATA[22], IORDATA[22]);  // ../RTL/cmsdk_ahb_to_iop.v(109)
  buf u3 (HRDATA[9], IORDATA[9]);  // ../RTL/cmsdk_ahb_to_iop.v(109)
  buf u30 (HRDATA[23], IORDATA[23]);  // ../RTL/cmsdk_ahb_to_iop.v(109)
  buf u31 (HRDATA[24], IORDATA[24]);  // ../RTL/cmsdk_ahb_to_iop.v(109)
  buf u32 (HRDATA[25], IORDATA[25]);  // ../RTL/cmsdk_ahb_to_iop.v(109)
  buf u33 (HRDATA[26], IORDATA[26]);  // ../RTL/cmsdk_ahb_to_iop.v(109)
  buf u34 (HRDATA[27], IORDATA[27]);  // ../RTL/cmsdk_ahb_to_iop.v(109)
  buf u35 (HRDATA[28], IORDATA[28]);  // ../RTL/cmsdk_ahb_to_iop.v(109)
  buf u36 (HRDATA[29], IORDATA[29]);  // ../RTL/cmsdk_ahb_to_iop.v(109)
  buf u37 (HRDATA[30], IORDATA[30]);  // ../RTL/cmsdk_ahb_to_iop.v(109)
  buf u38 (HRDATA[31], IORDATA[31]);  // ../RTL/cmsdk_ahb_to_iop.v(109)
  buf u39 (IOWDATA[1], HWDATA[1]);  // ../RTL/cmsdk_ahb_to_iop.v(108)
  buf u4 (HRDATA[8], IORDATA[8]);  // ../RTL/cmsdk_ahb_to_iop.v(109)
  buf u40 (IOWDATA[2], HWDATA[2]);  // ../RTL/cmsdk_ahb_to_iop.v(108)
  buf u41 (IOWDATA[3], HWDATA[3]);  // ../RTL/cmsdk_ahb_to_iop.v(108)
  buf u42 (IOWDATA[4], HWDATA[4]);  // ../RTL/cmsdk_ahb_to_iop.v(108)
  buf u43 (IOWDATA[5], HWDATA[5]);  // ../RTL/cmsdk_ahb_to_iop.v(108)
  buf u44 (IOWDATA[6], HWDATA[6]);  // ../RTL/cmsdk_ahb_to_iop.v(108)
  buf u45 (IOWDATA[7], HWDATA[7]);  // ../RTL/cmsdk_ahb_to_iop.v(108)
  buf u46 (IOWDATA[8], HWDATA[8]);  // ../RTL/cmsdk_ahb_to_iop.v(108)
  buf u47 (IOWDATA[9], HWDATA[9]);  // ../RTL/cmsdk_ahb_to_iop.v(108)
  buf u48 (IOWDATA[10], HWDATA[10]);  // ../RTL/cmsdk_ahb_to_iop.v(108)
  buf u49 (IOWDATA[11], HWDATA[11]);  // ../RTL/cmsdk_ahb_to_iop.v(108)
  not u5 (n1, HRESETn);  // ../RTL/cmsdk_ahb_to_iop.v(66)
  buf u50 (IOWDATA[12], HWDATA[12]);  // ../RTL/cmsdk_ahb_to_iop.v(108)
  buf u51 (IOWDATA[13], HWDATA[13]);  // ../RTL/cmsdk_ahb_to_iop.v(108)
  buf u52 (IOWDATA[14], HWDATA[14]);  // ../RTL/cmsdk_ahb_to_iop.v(108)
  buf u53 (IOWDATA[15], HWDATA[15]);  // ../RTL/cmsdk_ahb_to_iop.v(108)
  buf u54 (IOWDATA[16], HWDATA[16]);  // ../RTL/cmsdk_ahb_to_iop.v(108)
  buf u55 (IOWDATA[17], HWDATA[17]);  // ../RTL/cmsdk_ahb_to_iop.v(108)
  buf u56 (IOWDATA[18], HWDATA[18]);  // ../RTL/cmsdk_ahb_to_iop.v(108)
  buf u57 (IOWDATA[19], HWDATA[19]);  // ../RTL/cmsdk_ahb_to_iop.v(108)
  buf u58 (IOWDATA[20], HWDATA[20]);  // ../RTL/cmsdk_ahb_to_iop.v(108)
  buf u59 (IOWDATA[21], HWDATA[21]);  // ../RTL/cmsdk_ahb_to_iop.v(108)
  and u6 (n0, HSEL, HREADY);  // ../RTL/cmsdk_ahb_to_iop.v(69)
  buf u60 (IOWDATA[22], HWDATA[22]);  // ../RTL/cmsdk_ahb_to_iop.v(108)
  buf u61 (IOWDATA[23], HWDATA[23]);  // ../RTL/cmsdk_ahb_to_iop.v(108)
  buf u62 (IOWDATA[24], HWDATA[24]);  // ../RTL/cmsdk_ahb_to_iop.v(108)
  buf u63 (IOWDATA[25], HWDATA[25]);  // ../RTL/cmsdk_ahb_to_iop.v(108)
  buf u64 (IOWDATA[26], HWDATA[26]);  // ../RTL/cmsdk_ahb_to_iop.v(108)
  buf u65 (IOWDATA[27], HWDATA[27]);  // ../RTL/cmsdk_ahb_to_iop.v(108)
  buf u66 (IOWDATA[28], HWDATA[28]);  // ../RTL/cmsdk_ahb_to_iop.v(108)
  buf u67 (IOWDATA[29], HWDATA[29]);  // ../RTL/cmsdk_ahb_to_iop.v(108)
  buf u68 (IOWDATA[30], HWDATA[30]);  // ../RTL/cmsdk_ahb_to_iop.v(108)
  buf u69 (IOWDATA[31], HWDATA[31]);  // ../RTL/cmsdk_ahb_to_iop.v(108)
  buf u7 (HRDATA[7], IORDATA[7]);  // ../RTL/cmsdk_ahb_to_iop.v(109)
  buf u8 (HRDATA[3], IORDATA[3]);  // ../RTL/cmsdk_ahb_to_iop.v(109)
  buf u9 (HRDATA[6], IORDATA[6]);  // ../RTL/cmsdk_ahb_to_iop.v(109)

endmodule 

module cmsdk_iop_gpio  // ../RTL/cmsdk_iop_gpio.v(46)
  (
  ECOREVNUM,
  FCLK,
  HCLK,
  HRESETn,
  IOADDR,
  IOSEL,
  IOSIZE,
  IOTRANS,
  IOWDATA,
  IOWRITE,
  PORTIN,
  COMBINT,
  GPIOINT,
  IORDATA,
  PORTEN,
  PORTFUNC,
  PORTOUT
  );

  input [3:0] ECOREVNUM;  // ../RTL/cmsdk_iop_gpio.v(75)
  input FCLK;  // ../RTL/cmsdk_iop_gpio.v(65)
  input HCLK;  // ../RTL/cmsdk_iop_gpio.v(66)
  input HRESETn;  // ../RTL/cmsdk_iop_gpio.v(67)
  input [11:0] IOADDR;  // ../RTL/cmsdk_iop_gpio.v(69)
  input IOSEL;  // ../RTL/cmsdk_iop_gpio.v(68)
  input [1:0] IOSIZE;  // ../RTL/cmsdk_iop_gpio.v(71)
  input IOTRANS;  // ../RTL/cmsdk_iop_gpio.v(72)
  input [31:0] IOWDATA;  // ../RTL/cmsdk_iop_gpio.v(73)
  input IOWRITE;  // ../RTL/cmsdk_iop_gpio.v(70)
  input [15:0] PORTIN;  // ../RTL/cmsdk_iop_gpio.v(77)
  output COMBINT;  // ../RTL/cmsdk_iop_gpio.v(87)
  output [15:0] GPIOINT;  // ../RTL/cmsdk_iop_gpio.v(86)
  output [31:0] IORDATA;  // ../RTL/cmsdk_iop_gpio.v(80)
  output [15:0] PORTEN;  // ../RTL/cmsdk_iop_gpio.v(83)
  output [15:0] PORTFUNC;  // ../RTL/cmsdk_iop_gpio.v(84)
  output [15:0] PORTOUT;  // ../RTL/cmsdk_iop_gpio.v(82)

  parameter ALTERNATE_FUNC_DEFAULT = 16'b0000000000000000;
  parameter ALTERNATE_FUNC_MASK = 16'b1111111111111111;
  parameter BE = 0;
  // localparam ARM_CMSDK_IOP_GPIO_CID0 = 32'b00000000000000000000000000001101;
  // localparam ARM_CMSDK_IOP_GPIO_CID1 = 32'b00000000000000000000000011110000;
  // localparam ARM_CMSDK_IOP_GPIO_CID2 = 32'b00000000000000000000000000000101;
  // localparam ARM_CMSDK_IOP_GPIO_CID3 = 32'b00000000000000000000000010110001;
  // localparam ARM_CMSDK_IOP_GPIO_PID0 = 32'b00000000000000000000000000100000;
  // localparam ARM_CMSDK_IOP_GPIO_PID1 = 32'b00000000000000000000000010111000;
  // localparam ARM_CMSDK_IOP_GPIO_PID2 = 32'b00000000000000000000000000011011;
  // localparam ARM_CMSDK_IOP_GPIO_PID3 = 32'b00000000000000000000000000000000;
  // localparam ARM_CMSDK_IOP_GPIO_PID4 = 32'b00000000000000000000000000000100;
  // localparam ARM_CMSDK_IOP_GPIO_PID5 = 32'b00000000000000000000000000000000;
  // localparam ARM_CMSDK_IOP_GPIO_PID6 = 32'b00000000000000000000000000000000;
  // localparam ARM_CMSDK_IOP_GPIO_PID7 = 32'b00000000000000000000000000000000;
  // localparam PortWidth = 16;
  wire [31:0] IOWDATALE;  // ../RTL/cmsdk_iop_gpio.v(132)
  wire [32:0] current_dout_padded;  // ../RTL/cmsdk_iop_gpio.v(262)
  wire [15:0] fall_edge_int;  // ../RTL/cmsdk_iop_gpio.v(553)
  wire [15:0] high_level_int;  // ../RTL/cmsdk_iop_gpio.v(550)
  wire [1:0] iop_byte_strobe;  // ../RTL/cmsdk_iop_gpio.v(137)
  wire [15:0] low_level_int;  // ../RTL/cmsdk_iop_gpio.v(551)
  wire [7:0] n10;
  wire [7:0] n11;
  wire [31:0] n13;
  wire [31:0] n14;
  wire [31:0] n19;
  wire [1:0] n2;
  wire [31:0] n20;
  wire [1:0] n3;
  wire [7:0] n30;
  wire [15:0] n305;
  wire [15:0] n306;
  wire [15:0] n307;
  wire [15:0] n308;
  wire [15:0] n309;
  wire [7:0] n31;
  wire [15:0] n310;
  wire [7:0] n32;
  wire [15:0] n327;
  wire [15:0] n328;
  wire [15:0] n329;
  wire [7:0] n33;
  wire [15:0] n330;
  wire [15:0] n331;
  wire [15:0] n332;
  wire [15:0] n333;
  wire [15:0] n334;
  wire [15:0] n335;
  wire [7:0] n35;
  wire [7:0] n36;
  wire [7:0] n37;
  wire [7:0] n38;
  wire [1:0] n4;
  wire [7:0] n40;
  wire [1:0] n5;
  wire [31:0] n8;
  wire [31:0] n9;
  wire [15:0] new_masked_int;  // ../RTL/cmsdk_iop_gpio.v(517)
  wire [15:0] new_raw_int;  // ../RTL/cmsdk_iop_gpio.v(129)
  wire [15:0] nxt_dout_padded;  // ../RTL/cmsdk_iop_gpio.v(263)
  wire [31:0] read_mux;  // ../RTL/cmsdk_iop_gpio.v(114)
  wire [31:0] read_mux_le;  // ../RTL/cmsdk_iop_gpio.v(115)
  wire [15:0] reg_altfunc;  // ../RTL/cmsdk_iop_gpio.v(122)
  wire [15:0] reg_altfunc_padded;  // ../RTL/cmsdk_iop_gpio.v(359)
  wire [15:0] reg_altfuncclr;  // ../RTL/cmsdk_iop_gpio.v(362)
  wire [15:0] reg_altfuncset;  // ../RTL/cmsdk_iop_gpio.v(361)
  wire [15:0] reg_datain;  // ../RTL/cmsdk_iop_gpio.v(119)
  wire [31:0] reg_datain32;  // ../RTL/cmsdk_iop_gpio.v(118)
  wire [15:0] reg_dout;  // ../RTL/cmsdk_iop_gpio.v(120)
  wire [15:0] reg_dout_padded;  // ../RTL/cmsdk_iop_gpio.v(264)
  wire [15:0] reg_douten;  // ../RTL/cmsdk_iop_gpio.v(121)
  wire [15:0] reg_douten_padded;  // ../RTL/cmsdk_iop_gpio.v(319)
  wire [15:0] reg_doutenclr;  // ../RTL/cmsdk_iop_gpio.v(321)
  wire [15:0] reg_doutenset;  // ../RTL/cmsdk_iop_gpio.v(322)
  wire [15:0] reg_in_sync1;  // ../RTL/cmsdk_iop_gpio.v(238)
  wire [15:0] reg_in_sync2;  // ../RTL/cmsdk_iop_gpio.v(239)
  wire [15:0] reg_intclr_padded;  // ../RTL/cmsdk_iop_gpio.v(513)
  wire [15:0] reg_inten;  // ../RTL/cmsdk_iop_gpio.v(123)
  wire [15:0] reg_inten_padded;  // ../RTL/cmsdk_iop_gpio.v(397)
  wire [15:0] reg_intenclr;  // ../RTL/cmsdk_iop_gpio.v(400)
  wire [15:0] reg_intenset;  // ../RTL/cmsdk_iop_gpio.v(399)
  wire [15:0] reg_intpol;  // ../RTL/cmsdk_iop_gpio.v(125)
  wire [15:0] reg_intpol_padded;  // ../RTL/cmsdk_iop_gpio.v(474)
  wire [15:0] reg_intpolclr;  // ../RTL/cmsdk_iop_gpio.v(477)
  wire [15:0] reg_intpolset;  // ../RTL/cmsdk_iop_gpio.v(476)
  wire [15:0] reg_intstat;  // ../RTL/cmsdk_iop_gpio.v(126)
  wire [15:0] reg_intstat_padded;  // ../RTL/cmsdk_iop_gpio.v(511)
  wire [15:0] reg_inttype;  // ../RTL/cmsdk_iop_gpio.v(124)
  wire [15:0] reg_inttype_padded;  // ../RTL/cmsdk_iop_gpio.v(435)
  wire [15:0] reg_inttypeclr;  // ../RTL/cmsdk_iop_gpio.v(438)
  wire [15:0] reg_inttypeset;  // ../RTL/cmsdk_iop_gpio.v(437)
  wire [15:0] reg_last_datain;  // ../RTL/cmsdk_iop_gpio.v(549)
  wire [15:0] rise_edge_int;  // ../RTL/cmsdk_iop_gpio.v(552)
  wire bigendian;  // ../RTL/cmsdk_iop_gpio.v(131)
  wire n0;
  wire n1;
  wire n100;
  wire n101;
  wire n102;
  wire n103;
  wire n104;
  wire n105;
  wire n106;
  wire n107;
  wire n108;
  wire n109;
  wire n110;
  wire n111;
  wire n112;
  wire n113;
  wire n114;
  wire n115;
  wire n116;
  wire n117;
  wire n118;
  wire n119;
  wire n12;
  wire n120;
  wire n121;
  wire n122;
  wire n123;
  wire n124;
  wire n125;
  wire n126;
  wire n127;
  wire n128;
  wire n129;
  wire n130;
  wire n131;
  wire n132;
  wire n133;
  wire n134;
  wire n135;
  wire n136;
  wire n137;
  wire n138;
  wire n139;
  wire n140;
  wire n141;
  wire n142;
  wire n143;
  wire n144;
  wire n145;
  wire n146;
  wire n147;
  wire n148;
  wire n149;
  wire n15;
  wire n150;
  wire n151;
  wire n152;
  wire n153;
  wire n154;
  wire n155;
  wire n156;
  wire n157;
  wire n158;
  wire n159;
  wire n16;
  wire n160;
  wire n161;
  wire n162;
  wire n163;
  wire n164;
  wire n165;
  wire n166;
  wire n167;
  wire n168;
  wire n169;
  wire n17;
  wire n170;
  wire n171;
  wire n172;
  wire n173;
  wire n174;
  wire n175;
  wire n176;
  wire n177;
  wire n178;
  wire n179;
  wire n18;
  wire n180;
  wire n181;
  wire n182;
  wire n183;
  wire n184;
  wire n185;
  wire n186;
  wire n187;
  wire n188;
  wire n189;
  wire n190;
  wire n191;
  wire n192;
  wire n193;
  wire n194;
  wire n195;
  wire n196;
  wire n197;
  wire n198;
  wire n199;
  wire n200;
  wire n201;
  wire n202;
  wire n203;
  wire n204;
  wire n205;
  wire n206;
  wire n207;
  wire n208;
  wire n209;
  wire n21;
  wire n210;
  wire n211;
  wire n212;
  wire n213;
  wire n214;
  wire n215;
  wire n216;
  wire n217;
  wire n218;
  wire n219;
  wire n22;
  wire n220;
  wire n221;
  wire n222;
  wire n223;
  wire n224;
  wire n225;
  wire n226;
  wire n227;
  wire n228;
  wire n229;
  wire n23;
  wire n230;
  wire n231;
  wire n232;
  wire n233;
  wire n234;
  wire n235;
  wire n236;
  wire n237;
  wire n238;
  wire n239;
  wire n24;
  wire n240;
  wire n241;
  wire n242;
  wire n243;
  wire n244;
  wire n245;
  wire n246;
  wire n247;
  wire n248;
  wire n249;
  wire n25;
  wire n250;
  wire n251;
  wire n252;
  wire n253;
  wire n254;
  wire n255;
  wire n256;
  wire n257;
  wire n258;
  wire n259;
  wire n26;
  wire n260;
  wire n261;
  wire n262;
  wire n263;
  wire n264;
  wire n265;
  wire n266;
  wire n267;
  wire n268;
  wire n269;
  wire n27;
  wire n270;
  wire n271;
  wire n272;
  wire n273;
  wire n274;
  wire n275;
  wire n276;
  wire n277;
  wire n278;
  wire n279;
  wire n28;
  wire n280;
  wire n281;
  wire n282;
  wire n283;
  wire n284;
  wire n285;
  wire n286;
  wire n287;
  wire n288;
  wire n289;
  wire n29;
  wire n290;
  wire n291;
  wire n292;
  wire n293;
  wire n294;
  wire n295;
  wire n296;
  wire n297;
  wire n298;
  wire n299;
  wire n300;
  wire n301;
  wire n302;
  wire n303;
  wire n304;
  wire n311;
  wire n312;
  wire n313;
  wire n314;
  wire n315;
  wire n316;
  wire n317;
  wire n318;
  wire n319;
  wire n320;
  wire n321;
  wire n322;
  wire n323;
  wire n324;
  wire n325;
  wire n326;
  wire n34;
  wire n39;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n6;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n65;
  wire n66;
  wire n67;
  wire n68;
  wire n69;
  wire n7;
  wire n70;
  wire n71;
  wire n72;
  wire n73;
  wire n74;
  wire n75;
  wire n76;
  wire n77;
  wire n78;
  wire n79;
  wire n80;
  wire n81;
  wire n82;
  wire n83;
  wire n84;
  wire n85;
  wire n86;
  wire n87;
  wire n88;
  wire n89;
  wire n90;
  wire n91;
  wire n92;
  wire n93;
  wire n94;
  wire n95;
  wire n96;
  wire n97;
  wire n98;
  wire n99;
  wire reg_dout_masked_write0;  // ../RTL/cmsdk_iop_gpio.v(267)
  wire reg_dout_masked_write1;  // ../RTL/cmsdk_iop_gpio.v(268)
  wire reg_dout_normal_write0;  // ../RTL/cmsdk_iop_gpio.v(265)
  wire reg_dout_normal_write1;  // ../RTL/cmsdk_iop_gpio.v(266)
  wire reg_intclr_normal_write0;  // ../RTL/cmsdk_iop_gpio.v(514)
  wire reg_intclr_normal_write1;  // ../RTL/cmsdk_iop_gpio.v(515)
  wire write_trans;  // ../RTL/cmsdk_iop_gpio.v(135)

  eq_w2 eq0 (
    .i0(IOADDR[1:0]),
    .i1(2'b00),
    .o(n1));  // ../RTL/cmsdk_iop_gpio.v(142)
  eq_w2 eq1 (
    .i0(IOADDR[1:0]),
    .i1(2'b01),
    .o(n6));  // ../RTL/cmsdk_iop_gpio.v(143)
  eq_w10 eq10 (
    .i0(IOADDR[11:2]),
    .i1(10'b0000000100),
    .o(n41));  // ../RTL/cmsdk_iop_gpio.v(325)
  eq_w10 eq11 (
    .i0(IOADDR[11:2]),
    .i1(10'b0000000101),
    .o(n47));  // ../RTL/cmsdk_iop_gpio.v(331)
  eq_w10 eq12 (
    .i0(IOADDR[11:2]),
    .i1(10'b0000000110),
    .o(n86));  // ../RTL/cmsdk_iop_gpio.v(364)
  eq_w10 eq13 (
    .i0(IOADDR[11:2]),
    .i1(10'b0000000111),
    .o(n92));  // ../RTL/cmsdk_iop_gpio.v(370)
  eq_w10 eq14 (
    .i0(IOADDR[11:2]),
    .i1(10'b0000001000),
    .o(n131));  // ../RTL/cmsdk_iop_gpio.v(402)
  eq_w10 eq15 (
    .i0(IOADDR[11:2]),
    .i1(10'b0000001001),
    .o(n137));  // ../RTL/cmsdk_iop_gpio.v(408)
  eq_w10 eq16 (
    .i0(IOADDR[11:2]),
    .i1(10'b0000001010),
    .o(n176));  // ../RTL/cmsdk_iop_gpio.v(440)
  eq_w10 eq17 (
    .i0(IOADDR[11:2]),
    .i1(10'b0000001011),
    .o(n182));  // ../RTL/cmsdk_iop_gpio.v(446)
  eq_w10 eq18 (
    .i0(IOADDR[11:2]),
    .i1(10'b0000001100),
    .o(n221));  // ../RTL/cmsdk_iop_gpio.v(479)
  eq_w10 eq19 (
    .i0(IOADDR[11:2]),
    .i1(10'b0000001101),
    .o(n227));  // ../RTL/cmsdk_iop_gpio.v(485)
  eq_w4 eq2 (
    .i0(IOADDR[9:6]),
    .i1(4'b0000),
    .o(n7));  // ../RTL/cmsdk_iop_gpio.v(152)
  eq_w10 eq20 (
    .i0(IOADDR[11:2]),
    .i1(10'b0000001110),
    .o(n266));  // ../RTL/cmsdk_iop_gpio.v(520)
  eq_w4 eq3 (
    .i0(IOADDR[9:6]),
    .i1(4'b1111),
    .o(n12));  // ../RTL/cmsdk_iop_gpio.v(178)
  eq_w2 eq4 (
    .i0(IOSIZE),
    .i1(2'b10),
    .o(n15));  // ../RTL/cmsdk_iop_gpio.v(215)
  eq_w2 eq5 (
    .i0(IOSIZE),
    .i1(2'b01),
    .o(n17));  // ../RTL/cmsdk_iop_gpio.v(221)
  eq_w10 eq6 (
    .i0(IOADDR[11:2]),
    .i1(10'b0000000000),
    .o(n22));  // ../RTL/cmsdk_iop_gpio.v(271)
  eq_w10 eq7 (
    .i0(IOADDR[11:2]),
    .i1(10'b0000000001),
    .o(n23));  // ../RTL/cmsdk_iop_gpio.v(271)
  eq_w2 eq8 (
    .i0(IOADDR[11:10]),
    .i1(2'b01),
    .o(n26));  // ../RTL/cmsdk_iop_gpio.v(275)
  eq_w2 eq9 (
    .i0(IOADDR[11:10]),
    .i1(2'b10),
    .o(n28));  // ../RTL/cmsdk_iop_gpio.v(277)
  binary_mux_s4_w32 mux0 (
    .i0(reg_datain32),
    .i1({16'b0000000000000000,reg_dout}),
    .i10({16'b0000000000000000,reg_inttype}),
    .i11({16'b0000000000000000,reg_inttype}),
    .i12({16'b0000000000000000,reg_intpol}),
    .i13({16'b0000000000000000,reg_intpol}),
    .i14({16'b0000000000000000,reg_intstat}),
    .i15(32'b00000000000000000000000000000000),
    .i2(32'b00000000000000000000000000000000),
    .i3(32'b00000000000000000000000000000000),
    .i4({16'b0000000000000000,reg_douten}),
    .i5({16'b0000000000000000,reg_douten}),
    .i6({16'b0000000000000000,reg_altfunc}),
    .i7({16'b0000000000000000,reg_altfunc}),
    .i8({16'b0000000000000000,reg_inten}),
    .i9({16'b0000000000000000,reg_inten}),
    .sel(IOADDR[5:2]),
    .o(n8));  // ../RTL/cmsdk_iop_gpio.v(165)
  binary_mux_s1_w32 mux1 (
    .i0(32'b00000000000000000000000000000000),
    .i1(n8),
    .sel(n7),
    .o(n9));  // ../RTL/cmsdk_iop_gpio.v(167)
  binary_mux_s1_w8 mux10 (
    .i0(n33),
    .i1(IOWDATALE[7:0]),
    .sel(reg_dout_normal_write0),
    .o(nxt_dout_padded[7:0]));  // ../RTL/cmsdk_iop_gpio.v(286)
  binary_mux_s1_w8 mux11 (
    .i0(n38),
    .i1(IOWDATALE[15:8]),
    .sel(reg_dout_normal_write1),
    .o(nxt_dout_padded[15:8]));  // ../RTL/cmsdk_iop_gpio.v(301)
  binary_mux_s1_w8 mux12 (
    .i0(reg_dout_padded[7:0]),
    .i1(nxt_dout_padded[7:0]),
    .sel(n34),
    .o(n35));  // ../RTL/cmsdk_iop_gpio.v(294)
  binary_mux_s1_w8 mux13 (
    .i0(8'b00000000),
    .i1(IOWDATALE[7:0]),
    .sel(n43),
    .o(reg_doutenset[7:0]));  // ../RTL/cmsdk_iop_gpio.v(326)
  binary_mux_s1_w8 mux14 (
    .i0(8'b00000000),
    .i1(IOWDATALE[15:8]),
    .sel(n46),
    .o(reg_doutenset[15:8]));  // ../RTL/cmsdk_iop_gpio.v(329)
  binary_mux_s1_w8 mux15 (
    .i0(8'b00000000),
    .i1(IOWDATALE[7:0]),
    .sel(n49),
    .o(reg_doutenclr[7:0]));  // ../RTL/cmsdk_iop_gpio.v(332)
  binary_mux_s1_w8 mux16 (
    .i0(8'b00000000),
    .i1(IOWDATALE[15:8]),
    .sel(n52),
    .o(reg_doutenclr[15:8]));  // ../RTL/cmsdk_iop_gpio.v(335)
  binary_mux_s1_w8 mux17 (
    .i0(8'b00000000),
    .i1(IOWDATALE[7:0]),
    .sel(n88),
    .o(reg_altfuncset[7:0]));  // ../RTL/cmsdk_iop_gpio.v(365)
  binary_mux_s1_w8 mux18 (
    .i0(8'b00000000),
    .i1(IOWDATALE[15:8]),
    .sel(n91),
    .o(reg_altfuncset[15:8]));  // ../RTL/cmsdk_iop_gpio.v(368)
  binary_mux_s1_w8 mux19 (
    .i0(8'b00000000),
    .i1(IOWDATALE[7:0]),
    .sel(n94),
    .o(reg_altfuncclr[7:0]));  // ../RTL/cmsdk_iop_gpio.v(371)
  binary_mux_s4_w32 mux2 (
    .i0(32'b00000000000000000000000000000000),
    .i1(32'b00000000000000000000000000000000),
    .i10(32'b00000000000000000000000000011011),
    .i11({24'b000000000000000000000000,ECOREVNUM,4'b0000}),
    .i12(32'b00000000000000000000000000001101),
    .i13(32'b00000000000000000000000011110000),
    .i14(32'b00000000000000000000000000000101),
    .i15(32'b00000000000000000000000010110001),
    .i2(32'b00000000000000000000000000000000),
    .i3(32'b00000000000000000000000000000000),
    .i4(32'b00000000000000000000000000000100),
    .i5(32'b00000000000000000000000000000000),
    .i6(32'b00000000000000000000000000000000),
    .i7(32'b00000000000000000000000000000000),
    .i8(32'b00000000000000000000000000100000),
    .i9(32'b00000000000000000000000010111000),
    .sel(IOADDR[5:2]),
    .o(n13));  // ../RTL/cmsdk_iop_gpio.v(198)
  binary_mux_s1_w8 mux20 (
    .i0(8'b00000000),
    .i1(IOWDATALE[15:8]),
    .sel(n97),
    .o(reg_altfuncclr[15:8]));  // ../RTL/cmsdk_iop_gpio.v(374)
  binary_mux_s1_w8 mux21 (
    .i0(8'b00000000),
    .i1(IOWDATALE[7:0]),
    .sel(n133),
    .o(reg_intenset[7:0]));  // ../RTL/cmsdk_iop_gpio.v(403)
  binary_mux_s1_w8 mux22 (
    .i0(8'b00000000),
    .i1(IOWDATALE[15:8]),
    .sel(n136),
    .o(reg_intenset[15:8]));  // ../RTL/cmsdk_iop_gpio.v(406)
  binary_mux_s1_w8 mux23 (
    .i0(8'b00000000),
    .i1(IOWDATALE[7:0]),
    .sel(n139),
    .o(reg_intenclr[7:0]));  // ../RTL/cmsdk_iop_gpio.v(409)
  binary_mux_s1_w8 mux24 (
    .i0(8'b00000000),
    .i1(IOWDATALE[15:8]),
    .sel(n142),
    .o(reg_intenclr[15:8]));  // ../RTL/cmsdk_iop_gpio.v(412)
  binary_mux_s1_w8 mux25 (
    .i0(8'b00000000),
    .i1(IOWDATALE[7:0]),
    .sel(n178),
    .o(reg_inttypeset[7:0]));  // ../RTL/cmsdk_iop_gpio.v(441)
  binary_mux_s1_w8 mux26 (
    .i0(8'b00000000),
    .i1(IOWDATALE[15:8]),
    .sel(n181),
    .o(reg_inttypeset[15:8]));  // ../RTL/cmsdk_iop_gpio.v(444)
  binary_mux_s1_w8 mux27 (
    .i0(8'b00000000),
    .i1(IOWDATALE[7:0]),
    .sel(n184),
    .o(reg_inttypeclr[7:0]));  // ../RTL/cmsdk_iop_gpio.v(447)
  binary_mux_s1_w8 mux28 (
    .i0(8'b00000000),
    .i1(IOWDATALE[15:8]),
    .sel(n187),
    .o(reg_inttypeclr[15:8]));  // ../RTL/cmsdk_iop_gpio.v(450)
  binary_mux_s1_w8 mux29 (
    .i0(8'b00000000),
    .i1(IOWDATALE[7:0]),
    .sel(n223),
    .o(reg_intpolset[7:0]));  // ../RTL/cmsdk_iop_gpio.v(480)
  binary_mux_s1_w32 mux3 (
    .i0(32'b00000000000000000000000000000000),
    .i1(n13),
    .sel(n12),
    .o(n14));  // ../RTL/cmsdk_iop_gpio.v(204)
  binary_mux_s1_w8 mux30 (
    .i0(8'b00000000),
    .i1(IOWDATALE[15:8]),
    .sel(n226),
    .o(reg_intpolset[15:8]));  // ../RTL/cmsdk_iop_gpio.v(483)
  binary_mux_s1_w8 mux31 (
    .i0(8'b00000000),
    .i1(IOWDATALE[7:0]),
    .sel(n229),
    .o(reg_intpolclr[7:0]));  // ../RTL/cmsdk_iop_gpio.v(486)
  binary_mux_s1_w8 mux32 (
    .i0(8'b00000000),
    .i1(IOWDATALE[15:8]),
    .sel(n232),
    .o(reg_intpolclr[15:8]));  // ../RTL/cmsdk_iop_gpio.v(489)
  binary_mux_s1_w16 mux33 (
    .i0(reg_last_datain),
    .i1(reg_datain),
    .sel(n304),
    .o(n305));  // ../RTL/cmsdk_iop_gpio.v(561)
  binary_mux_s2_w32 mux4 (
    .i0(n9),
    .i1({24'b000000000000000000000000,n10}),
    .i2({16'b0000000000000000,n11,8'b00000000}),
    .i3(n14),
    .sel(IOADDR[11:10]),
    .o(read_mux_le));  // ../RTL/cmsdk_iop_gpio.v(209)
  binary_mux_s1_w32 mux5 (
    .i0(read_mux_le),
    .i1({read_mux_le[23:16],read_mux_le[31:24],read_mux_le[7:0],read_mux_le[15:8]}),
    .sel(n18),
    .o(n19));  // ../RTL/cmsdk_iop_gpio.v(231)
  binary_mux_s1_w32 mux6 (
    .i0(IOWDATA),
    .i1({IOWDATA[23:16],IOWDATA[31:24],IOWDATA[7:0],IOWDATA[15:8]}),
    .sel(n18),
    .o(n20));  // ../RTL/cmsdk_iop_gpio.v(231)
  binary_mux_s1_w32 mux7 (
    .i0(n19),
    .i1({read_mux_le[7:0],read_mux_le[15:8],read_mux_le[23:16],read_mux_le[31:24]}),
    .sel(n16),
    .o(read_mux));  // ../RTL/cmsdk_iop_gpio.v(231)
  binary_mux_s1_w32 mux8 (
    .i0(n20),
    .i1({IOWDATA[7:0],IOWDATA[15:8],IOWDATA[23:16],IOWDATA[31:24]}),
    .sel(n16),
    .o({open_n0,open_n1,open_n2,open_n3,open_n4,open_n5,open_n6,open_n7,open_n8,open_n9,open_n10,open_n11,open_n12,open_n13,open_n14,open_n15,IOWDATALE[15:0]}));  // ../RTL/cmsdk_iop_gpio.v(231)
  binary_mux_s1_w8 mux9 (
    .i0(reg_dout_padded[15:8]),
    .i1(nxt_dout_padded[15:8]),
    .sel(n39),
    .o(n40));  // ../RTL/cmsdk_iop_gpio.v(309)
  reg_ar_as_w16 reg0 (
    .clk(FCLK),
    .d(reg_in_sync1),
    .reset({n21,n21,n21,n21,n21,n21,n21,n21,n21,n21,n21,n21,n21,n21,n21,n21}),
    .set(16'b0000000000000000),
    .q(reg_in_sync2));  // ../RTL/cmsdk_iop_gpio.v(252)
  reg_ar_as_w16 reg1 (
    .clk(HCLK),
    .d({n40,n35}),
    .reset({n21,n21,n21,n21,n21,n21,n21,n21,n21,n21,n21,n21,n21,n21,n21,n21}),
    .set(16'b0000000000000000),
    .q(reg_dout_padded));  // ../RTL/cmsdk_iop_gpio.v(309)
  reg_ar_as_w16 reg2 (
    .clk(HCLK),
    .d({n85,n83,n81,n79,n77,n75,n73,n71,n69,n67,n65,n63,n61,n59,n57,n55}),
    .reset({n21,n21,n21,n21,n21,n21,n21,n21,n21,n21,n21,n21,n21,n21,n21,n21}),
    .set(16'b0000000000000000),
    .q(reg_douten_padded));  // ../RTL/cmsdk_iop_gpio.v(348)
  reg_ar_as_w16 reg3 (
    .clk(HCLK),
    .d({n130,n128,n126,n124,n122,n120,n118,n116,n114,n112,n110,n108,n106,n104,n102,n100}),
    .reset({n21,n21,n21,n21,n21,n21,n21,n21,n21,n21,n21,n21,n21,n21,n21,n21}),
    .set(16'b0000000000000000),
    .q(reg_altfunc_padded));  // ../RTL/cmsdk_iop_gpio.v(387)
  reg_ar_as_w16 reg4 (
    .clk(HCLK),
    .d({n175,n173,n171,n169,n167,n165,n163,n161,n159,n157,n155,n153,n151,n149,n147,n145}),
    .reset({n21,n21,n21,n21,n21,n21,n21,n21,n21,n21,n21,n21,n21,n21,n21,n21}),
    .set(16'b0000000000000000),
    .q(reg_inten_padded));  // ../RTL/cmsdk_iop_gpio.v(425)
  reg_ar_as_w16 reg5 (
    .clk(HCLK),
    .d({n220,n218,n216,n214,n212,n210,n208,n206,n204,n202,n200,n198,n196,n194,n192,n190}),
    .reset({n21,n21,n21,n21,n21,n21,n21,n21,n21,n21,n21,n21,n21,n21,n21,n21}),
    .set(16'b0000000000000000),
    .q(reg_inttype_padded));  // ../RTL/cmsdk_iop_gpio.v(463)
  reg_ar_as_w16 reg6 (
    .clk(HCLK),
    .d({n265,n263,n261,n259,n257,n255,n253,n251,n249,n247,n245,n243,n241,n239,n237,n235}),
    .reset({n21,n21,n21,n21,n21,n21,n21,n21,n21,n21,n21,n21,n21,n21,n21,n21}),
    .set(16'b0000000000000000),
    .q(reg_intpol_padded));  // ../RTL/cmsdk_iop_gpio.v(501)
  reg_ar_as_w16 reg7 (
    .clk(FCLK),
    .d({n302,n300,n298,n296,n294,n292,n290,n288,n286,n284,n282,n280,n278,n276,n274,n272}),
    .reset({n21,n21,n21,n21,n21,n21,n21,n21,n21,n21,n21,n21,n21,n21,n21,n21}),
    .set(16'b0000000000000000),
    .q(reg_intstat_padded));  // ../RTL/cmsdk_iop_gpio.v(539)
  reg_ar_as_w16 reg8 (
    .clk(FCLK),
    .d(n305),
    .reset({n21,n21,n21,n21,n21,n21,n21,n21,n21,n21,n21,n21,n21,n21,n21,n21}),
    .set(16'b0000000000000000),
    .q(reg_last_datain));  // ../RTL/cmsdk_iop_gpio.v(561)
  reg_ar_as_w16 reg9 (
    .clk(FCLK),
    .d(PORTIN),
    .reset({n21,n21,n21,n21,n21,n21,n21,n21,n21,n21,n21,n21,n21,n21,n21,n21}),
    .set(16'b0000000000000000),
    .q(reg_in_sync1));  // ../RTL/cmsdk_iop_gpio.v(252)
  or u10 (n335[6], n334[6], rise_edge_int[6]);  // ../RTL/cmsdk_iop_gpio.v(568)
  buf u100 (GPIOINT[11], reg_intstat[11]);  // ../RTL/cmsdk_iop_gpio.v(580)
  or u101 (n54, reg_doutenset[0], reg_doutenclr[0]);  // ../RTL/cmsdk_iop_gpio.v(346)
  AL_MUX u102 (
    .i0(reg_douten_padded[0]),
    .i1(reg_doutenset[0]),
    .sel(n54),
    .o(n55));  // ../RTL/cmsdk_iop_gpio.v(347)
  or u103 (n56, reg_doutenset[1], reg_doutenclr[1]);  // ../RTL/cmsdk_iop_gpio.v(346)
  AL_MUX u104 (
    .i0(reg_douten_padded[1]),
    .i1(reg_doutenset[1]),
    .sel(n56),
    .o(n57));  // ../RTL/cmsdk_iop_gpio.v(347)
  or u105 (n58, reg_doutenset[2], reg_doutenclr[2]);  // ../RTL/cmsdk_iop_gpio.v(346)
  AL_MUX u106 (
    .i0(reg_douten_padded[2]),
    .i1(reg_doutenset[2]),
    .sel(n58),
    .o(n59));  // ../RTL/cmsdk_iop_gpio.v(347)
  or u107 (n60, reg_doutenset[3], reg_doutenclr[3]);  // ../RTL/cmsdk_iop_gpio.v(346)
  AL_MUX u108 (
    .i0(reg_douten_padded[3]),
    .i1(reg_doutenset[3]),
    .sel(n60),
    .o(n61));  // ../RTL/cmsdk_iop_gpio.v(347)
  or u109 (n62, reg_doutenset[4], reg_doutenclr[4]);  // ../RTL/cmsdk_iop_gpio.v(346)
  or u11 (n335[7], n334[7], rise_edge_int[7]);  // ../RTL/cmsdk_iop_gpio.v(568)
  AL_MUX u110 (
    .i0(reg_douten_padded[4]),
    .i1(reg_doutenset[4]),
    .sel(n62),
    .o(n63));  // ../RTL/cmsdk_iop_gpio.v(347)
  or u111 (n64, reg_doutenset[5], reg_doutenclr[5]);  // ../RTL/cmsdk_iop_gpio.v(346)
  AL_MUX u112 (
    .i0(reg_douten_padded[5]),
    .i1(reg_doutenset[5]),
    .sel(n64),
    .o(n65));  // ../RTL/cmsdk_iop_gpio.v(347)
  or u113 (n66, reg_doutenset[6], reg_doutenclr[6]);  // ../RTL/cmsdk_iop_gpio.v(346)
  AL_MUX u114 (
    .i0(reg_douten_padded[6]),
    .i1(reg_doutenset[6]),
    .sel(n66),
    .o(n67));  // ../RTL/cmsdk_iop_gpio.v(347)
  or u115 (n68, reg_doutenset[7], reg_doutenclr[7]);  // ../RTL/cmsdk_iop_gpio.v(346)
  AL_MUX u116 (
    .i0(reg_douten_padded[7]),
    .i1(reg_doutenset[7]),
    .sel(n68),
    .o(n69));  // ../RTL/cmsdk_iop_gpio.v(347)
  or u117 (n70, reg_doutenset[8], reg_doutenclr[8]);  // ../RTL/cmsdk_iop_gpio.v(346)
  AL_MUX u118 (
    .i0(reg_douten_padded[8]),
    .i1(reg_doutenset[8]),
    .sel(n70),
    .o(n71));  // ../RTL/cmsdk_iop_gpio.v(347)
  or u119 (n72, reg_doutenset[9], reg_doutenclr[9]);  // ../RTL/cmsdk_iop_gpio.v(346)
  and u12 (n37[0], current_dout_padded[8], n31[0]);  // ../RTL/cmsdk_iop_gpio.v(301)
  AL_MUX u120 (
    .i0(reg_douten_padded[9]),
    .i1(reg_doutenset[9]),
    .sel(n72),
    .o(n73));  // ../RTL/cmsdk_iop_gpio.v(347)
  or u121 (n74, reg_doutenset[10], reg_doutenclr[10]);  // ../RTL/cmsdk_iop_gpio.v(346)
  AL_MUX u122 (
    .i0(reg_douten_padded[10]),
    .i1(reg_doutenset[10]),
    .sel(n74),
    .o(n75));  // ../RTL/cmsdk_iop_gpio.v(347)
  or u123 (n76, reg_doutenset[11], reg_doutenclr[11]);  // ../RTL/cmsdk_iop_gpio.v(346)
  AL_MUX u124 (
    .i0(reg_douten_padded[11]),
    .i1(reg_doutenset[11]),
    .sel(n76),
    .o(n77));  // ../RTL/cmsdk_iop_gpio.v(347)
  or u125 (n78, reg_doutenset[12], reg_doutenclr[12]);  // ../RTL/cmsdk_iop_gpio.v(346)
  AL_MUX u126 (
    .i0(reg_douten_padded[12]),
    .i1(reg_doutenset[12]),
    .sel(n78),
    .o(n79));  // ../RTL/cmsdk_iop_gpio.v(347)
  or u127 (n80, reg_doutenset[13], reg_doutenclr[13]);  // ../RTL/cmsdk_iop_gpio.v(346)
  AL_MUX u128 (
    .i0(reg_douten_padded[13]),
    .i1(reg_doutenset[13]),
    .sel(n80),
    .o(n81));  // ../RTL/cmsdk_iop_gpio.v(347)
  or u129 (n82, reg_doutenset[14], reg_doutenclr[14]);  // ../RTL/cmsdk_iop_gpio.v(346)
  and u13 (n4[1], n3[1], IOSIZE[0]);  // ../RTL/cmsdk_iop_gpio.v(143)
  AL_MUX u130 (
    .i0(reg_douten_padded[14]),
    .i1(reg_doutenset[14]),
    .sel(n82),
    .o(n83));  // ../RTL/cmsdk_iop_gpio.v(347)
  or u131 (n84, reg_doutenset[15], reg_doutenclr[15]);  // ../RTL/cmsdk_iop_gpio.v(346)
  AL_MUX u132 (
    .i0(reg_douten_padded[15]),
    .i1(reg_doutenset[15]),
    .sel(n84),
    .o(n85));  // ../RTL/cmsdk_iop_gpio.v(347)
  buf u133 (reg_dout[0], reg_dout_padded[0]);  // ../RTL/cmsdk_iop_gpio.v(312)
  buf u134 (PORTFUNC[14], reg_altfunc[14]);  // ../RTL/cmsdk_iop_gpio.v(575)
  and u135 (n87, write_trans, n86);  // ../RTL/cmsdk_iop_gpio.v(364)
  buf u136 (PORTFUNC[13], reg_altfunc[13]);  // ../RTL/cmsdk_iop_gpio.v(575)
  and u137 (n88, n87, iop_byte_strobe[0]);  // ../RTL/cmsdk_iop_gpio.v(365)
  buf u138 (PORTFUNC[12], reg_altfunc[12]);  // ../RTL/cmsdk_iop_gpio.v(575)
  buf u139 (GPIOINT[10], reg_intstat[10]);  // ../RTL/cmsdk_iop_gpio.v(580)
  buf u14 (IORDATA[8], read_mux[8]);  // ../RTL/cmsdk_iop_gpio.v(577)
  buf u140 (GPIOINT[9], reg_intstat[9]);  // ../RTL/cmsdk_iop_gpio.v(580)
  buf u141 (PORTFUNC[11], reg_altfunc[11]);  // ../RTL/cmsdk_iop_gpio.v(575)
  and u142 (n91, n87, iop_byte_strobe[1]);  // ../RTL/cmsdk_iop_gpio.v(368)
  buf u143 (PORTFUNC[10], reg_altfunc[10]);  // ../RTL/cmsdk_iop_gpio.v(575)
  and u144 (n93, write_trans, n92);  // ../RTL/cmsdk_iop_gpio.v(370)
  buf u145 (PORTFUNC[9], reg_altfunc[9]);  // ../RTL/cmsdk_iop_gpio.v(575)
  and u146 (n94, n93, iop_byte_strobe[0]);  // ../RTL/cmsdk_iop_gpio.v(371)
  buf u147 (PORTFUNC[8], reg_altfunc[8]);  // ../RTL/cmsdk_iop_gpio.v(575)
  buf u148 (GPIOINT[8], reg_intstat[8]);  // ../RTL/cmsdk_iop_gpio.v(580)
  buf u149 (GPIOINT[7], reg_intstat[7]);  // ../RTL/cmsdk_iop_gpio.v(580)
  or u15 (n5[1], IOSIZE[1], n4[1]);  // ../RTL/cmsdk_iop_gpio.v(143)
  buf u150 (PORTFUNC[7], reg_altfunc[7]);  // ../RTL/cmsdk_iop_gpio.v(575)
  and u151 (n97, n93, iop_byte_strobe[1]);  // ../RTL/cmsdk_iop_gpio.v(374)
  buf u152 (PORTFUNC[6], reg_altfunc[6]);  // ../RTL/cmsdk_iop_gpio.v(575)
  buf u153 (GPIOINT[6], reg_intstat[6]);  // ../RTL/cmsdk_iop_gpio.v(580)
  or u154 (n99, reg_altfuncset[0], reg_altfuncclr[0]);  // ../RTL/cmsdk_iop_gpio.v(385)
  AL_MUX u155 (
    .i0(reg_altfunc_padded[0]),
    .i1(reg_altfuncset[0]),
    .sel(n99),
    .o(n100));  // ../RTL/cmsdk_iop_gpio.v(386)
  or u156 (n101, reg_altfuncset[1], reg_altfuncclr[1]);  // ../RTL/cmsdk_iop_gpio.v(385)
  AL_MUX u157 (
    .i0(reg_altfunc_padded[1]),
    .i1(reg_altfuncset[1]),
    .sel(n101),
    .o(n102));  // ../RTL/cmsdk_iop_gpio.v(386)
  or u158 (n103, reg_altfuncset[2], reg_altfuncclr[2]);  // ../RTL/cmsdk_iop_gpio.v(385)
  AL_MUX u159 (
    .i0(reg_altfunc_padded[2]),
    .i1(reg_altfuncset[2]),
    .sel(n103),
    .o(n104));  // ../RTL/cmsdk_iop_gpio.v(386)
  or u16 (n335[8], n334[8], rise_edge_int[8]);  // ../RTL/cmsdk_iop_gpio.v(568)
  or u160 (n105, reg_altfuncset[3], reg_altfuncclr[3]);  // ../RTL/cmsdk_iop_gpio.v(385)
  AL_MUX u161 (
    .i0(reg_altfunc_padded[3]),
    .i1(reg_altfuncset[3]),
    .sel(n105),
    .o(n106));  // ../RTL/cmsdk_iop_gpio.v(386)
  or u162 (n107, reg_altfuncset[4], reg_altfuncclr[4]);  // ../RTL/cmsdk_iop_gpio.v(385)
  AL_MUX u163 (
    .i0(reg_altfunc_padded[4]),
    .i1(reg_altfuncset[4]),
    .sel(n107),
    .o(n108));  // ../RTL/cmsdk_iop_gpio.v(386)
  or u164 (n109, reg_altfuncset[5], reg_altfuncclr[5]);  // ../RTL/cmsdk_iop_gpio.v(385)
  AL_MUX u165 (
    .i0(reg_altfunc_padded[5]),
    .i1(reg_altfuncset[5]),
    .sel(n109),
    .o(n110));  // ../RTL/cmsdk_iop_gpio.v(386)
  or u166 (n111, reg_altfuncset[6], reg_altfuncclr[6]);  // ../RTL/cmsdk_iop_gpio.v(385)
  AL_MUX u167 (
    .i0(reg_altfunc_padded[6]),
    .i1(reg_altfuncset[6]),
    .sel(n111),
    .o(n112));  // ../RTL/cmsdk_iop_gpio.v(386)
  or u168 (n113, reg_altfuncset[7], reg_altfuncclr[7]);  // ../RTL/cmsdk_iop_gpio.v(385)
  AL_MUX u169 (
    .i0(reg_altfunc_padded[7]),
    .i1(reg_altfuncset[7]),
    .sel(n113),
    .o(n114));  // ../RTL/cmsdk_iop_gpio.v(386)
  or u17 (n2[0], n5[1], n1);  // ../RTL/cmsdk_iop_gpio.v(143)
  or u170 (n115, reg_altfuncset[8], reg_altfuncclr[8]);  // ../RTL/cmsdk_iop_gpio.v(385)
  AL_MUX u171 (
    .i0(reg_altfunc_padded[8]),
    .i1(reg_altfuncset[8]),
    .sel(n115),
    .o(n116));  // ../RTL/cmsdk_iop_gpio.v(386)
  or u172 (n117, reg_altfuncset[9], reg_altfuncclr[9]);  // ../RTL/cmsdk_iop_gpio.v(385)
  AL_MUX u173 (
    .i0(reg_altfunc_padded[9]),
    .i1(reg_altfuncset[9]),
    .sel(n117),
    .o(n118));  // ../RTL/cmsdk_iop_gpio.v(386)
  or u174 (n119, reg_altfuncset[10], reg_altfuncclr[10]);  // ../RTL/cmsdk_iop_gpio.v(385)
  AL_MUX u175 (
    .i0(reg_altfunc_padded[10]),
    .i1(reg_altfuncset[10]),
    .sel(n119),
    .o(n120));  // ../RTL/cmsdk_iop_gpio.v(386)
  or u176 (n121, reg_altfuncset[11], reg_altfuncclr[11]);  // ../RTL/cmsdk_iop_gpio.v(385)
  AL_MUX u177 (
    .i0(reg_altfunc_padded[11]),
    .i1(reg_altfuncset[11]),
    .sel(n121),
    .o(n122));  // ../RTL/cmsdk_iop_gpio.v(386)
  or u178 (n123, reg_altfuncset[12], reg_altfuncclr[12]);  // ../RTL/cmsdk_iop_gpio.v(385)
  AL_MUX u179 (
    .i0(reg_altfunc_padded[12]),
    .i1(reg_altfuncset[12]),
    .sel(n123),
    .o(n124));  // ../RTL/cmsdk_iop_gpio.v(386)
  and u18 (n16, bigendian, n15);  // ../RTL/cmsdk_iop_gpio.v(215)
  or u180 (n125, reg_altfuncset[13], reg_altfuncclr[13]);  // ../RTL/cmsdk_iop_gpio.v(385)
  AL_MUX u181 (
    .i0(reg_altfunc_padded[13]),
    .i1(reg_altfuncset[13]),
    .sel(n125),
    .o(n126));  // ../RTL/cmsdk_iop_gpio.v(386)
  or u182 (n127, reg_altfuncset[14], reg_altfuncclr[14]);  // ../RTL/cmsdk_iop_gpio.v(385)
  AL_MUX u183 (
    .i0(reg_altfunc_padded[14]),
    .i1(reg_altfuncset[14]),
    .sel(n127),
    .o(n128));  // ../RTL/cmsdk_iop_gpio.v(386)
  or u184 (n129, reg_altfuncset[15], reg_altfuncclr[15]);  // ../RTL/cmsdk_iop_gpio.v(385)
  AL_MUX u185 (
    .i0(reg_altfunc_padded[15]),
    .i1(reg_altfuncset[15]),
    .sel(n129),
    .o(n130));  // ../RTL/cmsdk_iop_gpio.v(386)
  buf u186 (reg_douten[0], reg_douten_padded[0]);  // ../RTL/cmsdk_iop_gpio.v(351)
  buf u187 (PORTFUNC[5], reg_altfunc[5]);  // ../RTL/cmsdk_iop_gpio.v(575)
  and u188 (n132, write_trans, n131);  // ../RTL/cmsdk_iop_gpio.v(402)
  buf u189 (PORTFUNC[4], reg_altfunc[4]);  // ../RTL/cmsdk_iop_gpio.v(575)
  and u19 (n18, bigendian, n17);  // ../RTL/cmsdk_iop_gpio.v(221)
  and u190 (n133, n132, iop_byte_strobe[0]);  // ../RTL/cmsdk_iop_gpio.v(403)
  buf u191 (PORTFUNC[3], reg_altfunc[3]);  // ../RTL/cmsdk_iop_gpio.v(575)
  buf u192 (GPIOINT[5], reg_intstat[5]);  // ../RTL/cmsdk_iop_gpio.v(580)
  buf u193 (GPIOINT[4], reg_intstat[4]);  // ../RTL/cmsdk_iop_gpio.v(580)
  buf u194 (PORTFUNC[2], reg_altfunc[2]);  // ../RTL/cmsdk_iop_gpio.v(575)
  and u195 (n136, n132, iop_byte_strobe[1]);  // ../RTL/cmsdk_iop_gpio.v(406)
  buf u196 (PORTFUNC[1], reg_altfunc[1]);  // ../RTL/cmsdk_iop_gpio.v(575)
  and u197 (n138, write_trans, n137);  // ../RTL/cmsdk_iop_gpio.v(408)
  buf u198 (IORDATA[31], read_mux[31]);  // ../RTL/cmsdk_iop_gpio.v(577)
  and u199 (n139, n138, iop_byte_strobe[0]);  // ../RTL/cmsdk_iop_gpio.v(409)
  buf u2 (PORTEN[13], reg_douten[13]);  // ../RTL/cmsdk_iop_gpio.v(574)
  buf u20 (PORTEN[11], reg_douten[11]);  // ../RTL/cmsdk_iop_gpio.v(574)
  buf u200 (IORDATA[30], read_mux[30]);  // ../RTL/cmsdk_iop_gpio.v(577)
  buf u201 (GPIOINT[3], reg_intstat[3]);  // ../RTL/cmsdk_iop_gpio.v(580)
  buf u202 (GPIOINT[2], reg_intstat[2]);  // ../RTL/cmsdk_iop_gpio.v(580)
  buf u203 (IORDATA[29], read_mux[29]);  // ../RTL/cmsdk_iop_gpio.v(577)
  and u204 (n142, n138, iop_byte_strobe[1]);  // ../RTL/cmsdk_iop_gpio.v(412)
  buf u205 (IORDATA[28], read_mux[28]);  // ../RTL/cmsdk_iop_gpio.v(577)
  buf u206 (GPIOINT[1], reg_intstat[1]);  // ../RTL/cmsdk_iop_gpio.v(580)
  or u207 (n144, reg_intenclr[0], reg_intenset[0]);  // ../RTL/cmsdk_iop_gpio.v(423)
  AL_MUX u208 (
    .i0(reg_inten_padded[0]),
    .i1(reg_intenset[0]),
    .sel(n144),
    .o(n145));  // ../RTL/cmsdk_iop_gpio.v(424)
  or u209 (n146, reg_intenclr[1], reg_intenset[1]);  // ../RTL/cmsdk_iop_gpio.v(423)
  not u21 (n21, HRESETn);  // ../RTL/cmsdk_iop_gpio.v(243)
  AL_MUX u210 (
    .i0(reg_inten_padded[1]),
    .i1(reg_intenset[1]),
    .sel(n146),
    .o(n147));  // ../RTL/cmsdk_iop_gpio.v(424)
  or u211 (n148, reg_intenclr[2], reg_intenset[2]);  // ../RTL/cmsdk_iop_gpio.v(423)
  AL_MUX u212 (
    .i0(reg_inten_padded[2]),
    .i1(reg_intenset[2]),
    .sel(n148),
    .o(n149));  // ../RTL/cmsdk_iop_gpio.v(424)
  or u213 (n150, reg_intenclr[3], reg_intenset[3]);  // ../RTL/cmsdk_iop_gpio.v(423)
  AL_MUX u214 (
    .i0(reg_inten_padded[3]),
    .i1(reg_intenset[3]),
    .sel(n150),
    .o(n151));  // ../RTL/cmsdk_iop_gpio.v(424)
  or u215 (n152, reg_intenclr[4], reg_intenset[4]);  // ../RTL/cmsdk_iop_gpio.v(423)
  AL_MUX u216 (
    .i0(reg_inten_padded[4]),
    .i1(reg_intenset[4]),
    .sel(n152),
    .o(n153));  // ../RTL/cmsdk_iop_gpio.v(424)
  or u217 (n154, reg_intenclr[5], reg_intenset[5]);  // ../RTL/cmsdk_iop_gpio.v(423)
  AL_MUX u218 (
    .i0(reg_inten_padded[5]),
    .i1(reg_intenset[5]),
    .sel(n154),
    .o(n155));  // ../RTL/cmsdk_iop_gpio.v(424)
  or u219 (n156, reg_intenclr[6], reg_intenset[6]);  // ../RTL/cmsdk_iop_gpio.v(423)
  buf u22 (PORTOUT[9], reg_dout[9]);  // ../RTL/cmsdk_iop_gpio.v(573)
  AL_MUX u220 (
    .i0(reg_inten_padded[6]),
    .i1(reg_intenset[6]),
    .sel(n156),
    .o(n157));  // ../RTL/cmsdk_iop_gpio.v(424)
  or u221 (n158, reg_intenclr[7], reg_intenset[7]);  // ../RTL/cmsdk_iop_gpio.v(423)
  AL_MUX u222 (
    .i0(reg_inten_padded[7]),
    .i1(reg_intenset[7]),
    .sel(n158),
    .o(n159));  // ../RTL/cmsdk_iop_gpio.v(424)
  or u223 (n160, reg_intenclr[8], reg_intenset[8]);  // ../RTL/cmsdk_iop_gpio.v(423)
  AL_MUX u224 (
    .i0(reg_inten_padded[8]),
    .i1(reg_intenset[8]),
    .sel(n160),
    .o(n161));  // ../RTL/cmsdk_iop_gpio.v(424)
  or u225 (n162, reg_intenclr[9], reg_intenset[9]);  // ../RTL/cmsdk_iop_gpio.v(423)
  AL_MUX u226 (
    .i0(reg_inten_padded[9]),
    .i1(reg_intenset[9]),
    .sel(n162),
    .o(n163));  // ../RTL/cmsdk_iop_gpio.v(424)
  or u227 (n164, reg_intenclr[10], reg_intenset[10]);  // ../RTL/cmsdk_iop_gpio.v(423)
  AL_MUX u228 (
    .i0(reg_inten_padded[10]),
    .i1(reg_intenset[10]),
    .sel(n164),
    .o(n165));  // ../RTL/cmsdk_iop_gpio.v(424)
  or u229 (n166, reg_intenclr[11], reg_intenset[11]);  // ../RTL/cmsdk_iop_gpio.v(423)
  and u23 (iop_byte_strobe[0], n2[0], IOSEL);  // ../RTL/cmsdk_iop_gpio.v(143)
  AL_MUX u230 (
    .i0(reg_inten_padded[11]),
    .i1(reg_intenset[11]),
    .sel(n166),
    .o(n167));  // ../RTL/cmsdk_iop_gpio.v(424)
  or u231 (n168, reg_intenclr[12], reg_intenset[12]);  // ../RTL/cmsdk_iop_gpio.v(423)
  AL_MUX u232 (
    .i0(reg_inten_padded[12]),
    .i1(reg_intenset[12]),
    .sel(n168),
    .o(n169));  // ../RTL/cmsdk_iop_gpio.v(424)
  or u233 (n170, reg_intenclr[13], reg_intenset[13]);  // ../RTL/cmsdk_iop_gpio.v(423)
  AL_MUX u234 (
    .i0(reg_inten_padded[13]),
    .i1(reg_intenset[13]),
    .sel(n170),
    .o(n171));  // ../RTL/cmsdk_iop_gpio.v(424)
  or u235 (n172, reg_intenclr[14], reg_intenset[14]);  // ../RTL/cmsdk_iop_gpio.v(423)
  AL_MUX u236 (
    .i0(reg_inten_padded[14]),
    .i1(reg_intenset[14]),
    .sel(n172),
    .o(n173));  // ../RTL/cmsdk_iop_gpio.v(424)
  or u237 (n174, reg_intenclr[15], reg_intenset[15]);  // ../RTL/cmsdk_iop_gpio.v(423)
  AL_MUX u238 (
    .i0(reg_inten_padded[15]),
    .i1(reg_intenset[15]),
    .sel(n174),
    .o(n175));  // ../RTL/cmsdk_iop_gpio.v(424)
  buf u239 (reg_altfunc[0], reg_altfunc_padded[0]);  // ../RTL/cmsdk_iop_gpio.v(390)
  buf u24 (reg_datain[0], reg_in_sync2[0]);  // ../RTL/cmsdk_iop_gpio.v(255)
  buf u240 (IORDATA[27], read_mux[27]);  // ../RTL/cmsdk_iop_gpio.v(577)
  and u241 (n177, write_trans, n176);  // ../RTL/cmsdk_iop_gpio.v(440)
  buf u242 (IORDATA[26], read_mux[26]);  // ../RTL/cmsdk_iop_gpio.v(577)
  and u243 (n178, n177, iop_byte_strobe[0]);  // ../RTL/cmsdk_iop_gpio.v(441)
  buf u244 (IORDATA[25], read_mux[25]);  // ../RTL/cmsdk_iop_gpio.v(577)
  or u245 (COMBINT, n320, n313);  // ../RTL/cmsdk_iop_gpio.v(581)
  or u246 (n313, n317, n314);  // ../RTL/cmsdk_iop_gpio.v(581)
  buf u247 (IORDATA[24], read_mux[24]);  // ../RTL/cmsdk_iop_gpio.v(577)
  and u248 (n181, n177, iop_byte_strobe[1]);  // ../RTL/cmsdk_iop_gpio.v(444)
  buf u249 (IORDATA[23], read_mux[23]);  // ../RTL/cmsdk_iop_gpio.v(577)
  or u25 (n24, n22, n23);  // ../RTL/cmsdk_iop_gpio.v(271)
  and u250 (n183, write_trans, n182);  // ../RTL/cmsdk_iop_gpio.v(446)
  buf u251 (IORDATA[22], read_mux[22]);  // ../RTL/cmsdk_iop_gpio.v(577)
  and u252 (n184, n183, iop_byte_strobe[0]);  // ../RTL/cmsdk_iop_gpio.v(447)
  buf u253 (IORDATA[21], read_mux[21]);  // ../RTL/cmsdk_iop_gpio.v(577)
  or u254 (n314, n316, n315);  // ../RTL/cmsdk_iop_gpio.v(581)
  or u255 (n315, reg_intstat[14], reg_intstat[15]);  // ../RTL/cmsdk_iop_gpio.v(581)
  buf u256 (IORDATA[20], read_mux[20]);  // ../RTL/cmsdk_iop_gpio.v(577)
  and u257 (n187, n183, iop_byte_strobe[1]);  // ../RTL/cmsdk_iop_gpio.v(450)
  buf u258 (IORDATA[19], read_mux[19]);  // ../RTL/cmsdk_iop_gpio.v(577)
  or u259 (n316, reg_intstat[12], reg_intstat[13]);  // ../RTL/cmsdk_iop_gpio.v(581)
  and u26 (n25, write_trans, n24);  // ../RTL/cmsdk_iop_gpio.v(271)
  or u260 (n189, reg_inttypeset[0], reg_inttypeclr[0]);  // ../RTL/cmsdk_iop_gpio.v(461)
  AL_MUX u261 (
    .i0(reg_inttype_padded[0]),
    .i1(reg_inttypeset[0]),
    .sel(n189),
    .o(n190));  // ../RTL/cmsdk_iop_gpio.v(462)
  or u262 (n191, reg_inttypeset[1], reg_inttypeclr[1]);  // ../RTL/cmsdk_iop_gpio.v(461)
  AL_MUX u263 (
    .i0(reg_inttype_padded[1]),
    .i1(reg_inttypeset[1]),
    .sel(n191),
    .o(n192));  // ../RTL/cmsdk_iop_gpio.v(462)
  or u264 (n193, reg_inttypeset[2], reg_inttypeclr[2]);  // ../RTL/cmsdk_iop_gpio.v(461)
  AL_MUX u265 (
    .i0(reg_inttype_padded[2]),
    .i1(reg_inttypeset[2]),
    .sel(n193),
    .o(n194));  // ../RTL/cmsdk_iop_gpio.v(462)
  or u266 (n195, reg_inttypeset[3], reg_inttypeclr[3]);  // ../RTL/cmsdk_iop_gpio.v(461)
  AL_MUX u267 (
    .i0(reg_inttype_padded[3]),
    .i1(reg_inttypeset[3]),
    .sel(n195),
    .o(n196));  // ../RTL/cmsdk_iop_gpio.v(462)
  or u268 (n197, reg_inttypeset[4], reg_inttypeclr[4]);  // ../RTL/cmsdk_iop_gpio.v(461)
  AL_MUX u269 (
    .i0(reg_inttype_padded[4]),
    .i1(reg_inttypeset[4]),
    .sel(n197),
    .o(n198));  // ../RTL/cmsdk_iop_gpio.v(462)
  and u27 (reg_dout_normal_write0, n25, iop_byte_strobe[0]);  // ../RTL/cmsdk_iop_gpio.v(271)
  or u270 (n199, reg_inttypeset[5], reg_inttypeclr[5]);  // ../RTL/cmsdk_iop_gpio.v(461)
  AL_MUX u271 (
    .i0(reg_inttype_padded[5]),
    .i1(reg_inttypeset[5]),
    .sel(n199),
    .o(n200));  // ../RTL/cmsdk_iop_gpio.v(462)
  or u272 (n201, reg_inttypeset[6], reg_inttypeclr[6]);  // ../RTL/cmsdk_iop_gpio.v(461)
  AL_MUX u273 (
    .i0(reg_inttype_padded[6]),
    .i1(reg_inttypeset[6]),
    .sel(n201),
    .o(n202));  // ../RTL/cmsdk_iop_gpio.v(462)
  or u274 (n203, reg_inttypeset[7], reg_inttypeclr[7]);  // ../RTL/cmsdk_iop_gpio.v(461)
  AL_MUX u275 (
    .i0(reg_inttype_padded[7]),
    .i1(reg_inttypeset[7]),
    .sel(n203),
    .o(n204));  // ../RTL/cmsdk_iop_gpio.v(462)
  or u276 (n205, reg_inttypeset[8], reg_inttypeclr[8]);  // ../RTL/cmsdk_iop_gpio.v(461)
  AL_MUX u277 (
    .i0(reg_inttype_padded[8]),
    .i1(reg_inttypeset[8]),
    .sel(n205),
    .o(n206));  // ../RTL/cmsdk_iop_gpio.v(462)
  or u278 (n207, reg_inttypeset[9], reg_inttypeclr[9]);  // ../RTL/cmsdk_iop_gpio.v(461)
  AL_MUX u279 (
    .i0(reg_inttype_padded[9]),
    .i1(reg_inttypeset[9]),
    .sel(n207),
    .o(n208));  // ../RTL/cmsdk_iop_gpio.v(462)
  buf u28 (IORDATA[7], read_mux[7]);  // ../RTL/cmsdk_iop_gpio.v(577)
  or u280 (n209, reg_inttypeset[10], reg_inttypeclr[10]);  // ../RTL/cmsdk_iop_gpio.v(461)
  AL_MUX u281 (
    .i0(reg_inttype_padded[10]),
    .i1(reg_inttypeset[10]),
    .sel(n209),
    .o(n210));  // ../RTL/cmsdk_iop_gpio.v(462)
  or u282 (n211, reg_inttypeset[11], reg_inttypeclr[11]);  // ../RTL/cmsdk_iop_gpio.v(461)
  AL_MUX u283 (
    .i0(reg_inttype_padded[11]),
    .i1(reg_inttypeset[11]),
    .sel(n211),
    .o(n212));  // ../RTL/cmsdk_iop_gpio.v(462)
  or u284 (n213, reg_inttypeset[12], reg_inttypeclr[12]);  // ../RTL/cmsdk_iop_gpio.v(461)
  AL_MUX u285 (
    .i0(reg_inttype_padded[12]),
    .i1(reg_inttypeset[12]),
    .sel(n213),
    .o(n214));  // ../RTL/cmsdk_iop_gpio.v(462)
  or u286 (n215, reg_inttypeset[13], reg_inttypeclr[13]);  // ../RTL/cmsdk_iop_gpio.v(461)
  AL_MUX u287 (
    .i0(reg_inttype_padded[13]),
    .i1(reg_inttypeset[13]),
    .sel(n215),
    .o(n216));  // ../RTL/cmsdk_iop_gpio.v(462)
  or u288 (n217, reg_inttypeset[14], reg_inttypeclr[14]);  // ../RTL/cmsdk_iop_gpio.v(461)
  AL_MUX u289 (
    .i0(reg_inttype_padded[14]),
    .i1(reg_inttypeset[14]),
    .sel(n217),
    .o(n218));  // ../RTL/cmsdk_iop_gpio.v(462)
  buf u29 (IORDATA[6], read_mux[6]);  // ../RTL/cmsdk_iop_gpio.v(577)
  or u290 (n219, reg_inttypeset[15], reg_inttypeclr[15]);  // ../RTL/cmsdk_iop_gpio.v(461)
  AL_MUX u291 (
    .i0(reg_inttype_padded[15]),
    .i1(reg_inttypeset[15]),
    .sel(n219),
    .o(n220));  // ../RTL/cmsdk_iop_gpio.v(462)
  buf u292 (reg_inten[0], reg_inten_padded[0]);  // ../RTL/cmsdk_iop_gpio.v(428)
  buf u293 (IORDATA[18], read_mux[18]);  // ../RTL/cmsdk_iop_gpio.v(577)
  and u294 (n222, write_trans, n221);  // ../RTL/cmsdk_iop_gpio.v(479)
  buf u295 (IORDATA[17], read_mux[17]);  // ../RTL/cmsdk_iop_gpio.v(577)
  and u296 (n223, n222, iop_byte_strobe[0]);  // ../RTL/cmsdk_iop_gpio.v(480)
  buf u297 (IORDATA[16], read_mux[16]);  // ../RTL/cmsdk_iop_gpio.v(577)
  or u298 (n317, n319, n318);  // ../RTL/cmsdk_iop_gpio.v(581)
  or u299 (n318, reg_intstat[10], reg_intstat[11]);  // ../RTL/cmsdk_iop_gpio.v(581)
  buf u3 (PORTEN[12], reg_douten[12]);  // ../RTL/cmsdk_iop_gpio.v(574)
  buf u30 (IORDATA[5], read_mux[5]);  // ../RTL/cmsdk_iop_gpio.v(577)
  buf u300 (IORDATA[15], read_mux[15]);  // ../RTL/cmsdk_iop_gpio.v(577)
  and u301 (n226, n222, iop_byte_strobe[1]);  // ../RTL/cmsdk_iop_gpio.v(483)
  buf u302 (IORDATA[14], read_mux[14]);  // ../RTL/cmsdk_iop_gpio.v(577)
  and u303 (n228, write_trans, n227);  // ../RTL/cmsdk_iop_gpio.v(485)
  buf u304 (IORDATA[13], read_mux[13]);  // ../RTL/cmsdk_iop_gpio.v(577)
  and u305 (n229, n228, iop_byte_strobe[0]);  // ../RTL/cmsdk_iop_gpio.v(486)
  buf u306 (IORDATA[12], read_mux[12]);  // ../RTL/cmsdk_iop_gpio.v(577)
  or u307 (n319, reg_intstat[8], reg_intstat[9]);  // ../RTL/cmsdk_iop_gpio.v(581)
  or u308 (n320, n324, n321);  // ../RTL/cmsdk_iop_gpio.v(581)
  buf u309 (IORDATA[11], read_mux[11]);  // ../RTL/cmsdk_iop_gpio.v(577)
  buf u31 (IORDATA[4], read_mux[4]);  // ../RTL/cmsdk_iop_gpio.v(577)
  and u310 (n232, n228, iop_byte_strobe[1]);  // ../RTL/cmsdk_iop_gpio.v(489)
  buf u311 (IORDATA[10], read_mux[10]);  // ../RTL/cmsdk_iop_gpio.v(577)
  or u312 (n321, n323, n322);  // ../RTL/cmsdk_iop_gpio.v(581)
  or u313 (n234, reg_intpolset[0], reg_intpolclr[0]);  // ../RTL/cmsdk_iop_gpio.v(499)
  AL_MUX u314 (
    .i0(reg_intpol_padded[0]),
    .i1(reg_intpolset[0]),
    .sel(n234),
    .o(n235));  // ../RTL/cmsdk_iop_gpio.v(500)
  or u315 (n236, reg_intpolset[1], reg_intpolclr[1]);  // ../RTL/cmsdk_iop_gpio.v(499)
  AL_MUX u316 (
    .i0(reg_intpol_padded[1]),
    .i1(reg_intpolset[1]),
    .sel(n236),
    .o(n237));  // ../RTL/cmsdk_iop_gpio.v(500)
  or u317 (n238, reg_intpolset[2], reg_intpolclr[2]);  // ../RTL/cmsdk_iop_gpio.v(499)
  AL_MUX u318 (
    .i0(reg_intpol_padded[2]),
    .i1(reg_intpolset[2]),
    .sel(n238),
    .o(n239));  // ../RTL/cmsdk_iop_gpio.v(500)
  or u319 (n240, reg_intpolset[3], reg_intpolclr[3]);  // ../RTL/cmsdk_iop_gpio.v(499)
  and u32 (reg_dout_normal_write1, n25, iop_byte_strobe[1]);  // ../RTL/cmsdk_iop_gpio.v(273)
  AL_MUX u320 (
    .i0(reg_intpol_padded[3]),
    .i1(reg_intpolset[3]),
    .sel(n240),
    .o(n241));  // ../RTL/cmsdk_iop_gpio.v(500)
  or u321 (n242, reg_intpolset[4], reg_intpolclr[4]);  // ../RTL/cmsdk_iop_gpio.v(499)
  AL_MUX u322 (
    .i0(reg_intpol_padded[4]),
    .i1(reg_intpolset[4]),
    .sel(n242),
    .o(n243));  // ../RTL/cmsdk_iop_gpio.v(500)
  or u323 (n244, reg_intpolset[5], reg_intpolclr[5]);  // ../RTL/cmsdk_iop_gpio.v(499)
  AL_MUX u324 (
    .i0(reg_intpol_padded[5]),
    .i1(reg_intpolset[5]),
    .sel(n244),
    .o(n245));  // ../RTL/cmsdk_iop_gpio.v(500)
  or u325 (n246, reg_intpolset[6], reg_intpolclr[6]);  // ../RTL/cmsdk_iop_gpio.v(499)
  AL_MUX u326 (
    .i0(reg_intpol_padded[6]),
    .i1(reg_intpolset[6]),
    .sel(n246),
    .o(n247));  // ../RTL/cmsdk_iop_gpio.v(500)
  or u327 (n248, reg_intpolset[7], reg_intpolclr[7]);  // ../RTL/cmsdk_iop_gpio.v(499)
  AL_MUX u328 (
    .i0(reg_intpol_padded[7]),
    .i1(reg_intpolset[7]),
    .sel(n248),
    .o(n249));  // ../RTL/cmsdk_iop_gpio.v(500)
  or u329 (n250, reg_intpolset[8], reg_intpolclr[8]);  // ../RTL/cmsdk_iop_gpio.v(499)
  and u33 (n27, write_trans, n26);  // ../RTL/cmsdk_iop_gpio.v(275)
  AL_MUX u330 (
    .i0(reg_intpol_padded[8]),
    .i1(reg_intpolset[8]),
    .sel(n250),
    .o(n251));  // ../RTL/cmsdk_iop_gpio.v(500)
  or u331 (n252, reg_intpolset[9], reg_intpolclr[9]);  // ../RTL/cmsdk_iop_gpio.v(499)
  AL_MUX u332 (
    .i0(reg_intpol_padded[9]),
    .i1(reg_intpolset[9]),
    .sel(n252),
    .o(n253));  // ../RTL/cmsdk_iop_gpio.v(500)
  or u333 (n254, reg_intpolset[10], reg_intpolclr[10]);  // ../RTL/cmsdk_iop_gpio.v(499)
  AL_MUX u334 (
    .i0(reg_intpol_padded[10]),
    .i1(reg_intpolset[10]),
    .sel(n254),
    .o(n255));  // ../RTL/cmsdk_iop_gpio.v(500)
  or u335 (n256, reg_intpolset[11], reg_intpolclr[11]);  // ../RTL/cmsdk_iop_gpio.v(499)
  AL_MUX u336 (
    .i0(reg_intpol_padded[11]),
    .i1(reg_intpolset[11]),
    .sel(n256),
    .o(n257));  // ../RTL/cmsdk_iop_gpio.v(500)
  or u337 (n258, reg_intpolset[12], reg_intpolclr[12]);  // ../RTL/cmsdk_iop_gpio.v(499)
  AL_MUX u338 (
    .i0(reg_intpol_padded[12]),
    .i1(reg_intpolset[12]),
    .sel(n258),
    .o(n259));  // ../RTL/cmsdk_iop_gpio.v(500)
  or u339 (n260, reg_intpolset[13], reg_intpolclr[13]);  // ../RTL/cmsdk_iop_gpio.v(499)
  and u34 (reg_dout_masked_write0, n27, iop_byte_strobe[0]);  // ../RTL/cmsdk_iop_gpio.v(275)
  AL_MUX u340 (
    .i0(reg_intpol_padded[13]),
    .i1(reg_intpolset[13]),
    .sel(n260),
    .o(n261));  // ../RTL/cmsdk_iop_gpio.v(500)
  or u341 (n262, reg_intpolset[14], reg_intpolclr[14]);  // ../RTL/cmsdk_iop_gpio.v(499)
  AL_MUX u342 (
    .i0(reg_intpol_padded[14]),
    .i1(reg_intpolset[14]),
    .sel(n262),
    .o(n263));  // ../RTL/cmsdk_iop_gpio.v(500)
  or u343 (n264, reg_intpolset[15], reg_intpolclr[15]);  // ../RTL/cmsdk_iop_gpio.v(499)
  AL_MUX u344 (
    .i0(reg_intpol_padded[15]),
    .i1(reg_intpolset[15]),
    .sel(n264),
    .o(n265));  // ../RTL/cmsdk_iop_gpio.v(500)
  buf u345 (reg_inttype[0], reg_inttype_padded[0]);  // ../RTL/cmsdk_iop_gpio.v(466)
  and u346 (n267, write_trans, n266);  // ../RTL/cmsdk_iop_gpio.v(520)
  and u347 (reg_intclr_normal_write0, n267, iop_byte_strobe[0]);  // ../RTL/cmsdk_iop_gpio.v(520)
  or u348 (n322, reg_intstat[6], reg_intstat[7]);  // ../RTL/cmsdk_iop_gpio.v(581)
  or u349 (n323, reg_intstat[4], reg_intstat[5]);  // ../RTL/cmsdk_iop_gpio.v(581)
  and u35 (n29, write_trans, n28);  // ../RTL/cmsdk_iop_gpio.v(277)
  and u350 (reg_intclr_normal_write1, n267, iop_byte_strobe[1]);  // ../RTL/cmsdk_iop_gpio.v(522)
  buf u351 (PORTOUT[1], reg_dout[1]);  // ../RTL/cmsdk_iop_gpio.v(573)
  buf u352 (reg_intpol[0], reg_intpol_padded[0]);  // ../RTL/cmsdk_iop_gpio.v(504)
  not u353 (n309[0], reg_intpol[0]);  // ../RTL/cmsdk_iop_gpio.v(565)
  buf u354 (IORDATA[9], read_mux[9]);  // ../RTL/cmsdk_iop_gpio.v(577)
  or u355 (n324, n326, n325);  // ../RTL/cmsdk_iop_gpio.v(581)
  or u356 (n271, new_masked_int[0], reg_intclr_padded[0]);  // ../RTL/cmsdk_iop_gpio.v(537)
  AL_MUX u357 (
    .i0(reg_intstat_padded[0]),
    .i1(new_masked_int[0]),
    .sel(n271),
    .o(n272));  // ../RTL/cmsdk_iop_gpio.v(538)
  or u358 (n273, new_masked_int[1], reg_intclr_padded[1]);  // ../RTL/cmsdk_iop_gpio.v(537)
  AL_MUX u359 (
    .i0(reg_intstat_padded[1]),
    .i1(new_masked_int[1]),
    .sel(n273),
    .o(n274));  // ../RTL/cmsdk_iop_gpio.v(538)
  and u36 (reg_dout_masked_write1, n29, iop_byte_strobe[1]);  // ../RTL/cmsdk_iop_gpio.v(277)
  or u360 (n275, new_masked_int[2], reg_intclr_padded[2]);  // ../RTL/cmsdk_iop_gpio.v(537)
  AL_MUX u361 (
    .i0(reg_intstat_padded[2]),
    .i1(new_masked_int[2]),
    .sel(n275),
    .o(n276));  // ../RTL/cmsdk_iop_gpio.v(538)
  or u362 (n277, new_masked_int[3], reg_intclr_padded[3]);  // ../RTL/cmsdk_iop_gpio.v(537)
  AL_MUX u363 (
    .i0(reg_intstat_padded[3]),
    .i1(new_masked_int[3]),
    .sel(n277),
    .o(n278));  // ../RTL/cmsdk_iop_gpio.v(538)
  or u364 (n279, new_masked_int[4], reg_intclr_padded[4]);  // ../RTL/cmsdk_iop_gpio.v(537)
  AL_MUX u365 (
    .i0(reg_intstat_padded[4]),
    .i1(new_masked_int[4]),
    .sel(n279),
    .o(n280));  // ../RTL/cmsdk_iop_gpio.v(538)
  or u366 (n281, new_masked_int[5], reg_intclr_padded[5]);  // ../RTL/cmsdk_iop_gpio.v(537)
  AL_MUX u367 (
    .i0(reg_intstat_padded[5]),
    .i1(new_masked_int[5]),
    .sel(n281),
    .o(n282));  // ../RTL/cmsdk_iop_gpio.v(538)
  or u368 (n283, new_masked_int[6], reg_intclr_padded[6]);  // ../RTL/cmsdk_iop_gpio.v(537)
  AL_MUX u369 (
    .i0(reg_intstat_padded[6]),
    .i1(new_masked_int[6]),
    .sel(n283),
    .o(n284));  // ../RTL/cmsdk_iop_gpio.v(538)
  buf u37 (reg_datain32[0], reg_datain[0]);  // ../RTL/cmsdk_iop_gpio.v(257)
  or u370 (n285, new_masked_int[7], reg_intclr_padded[7]);  // ../RTL/cmsdk_iop_gpio.v(537)
  AL_MUX u371 (
    .i0(reg_intstat_padded[7]),
    .i1(new_masked_int[7]),
    .sel(n285),
    .o(n286));  // ../RTL/cmsdk_iop_gpio.v(538)
  or u372 (n287, new_masked_int[8], reg_intclr_padded[8]);  // ../RTL/cmsdk_iop_gpio.v(537)
  AL_MUX u373 (
    .i0(reg_intstat_padded[8]),
    .i1(new_masked_int[8]),
    .sel(n287),
    .o(n288));  // ../RTL/cmsdk_iop_gpio.v(538)
  or u374 (n289, new_masked_int[9], reg_intclr_padded[9]);  // ../RTL/cmsdk_iop_gpio.v(537)
  AL_MUX u375 (
    .i0(reg_intstat_padded[9]),
    .i1(new_masked_int[9]),
    .sel(n289),
    .o(n290));  // ../RTL/cmsdk_iop_gpio.v(538)
  or u376 (n291, new_masked_int[10], reg_intclr_padded[10]);  // ../RTL/cmsdk_iop_gpio.v(537)
  AL_MUX u377 (
    .i0(reg_intstat_padded[10]),
    .i1(new_masked_int[10]),
    .sel(n291),
    .o(n292));  // ../RTL/cmsdk_iop_gpio.v(538)
  or u378 (n293, new_masked_int[11], reg_intclr_padded[11]);  // ../RTL/cmsdk_iop_gpio.v(537)
  AL_MUX u379 (
    .i0(reg_intstat_padded[11]),
    .i1(new_masked_int[11]),
    .sel(n293),
    .o(n294));  // ../RTL/cmsdk_iop_gpio.v(538)
  buf u38 (current_dout_padded[0], reg_dout[0]);  // ../RTL/cmsdk_iop_gpio.v(280)
  or u380 (n295, new_masked_int[12], reg_intclr_padded[12]);  // ../RTL/cmsdk_iop_gpio.v(537)
  AL_MUX u381 (
    .i0(reg_intstat_padded[12]),
    .i1(new_masked_int[12]),
    .sel(n295),
    .o(n296));  // ../RTL/cmsdk_iop_gpio.v(538)
  or u382 (n297, new_masked_int[13], reg_intclr_padded[13]);  // ../RTL/cmsdk_iop_gpio.v(537)
  AL_MUX u383 (
    .i0(reg_intstat_padded[13]),
    .i1(new_masked_int[13]),
    .sel(n297),
    .o(n298));  // ../RTL/cmsdk_iop_gpio.v(538)
  or u384 (n299, new_masked_int[14], reg_intclr_padded[14]);  // ../RTL/cmsdk_iop_gpio.v(537)
  AL_MUX u385 (
    .i0(reg_intstat_padded[14]),
    .i1(new_masked_int[14]),
    .sel(n299),
    .o(n300));  // ../RTL/cmsdk_iop_gpio.v(538)
  or u386 (n301, new_masked_int[15], reg_intclr_padded[15]);  // ../RTL/cmsdk_iop_gpio.v(537)
  AL_MUX u387 (
    .i0(reg_intstat_padded[15]),
    .i1(new_masked_int[15]),
    .sel(n301),
    .o(n302));  // ../RTL/cmsdk_iop_gpio.v(538)
  and u388 (new_masked_int[0], new_raw_int[0], reg_inten[0]);  // ../RTL/cmsdk_iop_gpio.v(527)
  buf u389 (reg_intstat[0], reg_intstat_padded[0]);  // ../RTL/cmsdk_iop_gpio.v(542)
  or u39 (n335[1], n334[1], rise_edge_int[1]);  // ../RTL/cmsdk_iop_gpio.v(568)
  or u390 (n325, reg_intstat[2], reg_intstat[3]);  // ../RTL/cmsdk_iop_gpio.v(581)
  not u391 (n3[1], IOADDR[1]);  // ../RTL/cmsdk_iop_gpio.v(143)
  or u392 (n312, reg_inttype[0], reg_inttype[1]);  // ../RTL/cmsdk_iop_gpio.v(560)
  and u393 (n10[0], reg_datain32[0], IOADDR[2]);  // ../RTL/cmsdk_iop_gpio.v(175)
  and u394 (n306[0], reg_datain[0], reg_intpol[0]);  // ../RTL/cmsdk_iop_gpio.v(564)
  not u395 (n307[0], reg_inttype[0]);  // ../RTL/cmsdk_iop_gpio.v(564)
  buf u396 (PORTEN[14], reg_douten[14]);  // ../RTL/cmsdk_iop_gpio.v(574)
  buf u397 (PORTEN[15], reg_douten[15]);  // ../RTL/cmsdk_iop_gpio.v(574)
  and u398 (high_level_int[0], n306[0], n307[0]);  // ../RTL/cmsdk_iop_gpio.v(564)
  or u399 (n326, reg_intstat[0], reg_intstat[1]);  // ../RTL/cmsdk_iop_gpio.v(581)
  and u4 (n0, IOSEL, IOWRITE);  // ../RTL/cmsdk_iop_gpio.v(135)
  not u40 (n31[0], IOADDR[2]);  // ../RTL/cmsdk_iop_gpio.v(286)
  and u400 (n310[0], n308[0], n309[0]);  // ../RTL/cmsdk_iop_gpio.v(565)
  and u401 (low_level_int[0], n310[0], n307[0]);  // ../RTL/cmsdk_iop_gpio.v(565)
  not u402 (n327[0], reg_last_datain[0]);  // ../RTL/cmsdk_iop_gpio.v(566)
  and u403 (n328[0], reg_datain[0], n327[0]);  // ../RTL/cmsdk_iop_gpio.v(566)
  and u404 (n329[0], n328[0], reg_intpol[0]);  // ../RTL/cmsdk_iop_gpio.v(566)
  and u405 (rise_edge_int[0], n329[0], reg_inttype[0]);  // ../RTL/cmsdk_iop_gpio.v(566)
  not u406 (n330[0], reg_datain[0]);  // ../RTL/cmsdk_iop_gpio.v(567)
  and u407 (n331[0], n330[0], reg_last_datain[0]);  // ../RTL/cmsdk_iop_gpio.v(567)
  not u408 (n332[0], reg_intpol[0]);  // ../RTL/cmsdk_iop_gpio.v(567)
  and u409 (n333[0], n331[0], n332[0]);  // ../RTL/cmsdk_iop_gpio.v(567)
  buf u41 (PORTEN[10], reg_douten[10]);  // ../RTL/cmsdk_iop_gpio.v(574)
  and u410 (fall_edge_int[0], n333[0], reg_inttype[0]);  // ../RTL/cmsdk_iop_gpio.v(567)
  or u411 (n334[0], high_level_int[0], low_level_int[0]);  // ../RTL/cmsdk_iop_gpio.v(568)
  or u412 (n335[0], n334[0], rise_edge_int[0]);  // ../RTL/cmsdk_iop_gpio.v(568)
  or u413 (new_raw_int[0], n335[0], fall_edge_int[0]);  // ../RTL/cmsdk_iop_gpio.v(568)
  buf u414 (PORTOUT[0], reg_dout[0]);  // ../RTL/cmsdk_iop_gpio.v(573)
  buf u415 (PORTEN[0], reg_douten[0]);  // ../RTL/cmsdk_iop_gpio.v(574)
  buf u416 (PORTFUNC[0], reg_altfunc[0]);  // ../RTL/cmsdk_iop_gpio.v(575)
  buf u417 (IORDATA[0], read_mux[0]);  // ../RTL/cmsdk_iop_gpio.v(577)
  buf u418 (GPIOINT[0], reg_intstat[0]);  // ../RTL/cmsdk_iop_gpio.v(580)
  or u419 (n335[9], n334[9], rise_edge_int[9]);  // ../RTL/cmsdk_iop_gpio.v(568)
  buf u42 (IORDATA[3], read_mux[3]);  // ../RTL/cmsdk_iop_gpio.v(577)
  or u420 (n335[10], n334[10], rise_edge_int[10]);  // ../RTL/cmsdk_iop_gpio.v(568)
  or u421 (n335[11], n334[11], rise_edge_int[11]);  // ../RTL/cmsdk_iop_gpio.v(568)
  or u422 (n335[12], n334[12], rise_edge_int[12]);  // ../RTL/cmsdk_iop_gpio.v(568)
  or u423 (n335[13], n334[13], rise_edge_int[13]);  // ../RTL/cmsdk_iop_gpio.v(568)
  or u424 (n335[14], n334[14], rise_edge_int[14]);  // ../RTL/cmsdk_iop_gpio.v(568)
  or u425 (n335[15], n334[15], rise_edge_int[15]);  // ../RTL/cmsdk_iop_gpio.v(568)
  or u426 (n334[1], high_level_int[1], low_level_int[1]);  // ../RTL/cmsdk_iop_gpio.v(568)
  or u427 (n334[2], high_level_int[2], low_level_int[2]);  // ../RTL/cmsdk_iop_gpio.v(568)
  or u428 (n334[3], high_level_int[3], low_level_int[3]);  // ../RTL/cmsdk_iop_gpio.v(568)
  or u429 (n334[4], high_level_int[4], low_level_int[4]);  // ../RTL/cmsdk_iop_gpio.v(568)
  or u43 (n34, reg_dout_normal_write0, reg_dout_masked_write0);  // ../RTL/cmsdk_iop_gpio.v(293)
  or u430 (n334[5], high_level_int[5], low_level_int[5]);  // ../RTL/cmsdk_iop_gpio.v(568)
  or u431 (n334[6], high_level_int[6], low_level_int[6]);  // ../RTL/cmsdk_iop_gpio.v(568)
  or u432 (n334[7], high_level_int[7], low_level_int[7]);  // ../RTL/cmsdk_iop_gpio.v(568)
  or u433 (n334[8], high_level_int[8], low_level_int[8]);  // ../RTL/cmsdk_iop_gpio.v(568)
  or u434 (n334[9], high_level_int[9], low_level_int[9]);  // ../RTL/cmsdk_iop_gpio.v(568)
  or u435 (n334[10], high_level_int[10], low_level_int[10]);  // ../RTL/cmsdk_iop_gpio.v(568)
  or u436 (n334[11], high_level_int[11], low_level_int[11]);  // ../RTL/cmsdk_iop_gpio.v(568)
  or u437 (n334[12], high_level_int[12], low_level_int[12]);  // ../RTL/cmsdk_iop_gpio.v(568)
  or u438 (n334[13], high_level_int[13], low_level_int[13]);  // ../RTL/cmsdk_iop_gpio.v(568)
  or u439 (n334[14], high_level_int[14], low_level_int[14]);  // ../RTL/cmsdk_iop_gpio.v(568)
  or u44 (new_raw_int[2], n335[2], fall_edge_int[2]);  // ../RTL/cmsdk_iop_gpio.v(568)
  or u440 (n334[15], high_level_int[15], low_level_int[15]);  // ../RTL/cmsdk_iop_gpio.v(568)
  and u441 (fall_edge_int[1], n333[1], reg_inttype[1]);  // ../RTL/cmsdk_iop_gpio.v(567)
  and u442 (fall_edge_int[2], n333[2], reg_inttype[2]);  // ../RTL/cmsdk_iop_gpio.v(567)
  and u443 (fall_edge_int[3], n333[3], reg_inttype[3]);  // ../RTL/cmsdk_iop_gpio.v(567)
  and u444 (fall_edge_int[4], n333[4], reg_inttype[4]);  // ../RTL/cmsdk_iop_gpio.v(567)
  and u445 (fall_edge_int[5], n333[5], reg_inttype[5]);  // ../RTL/cmsdk_iop_gpio.v(567)
  and u446 (fall_edge_int[6], n333[6], reg_inttype[6]);  // ../RTL/cmsdk_iop_gpio.v(567)
  and u447 (fall_edge_int[7], n333[7], reg_inttype[7]);  // ../RTL/cmsdk_iop_gpio.v(567)
  and u448 (fall_edge_int[8], n333[8], reg_inttype[8]);  // ../RTL/cmsdk_iop_gpio.v(567)
  and u449 (fall_edge_int[9], n333[9], reg_inttype[9]);  // ../RTL/cmsdk_iop_gpio.v(567)
  or u45 (new_raw_int[3], n335[3], fall_edge_int[3]);  // ../RTL/cmsdk_iop_gpio.v(568)
  and u450 (fall_edge_int[10], n333[10], reg_inttype[10]);  // ../RTL/cmsdk_iop_gpio.v(567)
  and u451 (fall_edge_int[11], n333[11], reg_inttype[11]);  // ../RTL/cmsdk_iop_gpio.v(567)
  and u452 (fall_edge_int[12], n333[12], reg_inttype[12]);  // ../RTL/cmsdk_iop_gpio.v(567)
  and u453 (fall_edge_int[13], n333[13], reg_inttype[13]);  // ../RTL/cmsdk_iop_gpio.v(567)
  and u454 (fall_edge_int[14], n333[14], reg_inttype[14]);  // ../RTL/cmsdk_iop_gpio.v(567)
  and u455 (fall_edge_int[15], n333[15], reg_inttype[15]);  // ../RTL/cmsdk_iop_gpio.v(567)
  and u456 (n333[1], n331[1], n332[1]);  // ../RTL/cmsdk_iop_gpio.v(567)
  and u457 (n333[2], n331[2], n332[2]);  // ../RTL/cmsdk_iop_gpio.v(567)
  and u458 (n333[3], n331[3], n332[3]);  // ../RTL/cmsdk_iop_gpio.v(567)
  and u459 (n333[4], n331[4], n332[4]);  // ../RTL/cmsdk_iop_gpio.v(567)
  or u46 (new_raw_int[4], n335[4], fall_edge_int[4]);  // ../RTL/cmsdk_iop_gpio.v(568)
  and u460 (n333[5], n331[5], n332[5]);  // ../RTL/cmsdk_iop_gpio.v(567)
  and u461 (n333[6], n331[6], n332[6]);  // ../RTL/cmsdk_iop_gpio.v(567)
  and u462 (n333[7], n331[7], n332[7]);  // ../RTL/cmsdk_iop_gpio.v(567)
  and u463 (n333[8], n331[8], n332[8]);  // ../RTL/cmsdk_iop_gpio.v(567)
  and u464 (n333[9], n331[9], n332[9]);  // ../RTL/cmsdk_iop_gpio.v(567)
  and u465 (n333[10], n331[10], n332[10]);  // ../RTL/cmsdk_iop_gpio.v(567)
  and u466 (n333[11], n331[11], n332[11]);  // ../RTL/cmsdk_iop_gpio.v(567)
  and u467 (n333[12], n331[12], n332[12]);  // ../RTL/cmsdk_iop_gpio.v(567)
  and u468 (n333[13], n331[13], n332[13]);  // ../RTL/cmsdk_iop_gpio.v(567)
  and u469 (n333[14], n331[14], n332[14]);  // ../RTL/cmsdk_iop_gpio.v(567)
  or u47 (new_raw_int[5], n335[5], fall_edge_int[5]);  // ../RTL/cmsdk_iop_gpio.v(568)
  and u470 (n333[15], n331[15], n332[15]);  // ../RTL/cmsdk_iop_gpio.v(567)
  not u471 (n332[1], reg_intpol[1]);  // ../RTL/cmsdk_iop_gpio.v(567)
  not u472 (n332[2], reg_intpol[2]);  // ../RTL/cmsdk_iop_gpio.v(567)
  not u473 (n332[3], reg_intpol[3]);  // ../RTL/cmsdk_iop_gpio.v(567)
  not u474 (n332[4], reg_intpol[4]);  // ../RTL/cmsdk_iop_gpio.v(567)
  not u475 (n332[5], reg_intpol[5]);  // ../RTL/cmsdk_iop_gpio.v(567)
  not u476 (n332[6], reg_intpol[6]);  // ../RTL/cmsdk_iop_gpio.v(567)
  not u477 (n332[7], reg_intpol[7]);  // ../RTL/cmsdk_iop_gpio.v(567)
  not u478 (n332[8], reg_intpol[8]);  // ../RTL/cmsdk_iop_gpio.v(567)
  not u479 (n332[9], reg_intpol[9]);  // ../RTL/cmsdk_iop_gpio.v(567)
  or u48 (new_raw_int[6], n335[6], fall_edge_int[6]);  // ../RTL/cmsdk_iop_gpio.v(568)
  not u480 (n332[10], reg_intpol[10]);  // ../RTL/cmsdk_iop_gpio.v(567)
  not u481 (n332[11], reg_intpol[11]);  // ../RTL/cmsdk_iop_gpio.v(567)
  not u482 (n332[12], reg_intpol[12]);  // ../RTL/cmsdk_iop_gpio.v(567)
  not u483 (n332[13], reg_intpol[13]);  // ../RTL/cmsdk_iop_gpio.v(567)
  not u484 (n332[14], reg_intpol[14]);  // ../RTL/cmsdk_iop_gpio.v(567)
  not u485 (n332[15], reg_intpol[15]);  // ../RTL/cmsdk_iop_gpio.v(567)
  and u486 (n331[1], n330[1], reg_last_datain[1]);  // ../RTL/cmsdk_iop_gpio.v(567)
  and u487 (n331[2], n330[2], reg_last_datain[2]);  // ../RTL/cmsdk_iop_gpio.v(567)
  and u488 (n331[3], n330[3], reg_last_datain[3]);  // ../RTL/cmsdk_iop_gpio.v(567)
  and u489 (n331[4], n330[4], reg_last_datain[4]);  // ../RTL/cmsdk_iop_gpio.v(567)
  or u49 (new_raw_int[7], n335[7], fall_edge_int[7]);  // ../RTL/cmsdk_iop_gpio.v(568)
  and u490 (n331[5], n330[5], reg_last_datain[5]);  // ../RTL/cmsdk_iop_gpio.v(567)
  and u491 (n331[6], n330[6], reg_last_datain[6]);  // ../RTL/cmsdk_iop_gpio.v(567)
  and u492 (n331[7], n330[7], reg_last_datain[7]);  // ../RTL/cmsdk_iop_gpio.v(567)
  and u493 (n331[8], n330[8], reg_last_datain[8]);  // ../RTL/cmsdk_iop_gpio.v(567)
  and u494 (n331[9], n330[9], reg_last_datain[9]);  // ../RTL/cmsdk_iop_gpio.v(567)
  and u495 (n331[10], n330[10], reg_last_datain[10]);  // ../RTL/cmsdk_iop_gpio.v(567)
  and u496 (n331[11], n330[11], reg_last_datain[11]);  // ../RTL/cmsdk_iop_gpio.v(567)
  and u497 (n331[12], n330[12], reg_last_datain[12]);  // ../RTL/cmsdk_iop_gpio.v(567)
  and u498 (n331[13], n330[13], reg_last_datain[13]);  // ../RTL/cmsdk_iop_gpio.v(567)
  and u499 (n331[14], n330[14], reg_last_datain[14]);  // ../RTL/cmsdk_iop_gpio.v(567)
  and u5 (write_trans, n0, IOTRANS);  // ../RTL/cmsdk_iop_gpio.v(135)
  or u50 (new_raw_int[8], n335[8], fall_edge_int[8]);  // ../RTL/cmsdk_iop_gpio.v(568)
  and u500 (n331[15], n330[15], reg_last_datain[15]);  // ../RTL/cmsdk_iop_gpio.v(567)
  not u501 (n330[1], reg_datain[1]);  // ../RTL/cmsdk_iop_gpio.v(567)
  not u502 (n330[2], reg_datain[2]);  // ../RTL/cmsdk_iop_gpio.v(567)
  not u503 (n330[3], reg_datain[3]);  // ../RTL/cmsdk_iop_gpio.v(567)
  not u504 (n330[4], reg_datain[4]);  // ../RTL/cmsdk_iop_gpio.v(567)
  not u505 (n330[5], reg_datain[5]);  // ../RTL/cmsdk_iop_gpio.v(567)
  not u506 (n330[6], reg_datain[6]);  // ../RTL/cmsdk_iop_gpio.v(567)
  not u507 (n330[7], reg_datain[7]);  // ../RTL/cmsdk_iop_gpio.v(567)
  not u508 (n330[8], reg_datain[8]);  // ../RTL/cmsdk_iop_gpio.v(567)
  not u509 (n330[9], reg_datain[9]);  // ../RTL/cmsdk_iop_gpio.v(567)
  buf u51 (PORTOUT[10], reg_dout[10]);  // ../RTL/cmsdk_iop_gpio.v(573)
  not u510 (n330[10], reg_datain[10]);  // ../RTL/cmsdk_iop_gpio.v(567)
  not u511 (n330[11], reg_datain[11]);  // ../RTL/cmsdk_iop_gpio.v(567)
  not u512 (n330[12], reg_datain[12]);  // ../RTL/cmsdk_iop_gpio.v(567)
  not u513 (n330[13], reg_datain[13]);  // ../RTL/cmsdk_iop_gpio.v(567)
  not u514 (n330[14], reg_datain[14]);  // ../RTL/cmsdk_iop_gpio.v(567)
  not u515 (n330[15], reg_datain[15]);  // ../RTL/cmsdk_iop_gpio.v(567)
  and u516 (rise_edge_int[1], n329[1], reg_inttype[1]);  // ../RTL/cmsdk_iop_gpio.v(566)
  and u517 (rise_edge_int[2], n329[2], reg_inttype[2]);  // ../RTL/cmsdk_iop_gpio.v(566)
  and u518 (rise_edge_int[3], n329[3], reg_inttype[3]);  // ../RTL/cmsdk_iop_gpio.v(566)
  and u519 (rise_edge_int[4], n329[4], reg_inttype[4]);  // ../RTL/cmsdk_iop_gpio.v(566)
  buf u52 (PORTOUT[11], reg_dout[11]);  // ../RTL/cmsdk_iop_gpio.v(573)
  and u520 (rise_edge_int[5], n329[5], reg_inttype[5]);  // ../RTL/cmsdk_iop_gpio.v(566)
  and u521 (rise_edge_int[6], n329[6], reg_inttype[6]);  // ../RTL/cmsdk_iop_gpio.v(566)
  and u522 (rise_edge_int[7], n329[7], reg_inttype[7]);  // ../RTL/cmsdk_iop_gpio.v(566)
  and u523 (rise_edge_int[8], n329[8], reg_inttype[8]);  // ../RTL/cmsdk_iop_gpio.v(566)
  and u524 (rise_edge_int[9], n329[9], reg_inttype[9]);  // ../RTL/cmsdk_iop_gpio.v(566)
  and u525 (rise_edge_int[10], n329[10], reg_inttype[10]);  // ../RTL/cmsdk_iop_gpio.v(566)
  and u526 (rise_edge_int[11], n329[11], reg_inttype[11]);  // ../RTL/cmsdk_iop_gpio.v(566)
  and u527 (rise_edge_int[12], n329[12], reg_inttype[12]);  // ../RTL/cmsdk_iop_gpio.v(566)
  and u528 (rise_edge_int[13], n329[13], reg_inttype[13]);  // ../RTL/cmsdk_iop_gpio.v(566)
  and u529 (rise_edge_int[14], n329[14], reg_inttype[14]);  // ../RTL/cmsdk_iop_gpio.v(566)
  buf u53 (PORTOUT[12], reg_dout[12]);  // ../RTL/cmsdk_iop_gpio.v(573)
  and u530 (rise_edge_int[15], n329[15], reg_inttype[15]);  // ../RTL/cmsdk_iop_gpio.v(566)
  and u531 (n329[1], n328[1], reg_intpol[1]);  // ../RTL/cmsdk_iop_gpio.v(566)
  and u532 (n329[2], n328[2], reg_intpol[2]);  // ../RTL/cmsdk_iop_gpio.v(566)
  and u533 (n329[3], n328[3], reg_intpol[3]);  // ../RTL/cmsdk_iop_gpio.v(566)
  and u534 (n329[4], n328[4], reg_intpol[4]);  // ../RTL/cmsdk_iop_gpio.v(566)
  and u535 (n329[5], n328[5], reg_intpol[5]);  // ../RTL/cmsdk_iop_gpio.v(566)
  and u536 (n329[6], n328[6], reg_intpol[6]);  // ../RTL/cmsdk_iop_gpio.v(566)
  and u537 (n329[7], n328[7], reg_intpol[7]);  // ../RTL/cmsdk_iop_gpio.v(566)
  and u538 (n329[8], n328[8], reg_intpol[8]);  // ../RTL/cmsdk_iop_gpio.v(566)
  and u539 (n329[9], n328[9], reg_intpol[9]);  // ../RTL/cmsdk_iop_gpio.v(566)
  buf u54 (PORTOUT[13], reg_dout[13]);  // ../RTL/cmsdk_iop_gpio.v(573)
  and u540 (n329[10], n328[10], reg_intpol[10]);  // ../RTL/cmsdk_iop_gpio.v(566)
  and u541 (n329[11], n328[11], reg_intpol[11]);  // ../RTL/cmsdk_iop_gpio.v(566)
  and u542 (n329[12], n328[12], reg_intpol[12]);  // ../RTL/cmsdk_iop_gpio.v(566)
  and u543 (n329[13], n328[13], reg_intpol[13]);  // ../RTL/cmsdk_iop_gpio.v(566)
  and u544 (n329[14], n328[14], reg_intpol[14]);  // ../RTL/cmsdk_iop_gpio.v(566)
  and u545 (n329[15], n328[15], reg_intpol[15]);  // ../RTL/cmsdk_iop_gpio.v(566)
  and u546 (n328[1], reg_datain[1], n327[1]);  // ../RTL/cmsdk_iop_gpio.v(566)
  and u547 (n328[2], reg_datain[2], n327[2]);  // ../RTL/cmsdk_iop_gpio.v(566)
  and u548 (n328[3], reg_datain[3], n327[3]);  // ../RTL/cmsdk_iop_gpio.v(566)
  and u549 (n328[4], reg_datain[4], n327[4]);  // ../RTL/cmsdk_iop_gpio.v(566)
  buf u55 (PORTOUT[14], reg_dout[14]);  // ../RTL/cmsdk_iop_gpio.v(573)
  and u550 (n328[5], reg_datain[5], n327[5]);  // ../RTL/cmsdk_iop_gpio.v(566)
  and u551 (n328[6], reg_datain[6], n327[6]);  // ../RTL/cmsdk_iop_gpio.v(566)
  and u552 (n328[7], reg_datain[7], n327[7]);  // ../RTL/cmsdk_iop_gpio.v(566)
  and u553 (n328[8], reg_datain[8], n327[8]);  // ../RTL/cmsdk_iop_gpio.v(566)
  and u554 (n328[9], reg_datain[9], n327[9]);  // ../RTL/cmsdk_iop_gpio.v(566)
  and u555 (n328[10], reg_datain[10], n327[10]);  // ../RTL/cmsdk_iop_gpio.v(566)
  and u556 (n328[11], reg_datain[11], n327[11]);  // ../RTL/cmsdk_iop_gpio.v(566)
  and u557 (n328[12], reg_datain[12], n327[12]);  // ../RTL/cmsdk_iop_gpio.v(566)
  and u558 (n328[13], reg_datain[13], n327[13]);  // ../RTL/cmsdk_iop_gpio.v(566)
  and u559 (n328[14], reg_datain[14], n327[14]);  // ../RTL/cmsdk_iop_gpio.v(566)
  buf u56 (PORTOUT[15], reg_dout[15]);  // ../RTL/cmsdk_iop_gpio.v(573)
  and u560 (n328[15], reg_datain[15], n327[15]);  // ../RTL/cmsdk_iop_gpio.v(566)
  not u561 (n327[1], reg_last_datain[1]);  // ../RTL/cmsdk_iop_gpio.v(566)
  not u562 (n327[2], reg_last_datain[2]);  // ../RTL/cmsdk_iop_gpio.v(566)
  not u563 (n327[3], reg_last_datain[3]);  // ../RTL/cmsdk_iop_gpio.v(566)
  not u564 (n327[4], reg_last_datain[4]);  // ../RTL/cmsdk_iop_gpio.v(566)
  not u565 (n327[5], reg_last_datain[5]);  // ../RTL/cmsdk_iop_gpio.v(566)
  not u566 (n327[6], reg_last_datain[6]);  // ../RTL/cmsdk_iop_gpio.v(566)
  not u567 (n327[7], reg_last_datain[7]);  // ../RTL/cmsdk_iop_gpio.v(566)
  not u568 (n327[8], reg_last_datain[8]);  // ../RTL/cmsdk_iop_gpio.v(566)
  not u569 (n327[9], reg_last_datain[9]);  // ../RTL/cmsdk_iop_gpio.v(566)
  or u57 (new_raw_int[1], n335[1], fall_edge_int[1]);  // ../RTL/cmsdk_iop_gpio.v(568)
  not u570 (n327[10], reg_last_datain[10]);  // ../RTL/cmsdk_iop_gpio.v(566)
  not u571 (n327[11], reg_last_datain[11]);  // ../RTL/cmsdk_iop_gpio.v(566)
  not u572 (n327[12], reg_last_datain[12]);  // ../RTL/cmsdk_iop_gpio.v(566)
  not u573 (n327[13], reg_last_datain[13]);  // ../RTL/cmsdk_iop_gpio.v(566)
  not u574 (n327[14], reg_last_datain[14]);  // ../RTL/cmsdk_iop_gpio.v(566)
  not u575 (n327[15], reg_last_datain[15]);  // ../RTL/cmsdk_iop_gpio.v(566)
  and u576 (low_level_int[1], n310[1], n307[1]);  // ../RTL/cmsdk_iop_gpio.v(565)
  and u577 (low_level_int[2], n310[2], n307[2]);  // ../RTL/cmsdk_iop_gpio.v(565)
  and u578 (low_level_int[3], n310[3], n307[3]);  // ../RTL/cmsdk_iop_gpio.v(565)
  and u579 (low_level_int[4], n310[4], n307[4]);  // ../RTL/cmsdk_iop_gpio.v(565)
  or u58 (n33[0], n30[0], n32[0]);  // ../RTL/cmsdk_iop_gpio.v(286)
  and u580 (low_level_int[5], n310[5], n307[5]);  // ../RTL/cmsdk_iop_gpio.v(565)
  and u581 (low_level_int[6], n310[6], n307[6]);  // ../RTL/cmsdk_iop_gpio.v(565)
  and u582 (low_level_int[7], n310[7], n307[7]);  // ../RTL/cmsdk_iop_gpio.v(565)
  and u583 (low_level_int[8], n310[8], n307[8]);  // ../RTL/cmsdk_iop_gpio.v(565)
  and u584 (low_level_int[9], n310[9], n307[9]);  // ../RTL/cmsdk_iop_gpio.v(565)
  and u585 (low_level_int[10], n310[10], n307[10]);  // ../RTL/cmsdk_iop_gpio.v(565)
  and u586 (low_level_int[11], n310[11], n307[11]);  // ../RTL/cmsdk_iop_gpio.v(565)
  and u587 (low_level_int[12], n310[12], n307[12]);  // ../RTL/cmsdk_iop_gpio.v(565)
  and u588 (low_level_int[13], n310[13], n307[13]);  // ../RTL/cmsdk_iop_gpio.v(565)
  and u589 (low_level_int[14], n310[14], n307[14]);  // ../RTL/cmsdk_iop_gpio.v(565)
  and u59 (reg_intclr_padded[0], reg_intclr_normal_write0, IOWDATALE[0]);  // ../RTL/cmsdk_iop_gpio.v(525)
  and u590 (low_level_int[15], n310[15], n307[15]);  // ../RTL/cmsdk_iop_gpio.v(565)
  and u591 (n310[1], n308[1], n309[1]);  // ../RTL/cmsdk_iop_gpio.v(565)
  and u592 (n310[2], n308[2], n309[2]);  // ../RTL/cmsdk_iop_gpio.v(565)
  and u593 (n310[3], n308[3], n309[3]);  // ../RTL/cmsdk_iop_gpio.v(565)
  and u594 (n310[4], n308[4], n309[4]);  // ../RTL/cmsdk_iop_gpio.v(565)
  and u595 (n310[5], n308[5], n309[5]);  // ../RTL/cmsdk_iop_gpio.v(565)
  and u596 (n310[6], n308[6], n309[6]);  // ../RTL/cmsdk_iop_gpio.v(565)
  and u597 (n310[7], n308[7], n309[7]);  // ../RTL/cmsdk_iop_gpio.v(565)
  and u598 (n310[8], n308[8], n309[8]);  // ../RTL/cmsdk_iop_gpio.v(565)
  and u599 (n310[9], n308[9], n309[9]);  // ../RTL/cmsdk_iop_gpio.v(565)
  buf u6 (bigendian, 1'b0);  // ../RTL/cmsdk_iop_gpio.v(139)
  buf u60 (IORDATA[2], read_mux[2]);  // ../RTL/cmsdk_iop_gpio.v(577)
  and u600 (n310[10], n308[10], n309[10]);  // ../RTL/cmsdk_iop_gpio.v(565)
  and u601 (n310[11], n308[11], n309[11]);  // ../RTL/cmsdk_iop_gpio.v(565)
  and u602 (n310[12], n308[12], n309[12]);  // ../RTL/cmsdk_iop_gpio.v(565)
  and u603 (n310[13], n308[13], n309[13]);  // ../RTL/cmsdk_iop_gpio.v(565)
  and u604 (n310[14], n308[14], n309[14]);  // ../RTL/cmsdk_iop_gpio.v(565)
  and u605 (n310[15], n308[15], n309[15]);  // ../RTL/cmsdk_iop_gpio.v(565)
  and u606 (high_level_int[1], n306[1], n307[1]);  // ../RTL/cmsdk_iop_gpio.v(564)
  and u607 (high_level_int[2], n306[2], n307[2]);  // ../RTL/cmsdk_iop_gpio.v(564)
  and u608 (high_level_int[3], n306[3], n307[3]);  // ../RTL/cmsdk_iop_gpio.v(564)
  and u609 (high_level_int[4], n306[4], n307[4]);  // ../RTL/cmsdk_iop_gpio.v(564)
  or u61 (n335[2], n334[2], rise_edge_int[2]);  // ../RTL/cmsdk_iop_gpio.v(568)
  and u610 (high_level_int[5], n306[5], n307[5]);  // ../RTL/cmsdk_iop_gpio.v(564)
  and u611 (high_level_int[6], n306[6], n307[6]);  // ../RTL/cmsdk_iop_gpio.v(564)
  and u612 (high_level_int[7], n306[7], n307[7]);  // ../RTL/cmsdk_iop_gpio.v(564)
  and u613 (high_level_int[8], n306[8], n307[8]);  // ../RTL/cmsdk_iop_gpio.v(564)
  and u614 (high_level_int[9], n306[9], n307[9]);  // ../RTL/cmsdk_iop_gpio.v(564)
  and u615 (high_level_int[10], n306[10], n307[10]);  // ../RTL/cmsdk_iop_gpio.v(564)
  and u616 (high_level_int[11], n306[11], n307[11]);  // ../RTL/cmsdk_iop_gpio.v(564)
  and u617 (high_level_int[12], n306[12], n307[12]);  // ../RTL/cmsdk_iop_gpio.v(564)
  and u618 (high_level_int[13], n306[13], n307[13]);  // ../RTL/cmsdk_iop_gpio.v(564)
  and u619 (high_level_int[14], n306[14], n307[14]);  // ../RTL/cmsdk_iop_gpio.v(564)
  and u62 (n32[0], current_dout_padded[0], n31[0]);  // ../RTL/cmsdk_iop_gpio.v(286)
  and u620 (high_level_int[15], n306[15], n307[15]);  // ../RTL/cmsdk_iop_gpio.v(564)
  not u621 (n307[1], reg_inttype[1]);  // ../RTL/cmsdk_iop_gpio.v(564)
  not u622 (n307[2], reg_inttype[2]);  // ../RTL/cmsdk_iop_gpio.v(564)
  not u623 (n307[3], reg_inttype[3]);  // ../RTL/cmsdk_iop_gpio.v(564)
  not u624 (n307[4], reg_inttype[4]);  // ../RTL/cmsdk_iop_gpio.v(564)
  not u625 (n307[5], reg_inttype[5]);  // ../RTL/cmsdk_iop_gpio.v(564)
  not u626 (n307[6], reg_inttype[6]);  // ../RTL/cmsdk_iop_gpio.v(564)
  not u627 (n307[7], reg_inttype[7]);  // ../RTL/cmsdk_iop_gpio.v(564)
  not u628 (n307[8], reg_inttype[8]);  // ../RTL/cmsdk_iop_gpio.v(564)
  not u629 (n307[9], reg_inttype[9]);  // ../RTL/cmsdk_iop_gpio.v(564)
  buf u63 (PORTEN[9], reg_douten[9]);  // ../RTL/cmsdk_iop_gpio.v(574)
  not u630 (n307[10], reg_inttype[10]);  // ../RTL/cmsdk_iop_gpio.v(564)
  not u631 (n307[11], reg_inttype[11]);  // ../RTL/cmsdk_iop_gpio.v(564)
  not u632 (n307[12], reg_inttype[12]);  // ../RTL/cmsdk_iop_gpio.v(564)
  not u633 (n307[13], reg_inttype[13]);  // ../RTL/cmsdk_iop_gpio.v(564)
  not u634 (n307[14], reg_inttype[14]);  // ../RTL/cmsdk_iop_gpio.v(564)
  not u635 (n307[15], reg_inttype[15]);  // ../RTL/cmsdk_iop_gpio.v(564)
  and u636 (n306[1], reg_datain[1], reg_intpol[1]);  // ../RTL/cmsdk_iop_gpio.v(564)
  and u637 (n306[2], reg_datain[2], reg_intpol[2]);  // ../RTL/cmsdk_iop_gpio.v(564)
  and u638 (n306[3], reg_datain[3], reg_intpol[3]);  // ../RTL/cmsdk_iop_gpio.v(564)
  and u639 (n306[4], reg_datain[4], reg_intpol[4]);  // ../RTL/cmsdk_iop_gpio.v(564)
  buf u64 (IORDATA[1], read_mux[1]);  // ../RTL/cmsdk_iop_gpio.v(577)
  and u640 (n306[5], reg_datain[5], reg_intpol[5]);  // ../RTL/cmsdk_iop_gpio.v(564)
  and u641 (n306[6], reg_datain[6], reg_intpol[6]);  // ../RTL/cmsdk_iop_gpio.v(564)
  and u642 (n306[7], reg_datain[7], reg_intpol[7]);  // ../RTL/cmsdk_iop_gpio.v(564)
  and u643 (n306[8], reg_datain[8], reg_intpol[8]);  // ../RTL/cmsdk_iop_gpio.v(564)
  and u644 (n306[9], reg_datain[9], reg_intpol[9]);  // ../RTL/cmsdk_iop_gpio.v(564)
  and u645 (n306[10], reg_datain[10], reg_intpol[10]);  // ../RTL/cmsdk_iop_gpio.v(564)
  and u646 (n306[11], reg_datain[11], reg_intpol[11]);  // ../RTL/cmsdk_iop_gpio.v(564)
  and u647 (n306[12], reg_datain[12], reg_intpol[12]);  // ../RTL/cmsdk_iop_gpio.v(564)
  and u648 (n306[13], reg_datain[13], reg_intpol[13]);  // ../RTL/cmsdk_iop_gpio.v(564)
  and u649 (n306[14], reg_datain[14], reg_intpol[14]);  // ../RTL/cmsdk_iop_gpio.v(564)
  or u65 (n39, reg_dout_normal_write1, reg_dout_masked_write1);  // ../RTL/cmsdk_iop_gpio.v(308)
  and u650 (n306[15], reg_datain[15], reg_intpol[15]);  // ../RTL/cmsdk_iop_gpio.v(564)
  and u651 (n10[1], reg_datain32[1], IOADDR[3]);  // ../RTL/cmsdk_iop_gpio.v(175)
  and u652 (n10[2], reg_datain32[2], IOADDR[4]);  // ../RTL/cmsdk_iop_gpio.v(175)
  and u653 (n10[3], reg_datain32[3], IOADDR[5]);  // ../RTL/cmsdk_iop_gpio.v(175)
  and u654 (n10[4], reg_datain32[4], IOADDR[6]);  // ../RTL/cmsdk_iop_gpio.v(175)
  and u655 (n10[5], reg_datain32[5], IOADDR[7]);  // ../RTL/cmsdk_iop_gpio.v(175)
  and u656 (n10[6], reg_datain32[6], IOADDR[8]);  // ../RTL/cmsdk_iop_gpio.v(175)
  and u657 (n10[7], reg_datain32[7], IOADDR[9]);  // ../RTL/cmsdk_iop_gpio.v(175)
  and u658 (n11[0], reg_datain32[8], IOADDR[2]);  // ../RTL/cmsdk_iop_gpio.v(175)
  and u659 (n11[1], reg_datain32[9], IOADDR[3]);  // ../RTL/cmsdk_iop_gpio.v(175)
  or u66 (new_raw_int[9], n335[9], fall_edge_int[9]);  // ../RTL/cmsdk_iop_gpio.v(568)
  and u660 (n11[2], reg_datain32[10], IOADDR[4]);  // ../RTL/cmsdk_iop_gpio.v(175)
  and u661 (n11[3], reg_datain32[11], IOADDR[5]);  // ../RTL/cmsdk_iop_gpio.v(175)
  and u662 (n11[4], reg_datain32[12], IOADDR[6]);  // ../RTL/cmsdk_iop_gpio.v(175)
  and u663 (n11[5], reg_datain32[13], IOADDR[7]);  // ../RTL/cmsdk_iop_gpio.v(175)
  and u664 (n11[6], reg_datain32[14], IOADDR[8]);  // ../RTL/cmsdk_iop_gpio.v(175)
  and u665 (n11[7], reg_datain32[15], IOADDR[9]);  // ../RTL/cmsdk_iop_gpio.v(175)
  or u666 (n311, reg_inttype[2], reg_inttype[3]);  // ../RTL/cmsdk_iop_gpio.v(560)
  or u667 (n303, n312, n311);  // ../RTL/cmsdk_iop_gpio.v(560)
  or u668 (n270, reg_inttype[4], reg_inttype[5]);  // ../RTL/cmsdk_iop_gpio.v(560)
  or u669 (n269, reg_inttype[6], reg_inttype[7]);  // ../RTL/cmsdk_iop_gpio.v(560)
  or u67 (new_raw_int[10], n335[10], fall_edge_int[10]);  // ../RTL/cmsdk_iop_gpio.v(568)
  or u670 (n268, n270, n269);  // ../RTL/cmsdk_iop_gpio.v(560)
  or u671 (n233, n303, n268);  // ../RTL/cmsdk_iop_gpio.v(560)
  or u672 (n231, reg_inttype[8], reg_inttype[9]);  // ../RTL/cmsdk_iop_gpio.v(560)
  or u673 (n230, reg_inttype[10], reg_inttype[11]);  // ../RTL/cmsdk_iop_gpio.v(560)
  or u674 (n225, n231, n230);  // ../RTL/cmsdk_iop_gpio.v(560)
  or u675 (n224, reg_inttype[12], reg_inttype[13]);  // ../RTL/cmsdk_iop_gpio.v(560)
  or u676 (n188, reg_inttype[14], reg_inttype[15]);  // ../RTL/cmsdk_iop_gpio.v(560)
  or u677 (n186, n224, n188);  // ../RTL/cmsdk_iop_gpio.v(560)
  or u678 (n185, n225, n186);  // ../RTL/cmsdk_iop_gpio.v(560)
  or u679 (n304, n233, n185);  // ../RTL/cmsdk_iop_gpio.v(560)
  or u68 (new_raw_int[11], n335[11], fall_edge_int[11]);  // ../RTL/cmsdk_iop_gpio.v(568)
  buf u680 (reg_intstat[1], reg_intstat_padded[1]);  // ../RTL/cmsdk_iop_gpio.v(542)
  buf u681 (reg_intstat[2], reg_intstat_padded[2]);  // ../RTL/cmsdk_iop_gpio.v(542)
  buf u682 (reg_intstat[3], reg_intstat_padded[3]);  // ../RTL/cmsdk_iop_gpio.v(542)
  buf u683 (reg_intstat[4], reg_intstat_padded[4]);  // ../RTL/cmsdk_iop_gpio.v(542)
  buf u684 (reg_intstat[5], reg_intstat_padded[5]);  // ../RTL/cmsdk_iop_gpio.v(542)
  buf u685 (reg_intstat[6], reg_intstat_padded[6]);  // ../RTL/cmsdk_iop_gpio.v(542)
  buf u686 (reg_intstat[7], reg_intstat_padded[7]);  // ../RTL/cmsdk_iop_gpio.v(542)
  buf u687 (reg_intstat[8], reg_intstat_padded[8]);  // ../RTL/cmsdk_iop_gpio.v(542)
  buf u688 (reg_intstat[9], reg_intstat_padded[9]);  // ../RTL/cmsdk_iop_gpio.v(542)
  buf u689 (reg_intstat[10], reg_intstat_padded[10]);  // ../RTL/cmsdk_iop_gpio.v(542)
  or u69 (new_raw_int[12], n335[12], fall_edge_int[12]);  // ../RTL/cmsdk_iop_gpio.v(568)
  buf u690 (reg_intstat[11], reg_intstat_padded[11]);  // ../RTL/cmsdk_iop_gpio.v(542)
  buf u691 (reg_intstat[12], reg_intstat_padded[12]);  // ../RTL/cmsdk_iop_gpio.v(542)
  buf u692 (reg_intstat[13], reg_intstat_padded[13]);  // ../RTL/cmsdk_iop_gpio.v(542)
  buf u693 (reg_intstat[14], reg_intstat_padded[14]);  // ../RTL/cmsdk_iop_gpio.v(542)
  buf u694 (reg_intstat[15], reg_intstat_padded[15]);  // ../RTL/cmsdk_iop_gpio.v(542)
  and u695 (new_masked_int[1], new_raw_int[1], reg_inten[1]);  // ../RTL/cmsdk_iop_gpio.v(527)
  and u696 (new_masked_int[2], new_raw_int[2], reg_inten[2]);  // ../RTL/cmsdk_iop_gpio.v(527)
  and u697 (new_masked_int[3], new_raw_int[3], reg_inten[3]);  // ../RTL/cmsdk_iop_gpio.v(527)
  and u698 (new_masked_int[4], new_raw_int[4], reg_inten[4]);  // ../RTL/cmsdk_iop_gpio.v(527)
  and u699 (new_masked_int[5], new_raw_int[5], reg_inten[5]);  // ../RTL/cmsdk_iop_gpio.v(527)
  or u7 (n335[3], n334[3], rise_edge_int[3]);  // ../RTL/cmsdk_iop_gpio.v(568)
  or u70 (new_raw_int[13], n335[13], fall_edge_int[13]);  // ../RTL/cmsdk_iop_gpio.v(568)
  and u700 (new_masked_int[6], new_raw_int[6], reg_inten[6]);  // ../RTL/cmsdk_iop_gpio.v(527)
  and u701 (new_masked_int[7], new_raw_int[7], reg_inten[7]);  // ../RTL/cmsdk_iop_gpio.v(527)
  and u702 (new_masked_int[8], new_raw_int[8], reg_inten[8]);  // ../RTL/cmsdk_iop_gpio.v(527)
  and u703 (new_masked_int[9], new_raw_int[9], reg_inten[9]);  // ../RTL/cmsdk_iop_gpio.v(527)
  and u704 (new_masked_int[10], new_raw_int[10], reg_inten[10]);  // ../RTL/cmsdk_iop_gpio.v(527)
  and u705 (new_masked_int[11], new_raw_int[11], reg_inten[11]);  // ../RTL/cmsdk_iop_gpio.v(527)
  and u706 (new_masked_int[12], new_raw_int[12], reg_inten[12]);  // ../RTL/cmsdk_iop_gpio.v(527)
  and u707 (new_masked_int[13], new_raw_int[13], reg_inten[13]);  // ../RTL/cmsdk_iop_gpio.v(527)
  and u708 (new_masked_int[14], new_raw_int[14], reg_inten[14]);  // ../RTL/cmsdk_iop_gpio.v(527)
  and u709 (new_masked_int[15], new_raw_int[15], reg_inten[15]);  // ../RTL/cmsdk_iop_gpio.v(527)
  or u71 (new_raw_int[14], n335[14], fall_edge_int[14]);  // ../RTL/cmsdk_iop_gpio.v(568)
  not u710 (n309[1], reg_intpol[1]);  // ../RTL/cmsdk_iop_gpio.v(565)
  not u711 (n309[2], reg_intpol[2]);  // ../RTL/cmsdk_iop_gpio.v(565)
  not u712 (n309[3], reg_intpol[3]);  // ../RTL/cmsdk_iop_gpio.v(565)
  not u713 (n309[4], reg_intpol[4]);  // ../RTL/cmsdk_iop_gpio.v(565)
  not u714 (n309[5], reg_intpol[5]);  // ../RTL/cmsdk_iop_gpio.v(565)
  not u715 (n309[6], reg_intpol[6]);  // ../RTL/cmsdk_iop_gpio.v(565)
  not u716 (n309[7], reg_intpol[7]);  // ../RTL/cmsdk_iop_gpio.v(565)
  not u717 (n309[8], reg_intpol[8]);  // ../RTL/cmsdk_iop_gpio.v(565)
  not u718 (n309[9], reg_intpol[9]);  // ../RTL/cmsdk_iop_gpio.v(565)
  not u719 (n309[10], reg_intpol[10]);  // ../RTL/cmsdk_iop_gpio.v(565)
  or u72 (new_raw_int[15], n335[15], fall_edge_int[15]);  // ../RTL/cmsdk_iop_gpio.v(568)
  not u720 (n309[11], reg_intpol[11]);  // ../RTL/cmsdk_iop_gpio.v(565)
  not u721 (n309[12], reg_intpol[12]);  // ../RTL/cmsdk_iop_gpio.v(565)
  not u722 (n309[13], reg_intpol[13]);  // ../RTL/cmsdk_iop_gpio.v(565)
  not u723 (n309[14], reg_intpol[14]);  // ../RTL/cmsdk_iop_gpio.v(565)
  not u724 (n309[15], reg_intpol[15]);  // ../RTL/cmsdk_iop_gpio.v(565)
  not u725 (n308[0], reg_datain[0]);  // ../RTL/cmsdk_iop_gpio.v(565)
  not u726 (n308[1], reg_datain[1]);  // ../RTL/cmsdk_iop_gpio.v(565)
  not u727 (n308[2], reg_datain[2]);  // ../RTL/cmsdk_iop_gpio.v(565)
  not u728 (n308[3], reg_datain[3]);  // ../RTL/cmsdk_iop_gpio.v(565)
  not u729 (n308[4], reg_datain[4]);  // ../RTL/cmsdk_iop_gpio.v(565)
  buf u73 (PORTOUT[2], reg_dout[2]);  // ../RTL/cmsdk_iop_gpio.v(573)
  not u730 (n308[5], reg_datain[5]);  // ../RTL/cmsdk_iop_gpio.v(565)
  not u731 (n308[6], reg_datain[6]);  // ../RTL/cmsdk_iop_gpio.v(565)
  not u732 (n308[7], reg_datain[7]);  // ../RTL/cmsdk_iop_gpio.v(565)
  not u733 (n308[8], reg_datain[8]);  // ../RTL/cmsdk_iop_gpio.v(565)
  not u734 (n308[9], reg_datain[9]);  // ../RTL/cmsdk_iop_gpio.v(565)
  not u735 (n308[10], reg_datain[10]);  // ../RTL/cmsdk_iop_gpio.v(565)
  not u736 (n308[11], reg_datain[11]);  // ../RTL/cmsdk_iop_gpio.v(565)
  not u737 (n308[12], reg_datain[12]);  // ../RTL/cmsdk_iop_gpio.v(565)
  not u738 (n308[13], reg_datain[13]);  // ../RTL/cmsdk_iop_gpio.v(565)
  not u739 (n308[14], reg_datain[14]);  // ../RTL/cmsdk_iop_gpio.v(565)
  buf u74 (PORTOUT[3], reg_dout[3]);  // ../RTL/cmsdk_iop_gpio.v(573)
  not u740 (n308[15], reg_datain[15]);  // ../RTL/cmsdk_iop_gpio.v(565)
  buf u741 (reg_intpol[1], reg_intpol_padded[1]);  // ../RTL/cmsdk_iop_gpio.v(504)
  buf u742 (reg_intpol[2], reg_intpol_padded[2]);  // ../RTL/cmsdk_iop_gpio.v(504)
  buf u743 (reg_intpol[3], reg_intpol_padded[3]);  // ../RTL/cmsdk_iop_gpio.v(504)
  buf u744 (reg_intpol[4], reg_intpol_padded[4]);  // ../RTL/cmsdk_iop_gpio.v(504)
  buf u745 (reg_intpol[5], reg_intpol_padded[5]);  // ../RTL/cmsdk_iop_gpio.v(504)
  buf u746 (reg_intpol[6], reg_intpol_padded[6]);  // ../RTL/cmsdk_iop_gpio.v(504)
  buf u747 (reg_intpol[7], reg_intpol_padded[7]);  // ../RTL/cmsdk_iop_gpio.v(504)
  buf u748 (reg_intpol[8], reg_intpol_padded[8]);  // ../RTL/cmsdk_iop_gpio.v(504)
  buf u749 (reg_intpol[9], reg_intpol_padded[9]);  // ../RTL/cmsdk_iop_gpio.v(504)
  buf u75 (PORTOUT[4], reg_dout[4]);  // ../RTL/cmsdk_iop_gpio.v(573)
  buf u750 (reg_intpol[10], reg_intpol_padded[10]);  // ../RTL/cmsdk_iop_gpio.v(504)
  buf u751 (reg_intpol[11], reg_intpol_padded[11]);  // ../RTL/cmsdk_iop_gpio.v(504)
  buf u752 (reg_intpol[12], reg_intpol_padded[12]);  // ../RTL/cmsdk_iop_gpio.v(504)
  buf u753 (reg_intpol[13], reg_intpol_padded[13]);  // ../RTL/cmsdk_iop_gpio.v(504)
  buf u754 (reg_intpol[14], reg_intpol_padded[14]);  // ../RTL/cmsdk_iop_gpio.v(504)
  buf u755 (reg_intpol[15], reg_intpol_padded[15]);  // ../RTL/cmsdk_iop_gpio.v(504)
  buf u756 (reg_inttype[1], reg_inttype_padded[1]);  // ../RTL/cmsdk_iop_gpio.v(466)
  buf u757 (reg_inttype[2], reg_inttype_padded[2]);  // ../RTL/cmsdk_iop_gpio.v(466)
  buf u758 (reg_inttype[3], reg_inttype_padded[3]);  // ../RTL/cmsdk_iop_gpio.v(466)
  buf u759 (reg_inttype[4], reg_inttype_padded[4]);  // ../RTL/cmsdk_iop_gpio.v(466)
  buf u76 (PORTOUT[5], reg_dout[5]);  // ../RTL/cmsdk_iop_gpio.v(573)
  buf u760 (reg_inttype[5], reg_inttype_padded[5]);  // ../RTL/cmsdk_iop_gpio.v(466)
  buf u761 (reg_inttype[6], reg_inttype_padded[6]);  // ../RTL/cmsdk_iop_gpio.v(466)
  buf u762 (reg_inttype[7], reg_inttype_padded[7]);  // ../RTL/cmsdk_iop_gpio.v(466)
  buf u763 (reg_inttype[8], reg_inttype_padded[8]);  // ../RTL/cmsdk_iop_gpio.v(466)
  buf u764 (reg_inttype[9], reg_inttype_padded[9]);  // ../RTL/cmsdk_iop_gpio.v(466)
  buf u765 (reg_inttype[10], reg_inttype_padded[10]);  // ../RTL/cmsdk_iop_gpio.v(466)
  buf u766 (reg_inttype[11], reg_inttype_padded[11]);  // ../RTL/cmsdk_iop_gpio.v(466)
  buf u767 (reg_inttype[12], reg_inttype_padded[12]);  // ../RTL/cmsdk_iop_gpio.v(466)
  buf u768 (reg_inttype[13], reg_inttype_padded[13]);  // ../RTL/cmsdk_iop_gpio.v(466)
  buf u769 (reg_inttype[14], reg_inttype_padded[14]);  // ../RTL/cmsdk_iop_gpio.v(466)
  buf u77 (PORTOUT[6], reg_dout[6]);  // ../RTL/cmsdk_iop_gpio.v(573)
  buf u770 (reg_inttype[15], reg_inttype_padded[15]);  // ../RTL/cmsdk_iop_gpio.v(466)
  buf u771 (reg_inten[1], reg_inten_padded[1]);  // ../RTL/cmsdk_iop_gpio.v(428)
  buf u772 (reg_inten[2], reg_inten_padded[2]);  // ../RTL/cmsdk_iop_gpio.v(428)
  buf u773 (reg_inten[3], reg_inten_padded[3]);  // ../RTL/cmsdk_iop_gpio.v(428)
  buf u774 (reg_inten[4], reg_inten_padded[4]);  // ../RTL/cmsdk_iop_gpio.v(428)
  buf u775 (reg_inten[5], reg_inten_padded[5]);  // ../RTL/cmsdk_iop_gpio.v(428)
  buf u776 (reg_inten[6], reg_inten_padded[6]);  // ../RTL/cmsdk_iop_gpio.v(428)
  buf u777 (reg_inten[7], reg_inten_padded[7]);  // ../RTL/cmsdk_iop_gpio.v(428)
  buf u778 (reg_inten[8], reg_inten_padded[8]);  // ../RTL/cmsdk_iop_gpio.v(428)
  buf u779 (reg_inten[9], reg_inten_padded[9]);  // ../RTL/cmsdk_iop_gpio.v(428)
  buf u78 (PORTOUT[7], reg_dout[7]);  // ../RTL/cmsdk_iop_gpio.v(573)
  buf u780 (reg_inten[10], reg_inten_padded[10]);  // ../RTL/cmsdk_iop_gpio.v(428)
  buf u781 (reg_inten[11], reg_inten_padded[11]);  // ../RTL/cmsdk_iop_gpio.v(428)
  buf u782 (reg_inten[12], reg_inten_padded[12]);  // ../RTL/cmsdk_iop_gpio.v(428)
  buf u783 (reg_inten[13], reg_inten_padded[13]);  // ../RTL/cmsdk_iop_gpio.v(428)
  buf u784 (reg_inten[14], reg_inten_padded[14]);  // ../RTL/cmsdk_iop_gpio.v(428)
  buf u785 (reg_inten[15], reg_inten_padded[15]);  // ../RTL/cmsdk_iop_gpio.v(428)
  buf u786 (reg_altfunc[1], reg_altfunc_padded[1]);  // ../RTL/cmsdk_iop_gpio.v(390)
  buf u787 (reg_altfunc[2], reg_altfunc_padded[2]);  // ../RTL/cmsdk_iop_gpio.v(390)
  buf u788 (reg_altfunc[3], reg_altfunc_padded[3]);  // ../RTL/cmsdk_iop_gpio.v(390)
  buf u789 (reg_altfunc[4], reg_altfunc_padded[4]);  // ../RTL/cmsdk_iop_gpio.v(390)
  buf u79 (PORTOUT[8], reg_dout[8]);  // ../RTL/cmsdk_iop_gpio.v(573)
  buf u790 (reg_altfunc[5], reg_altfunc_padded[5]);  // ../RTL/cmsdk_iop_gpio.v(390)
  buf u791 (reg_altfunc[6], reg_altfunc_padded[6]);  // ../RTL/cmsdk_iop_gpio.v(390)
  buf u792 (reg_altfunc[7], reg_altfunc_padded[7]);  // ../RTL/cmsdk_iop_gpio.v(390)
  buf u793 (reg_altfunc[8], reg_altfunc_padded[8]);  // ../RTL/cmsdk_iop_gpio.v(390)
  buf u794 (reg_altfunc[9], reg_altfunc_padded[9]);  // ../RTL/cmsdk_iop_gpio.v(390)
  buf u795 (reg_altfunc[10], reg_altfunc_padded[10]);  // ../RTL/cmsdk_iop_gpio.v(390)
  buf u796 (reg_altfunc[11], reg_altfunc_padded[11]);  // ../RTL/cmsdk_iop_gpio.v(390)
  buf u797 (reg_altfunc[12], reg_altfunc_padded[12]);  // ../RTL/cmsdk_iop_gpio.v(390)
  buf u798 (reg_altfunc[13], reg_altfunc_padded[13]);  // ../RTL/cmsdk_iop_gpio.v(390)
  buf u799 (reg_altfunc[14], reg_altfunc_padded[14]);  // ../RTL/cmsdk_iop_gpio.v(390)
  or u8 (n335[4], n334[4], rise_edge_int[4]);  // ../RTL/cmsdk_iop_gpio.v(568)
  or u80 (n38[0], n36[0], n37[0]);  // ../RTL/cmsdk_iop_gpio.v(301)
  buf u800 (reg_altfunc[15], reg_altfunc_padded[15]);  // ../RTL/cmsdk_iop_gpio.v(390)
  buf u801 (reg_douten[1], reg_douten_padded[1]);  // ../RTL/cmsdk_iop_gpio.v(351)
  buf u802 (reg_douten[2], reg_douten_padded[2]);  // ../RTL/cmsdk_iop_gpio.v(351)
  buf u803 (reg_douten[3], reg_douten_padded[3]);  // ../RTL/cmsdk_iop_gpio.v(351)
  buf u804 (reg_douten[4], reg_douten_padded[4]);  // ../RTL/cmsdk_iop_gpio.v(351)
  buf u805 (reg_douten[5], reg_douten_padded[5]);  // ../RTL/cmsdk_iop_gpio.v(351)
  buf u806 (reg_douten[6], reg_douten_padded[6]);  // ../RTL/cmsdk_iop_gpio.v(351)
  buf u807 (reg_douten[7], reg_douten_padded[7]);  // ../RTL/cmsdk_iop_gpio.v(351)
  buf u808 (reg_douten[8], reg_douten_padded[8]);  // ../RTL/cmsdk_iop_gpio.v(351)
  buf u809 (reg_douten[9], reg_douten_padded[9]);  // ../RTL/cmsdk_iop_gpio.v(351)
  buf u81 (PORTEN[8], reg_douten[8]);  // ../RTL/cmsdk_iop_gpio.v(574)
  buf u810 (reg_douten[10], reg_douten_padded[10]);  // ../RTL/cmsdk_iop_gpio.v(351)
  buf u811 (reg_douten[11], reg_douten_padded[11]);  // ../RTL/cmsdk_iop_gpio.v(351)
  buf u812 (reg_douten[12], reg_douten_padded[12]);  // ../RTL/cmsdk_iop_gpio.v(351)
  buf u813 (reg_douten[13], reg_douten_padded[13]);  // ../RTL/cmsdk_iop_gpio.v(351)
  buf u814 (reg_douten[14], reg_douten_padded[14]);  // ../RTL/cmsdk_iop_gpio.v(351)
  buf u815 (reg_douten[15], reg_douten_padded[15]);  // ../RTL/cmsdk_iop_gpio.v(351)
  buf u816 (reg_dout[1], reg_dout_padded[1]);  // ../RTL/cmsdk_iop_gpio.v(312)
  buf u817 (reg_dout[2], reg_dout_padded[2]);  // ../RTL/cmsdk_iop_gpio.v(312)
  buf u818 (reg_dout[3], reg_dout_padded[3]);  // ../RTL/cmsdk_iop_gpio.v(312)
  buf u819 (reg_dout[4], reg_dout_padded[4]);  // ../RTL/cmsdk_iop_gpio.v(312)
  and u82 (n42, write_trans, n41);  // ../RTL/cmsdk_iop_gpio.v(325)
  buf u820 (reg_dout[5], reg_dout_padded[5]);  // ../RTL/cmsdk_iop_gpio.v(312)
  buf u821 (reg_dout[6], reg_dout_padded[6]);  // ../RTL/cmsdk_iop_gpio.v(312)
  buf u822 (reg_dout[7], reg_dout_padded[7]);  // ../RTL/cmsdk_iop_gpio.v(312)
  buf u823 (reg_dout[8], reg_dout_padded[8]);  // ../RTL/cmsdk_iop_gpio.v(312)
  buf u824 (reg_dout[9], reg_dout_padded[9]);  // ../RTL/cmsdk_iop_gpio.v(312)
  buf u825 (reg_dout[10], reg_dout_padded[10]);  // ../RTL/cmsdk_iop_gpio.v(312)
  buf u826 (reg_dout[11], reg_dout_padded[11]);  // ../RTL/cmsdk_iop_gpio.v(312)
  buf u827 (reg_dout[12], reg_dout_padded[12]);  // ../RTL/cmsdk_iop_gpio.v(312)
  buf u828 (reg_dout[13], reg_dout_padded[13]);  // ../RTL/cmsdk_iop_gpio.v(312)
  buf u829 (reg_dout[14], reg_dout_padded[14]);  // ../RTL/cmsdk_iop_gpio.v(312)
  buf u83 (PORTEN[7], reg_douten[7]);  // ../RTL/cmsdk_iop_gpio.v(574)
  buf u830 (reg_dout[15], reg_dout_padded[15]);  // ../RTL/cmsdk_iop_gpio.v(312)
  or u831 (n38[1], n36[1], n37[1]);  // ../RTL/cmsdk_iop_gpio.v(301)
  or u832 (n38[2], n36[2], n37[2]);  // ../RTL/cmsdk_iop_gpio.v(301)
  or u833 (n38[3], n36[3], n37[3]);  // ../RTL/cmsdk_iop_gpio.v(301)
  or u834 (n38[4], n36[4], n37[4]);  // ../RTL/cmsdk_iop_gpio.v(301)
  or u835 (n38[5], n36[5], n37[5]);  // ../RTL/cmsdk_iop_gpio.v(301)
  or u836 (n38[6], n36[6], n37[6]);  // ../RTL/cmsdk_iop_gpio.v(301)
  or u837 (n38[7], n36[7], n37[7]);  // ../RTL/cmsdk_iop_gpio.v(301)
  and u838 (n32[1], current_dout_padded[1], n31[1]);  // ../RTL/cmsdk_iop_gpio.v(286)
  and u839 (n32[2], current_dout_padded[2], n31[2]);  // ../RTL/cmsdk_iop_gpio.v(286)
  and u84 (n43, n42, iop_byte_strobe[0]);  // ../RTL/cmsdk_iop_gpio.v(326)
  and u840 (n32[3], current_dout_padded[3], n31[3]);  // ../RTL/cmsdk_iop_gpio.v(286)
  and u841 (n32[4], current_dout_padded[4], n31[4]);  // ../RTL/cmsdk_iop_gpio.v(286)
  and u842 (n32[5], current_dout_padded[5], n31[5]);  // ../RTL/cmsdk_iop_gpio.v(286)
  and u843 (n32[6], current_dout_padded[6], n31[6]);  // ../RTL/cmsdk_iop_gpio.v(286)
  and u844 (n32[7], current_dout_padded[7], n31[7]);  // ../RTL/cmsdk_iop_gpio.v(286)
  and u845 (n30[0], IOWDATALE[0], IOADDR[2]);  // ../RTL/cmsdk_iop_gpio.v(286)
  and u846 (n30[1], IOWDATALE[1], IOADDR[3]);  // ../RTL/cmsdk_iop_gpio.v(286)
  and u847 (n30[2], IOWDATALE[2], IOADDR[4]);  // ../RTL/cmsdk_iop_gpio.v(286)
  and u848 (n30[3], IOWDATALE[3], IOADDR[5]);  // ../RTL/cmsdk_iop_gpio.v(286)
  and u849 (n30[4], IOWDATALE[4], IOADDR[6]);  // ../RTL/cmsdk_iop_gpio.v(286)
  buf u85 (PORTEN[6], reg_douten[6]);  // ../RTL/cmsdk_iop_gpio.v(574)
  and u850 (n30[5], IOWDATALE[5], IOADDR[7]);  // ../RTL/cmsdk_iop_gpio.v(286)
  and u851 (n30[6], IOWDATALE[6], IOADDR[8]);  // ../RTL/cmsdk_iop_gpio.v(286)
  and u852 (n30[7], IOWDATALE[7], IOADDR[9]);  // ../RTL/cmsdk_iop_gpio.v(286)
  and u853 (reg_intclr_padded[1], reg_intclr_normal_write0, IOWDATALE[1]);  // ../RTL/cmsdk_iop_gpio.v(525)
  and u854 (reg_intclr_padded[2], reg_intclr_normal_write0, IOWDATALE[2]);  // ../RTL/cmsdk_iop_gpio.v(525)
  and u855 (reg_intclr_padded[3], reg_intclr_normal_write0, IOWDATALE[3]);  // ../RTL/cmsdk_iop_gpio.v(525)
  and u856 (reg_intclr_padded[4], reg_intclr_normal_write0, IOWDATALE[4]);  // ../RTL/cmsdk_iop_gpio.v(525)
  and u857 (reg_intclr_padded[5], reg_intclr_normal_write0, IOWDATALE[5]);  // ../RTL/cmsdk_iop_gpio.v(525)
  and u858 (reg_intclr_padded[6], reg_intclr_normal_write0, IOWDATALE[6]);  // ../RTL/cmsdk_iop_gpio.v(525)
  and u859 (reg_intclr_padded[7], reg_intclr_normal_write0, IOWDATALE[7]);  // ../RTL/cmsdk_iop_gpio.v(525)
  buf u86 (GPIOINT[15], reg_intstat[15]);  // ../RTL/cmsdk_iop_gpio.v(580)
  and u860 (reg_intclr_padded[8], reg_intclr_normal_write1, IOWDATALE[8]);  // ../RTL/cmsdk_iop_gpio.v(525)
  and u861 (reg_intclr_padded[9], reg_intclr_normal_write1, IOWDATALE[9]);  // ../RTL/cmsdk_iop_gpio.v(525)
  and u862 (reg_intclr_padded[10], reg_intclr_normal_write1, IOWDATALE[10]);  // ../RTL/cmsdk_iop_gpio.v(525)
  and u863 (reg_intclr_padded[11], reg_intclr_normal_write1, IOWDATALE[11]);  // ../RTL/cmsdk_iop_gpio.v(525)
  and u864 (reg_intclr_padded[12], reg_intclr_normal_write1, IOWDATALE[12]);  // ../RTL/cmsdk_iop_gpio.v(525)
  and u865 (reg_intclr_padded[13], reg_intclr_normal_write1, IOWDATALE[13]);  // ../RTL/cmsdk_iop_gpio.v(525)
  and u866 (reg_intclr_padded[14], reg_intclr_normal_write1, IOWDATALE[14]);  // ../RTL/cmsdk_iop_gpio.v(525)
  and u867 (reg_intclr_padded[15], reg_intclr_normal_write1, IOWDATALE[15]);  // ../RTL/cmsdk_iop_gpio.v(525)
  or u868 (n33[1], n30[1], n32[1]);  // ../RTL/cmsdk_iop_gpio.v(286)
  or u869 (n33[2], n30[2], n32[2]);  // ../RTL/cmsdk_iop_gpio.v(286)
  buf u87 (GPIOINT[14], reg_intstat[14]);  // ../RTL/cmsdk_iop_gpio.v(580)
  or u870 (n33[3], n30[3], n32[3]);  // ../RTL/cmsdk_iop_gpio.v(286)
  or u871 (n33[4], n30[4], n32[4]);  // ../RTL/cmsdk_iop_gpio.v(286)
  or u872 (n33[5], n30[5], n32[5]);  // ../RTL/cmsdk_iop_gpio.v(286)
  or u873 (n33[6], n30[6], n32[6]);  // ../RTL/cmsdk_iop_gpio.v(286)
  or u874 (n33[7], n30[7], n32[7]);  // ../RTL/cmsdk_iop_gpio.v(286)
  not u875 (n31[1], IOADDR[3]);  // ../RTL/cmsdk_iop_gpio.v(286)
  not u876 (n31[2], IOADDR[4]);  // ../RTL/cmsdk_iop_gpio.v(286)
  not u877 (n31[3], IOADDR[5]);  // ../RTL/cmsdk_iop_gpio.v(286)
  not u878 (n31[4], IOADDR[6]);  // ../RTL/cmsdk_iop_gpio.v(286)
  not u879 (n31[5], IOADDR[7]);  // ../RTL/cmsdk_iop_gpio.v(286)
  buf u88 (PORTEN[5], reg_douten[5]);  // ../RTL/cmsdk_iop_gpio.v(574)
  not u880 (n31[6], IOADDR[8]);  // ../RTL/cmsdk_iop_gpio.v(286)
  not u881 (n31[7], IOADDR[9]);  // ../RTL/cmsdk_iop_gpio.v(286)
  buf u882 (current_dout_padded[1], reg_dout[1]);  // ../RTL/cmsdk_iop_gpio.v(280)
  buf u883 (current_dout_padded[2], reg_dout[2]);  // ../RTL/cmsdk_iop_gpio.v(280)
  buf u884 (current_dout_padded[3], reg_dout[3]);  // ../RTL/cmsdk_iop_gpio.v(280)
  buf u885 (current_dout_padded[4], reg_dout[4]);  // ../RTL/cmsdk_iop_gpio.v(280)
  buf u886 (current_dout_padded[5], reg_dout[5]);  // ../RTL/cmsdk_iop_gpio.v(280)
  buf u887 (current_dout_padded[6], reg_dout[6]);  // ../RTL/cmsdk_iop_gpio.v(280)
  buf u888 (current_dout_padded[7], reg_dout[7]);  // ../RTL/cmsdk_iop_gpio.v(280)
  buf u889 (current_dout_padded[8], reg_dout[8]);  // ../RTL/cmsdk_iop_gpio.v(280)
  and u89 (n46, n42, iop_byte_strobe[1]);  // ../RTL/cmsdk_iop_gpio.v(329)
  buf u890 (current_dout_padded[9], reg_dout[9]);  // ../RTL/cmsdk_iop_gpio.v(280)
  buf u891 (current_dout_padded[10], reg_dout[10]);  // ../RTL/cmsdk_iop_gpio.v(280)
  buf u892 (current_dout_padded[11], reg_dout[11]);  // ../RTL/cmsdk_iop_gpio.v(280)
  buf u893 (current_dout_padded[12], reg_dout[12]);  // ../RTL/cmsdk_iop_gpio.v(280)
  buf u894 (current_dout_padded[13], reg_dout[13]);  // ../RTL/cmsdk_iop_gpio.v(280)
  buf u895 (current_dout_padded[14], reg_dout[14]);  // ../RTL/cmsdk_iop_gpio.v(280)
  buf u896 (current_dout_padded[15], reg_dout[15]);  // ../RTL/cmsdk_iop_gpio.v(280)
  buf u897 (n180, 1'b0);  // ../RTL/cmsdk_iop_gpio.v(280)
  buf u898 (n179, 1'b0);  // ../RTL/cmsdk_iop_gpio.v(280)
  buf u899 (n143, 1'b0);  // ../RTL/cmsdk_iop_gpio.v(280)
  or u9 (n335[5], n334[5], rise_edge_int[5]);  // ../RTL/cmsdk_iop_gpio.v(568)
  buf u90 (PORTEN[4], reg_douten[4]);  // ../RTL/cmsdk_iop_gpio.v(574)
  buf u900 (n141, 1'b0);  // ../RTL/cmsdk_iop_gpio.v(280)
  buf u901 (n140, 1'b0);  // ../RTL/cmsdk_iop_gpio.v(280)
  buf u902 (n135, 1'b0);  // ../RTL/cmsdk_iop_gpio.v(280)
  buf u903 (n134, 1'b0);  // ../RTL/cmsdk_iop_gpio.v(280)
  buf u904 (n98, 1'b0);  // ../RTL/cmsdk_iop_gpio.v(280)
  buf u905 (n96, 1'b0);  // ../RTL/cmsdk_iop_gpio.v(280)
  buf u906 (n95, 1'b0);  // ../RTL/cmsdk_iop_gpio.v(280)
  buf u907 (n90, 1'b0);  // ../RTL/cmsdk_iop_gpio.v(280)
  buf u908 (n89, 1'b0);  // ../RTL/cmsdk_iop_gpio.v(280)
  buf u909 (n53, 1'b0);  // ../RTL/cmsdk_iop_gpio.v(280)
  and u91 (n48, write_trans, n47);  // ../RTL/cmsdk_iop_gpio.v(331)
  buf u910 (n51, 1'b0);  // ../RTL/cmsdk_iop_gpio.v(280)
  buf u911 (n50, 1'b0);  // ../RTL/cmsdk_iop_gpio.v(280)
  buf u912 (n45, 1'b0);  // ../RTL/cmsdk_iop_gpio.v(280)
  buf u913 (n44, 1'b0);  // ../RTL/cmsdk_iop_gpio.v(280)
  buf u914 (reg_datain32[1], reg_datain[1]);  // ../RTL/cmsdk_iop_gpio.v(257)
  buf u915 (reg_datain32[2], reg_datain[2]);  // ../RTL/cmsdk_iop_gpio.v(257)
  buf u916 (reg_datain32[3], reg_datain[3]);  // ../RTL/cmsdk_iop_gpio.v(257)
  buf u917 (reg_datain32[4], reg_datain[4]);  // ../RTL/cmsdk_iop_gpio.v(257)
  buf u918 (reg_datain32[5], reg_datain[5]);  // ../RTL/cmsdk_iop_gpio.v(257)
  buf u919 (reg_datain32[6], reg_datain[6]);  // ../RTL/cmsdk_iop_gpio.v(257)
  buf u92 (PORTEN[3], reg_douten[3]);  // ../RTL/cmsdk_iop_gpio.v(574)
  buf u920 (reg_datain32[7], reg_datain[7]);  // ../RTL/cmsdk_iop_gpio.v(257)
  buf u921 (reg_datain32[8], reg_datain[8]);  // ../RTL/cmsdk_iop_gpio.v(257)
  buf u922 (reg_datain32[9], reg_datain[9]);  // ../RTL/cmsdk_iop_gpio.v(257)
  buf u923 (reg_datain32[10], reg_datain[10]);  // ../RTL/cmsdk_iop_gpio.v(257)
  buf u924 (reg_datain32[11], reg_datain[11]);  // ../RTL/cmsdk_iop_gpio.v(257)
  buf u925 (reg_datain32[12], reg_datain[12]);  // ../RTL/cmsdk_iop_gpio.v(257)
  buf u926 (reg_datain32[13], reg_datain[13]);  // ../RTL/cmsdk_iop_gpio.v(257)
  buf u927 (reg_datain32[14], reg_datain[14]);  // ../RTL/cmsdk_iop_gpio.v(257)
  buf u928 (reg_datain32[15], reg_datain[15]);  // ../RTL/cmsdk_iop_gpio.v(257)
  buf u929 (reg_datain32[16], 1'b0);  // ../RTL/cmsdk_iop_gpio.v(257)
  and u93 (n49, n48, iop_byte_strobe[0]);  // ../RTL/cmsdk_iop_gpio.v(332)
  buf u930 (reg_datain32[17], 1'b0);  // ../RTL/cmsdk_iop_gpio.v(257)
  buf u931 (reg_datain32[18], 1'b0);  // ../RTL/cmsdk_iop_gpio.v(257)
  buf u932 (reg_datain32[19], 1'b0);  // ../RTL/cmsdk_iop_gpio.v(257)
  buf u933 (reg_datain32[20], 1'b0);  // ../RTL/cmsdk_iop_gpio.v(257)
  buf u934 (reg_datain32[21], 1'b0);  // ../RTL/cmsdk_iop_gpio.v(257)
  buf u935 (reg_datain32[22], 1'b0);  // ../RTL/cmsdk_iop_gpio.v(257)
  buf u936 (reg_datain32[23], 1'b0);  // ../RTL/cmsdk_iop_gpio.v(257)
  buf u937 (reg_datain32[24], 1'b0);  // ../RTL/cmsdk_iop_gpio.v(257)
  buf u938 (reg_datain32[25], 1'b0);  // ../RTL/cmsdk_iop_gpio.v(257)
  buf u939 (reg_datain32[26], 1'b0);  // ../RTL/cmsdk_iop_gpio.v(257)
  buf u94 (PORTEN[2], reg_douten[2]);  // ../RTL/cmsdk_iop_gpio.v(574)
  buf u940 (reg_datain32[27], 1'b0);  // ../RTL/cmsdk_iop_gpio.v(257)
  buf u941 (reg_datain32[28], 1'b0);  // ../RTL/cmsdk_iop_gpio.v(257)
  buf u942 (reg_datain32[29], 1'b0);  // ../RTL/cmsdk_iop_gpio.v(257)
  buf u943 (reg_datain32[30], 1'b0);  // ../RTL/cmsdk_iop_gpio.v(257)
  buf u944 (reg_datain32[31], 1'b0);  // ../RTL/cmsdk_iop_gpio.v(257)
  buf u945 (reg_datain[1], reg_in_sync2[1]);  // ../RTL/cmsdk_iop_gpio.v(255)
  buf u946 (reg_datain[2], reg_in_sync2[2]);  // ../RTL/cmsdk_iop_gpio.v(255)
  buf u947 (reg_datain[3], reg_in_sync2[3]);  // ../RTL/cmsdk_iop_gpio.v(255)
  buf u948 (reg_datain[4], reg_in_sync2[4]);  // ../RTL/cmsdk_iop_gpio.v(255)
  buf u949 (reg_datain[5], reg_in_sync2[5]);  // ../RTL/cmsdk_iop_gpio.v(255)
  buf u95 (GPIOINT[13], reg_intstat[13]);  // ../RTL/cmsdk_iop_gpio.v(580)
  buf u950 (reg_datain[6], reg_in_sync2[6]);  // ../RTL/cmsdk_iop_gpio.v(255)
  buf u951 (reg_datain[7], reg_in_sync2[7]);  // ../RTL/cmsdk_iop_gpio.v(255)
  buf u952 (reg_datain[8], reg_in_sync2[8]);  // ../RTL/cmsdk_iop_gpio.v(255)
  buf u953 (reg_datain[9], reg_in_sync2[9]);  // ../RTL/cmsdk_iop_gpio.v(255)
  buf u954 (reg_datain[10], reg_in_sync2[10]);  // ../RTL/cmsdk_iop_gpio.v(255)
  buf u955 (reg_datain[11], reg_in_sync2[11]);  // ../RTL/cmsdk_iop_gpio.v(255)
  buf u956 (reg_datain[12], reg_in_sync2[12]);  // ../RTL/cmsdk_iop_gpio.v(255)
  buf u957 (reg_datain[13], reg_in_sync2[13]);  // ../RTL/cmsdk_iop_gpio.v(255)
  buf u958 (reg_datain[14], reg_in_sync2[14]);  // ../RTL/cmsdk_iop_gpio.v(255)
  buf u959 (reg_datain[15], reg_in_sync2[15]);  // ../RTL/cmsdk_iop_gpio.v(255)
  buf u96 (GPIOINT[12], reg_intstat[12]);  // ../RTL/cmsdk_iop_gpio.v(580)
  and u960 (iop_byte_strobe[1], n2[1], IOSEL);  // ../RTL/cmsdk_iop_gpio.v(143)
  or u961 (n2[1], n5[1], n6);  // ../RTL/cmsdk_iop_gpio.v(143)
  and u962 (n37[1], current_dout_padded[9], n31[1]);  // ../RTL/cmsdk_iop_gpio.v(301)
  and u963 (n37[2], current_dout_padded[10], n31[2]);  // ../RTL/cmsdk_iop_gpio.v(301)
  and u964 (n37[3], current_dout_padded[11], n31[3]);  // ../RTL/cmsdk_iop_gpio.v(301)
  and u965 (n37[4], current_dout_padded[12], n31[4]);  // ../RTL/cmsdk_iop_gpio.v(301)
  and u966 (n37[5], current_dout_padded[13], n31[5]);  // ../RTL/cmsdk_iop_gpio.v(301)
  and u967 (n37[6], current_dout_padded[14], n31[6]);  // ../RTL/cmsdk_iop_gpio.v(301)
  and u968 (n37[7], current_dout_padded[15], n31[7]);  // ../RTL/cmsdk_iop_gpio.v(301)
  and u969 (n36[0], IOWDATALE[8], IOADDR[2]);  // ../RTL/cmsdk_iop_gpio.v(301)
  buf u97 (PORTEN[1], reg_douten[1]);  // ../RTL/cmsdk_iop_gpio.v(574)
  and u970 (n36[1], IOWDATALE[9], IOADDR[3]);  // ../RTL/cmsdk_iop_gpio.v(301)
  and u971 (n36[2], IOWDATALE[10], IOADDR[4]);  // ../RTL/cmsdk_iop_gpio.v(301)
  and u972 (n36[3], IOWDATALE[11], IOADDR[5]);  // ../RTL/cmsdk_iop_gpio.v(301)
  and u973 (n36[4], IOWDATALE[12], IOADDR[6]);  // ../RTL/cmsdk_iop_gpio.v(301)
  and u974 (n36[5], IOWDATALE[13], IOADDR[7]);  // ../RTL/cmsdk_iop_gpio.v(301)
  and u975 (n36[6], IOWDATALE[14], IOADDR[8]);  // ../RTL/cmsdk_iop_gpio.v(301)
  and u976 (n36[7], IOWDATALE[15], IOADDR[9]);  // ../RTL/cmsdk_iop_gpio.v(301)
  and u98 (n52, n48, iop_byte_strobe[1]);  // ../RTL/cmsdk_iop_gpio.v(335)
  buf u99 (PORTFUNC[15], reg_altfunc[15]);  // ../RTL/cmsdk_iop_gpio.v(575)

endmodule 

module binary_mux_s1_w10
  (
  i0,
  i1,
  sel,
  o
  );

  input [9:0] i0;
  input [9:0] i1;
  input sel;
  output [9:0] o;



endmodule 

module reg_ar_as_w10
  (
  clk,
  d,
  en,
  reset,
  set,
  q
  );

  input clk;
  input [9:0] d;
  input en;
  input [9:0] reset;
  input [9:0] set;
  output [9:0] q;



endmodule 

module eq_w2
  (
  i0,
  i1,
  o
  );

  input [1:0] i0;
  input [1:0] i1;
  output o;



endmodule 

module gpio  // ../RTL/gpio.v(23)
  (
  paddr,
  pclk,
  pclk_intr,
  penable,
  presetn,
  psel,
  pwdata,
  pwrite,
  gpio_intr,
  prdata,
  pready,
  pslverr,
  b_pad_gpio_porta
  );

  input [6:2] paddr;  // ../RTL/gpio.v(40)
  input pclk;  // ../RTL/gpio.v(41)
  input pclk_intr;  // ../RTL/gpio.v(42)
  input penable;  // ../RTL/gpio.v(43)
  input presetn;  // ../RTL/gpio.v(44)
  input psel;  // ../RTL/gpio.v(45)
  input [31:0] pwdata;  // ../RTL/gpio.v(46)
  input pwrite;  // ../RTL/gpio.v(47)
  output [7:0] gpio_intr;  // ../RTL/gpio.v(48)
  output [31:0] prdata;  // ../RTL/gpio.v(49)
  output pready;  // ../RTL/gpio.v(50)
  output pslverr;  // ../RTL/gpio.v(51)
  inout [7:0] b_pad_gpio_porta;  // ../RTL/gpio.v(52)

  wire [7:0] gpio_ext_porta;  // ../RTL/gpio.v(58)
  wire [7:0] gpio_ext_porta_rb;  // ../RTL/gpio.v(59)
  wire [7:0] gpio_int_polarity;  // ../RTL/gpio.v(60)
  wire [7:0] gpio_inten;  // ../RTL/gpio.v(61)
  wire [7:0] gpio_intmask;  // ../RTL/gpio.v(62)
  wire [7:0] gpio_intstatus;  // ../RTL/gpio.v(66)
  wire [7:0] gpio_inttype_level;  // ../RTL/gpio.v(67)
  wire [7:0] gpio_porta_ddr;  // ../RTL/gpio.v(69)
  wire [7:0] gpio_porta_dr;  // ../RTL/gpio.v(70)
  wire [7:0] gpio_porta_eoi;  // ../RTL/gpio.v(71)
  wire [7:0] gpio_porta_oe;  // ../RTL/gpio.v(72)
  wire [7:0] gpio_raw_intstatus;  // ../RTL/gpio.v(73)
  wire [7:0] gpio_swporta_ctl;  // ../RTL/gpio.v(74)
  wire [7:0] gpio_swporta_ddr;  // ../RTL/gpio.v(75)
  wire [7:0] gpio_swporta_dr;  // ../RTL/gpio.v(76)
  wire gpio_ls_sync;  // ../RTL/gpio.v(68)

  bufif1 u10 (b_pad_gpio_porta[3], gpio_porta_dr[3], gpio_porta_oe[3]);  // ../RTL/gpio.v(166)
  buf u11 (gpio_porta_oe[4], gpio_porta_ddr[4]);  // ../RTL/gpio.v(180)
  buf u12 (gpio_porta_oe[3], gpio_porta_ddr[3]);  // ../RTL/gpio.v(180)
  buf u13 (gpio_porta_oe[2], gpio_porta_ddr[2]);  // ../RTL/gpio.v(180)
  bufif1 u14 (b_pad_gpio_porta[4], gpio_porta_dr[4], gpio_porta_oe[4]);  // ../RTL/gpio.v(170)
  buf u15 (gpio_porta_oe[1], gpio_porta_ddr[1]);  // ../RTL/gpio.v(180)
  buf u16 (gpio_ext_porta[7], b_pad_gpio_porta[7]);  // ../RTL/gpio.v(181)
  buf u17 (gpio_ext_porta[6], b_pad_gpio_porta[6]);  // ../RTL/gpio.v(181)
  bufif1 u18 (b_pad_gpio_porta[5], gpio_porta_dr[5], gpio_porta_oe[5]);  // ../RTL/gpio.v(174)
  buf u19 (gpio_ext_porta[5], b_pad_gpio_porta[5]);  // ../RTL/gpio.v(181)
  buf u2 (pready, 1'b1);  // ../RTL/gpio.v(148)
  buf u20 (gpio_ext_porta[4], b_pad_gpio_porta[4]);  // ../RTL/gpio.v(181)
  buf u21 (gpio_ext_porta[3], b_pad_gpio_porta[3]);  // ../RTL/gpio.v(181)
  bufif1 u22 (b_pad_gpio_porta[6], gpio_porta_dr[6], gpio_porta_oe[6]);  // ../RTL/gpio.v(178)
  buf u23 (gpio_ext_porta[2], b_pad_gpio_porta[2]);  // ../RTL/gpio.v(181)
  buf u24 (gpio_ext_porta[1], b_pad_gpio_porta[1]);  // ../RTL/gpio.v(181)
  buf u25 (gpio_ext_porta[0], b_pad_gpio_porta[0]);  // ../RTL/gpio.v(181)
  bufif1 u26 (b_pad_gpio_porta[7], gpio_porta_dr[7], gpio_porta_oe[7]);  // ../RTL/gpio.v(182)
  buf u27 (gpio_porta_oe[0], gpio_porta_ddr[0]);  // ../RTL/gpio.v(180)
  buf u3 (pslverr, 1'b0);  // ../RTL/gpio.v(149)
  bufif1 u4 (b_pad_gpio_porta[0], gpio_porta_dr[0], gpio_porta_oe[0]);  // ../RTL/gpio.v(154)
  bufif1 u5 (b_pad_gpio_porta[1], gpio_porta_dr[1], gpio_porta_oe[1]);  // ../RTL/gpio.v(158)
  bufif1 u6 (b_pad_gpio_porta[2], gpio_porta_dr[2], gpio_porta_oe[2]);  // ../RTL/gpio.v(162)
  buf u7 (gpio_porta_oe[7], gpio_porta_ddr[7]);  // ../RTL/gpio.v(180)
  buf u8 (gpio_porta_oe[6], gpio_porta_ddr[6]);  // ../RTL/gpio.v(180)
  buf u9 (gpio_porta_oe[5], gpio_porta_ddr[5]);  // ../RTL/gpio.v(180)
  gpio_apbif x_gpio_apbif (
    .gpio_ext_porta_rb(gpio_ext_porta_rb),
    .gpio_intstatus(gpio_intstatus),
    .gpio_raw_intstatus(gpio_raw_intstatus),
    .paddr(paddr),
    .pclk(pclk),
    .penable(penable),
    .presetn(presetn),
    .psel(psel),
    .pwdata(pwdata),
    .pwrite(pwrite),
    .gpio_int_polarity(gpio_int_polarity),
    .gpio_inten(gpio_inten),
    .gpio_intmask(gpio_intmask),
    .gpio_inttype_level(gpio_inttype_level),
    .gpio_ls_sync(gpio_ls_sync),
    .gpio_porta_eoi(gpio_porta_eoi),
    .gpio_swporta_ctl(gpio_swporta_ctl),
    .gpio_swporta_ddr(gpio_swporta_ddr),
    .gpio_swporta_dr(gpio_swporta_dr),
    .prdata(prdata));  // ../RTL/gpio.v(98)
  gpio_ctrl x_gpio_ctrl (
    .gpio_ext_porta(gpio_ext_porta),
    .gpio_int_polarity(gpio_int_polarity),
    .gpio_inten(gpio_inten),
    .gpio_intmask(gpio_intmask),
    .gpio_inttype_level(gpio_inttype_level),
    .gpio_ls_sync(gpio_ls_sync),
    .gpio_porta_eoi(gpio_porta_eoi),
    .gpio_swporta_ctl(gpio_swporta_ctl),
    .gpio_swporta_ddr(gpio_swporta_ddr),
    .gpio_swporta_dr(gpio_swporta_dr),
    .pclk(pclk),
    .pclk_intr(pclk_intr),
    .presetn(presetn),
    .gpio_ext_porta_rb(gpio_ext_porta_rb),
    .gpio_intr(gpio_intr),
    .gpio_intr_int(gpio_intstatus),
    .gpio_porta_ddr(gpio_porta_ddr),
    .gpio_porta_dr(gpio_porta_dr),
    .gpio_raw_intstatus(gpio_raw_intstatus));  // ../RTL/gpio.v(122)

endmodule 

module cmsdk_apb_uart  // ../RTL/cmsdk_apb_uart.v(53)
  (
  ECOREVNUM,
  PADDR,
  PCLK,
  PCLKG,
  PENABLE,
  PRESETn,
  PSEL,
  PWDATA,
  PWRITE,
  RXD,
  BAUDTICK,
  PRDATA,
  PREADY,
  PSLVERR,
  RXINT,
  RXOVRINT,
  TXD,
  TXEN,
  TXINT,
  TXOVRINT,
  UARTINT
  );

  input [3:0] ECOREVNUM;  // ../RTL/cmsdk_apb_uart.v(67)
  input [11:2] PADDR;  // ../RTL/cmsdk_apb_uart.v(62)
  input PCLK;  // ../RTL/cmsdk_apb_uart.v(57)
  input PCLKG;  // ../RTL/cmsdk_apb_uart.v(58)
  input PENABLE;  // ../RTL/cmsdk_apb_uart.v(63)
  input PRESETn;  // ../RTL/cmsdk_apb_uart.v(59)
  input PSEL;  // ../RTL/cmsdk_apb_uart.v(61)
  input [31:0] PWDATA;  // ../RTL/cmsdk_apb_uart.v(65)
  input PWRITE;  // ../RTL/cmsdk_apb_uart.v(64)
  input RXD;  // ../RTL/cmsdk_apb_uart.v(73)
  output BAUDTICK;  // ../RTL/cmsdk_apb_uart.v(76)
  output [31:0] PRDATA;  // ../RTL/cmsdk_apb_uart.v(69)
  output PREADY;  // ../RTL/cmsdk_apb_uart.v(70)
  output PSLVERR;  // ../RTL/cmsdk_apb_uart.v(71)
  output RXINT;  // ../RTL/cmsdk_apb_uart.v(79)
  output RXOVRINT;  // ../RTL/cmsdk_apb_uart.v(81)
  output TXD;  // ../RTL/cmsdk_apb_uart.v(74)
  output TXEN;  // ../RTL/cmsdk_apb_uart.v(75)
  output TXINT;  // ../RTL/cmsdk_apb_uart.v(78)
  output TXOVRINT;  // ../RTL/cmsdk_apb_uart.v(80)
  output UARTINT;  // ../RTL/cmsdk_apb_uart.v(82)

  // localparam ARM_CMSDK_APB_UART_CID0 = 8'b00001101;
  // localparam ARM_CMSDK_APB_UART_CID1 = 8'b11110000;
  // localparam ARM_CMSDK_APB_UART_CID2 = 8'b00000101;
  // localparam ARM_CMSDK_APB_UART_CID3 = 8'b10110001;
  // localparam ARM_CMSDK_APB_UART_PID0 = 8'b00100001;
  // localparam ARM_CMSDK_APB_UART_PID1 = 8'b10111000;
  // localparam ARM_CMSDK_APB_UART_PID2 = 8'b00011011;
  // localparam ARM_CMSDK_APB_UART_PID3 = 4'b0000;
  // localparam ARM_CMSDK_APB_UART_PID4 = 8'b00000100;
  // localparam ARM_CMSDK_APB_UART_PID5 = 8'b00000000;
  // localparam ARM_CMSDK_APB_UART_PID6 = 8'b00000000;
  // localparam ARM_CMSDK_APB_UART_PID7 = 8'b00000000;
  wire [1:0] intr_stat_clear;  // ../RTL/cmsdk_apb_uart.v(148)
  wire [1:0] intr_stat_set;  // ../RTL/cmsdk_apb_uart.v(147)
  wire [3:0] intr_state;  // ../RTL/cmsdk_apb_uart.v(146)
  wire [3:0] mapped_cntr_f;  // ../RTL/cmsdk_apb_uart.v(126)
  wire [3:0] n102;
  wire [3:0] n103;
  wire [3:0] n105;
  wire [7:0] n108;
  wire [6:0] n110;
  wire [6:0] n22;
  wire [19:0] n24;
  wire [7:0] n26;
  wire [7:0] n28;
  wire [7:0] n29;
  wire [7:0] n30;
  wire [15:0] n37;
  wire [15:0] n39;
  wire [3:0] n43;
  wire [3:0] n45;
  wire [3:0] n55;
  wire [3:0] n56;
  wire [3:0] n67;
  wire [3:0] n68;
  wire [3:0] n72;
  wire [7:0] n75;
  wire [7:0] n8;
  wire [2:0] n83;
  wire [3:0] n92;
  wire [3:0] n93;
  wire [3:0] nxt_baud_cntr_f;  // ../RTL/cmsdk_apb_uart.v(125)
  wire [15:0] nxt_baud_cntr_i;  // ../RTL/cmsdk_apb_uart.v(123)
  wire [7:0] nxt_rx_buf;  // ../RTL/cmsdk_apb_uart.v(188)
  wire [6:0] nxt_rx_shift_buf;  // ../RTL/cmsdk_apb_uart.v(183)
  wire [4:0] nxt_rx_state;  // ../RTL/cmsdk_apb_uart.v(176)
  wire [4:0] nxt_rx_tick_cnt;  // ../RTL/cmsdk_apb_uart.v(179)
  wire [2:0] nxt_rxd_lpf;  // ../RTL/cmsdk_apb_uart.v(171)
  wire [7:0] nxt_tx_shift_buf;  // ../RTL/cmsdk_apb_uart.v(158)
  wire [4:0] nxt_tx_state;  // ../RTL/cmsdk_apb_uart.v(152)
  wire [4:0] nxt_tx_tick_cnt;  // ../RTL/cmsdk_apb_uart.v(156)
  wire [3:0] pid3_value;  // ../RTL/cmsdk_apb_uart.v(112)
  wire [7:0] read_mux_byte0;  // ../RTL/cmsdk_apb_uart.v(109)
  wire [7:0] read_mux_byte0_reg;  // ../RTL/cmsdk_apb_uart.v(110)
  wire [31:0] read_mux_word;  // ../RTL/cmsdk_apb_uart.v(111)
  wire [3:0] reg_baud_cntr_f;  // ../RTL/cmsdk_apb_uart.v(124)
  wire [15:0] reg_baud_cntr_i;  // ../RTL/cmsdk_apb_uart.v(122)
  wire [19:0] reg_baud_div;  // ../RTL/cmsdk_apb_uart.v(118)
  wire [6:0] reg_ctrl;  // ../RTL/cmsdk_apb_uart.v(115)
  wire [7:0] reg_rx_buf;  // ../RTL/cmsdk_apb_uart.v(117)
  wire [7:0] reg_tx_buf;  // ../RTL/cmsdk_apb_uart.v(116)
  wire [6:0] rx_shift_buf;  // ../RTL/cmsdk_apb_uart.v(182)
  wire [3:0] rx_state;  // ../RTL/cmsdk_apb_uart.v(175)
  wire [3:0] rx_tick_cnt;  // ../RTL/cmsdk_apb_uart.v(178)
  wire [2:0] rxd_lpf;  // ../RTL/cmsdk_apb_uart.v(170)
  wire [7:0] tx_shift_buf;  // ../RTL/cmsdk_apb_uart.v(157)
  wire [3:0] tx_state;  // ../RTL/cmsdk_apb_uart.v(151)
  wire [3:0] tx_tick_cnt;  // ../RTL/cmsdk_apb_uart.v(155)
  wire [3:0] uart_status;  // ../RTL/cmsdk_apb_uart.v(134)
  wire baud_div_en;  // ../RTL/cmsdk_apb_uart.v(131)
  wire baud_updated;  // ../RTL/cmsdk_apb_uart.v(128)
  wire n0;
  wire n1;
  wire n10;
  wire n100;
  wire n101;
  wire n104;
  wire n106;
  wire n107;
  wire n109;
  wire n11;
  wire n111;
  wire n112;
  wire n113;
  wire n114;
  wire n115;
  wire n116;
  wire n117;
  wire n118;
  wire n119;
  wire n12;
  wire n120;
  wire n13;
  wire n14;
  wire n15;
  wire n16;
  wire n17;
  wire n18;
  wire n19;
  wire n2;
  wire n20;
  wire n21;
  wire n23;
  wire n25;
  wire n27;
  wire n3;
  wire n31;
  wire n32;
  wire n33;
  wire n34;
  wire n35;
  wire n36;
  wire n38;
  wire n4;
  wire n40;
  wire n41;
  wire n42;
  wire n44;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n5;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n57;
  wire n58;
  wire n59;
  wire n6;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n65;
  wire n66;
  wire n69;
  wire n7;
  wire n70;
  wire n71;
  wire n73;
  wire n74;
  wire n76;
  wire n77;
  wire n78;
  wire n79;
  wire n80;
  wire n81;
  wire n82;
  wire n84;
  wire n85;
  wire n86;
  wire n87;
  wire n88;
  wire n89;
  wire n9;
  wire n90;
  wire n91;
  wire n94;
  wire n95;
  wire n96;
  wire n97;
  wire n98;
  wire n99;
  wire nxt_rx_buf_full;  // ../RTL/cmsdk_apb_uart.v(185)
  wire nxt_rx_overrun;  // ../RTL/cmsdk_apb_uart.v(139)
  wire nxt_tx_overrun;  // ../RTL/cmsdk_apb_uart.v(140)
  wire nxt_txd;  // ../RTL/cmsdk_apb_uart.v(163)
  wire read_enable;  // ../RTL/cmsdk_apb_uart.v(102)
  wire reg_baud_tick;  // ../RTL/cmsdk_apb_uart.v(127)
  wire reg_rx_overrun;  // ../RTL/cmsdk_apb_uart.v(135)
  wire reg_rxintr;  // ../RTL/cmsdk_apb_uart.v(143)
  wire reg_tx_overrun;  // ../RTL/cmsdk_apb_uart.v(137)
  wire reg_txd;  // ../RTL/cmsdk_apb_uart.v(162)
  wire reg_txintr;  // ../RTL/cmsdk_apb_uart.v(142)
  wire reload_f;  // ../RTL/cmsdk_apb_uart.v(130)
  wire reload_i;  // ../RTL/cmsdk_apb_uart.v(129)
  wire rx_buf_full;  // ../RTL/cmsdk_apb_uart.v(184)
  wire rx_data_read;  // ../RTL/cmsdk_apb_uart.v(187)
  wire rx_overflow_intr;  // ../RTL/cmsdk_apb_uart.v(145)
  wire rx_overrun;  // ../RTL/cmsdk_apb_uart.v(136)
  wire rx_shift_in;  // ../RTL/cmsdk_apb_uart.v(172)
  wire rx_state_inc;  // ../RTL/cmsdk_apb_uart.v(181)
  wire rx_state_update;  // ../RTL/cmsdk_apb_uart.v(177)
  wire rxbuf_sample;  // ../RTL/cmsdk_apb_uart.v(186)
  wire rxd_sync_1;  // ../RTL/cmsdk_apb_uart.v(168)
  wire rxd_sync_2;  // ../RTL/cmsdk_apb_uart.v(169)
  wire tx_buf_clear;  // ../RTL/cmsdk_apb_uart.v(165)
  wire tx_buf_ctrl_shift;  // ../RTL/cmsdk_apb_uart.v(159)
  wire tx_buf_full;  // ../RTL/cmsdk_apb_uart.v(161)
  wire tx_overflow_intr;  // ../RTL/cmsdk_apb_uart.v(144)
  wire tx_overrun;  // ../RTL/cmsdk_apb_uart.v(138)
  wire tx_state_inc;  // ../RTL/cmsdk_apb_uart.v(154)
  wire tx_state_update;  // ../RTL/cmsdk_apb_uart.v(153)
  wire update_reg_txd;  // ../RTL/cmsdk_apb_uart.v(164)
  wire update_rx_tick_cnt;  // ../RTL/cmsdk_apb_uart.v(180)
  wire write_enable;  // ../RTL/cmsdk_apb_uart.v(103)
  wire write_enable00;  // ../RTL/cmsdk_apb_uart.v(104)
  wire write_enable04;  // ../RTL/cmsdk_apb_uart.v(105)
  wire write_enable08;  // ../RTL/cmsdk_apb_uart.v(106)
  wire write_enable0c;  // ../RTL/cmsdk_apb_uart.v(107)
  wire write_enable10;  // ../RTL/cmsdk_apb_uart.v(108)

  add_pu4_pu4_o5 add0 (
    .i0(tx_tick_cnt),
    .i1({3'b000,reg_baud_tick}),
    .o({n54,n55}));  // ../RTL/cmsdk_apb_uart.v(397)
  add_pu4_pu4_o5 add1 (
    .i0(tx_state),
    .i1({3'b000,tx_state_inc}),
    .o({n66,n67}));  // ../RTL/cmsdk_apb_uart.v(427)
  add_pu4_pu4_o5 add2 (
    .i0(rx_tick_cnt),
    .i1({3'b000,reg_baud_tick}),
    .o({n91,n92}));  // ../RTL/cmsdk_apb_uart.v(525)
  add_pu4_pu4_o5 add3 (
    .i0(rx_state),
    .i1({3'b000,rx_state_inc}),
    .o({n101,n102}));  // ../RTL/cmsdk_apb_uart.v(565)
  AL_DFF baud_updated_reg (
    .clk(PCLK),
    .d(n47),
    .reset(n23),
    .set(1'b0),
    .q(baud_updated));  // ../RTL/cmsdk_apb_uart.v(368)
  eq_w10 eq0 (
    .i0(PADDR),
    .i1(10'b0000000000),
    .o(n3));  // ../RTL/cmsdk_apb_uart.v(194)
  eq_w10 eq1 (
    .i0(PADDR),
    .i1(10'b0000000001),
    .o(n4));  // ../RTL/cmsdk_apb_uart.v(195)
  eq_w4 eq10 (
    .i0(tx_state),
    .i1(4'b0001),
    .o(n52));  // ../RTL/cmsdk_apb_uart.v(396)
  eq_w4 eq11 (
    .i0(tx_state),
    .i1(4'b0000),
    .o(n60));  // ../RTL/cmsdk_apb_uart.v(412)
  eq_w4 eq12 (
    .i0(tx_state),
    .i1(4'b1011),
    .o(n62));  // ../RTL/cmsdk_apb_uart.v(413)
  eq_w4 eq13 (
    .i0(tx_state),
    .i1(4'b0010),
    .o(n76));  // ../RTL/cmsdk_apb_uart.v(465)
  eq_w4 eq14 (
    .i0(rx_state),
    .i1(4'b0000),
    .o(n88));  // ../RTL/cmsdk_apb_uart.v(524)
  eq_w4 eq15 (
    .i0(rx_state),
    .i1(4'b1001),
    .o(n97));  // ../RTL/cmsdk_apb_uart.v(544)
  eq_w10 eq2 (
    .i0(PADDR),
    .i1(10'b0000000010),
    .o(n5));  // ../RTL/cmsdk_apb_uart.v(196)
  eq_w10 eq3 (
    .i0(PADDR),
    .i1(10'b0000000011),
    .o(n6));  // ../RTL/cmsdk_apb_uart.v(197)
  eq_w10 eq4 (
    .i0(PADDR),
    .i1(10'b0000000100),
    .o(n7));  // ../RTL/cmsdk_apb_uart.v(198)
  eq_w7 eq5 (
    .i0(PADDR[11:5]),
    .i1(7'b0000000),
    .o(n25));  // ../RTL/cmsdk_apb_uart.v(259)
  eq_w6 eq6 (
    .i0(PADDR[11:6]),
    .i1(6'b111111),
    .o(n27));  // ../RTL/cmsdk_apb_uart.v(270)
  eq_w15 eq7 (
    .i0(reg_baud_cntr_i[15:1]),
    .i1(15'b000000000000000),
    .o(n32));  // ../RTL/cmsdk_apb_uart.v(329)
  eq_w16 eq8 (
    .i0(reg_baud_cntr_i),
    .i1(16'b0000000000000000),
    .o(n34));  // ../RTL/cmsdk_apb_uart.v(330)
  eq_w4 eq9 (
    .i0(reg_baud_cntr_f),
    .i1(4'b0000),
    .o(n40));  // ../RTL/cmsdk_apb_uart.v(345)
  lt_u4_u4 lt0 (
    .ci(1'b1),
    .i0(reg_baud_div[3:0]),
    .i1(mapped_cntr_f),
    .o(n31));  // ../RTL/cmsdk_apb_uart.v(328)
  lt_u4_u4 lt1 (
    .ci(1'b0),
    .i0(4'b1011),
    .i1(tx_state),
    .o(n71));  // ../RTL/cmsdk_apb_uart.v(437)
  lt_u4_u4 lt2 (
    .ci(1'b0),
    .i0(4'b0010),
    .i1(tx_state),
    .o(n73));  // ../RTL/cmsdk_apb_uart.v(451)
  binary_mux_s1_w8 mux0 (
    .i0(reg_tx_buf),
    .i1(PWDATA[7:0]),
    .sel(write_enable00),
    .o(n8));  // ../RTL/cmsdk_apb_uart.v(207)
  binary_mux_s1_w7 mux1 (
    .i0(reg_ctrl),
    .i1(PWDATA[6:0]),
    .sel(write_enable08),
    .o(n22));  // ../RTL/cmsdk_apb_uart.v(238)
  binary_mux_s1_w16 mux10 (
    .i0(n37),
    .i1(reg_baud_div[19:4]),
    .sel(n36),
    .o(nxt_baud_cntr_i));  // ../RTL/cmsdk_apb_uart.v(334)
  binary_mux_s1_w16 mux11 (
    .i0(reg_baud_cntr_i),
    .i1(nxt_baud_cntr_i),
    .sel(n38),
    .o(n39));  // ../RTL/cmsdk_apb_uart.v(341)
  binary_mux_s1_w4 mux12 (
    .i0(n43),
    .i1(4'b1111),
    .sel(n42),
    .o(nxt_baud_cntr_f));  // ../RTL/cmsdk_apb_uart.v(350)
  binary_mux_s1_w4 mux13 (
    .i0(reg_baud_cntr_f),
    .i1(nxt_baud_cntr_f),
    .sel(n44),
    .o(n45));  // ../RTL/cmsdk_apb_uart.v(358)
  binary_mux_s1_w5 mux14 (
    .i0({n54,n55}),
    .i1(5'b00000),
    .sel(n53),
    .o({open_n0,nxt_tx_tick_cnt[3:0]}));  // ../RTL/cmsdk_apb_uart.v(397)
  binary_mux_s1_w4 mux15 (
    .i0(tx_tick_cnt),
    .i1(nxt_tx_tick_cnt[3:0]),
    .sel(reg_baud_tick),
    .o(n56));  // ../RTL/cmsdk_apb_uart.v(405)
  binary_mux_s1_w4 mux16 (
    .i0(tx_state),
    .i1({2'b00,tx_buf_full,1'b0}),
    .sel(tx_state_inc),
    .o(n68));  // ../RTL/cmsdk_apb_uart.v(430)
  binary_mux_s4_w5 mux17 (
    .i0({4'b0000,n65}),
    .i1({n66,n67}),
    .i10({n66,n67}),
    .i11({1'b0,n68}),
    .i12(5'bxxxxx),
    .i13(5'bxxxxx),
    .i14(5'bxxxxx),
    .i15(5'bxxxxx),
    .i2({n66,n67}),
    .i3({n66,n67}),
    .i4({n66,n67}),
    .i5({n66,n67}),
    .i6({n66,n67}),
    .i7({n66,n67}),
    .i8({n66,n67}),
    .i9({n66,n67}),
    .sel(tx_state),
    .o({open_n1,nxt_tx_state[3:0]}));  // ../RTL/cmsdk_apb_uart.v(434)
  binary_mux_s1_w4 mux18 (
    .i0(tx_state),
    .i1(nxt_tx_state[3:0]),
    .sel(tx_state_update),
    .o(n72));  // ../RTL/cmsdk_apb_uart.v(445)
  binary_mux_s1_w8 mux19 (
    .i0({1'b1,tx_shift_buf[7:1]}),
    .i1(reg_tx_buf),
    .sel(tx_buf_clear),
    .o(nxt_tx_shift_buf));  // ../RTL/cmsdk_apb_uart.v(453)
  binary_mux_s1_w20 mux2 (
    .i0(reg_baud_div),
    .i1(PWDATA[19:0]),
    .sel(write_enable10),
    .o(n24));  // ../RTL/cmsdk_apb_uart.v(247)
  binary_mux_s1_w8 mux20 (
    .i0(tx_shift_buf),
    .i1(nxt_tx_shift_buf),
    .sel(n74),
    .o(n75));  // ../RTL/cmsdk_apb_uart.v(461)
  binary_mux_s1_w3 mux21 (
    .i0(rxd_lpf),
    .i1(nxt_rxd_lpf),
    .sel(reg_baud_tick),
    .o(n83));  // ../RTL/cmsdk_apb_uart.v(512)
  binary_mux_s1_w5 mux22 (
    .i0({n91,n92}),
    .i1(5'b01000),
    .sel(n90),
    .o({open_n2,nxt_rx_tick_cnt[3:0]}));  // ../RTL/cmsdk_apb_uart.v(525)
  binary_mux_s1_w4 mux23 (
    .i0(rx_tick_cnt),
    .i1(nxt_rx_tick_cnt[3:0]),
    .sel(update_rx_tick_cnt),
    .o(n93));  // ../RTL/cmsdk_apb_uart.v(535)
  binary_mux_s4_w5 mux24 (
    .i0({4'b0000,n100}),
    .i1({n101,n102}),
    .i10({1'b0,n103[3],1'b0,n103[3],1'b0}),
    .i11(5'bxxxxx),
    .i12(5'bxxxxx),
    .i13(5'bxxxxx),
    .i14(5'bxxxxx),
    .i15(5'bxxxxx),
    .i2({n101,n102}),
    .i3({n101,n102}),
    .i4({n101,n102}),
    .i5({n101,n102}),
    .i6({n101,n102}),
    .i7({n101,n102}),
    .i8({n101,n102}),
    .i9({n101,n102}),
    .sel(rx_state),
    .o({open_n3,nxt_rx_state[3:0]}));  // ../RTL/cmsdk_apb_uart.v(572)
  binary_mux_s1_w4 mux25 (
    .i0(rx_state),
    .i1(nxt_rx_state[3:0]),
    .sel(rx_state_update),
    .o(n105));  // ../RTL/cmsdk_apb_uart.v(583)
  binary_mux_s1_w8 mux26 (
    .i0(reg_rx_buf),
    .i1(nxt_rx_buf),
    .sel(rxbuf_sample),
    .o(n108));  // ../RTL/cmsdk_apb_uart.v(603)
  binary_mux_s1_w7 mux27 (
    .i0(rx_shift_buf),
    .i1(nxt_rx_shift_buf),
    .sel(rx_state_inc),
    .o(n110));  // ../RTL/cmsdk_apb_uart.v(614)
  binary_mux_s3_w8 mux3 (
    .i0(reg_rx_buf),
    .i1({4'b0000,uart_status}),
    .i2({1'b0,reg_ctrl}),
    .i3({4'b0000,intr_state}),
    .i4(reg_baud_div[7:0]),
    .i5(8'b00000000),
    .i6(8'b00000000),
    .i7(8'b00000000),
    .sel(PADDR[4:2]),
    .o(n26));  // ../RTL/cmsdk_apb_uart.v(268)
  binary_mux_s4_w8 mux4 (
    .i0(8'b00000000),
    .i1(8'b00000000),
    .i10(8'b00011011),
    .i11({ECOREVNUM,pid3_value}),
    .i12(8'b00001101),
    .i13(8'b11110000),
    .i14(8'b00000101),
    .i15(8'b10110001),
    .i2(8'b00000000),
    .i3(8'b00000000),
    .i4(8'b00000100),
    .i5(8'b00000000),
    .i6(8'b00000000),
    .i7(8'b00000000),
    .i8(8'b00100001),
    .i9(8'b10111000),
    .sel(PADDR[5:2]),
    .o(n28));  // ../RTL/cmsdk_apb_uart.v(288)
  binary_mux_s1_w8 mux5 (
    .i0(8'b00000000),
    .i1(n28),
    .sel(n27),
    .o(n29));  // ../RTL/cmsdk_apb_uart.v(292)
  binary_mux_s1_w8 mux6 (
    .i0(n29),
    .i1(n26),
    .sel(n25),
    .o(read_mux_byte0));  // ../RTL/cmsdk_apb_uart.v(292)
  binary_mux_s1_w8 mux7 (
    .i0(read_mux_byte0_reg),
    .i1(read_mux_byte0),
    .sel(read_enable),
    .o(n30));  // ../RTL/cmsdk_apb_uart.v(303)
  binary_mux_s1_w12 mux8 (
    .i0(12'b000000000000),
    .i1(reg_baud_div[19:8]),
    .sel(n7),
    .o(read_mux_word[19:8]));  // ../RTL/cmsdk_apb_uart.v(308)
  binary_mux_s1_w32 mux9 (
    .i0(32'b00000000000000000000000000000000),
    .i1(read_mux_word),
    .sel(read_enable),
    .o(PRDATA));  // ../RTL/cmsdk_apb_uart.v(313)
  ne_w2 neq0 (
    .i0(reg_ctrl[1:0]),
    .i1(2'b00),
    .o(baud_div_en));  // ../RTL/cmsdk_apb_uart.v(320)
  reg_ar_as_w7 reg0 (
    .clk(PCLKG),
    .d(n22),
    .reset({n23,n23,n23,n23,n23,n23,n23}),
    .set(7'b0000000),
    .q(reg_ctrl));  // ../RTL/cmsdk_apb_uart.v(238)
  reg_ar_as_w20 reg1 (
    .clk(PCLKG),
    .d(n24),
    .reset({n23,n23,n23,n23,n23,n23,n23,n23,n23,n23,n23,n23,n23,n23,n23,n23,n23,n23,n23,n23}),
    .set(20'b00000000000000000000),
    .q(reg_baud_div));  // ../RTL/cmsdk_apb_uart.v(247)
  reg_ar_as_w4 reg10 (
    .clk(PCLK),
    .d(n105),
    .reset({n23,n23,n23,n23}),
    .set(4'b0000),
    .q(rx_state));  // ../RTL/cmsdk_apb_uart.v(583)
  reg_ar_as_w8 reg11 (
    .clk(PCLK),
    .d(n108),
    .reset({n23,n23,n23,n23,n23,n23,n23,n23}),
    .set(8'b00000000),
    .q(reg_rx_buf));  // ../RTL/cmsdk_apb_uart.v(603)
  reg_ar_as_w7 reg12 (
    .clk(PCLK),
    .d(n110),
    .reset({n23,n23,n23,n23,n23,n23,n23}),
    .set(7'b0000000),
    .q(rx_shift_buf));  // ../RTL/cmsdk_apb_uart.v(614)
  reg_ar_as_w8 reg13 (
    .clk(PCLKG),
    .d(n8),
    .reset({n23,n23,n23,n23,n23,n23,n23,n23}),
    .set(8'b00000000),
    .q(reg_tx_buf));  // ../RTL/cmsdk_apb_uart.v(207)
  reg_ar_as_w8 reg2 (
    .clk(PCLKG),
    .d(n30),
    .reset({n23,n23,n23,n23,n23,n23,n23,n23}),
    .set(8'b00000000),
    .q(read_mux_byte0_reg));  // ../RTL/cmsdk_apb_uart.v(303)
  reg_ar_as_w16 reg3 (
    .clk(PCLK),
    .d(n39),
    .reset({n23,n23,n23,n23,n23,n23,n23,n23,n23,n23,n23,n23,n23,n23,n23,n23}),
    .set(16'b0000000000000000),
    .q(reg_baud_cntr_i));  // ../RTL/cmsdk_apb_uart.v(341)
  reg_ar_as_w4 reg4 (
    .clk(PCLK),
    .d(n45),
    .reset({n23,n23,n23,n23}),
    .set(4'b0000),
    .q(reg_baud_cntr_f));  // ../RTL/cmsdk_apb_uart.v(358)
  reg_ar_as_w4 reg5 (
    .clk(PCLK),
    .d(n56),
    .reset({n23,n23,n23,n23}),
    .set(4'b0000),
    .q(tx_tick_cnt));  // ../RTL/cmsdk_apb_uart.v(405)
  reg_ar_as_w4 reg6 (
    .clk(PCLK),
    .d(n72),
    .reset({n23,n23,n23,n23}),
    .set(4'b0000),
    .q(tx_state));  // ../RTL/cmsdk_apb_uart.v(445)
  reg_ar_as_w8 reg7 (
    .clk(PCLK),
    .d(n75),
    .reset({n23,n23,n23,n23,n23,n23,n23,n23}),
    .set(8'b00000000),
    .q(tx_shift_buf));  // ../RTL/cmsdk_apb_uart.v(461)
  reg_ar_as_w3 reg8 (
    .clk(PCLK),
    .d(n83),
    .reset(3'b000),
    .set({n23,n23,n23}),
    .q(rxd_lpf));  // ../RTL/cmsdk_apb_uart.v(512)
  reg_ar_as_w4 reg9 (
    .clk(PCLK),
    .d(n93),
    .reset({n23,n23,n23,n23}),
    .set(4'b0000),
    .q(rx_tick_cnt));  // ../RTL/cmsdk_apb_uart.v(535)
  AL_DFF reg_baud_tick_reg (
    .clk(PCLK),
    .d(n49),
    .reset(n23),
    .set(1'b0),
    .q(reg_baud_tick));  // ../RTL/cmsdk_apb_uart.v(377)
  AL_DFF reg_rx_overrun_reg (
    .clk(PCLK),
    .d(n18),
    .reset(n23),
    .set(1'b0),
    .q(reg_rx_overrun));  // ../RTL/cmsdk_apb_uart.v(220)
  AL_DFF reg_rxintr_reg (
    .clk(PCLK),
    .d(n118),
    .reset(n23),
    .set(1'b0),
    .q(reg_rxintr));  // ../RTL/cmsdk_apb_uart.v(642)
  AL_DFF reg_tx_overrun_reg (
    .clk(PCLK),
    .d(n21),
    .reset(n23),
    .set(1'b0),
    .q(reg_tx_overrun));  // ../RTL/cmsdk_apb_uart.v(229)
  AL_DFF reg_txd_reg (
    .clk(PCLK),
    .d(n78),
    .reset(1'b0),
    .set(n23),
    .q(reg_txd));  // ../RTL/cmsdk_apb_uart.v(476)
  AL_DFF reg_txintr_reg (
    .clk(PCLK),
    .d(n115),
    .reset(n23),
    .set(1'b0),
    .q(reg_txintr));  // ../RTL/cmsdk_apb_uart.v(634)
  AL_DFF rx_buf_full_reg (
    .clk(PCLK),
    .d(n107),
    .reset(n23),
    .set(1'b0),
    .q(rx_buf_full));  // ../RTL/cmsdk_apb_uart.v(592)
  AL_DFF rxd_sync_1_reg (
    .clk(PCLK),
    .d(n81),
    .reset(1'b0),
    .set(n23),
    .q(rxd_sync_1));  // ../RTL/cmsdk_apb_uart.v(501)
  AL_DFF rxd_sync_2_reg (
    .clk(PCLK),
    .d(n82),
    .reset(1'b0),
    .set(n23),
    .q(rxd_sync_2));  // ../RTL/cmsdk_apb_uart.v(501)
  add_pu16_mu16_o16 sub0 (
    .i0(reg_baud_cntr_i),
    .i1(16'b0000000000000001),
    .o(n37));  // ../RTL/cmsdk_apb_uart.v(334)
  add_pu4_mu4_o4 sub1 (
    .i0(reg_baud_cntr_f),
    .i1(4'b0001),
    .o(n43));  // ../RTL/cmsdk_apb_uart.v(350)
  AL_DFF tx_buf_full_reg (
    .clk(PCLK),
    .d(n51),
    .reset(n23),
    .set(1'b0),
    .q(tx_buf_full));  // ../RTL/cmsdk_apb_uart.v(392)
  and u10 (write_enable08, write_enable, n5);  // ../RTL/cmsdk_apb_uart.v(196)
  and u100 (tx_overrun, n80, write_enable00);  // ../RTL/cmsdk_apb_uart.v(480)
  buf u101 (TXD, reg_txd);  // ../RTL/cmsdk_apb_uart.v(483)
  buf u102 (TXEN, reg_ctrl[0]);  // ../RTL/cmsdk_apb_uart.v(484)
  buf u103 (read_mux_word[29], 1'b0);  // ../RTL/cmsdk_apb_uart.v(309)
  AL_MUX u104 (
    .i0(rxd_sync_1),
    .i1(RXD),
    .sel(reg_ctrl[1]),
    .o(n81));  // ../RTL/cmsdk_apb_uart.v(501)
  AL_MUX u105 (
    .i0(rxd_sync_2),
    .i1(rxd_sync_1),
    .sel(reg_ctrl[1]),
    .o(n82));  // ../RTL/cmsdk_apb_uart.v(501)
  and u106 (n113, tx_tick_cnt[0], tx_tick_cnt[1]);  // ../RTL/cmsdk_apb_uart.v(409)
  buf u107 (read_mux_word[28], 1'b0);  // ../RTL/cmsdk_apb_uart.v(309)
  and u108 (n84, rxd_lpf[1], rxd_lpf[0]);  // ../RTL/cmsdk_apb_uart.v(516)
  and u109 (n85, rxd_lpf[1], rxd_lpf[2]);  // ../RTL/cmsdk_apb_uart.v(517)
  and u11 (write_enable0c, write_enable, n6);  // ../RTL/cmsdk_apb_uart.v(197)
  or u110 (n86, n84, n85);  // ../RTL/cmsdk_apb_uart.v(517)
  and u111 (n87, rxd_lpf[0], rxd_lpf[2]);  // ../RTL/cmsdk_apb_uart.v(518)
  or u112 (rx_shift_in, n86, n87);  // ../RTL/cmsdk_apb_uart.v(518)
  not u113 (n89, rx_shift_in);  // ../RTL/cmsdk_apb_uart.v(524)
  and u114 (n90, n88, n89);  // ../RTL/cmsdk_apb_uart.v(524)
  buf u115 (read_mux_word[27], 1'b0);  // ../RTL/cmsdk_apb_uart.v(309)
  buf u116 (read_mux_word[26], 1'b0);  // ../RTL/cmsdk_apb_uart.v(309)
  buf u117 (read_mux_word[25], 1'b0);  // ../RTL/cmsdk_apb_uart.v(309)
  or u118 (update_rx_tick_cnt, n90, reg_baud_tick);  // ../RTL/cmsdk_apb_uart.v(527)
  buf u119 (read_mux_word[24], 1'b0);  // ../RTL/cmsdk_apb_uart.v(309)
  and u12 (write_enable10, write_enable, n7);  // ../RTL/cmsdk_apb_uart.v(198)
  buf u120 (nxt_rxd_lpf[0], rxd_sync_2);  // ../RTL/cmsdk_apb_uart.v(505)
  and u121 (rx_state_inc, n94, reg_baud_tick);  // ../RTL/cmsdk_apb_uart.v(539)
  not u122 (n95, rx_data_read);  // ../RTL/cmsdk_apb_uart.v(541)
  and u123 (n96, rx_buf_full, n95);  // ../RTL/cmsdk_apb_uart.v(541)
  or u124 (nxt_rx_buf_full, rxbuf_sample, n96);  // ../RTL/cmsdk_apb_uart.v(541)
  and u125 (rxbuf_sample, n97, rx_state_inc);  // ../RTL/cmsdk_apb_uart.v(544)
  buf u126 (read_mux_word[23], 1'b0);  // ../RTL/cmsdk_apb_uart.v(309)
  buf u127 (read_mux_word[22], 1'b0);  // ../RTL/cmsdk_apb_uart.v(309)
  buf u128 (read_mux_word[21], 1'b0);  // ../RTL/cmsdk_apb_uart.v(309)
  and u129 (n98, n2, n3);  // ../RTL/cmsdk_apb_uart.v(548)
  not u13 (n23, PRESETn);  // ../RTL/cmsdk_apb_uart.v(204)
  buf u130 (read_mux_word[20], 1'b0);  // ../RTL/cmsdk_apb_uart.v(309)
  and u131 (rx_data_read, n98, n0);  // ../RTL/cmsdk_apb_uart.v(548)
  and u132 (n99, rx_buf_full, rxbuf_sample);  // ../RTL/cmsdk_apb_uart.v(550)
  buf u133 (read_mux_word[7], read_mux_byte0_reg[7]);  // ../RTL/cmsdk_apb_uart.v(309)
  and u134 (rx_overrun, n99, n95);  // ../RTL/cmsdk_apb_uart.v(550)
  buf u135 (read_mux_word[6], read_mux_byte0_reg[6]);  // ../RTL/cmsdk_apb_uart.v(309)
  and u136 (n100, n89, reg_ctrl[1]);  // ../RTL/cmsdk_apb_uart.v(561)
  buf u137 (pid3_value[3], 1'b0);  // ../RTL/cmsdk_apb_uart.v(253)
  buf u138 (read_mux_word[5], read_mux_byte0_reg[5]);  // ../RTL/cmsdk_apb_uart.v(309)
  buf u139 (read_mux_word[4], read_mux_byte0_reg[4]);  // ../RTL/cmsdk_apb_uart.v(309)
  or u14 (n9, write_enable04, write_enable0c);  // ../RTL/cmsdk_apb_uart.v(211)
  or u140 (rx_state_update, rx_state_inc, n100);  // ../RTL/cmsdk_apb_uart.v(575)
  buf u141 (read_mux_word[3], read_mux_byte0_reg[3]);  // ../RTL/cmsdk_apb_uart.v(309)
  buf u142 (read_mux_word[2], read_mux_byte0_reg[2]);  // ../RTL/cmsdk_apb_uart.v(309)
  or u143 (n106, rxbuf_sample, rx_data_read);  // ../RTL/cmsdk_apb_uart.v(591)
  AL_MUX u144 (
    .i0(rx_buf_full),
    .i1(nxt_rx_buf_full),
    .sel(n106),
    .o(n107));  // ../RTL/cmsdk_apb_uart.v(592)
  and u145 (n116, rx_tick_cnt[0], rx_tick_cnt[1]);  // ../RTL/cmsdk_apb_uart.v(539)
  buf u146 (uart_status[3], reg_rx_overrun);  // ../RTL/cmsdk_apb_uart.v(251)
  buf u147 (read_mux_word[1], read_mux_byte0_reg[1]);  // ../RTL/cmsdk_apb_uart.v(309)
  buf u148 (nxt_rx_buf[0], rx_shift_buf[0]);  // ../RTL/cmsdk_apb_uart.v(596)
  buf u149 (uart_status[2], reg_tx_overrun);  // ../RTL/cmsdk_apb_uart.v(251)
  and u15 (n10, n9, PWDATA[3]);  // ../RTL/cmsdk_apb_uart.v(211)
  buf u150 (intr_state[3], rx_overflow_intr);  // ../RTL/cmsdk_apb_uart.v(649)
  and u151 (n111, reg_ctrl[2], reg_ctrl[0]);  // ../RTL/cmsdk_apb_uart.v(623)
  and u152 (n112, n111, tx_buf_full);  // ../RTL/cmsdk_apb_uart.v(623)
  buf u153 (nxt_rx_shift_buf[0], rx_shift_buf[1]);  // ../RTL/cmsdk_apb_uart.v(607)
  buf u154 (uart_status[1], rx_buf_full);  // ../RTL/cmsdk_apb_uart.v(251)
  buf u155 (intr_state[2], tx_overflow_intr);  // ../RTL/cmsdk_apb_uart.v(649)
  or u156 (n114, intr_stat_set[0], intr_stat_clear[0]);  // ../RTL/cmsdk_apb_uart.v(633)
  AL_MUX u157 (
    .i0(reg_txintr),
    .i1(intr_stat_set[0]),
    .sel(n114),
    .o(n115));  // ../RTL/cmsdk_apb_uart.v(634)
  buf u158 (intr_state[1], reg_rxintr);  // ../RTL/cmsdk_apb_uart.v(649)
  buf u159 (intr_state[0], reg_txintr);  // ../RTL/cmsdk_apb_uart.v(649)
  not u16 (n11, n10);  // ../RTL/cmsdk_apb_uart.v(211)
  or u160 (n117, intr_stat_set[1], intr_stat_clear[1]);  // ../RTL/cmsdk_apb_uart.v(641)
  AL_MUX u161 (
    .i0(reg_rxintr),
    .i1(intr_stat_set[1]),
    .sel(n117),
    .o(n118));  // ../RTL/cmsdk_apb_uart.v(642)
  and u162 (intr_stat_clear[0], write_enable0c, PWDATA[0]);  // ../RTL/cmsdk_apb_uart.v(626)
  and u163 (rx_overflow_intr, reg_rx_overrun, reg_ctrl[5]);  // ../RTL/cmsdk_apb_uart.v(645)
  and u164 (tx_overflow_intr, reg_tx_overrun, reg_ctrl[4]);  // ../RTL/cmsdk_apb_uart.v(646)
  buf u165 (read_mux_word[0], read_mux_byte0_reg[0]);  // ../RTL/cmsdk_apb_uart.v(309)
  buf u166 (TXINT, reg_txintr);  // ../RTL/cmsdk_apb_uart.v(652)
  buf u167 (RXINT, reg_rxintr);  // ../RTL/cmsdk_apb_uart.v(653)
  buf u168 (TXOVRINT, tx_overflow_intr);  // ../RTL/cmsdk_apb_uart.v(654)
  buf u169 (RXOVRINT, rx_overflow_intr);  // ../RTL/cmsdk_apb_uart.v(655)
  and u17 (n12, reg_rx_overrun, n11);  // ../RTL/cmsdk_apb_uart.v(211)
  or u170 (n119, reg_txintr, reg_rxintr);  // ../RTL/cmsdk_apb_uart.v(656)
  or u171 (n120, n119, tx_overflow_intr);  // ../RTL/cmsdk_apb_uart.v(656)
  or u172 (UARTINT, n120, rx_overflow_intr);  // ../RTL/cmsdk_apb_uart.v(656)
  or u18 (nxt_rx_overrun, n12, rx_overrun);  // ../RTL/cmsdk_apb_uart.v(211)
  buf u19 (pid3_value[2], 1'b0);  // ../RTL/cmsdk_apb_uart.v(253)
  and u20 (n13, n9, PWDATA[2]);  // ../RTL/cmsdk_apb_uart.v(212)
  not u21 (n14, n13);  // ../RTL/cmsdk_apb_uart.v(212)
  and u22 (n15, reg_tx_overrun, n14);  // ../RTL/cmsdk_apb_uart.v(212)
  or u23 (nxt_tx_overrun, n15, tx_overrun);  // ../RTL/cmsdk_apb_uart.v(212)
  buf u24 (pid3_value[1], 1'b0);  // ../RTL/cmsdk_apb_uart.v(253)
  or u25 (n16, rx_overrun, write_enable04);  // ../RTL/cmsdk_apb_uart.v(219)
  or u26 (n17, n16, write_enable0c);  // ../RTL/cmsdk_apb_uart.v(219)
  AL_MUX u27 (
    .i0(reg_rx_overrun),
    .i1(nxt_rx_overrun),
    .sel(n17),
    .o(n18));  // ../RTL/cmsdk_apb_uart.v(220)
  and u28 (intr_stat_set[1], reg_ctrl[3], rxbuf_sample);  // ../RTL/cmsdk_apb_uart.v(622)
  or u29 (n19, tx_overrun, write_enable04);  // ../RTL/cmsdk_apb_uart.v(228)
  not u3 (n0, PWRITE);  // ../RTL/cmsdk_apb_uart.v(192)
  or u30 (n20, n19, write_enable0c);  // ../RTL/cmsdk_apb_uart.v(228)
  AL_MUX u31 (
    .i0(reg_tx_overrun),
    .i1(nxt_tx_overrun),
    .sel(n20),
    .o(n21));  // ../RTL/cmsdk_apb_uart.v(229)
  buf u32 (mapped_cntr_f[3], reg_baud_cntr_f[0]);  // ../RTL/cmsdk_apb_uart.v(322)
  buf u33 (mapped_cntr_f[2], reg_baud_cntr_f[1]);  // ../RTL/cmsdk_apb_uart.v(322)
  buf u34 (uart_status[0], tx_buf_full);  // ../RTL/cmsdk_apb_uart.v(251)
  buf u35 (mapped_cntr_f[1], reg_baud_cntr_f[2]);  // ../RTL/cmsdk_apb_uart.v(322)
  and u36 (n57, n113, n109);  // ../RTL/cmsdk_apb_uart.v(409)
  buf u37 (pid3_value[0], 1'b0);  // ../RTL/cmsdk_apb_uart.v(253)
  buf u38 (PREADY, 1'b1);  // ../RTL/cmsdk_apb_uart.v(314)
  buf u39 (PSLVERR, 1'b0);  // ../RTL/cmsdk_apb_uart.v(315)
  and u4 (read_enable, PSEL, n0);  // ../RTL/cmsdk_apb_uart.v(192)
  and u40 (intr_stat_set[0], n112, tx_buf_clear);  // ../RTL/cmsdk_apb_uart.v(622)
  and u41 (n33, n31, n32);  // ../RTL/cmsdk_apb_uart.v(329)
  or u42 (n35, n33, n34);  // ../RTL/cmsdk_apb_uart.v(330)
  and u43 (reload_i, baud_div_en, n35);  // ../RTL/cmsdk_apb_uart.v(330)
  or u44 (n36, baud_updated, reload_i);  // ../RTL/cmsdk_apb_uart.v(333)
  and u45 (n109, tx_tick_cnt[2], tx_tick_cnt[3]);  // ../RTL/cmsdk_apb_uart.v(409)
  or u46 (n38, baud_updated, baud_div_en);  // ../RTL/cmsdk_apb_uart.v(340)
  and u47 (n41, baud_div_en, n40);  // ../RTL/cmsdk_apb_uart.v(345)
  and u48 (reload_f, n41, reload_i);  // ../RTL/cmsdk_apb_uart.v(346)
  or u49 (n42, reload_f, baud_updated);  // ../RTL/cmsdk_apb_uart.v(349)
  not u5 (n1, PENABLE);  // ../RTL/cmsdk_apb_uart.v(193)
  buf u50 (nxt_rxd_lpf[2], rxd_lpf[1]);  // ../RTL/cmsdk_apb_uart.v(505)
  buf u51 (nxt_rxd_lpf[1], rxd_lpf[0]);  // ../RTL/cmsdk_apb_uart.v(505)
  or u52 (n44, n42, reload_i);  // ../RTL/cmsdk_apb_uart.v(357)
  and u53 (n94, n116, n104);  // ../RTL/cmsdk_apb_uart.v(539)
  or u54 (n46, write_enable10, baud_updated);  // ../RTL/cmsdk_apb_uart.v(366)
  AL_MUX u55 (
    .i0(baud_updated),
    .i1(write_enable10),
    .sel(n46),
    .o(n47));  // ../RTL/cmsdk_apb_uart.v(368)
  and u56 (n104, rx_tick_cnt[2], rx_tick_cnt[3]);  // ../RTL/cmsdk_apb_uart.v(539)
  or u57 (n48, reload_i, reg_baud_tick);  // ../RTL/cmsdk_apb_uart.v(376)
  AL_MUX u58 (
    .i0(reg_baud_tick),
    .i1(reload_i),
    .sel(n48),
    .o(n49));  // ../RTL/cmsdk_apb_uart.v(377)
  buf u59 (BAUDTICK, reg_baud_tick);  // ../RTL/cmsdk_apb_uart.v(381)
  and u6 (n2, PSEL, n1);  // ../RTL/cmsdk_apb_uart.v(193)
  buf u60 (nxt_rx_buf[7], rx_shift_in);  // ../RTL/cmsdk_apb_uart.v(596)
  or u61 (n50, write_enable00, tx_buf_clear);  // ../RTL/cmsdk_apb_uart.v(391)
  AL_MUX u62 (
    .i0(tx_buf_full),
    .i1(write_enable00),
    .sel(n50),
    .o(n51));  // ../RTL/cmsdk_apb_uart.v(392)
  and u63 (n53, n52, reg_baud_tick);  // ../RTL/cmsdk_apb_uart.v(396)
  buf u64 (nxt_rx_buf[6], rx_shift_buf[6]);  // ../RTL/cmsdk_apb_uart.v(596)
  buf u65 (mapped_cntr_f[0], reg_baud_cntr_f[3]);  // ../RTL/cmsdk_apb_uart.v(322)
  buf u66 (nxt_rx_buf[5], rx_shift_buf[5]);  // ../RTL/cmsdk_apb_uart.v(596)
  or u67 (n58, n57, n52);  // ../RTL/cmsdk_apb_uart.v(409)
  and u68 (n59, n58, reg_baud_tick);  // ../RTL/cmsdk_apb_uart.v(409)
  or u69 (tx_state_inc, n59, reg_ctrl[6]);  // ../RTL/cmsdk_apb_uart.v(409)
  and u7 (write_enable, n2, PWRITE);  // ../RTL/cmsdk_apb_uart.v(193)
  and u70 (n61, n60, tx_buf_full);  // ../RTL/cmsdk_apb_uart.v(412)
  and u71 (n63, n62, tx_buf_full);  // ../RTL/cmsdk_apb_uart.v(413)
  and u72 (n64, n63, tx_state_inc);  // ../RTL/cmsdk_apb_uart.v(413)
  or u73 (tx_buf_clear, n61, n64);  // ../RTL/cmsdk_apb_uart.v(413)
  and u74 (n65, tx_buf_full, reg_ctrl[0]);  // ../RTL/cmsdk_apb_uart.v(423)
  not u75 (n103[3], rx_state_inc);  // ../RTL/cmsdk_apb_uart.v(568)
  buf u76 (nxt_rx_buf[4], rx_shift_buf[4]);  // ../RTL/cmsdk_apb_uart.v(596)
  buf u77 (nxt_rx_buf[3], rx_shift_buf[3]);  // ../RTL/cmsdk_apb_uart.v(596)
  and u78 (n69, n61, reg_ctrl[0]);  // ../RTL/cmsdk_apb_uart.v(437)
  or u79 (n70, tx_state_inc, n69);  // ../RTL/cmsdk_apb_uart.v(437)
  and u8 (write_enable00, write_enable, n3);  // ../RTL/cmsdk_apb_uart.v(194)
  or u80 (tx_state_update, n70, n71);  // ../RTL/cmsdk_apb_uart.v(437)
  buf u81 (nxt_rx_buf[2], rx_shift_buf[2]);  // ../RTL/cmsdk_apb_uart.v(596)
  buf u82 (nxt_rx_buf[1], rx_shift_buf[1]);  // ../RTL/cmsdk_apb_uart.v(596)
  buf u83 (nxt_rx_shift_buf[6], rx_shift_in);  // ../RTL/cmsdk_apb_uart.v(607)
  buf u84 (nxt_rx_shift_buf[5], rx_shift_buf[6]);  // ../RTL/cmsdk_apb_uart.v(607)
  buf u85 (nxt_rx_shift_buf[4], rx_shift_buf[5]);  // ../RTL/cmsdk_apb_uart.v(607)
  buf u86 (nxt_rx_shift_buf[3], rx_shift_buf[4]);  // ../RTL/cmsdk_apb_uart.v(607)
  buf u87 (nxt_rx_shift_buf[2], rx_shift_buf[3]);  // ../RTL/cmsdk_apb_uart.v(607)
  and u88 (tx_buf_ctrl_shift, n73, tx_state_inc);  // ../RTL/cmsdk_apb_uart.v(451)
  buf u89 (nxt_rx_shift_buf[1], rx_shift_buf[2]);  // ../RTL/cmsdk_apb_uart.v(607)
  and u9 (write_enable04, write_enable, n4);  // ../RTL/cmsdk_apb_uart.v(195)
  or u90 (n74, tx_buf_ctrl_shift, tx_buf_clear);  // ../RTL/cmsdk_apb_uart.v(460)
  and u91 (intr_stat_clear[1], write_enable0c, PWDATA[1]);  // ../RTL/cmsdk_apb_uart.v(626)
  buf u92 (read_mux_word[31], 1'b0);  // ../RTL/cmsdk_apb_uart.v(309)
  AL_MUX u93 (
    .i0(1'b1),
    .i1(tx_shift_buf[0]),
    .sel(n73),
    .o(n77));  // ../RTL/cmsdk_apb_uart.v(466)
  AL_MUX u94 (
    .i0(n77),
    .i1(1'b0),
    .sel(n76),
    .o(nxt_txd));  // ../RTL/cmsdk_apb_uart.v(466)
  xor u95 (update_reg_txd, nxt_txd, reg_txd);  // ../RTL/cmsdk_apb_uart.v(468)
  buf u96 (read_mux_word[30], 1'b0);  // ../RTL/cmsdk_apb_uart.v(309)
  AL_MUX u97 (
    .i0(reg_txd),
    .i1(nxt_txd),
    .sel(update_reg_txd),
    .o(n78));  // ../RTL/cmsdk_apb_uart.v(476)
  not u98 (n79, tx_buf_clear);  // ../RTL/cmsdk_apb_uart.v(480)
  and u99 (n80, tx_buf_full, n79);  // ../RTL/cmsdk_apb_uart.v(480)

endmodule 

module binary_mux_s1_w2
  (
  i0,
  i1,
  sel,
  o
  );

  input [1:0] i0;
  input [1:0] i1;
  input sel;
  output [1:0] o;



endmodule 

module ne_w2
  (
  i0,
  i1,
  o
  );

  input [1:0] i0;
  input [1:0] i1;
  output o;



endmodule 

module cmsdk_ahb_to_apb  // ../RTL/cmsdk_ahb_to_apb.v(31)
  (
  HADDR,
  HCLK,
  HPROT,
  HREADY,
  HRESETn,
  HSEL,
  HSIZE,
  HTRANS,
  HWDATA,
  HWRITE,
  PCLKEN,
  PRDATA,
  PREADY,
  PSLVERR,
  APBACTIVE,
  HRDATA,
  HREADYOUT,
  HRESP,
  PADDR,
  PENABLE,
  PPROT,
  PSEL,
  PSTRB,
  PWDATA,
  PWRITE
  );

  input [15:0] HADDR;  // ../RTL/cmsdk_ahb_to_apb.v(46)
  input HCLK;  // ../RTL/cmsdk_ahb_to_apb.v(41)
  input [3:0] HPROT;  // ../RTL/cmsdk_ahb_to_apb.v(49)
  input HREADY;  // ../RTL/cmsdk_ahb_to_apb.v(51)
  input HRESETn;  // ../RTL/cmsdk_ahb_to_apb.v(42)
  input HSEL;  // ../RTL/cmsdk_ahb_to_apb.v(45)
  input [2:0] HSIZE;  // ../RTL/cmsdk_ahb_to_apb.v(48)
  input [1:0] HTRANS;  // ../RTL/cmsdk_ahb_to_apb.v(47)
  input [31:0] HWDATA;  // ../RTL/cmsdk_ahb_to_apb.v(52)
  input HWRITE;  // ../RTL/cmsdk_ahb_to_apb.v(50)
  input PCLKEN;  // ../RTL/cmsdk_ahb_to_apb.v(43)
  input [31:0] PRDATA;  // ../RTL/cmsdk_ahb_to_apb.v(70)
  input PREADY;  // ../RTL/cmsdk_ahb_to_apb.v(71)
  input PSLVERR;  // ../RTL/cmsdk_ahb_to_apb.v(72)
  output APBACTIVE;  // ../RTL/cmsdk_ahb_to_apb.v(66)
  output [31:0] HRDATA;  // ../RTL/cmsdk_ahb_to_apb.v(55)
  output HREADYOUT;  // ../RTL/cmsdk_ahb_to_apb.v(54)
  output HRESP;  // ../RTL/cmsdk_ahb_to_apb.v(56)
  output [15:0] PADDR;  // ../RTL/cmsdk_ahb_to_apb.v(58)
  output PENABLE;  // ../RTL/cmsdk_ahb_to_apb.v(59)
  output [2:0] PPROT;  // ../RTL/cmsdk_ahb_to_apb.v(62)
  output PSEL;  // ../RTL/cmsdk_ahb_to_apb.v(64)
  output [3:0] PSTRB;  // ../RTL/cmsdk_ahb_to_apb.v(61)
  output [31:0] PWDATA;  // ../RTL/cmsdk_ahb_to_apb.v(63)
  output PWRITE;  // ../RTL/cmsdk_ahb_to_apb.v(60)

  parameter ADDRWIDTH = 16;
  parameter REGISTER_RDATA = 1;
  parameter REGISTER_WDATA = 0;
  // localparam ST_APB_ENDOK = 3'b100;
  // localparam ST_APB_ERR1 = 3'b101;
  // localparam ST_APB_ERR2 = 3'b110;
  // localparam ST_APB_TRNF = 3'b010;
  // localparam ST_APB_TRNF2 = 3'b011;
  // localparam ST_APB_WAIT = 3'b001;
  // localparam ST_BITS = 3;
  // localparam ST_IDLE = 3'b000;
  // localparam ST_ILLEGAL = 3'b111;
  wire [13:0] addr_reg;  // ../RTL/cmsdk_ahb_to_apb.v(78)
  wire [13:0] n10;
  wire [1:0] n12;
  wire [3:0] n13;
  wire [1:0] n21;
  wire [1:0] n22;
  wire [2:0] n28;
  wire [2:0] n29;
  wire [2:0] n30;
  wire [31:0] n36;
  wire [31:0] n37;
  wire [3:0] n4;
  wire [3:0] n5;
  wire [3:0] n6;
  wire [2:0] next_state;  // ../RTL/cmsdk_ahb_to_apb.v(89)
  wire [1:0] pprot_nxt;  // ../RTL/cmsdk_ahb_to_apb.v(85)
  wire [1:0] pprot_reg;  // ../RTL/cmsdk_ahb_to_apb.v(84)
  wire [3:0] pstrb_nxt;  // ../RTL/cmsdk_ahb_to_apb.v(83)
  wire [3:0] pstrb_reg;  // ../RTL/cmsdk_ahb_to_apb.v(82)
  wire [31:0] rwdata_reg;  // ../RTL/cmsdk_ahb_to_apb.v(90)
  wire [2:0] state_reg;  // ../RTL/cmsdk_ahb_to_apb.v(80)
  wire apb_select;  // ../RTL/cmsdk_ahb_to_apb.v(87)
  wire apb_tran_end;  // ../RTL/cmsdk_ahb_to_apb.v(88)
  wire n0;
  wire n1;
  wire n11;
  wire n14;
  wire n15;
  wire n16;
  wire n17;
  wire n18;
  wire n19;
  wire n2;
  wire n20;
  wire n23;
  wire n24;
  wire n25;
  wire n26;
  wire n27;
  wire n3;
  wire n31;
  wire n32;
  wire n33;
  wire n34;
  wire n35;
  wire n38;
  wire n39;
  wire n40;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n7;
  wire n8;
  wire n9;
  wire reg_rdata_cfg;  // ../RTL/cmsdk_ahb_to_apb.v(92)
  wire reg_wdata_cfg;  // ../RTL/cmsdk_ahb_to_apb.v(93)
  wire sample_wdata_clr;  // ../RTL/cmsdk_ahb_to_apb.v(159)
  wire sample_wdata_reg;  // ../RTL/cmsdk_ahb_to_apb.v(95)
  wire sample_wdata_set;  // ../RTL/cmsdk_ahb_to_apb.v(158)
  wire wr_reg;  // ../RTL/cmsdk_ahb_to_apb.v(79)

  eq_w3 eq0 (
    .i0(state_reg),
    .i1(3'b011),
    .o(PENABLE));  // ../RTL/cmsdk_ahb_to_apb.v(122)
  eq_w2 eq1 (
    .i0(HADDR[1:0]),
    .i1(2'b00),
    .o(n3));  // ../RTL/cmsdk_ahb_to_apb.v(132)
  eq_w2 eq2 (
    .i0(HADDR[1:0]),
    .i1(2'b01),
    .o(n7));  // ../RTL/cmsdk_ahb_to_apb.v(133)
  eq_w2 eq3 (
    .i0(HADDR[1:0]),
    .i1(2'b10),
    .o(n8));  // ../RTL/cmsdk_ahb_to_apb.v(134)
  eq_w2 eq4 (
    .i0(HADDR[1:0]),
    .i1(2'b11),
    .o(n9));  // ../RTL/cmsdk_ahb_to_apb.v(135)
  eq_w3 eq5 (
    .i0(state_reg),
    .i1(3'b010),
    .o(n38));  // ../RTL/cmsdk_ahb_to_apb.v(273)
  eq_w3 eq6 (
    .i0(state_reg),
    .i1(3'b101),
    .o(n43));  // ../RTL/cmsdk_ahb_to_apb.v(299)
  eq_w3 eq7 (
    .i0(state_reg),
    .i1(3'b110),
    .o(n44));  // ../RTL/cmsdk_ahb_to_apb.v(299)
  binary_mux_s1_w14 mux0 (
    .i0(addr_reg),
    .i1(HADDR[15:2]),
    .sel(apb_select),
    .o(n10));  // ../RTL/cmsdk_ahb_to_apb.v(153)
  binary_mux_s1_w2 mux1 (
    .i0(pprot_reg),
    .i1(pprot_nxt),
    .sel(apb_select),
    .o(n12));  // ../RTL/cmsdk_ahb_to_apb.v(153)
  binary_mux_s1_w32 mux10 (
    .i0(HWDATA),
    .i1(rwdata_reg),
    .sel(reg_wdata_cfg),
    .o(PWDATA));  // ../RTL/cmsdk_ahb_to_apb.v(272)
  binary_mux_s3_w1 mux11 (
    .i0(1'b1),
    .i1(1'b0),
    .i2(1'b0),
    .i3(n42),
    .i4(reg_rdata_cfg),
    .i5(1'b0),
    .i6(1'b1),
    .i7(1'bx),
    .sel(state_reg),
    .o(HREADYOUT));  // ../RTL/cmsdk_ahb_to_apb.v(294)
  binary_mux_s1_w32 mux12 (
    .i0(PRDATA),
    .i1(rwdata_reg),
    .sel(reg_rdata_cfg),
    .o(HRDATA));  // ../RTL/cmsdk_ahb_to_apb.v(298)
  binary_mux_s1_w4 mux2 (
    .i0(pstrb_reg),
    .i1(pstrb_nxt),
    .sel(apb_select),
    .o(n13));  // ../RTL/cmsdk_ahb_to_apb.v(153)
  binary_mux_s1_w2 mux3 (
    .i0({1'b0,apb_select}),
    .i1(2'b10),
    .sel(n20),
    .o(n21));  // ../RTL/cmsdk_ahb_to_apb.v(184)
  binary_mux_s1_w3 mux4 (
    .i0({2'b00,apb_select}),
    .i1(3'b100),
    .sel(reg_rdata_cfg),
    .o(n28));  // ../RTL/cmsdk_ahb_to_apb.v(215)
  binary_mux_s1_w3 mux5 (
    .i0(3'b011),
    .i1(n28),
    .sel(n27),
    .o(n29));  // ../RTL/cmsdk_ahb_to_apb.v(218)
  binary_mux_s1_w3 mux6 (
    .i0(n29),
    .i1(3'b101),
    .sel(n24),
    .o(n30));  // ../RTL/cmsdk_ahb_to_apb.v(218)
  binary_mux_s3_w3 mux7 (
    .i0({1'b0,n21}),
    .i1({1'b0,PCLKEN,n22[0]}),
    .i2({2'b01,PCLKEN}),
    .i3(n30),
    .i4({1'b0,n21}),
    .i5(3'b110),
    .i6({1'b0,n21}),
    .i7(3'bxxx),
    .sel(state_reg),
    .o(next_state));  // ../RTL/cmsdk_ahb_to_apb.v(244)
  binary_mux_s1_w32 mux8 (
    .i0(rwdata_reg),
    .i1(PRDATA),
    .sel(n35),
    .o(n36));  // ../RTL/cmsdk_ahb_to_apb.v(265)
  binary_mux_s1_w32 mux9 (
    .i0(n36),
    .i1(HWDATA),
    .sel(n33),
    .o(n37));  // ../RTL/cmsdk_ahb_to_apb.v(265)
  reg_ar_as_w2 reg0 (
    .clk(HCLK),
    .d(n12),
    .reset({n31,n31}),
    .set(2'b00),
    .q(pprot_reg));  // ../RTL/cmsdk_ahb_to_apb.v(153)
  reg_ar_as_w4 reg1 (
    .clk(HCLK),
    .d(n13),
    .reset({n31,n31,n31,n31}),
    .set(4'b0000),
    .q(pstrb_reg));  // ../RTL/cmsdk_ahb_to_apb.v(153)
  reg_ar_as_w3 reg2 (
    .clk(HCLK),
    .d(next_state),
    .reset({n31,n31,n31}),
    .set(3'b000),
    .q(state_reg));  // ../RTL/cmsdk_ahb_to_apb.v(253)
  reg_ar_as_w32 reg3 (
    .clk(HCLK),
    .d(n37),
    .reset({n31,n31,n31,n31,n31,n31,n31,n31,n31,n31,n31,n31,n31,n31,n31,n31,n31,n31,n31,n31,n31,n31,n31,n31,n31,n31,n31,n31,n31,n31,n31,n31}),
    .set(32'b00000000000000000000000000000000),
    .q(rwdata_reg));  // ../RTL/cmsdk_ahb_to_apb.v(265)
  reg_ar_as_w14 reg4 (
    .clk(HCLK),
    .d(n10),
    .reset({n31,n31,n31,n31,n31,n31,n31,n31,n31,n31,n31,n31,n31,n31}),
    .set(14'b00000000000000),
    .q(addr_reg));  // ../RTL/cmsdk_ahb_to_apb.v(153)
  AL_DFF sample_wdata_reg_reg (
    .clk(HCLK),
    .d(n16),
    .reset(n31),
    .set(1'b0),
    .q(sample_wdata_reg));  // ../RTL/cmsdk_ahb_to_apb.v(166)
  not u10 (pprot_nxt[1], HPROT[0]);  // ../RTL/cmsdk_ahb_to_apb.v(125)
  not u11 (n1, HADDR[1]);  // ../RTL/cmsdk_ahb_to_apb.v(132)
  or u12 (n6[3], HSIZE[1], n5[3]);  // ../RTL/cmsdk_ahb_to_apb.v(135)
  or u13 (n4[3], n6[3], n9);  // ../RTL/cmsdk_ahb_to_apb.v(135)
  buf u14 (PADDR[10], addr_reg[8]);  // ../RTL/cmsdk_ahb_to_apb.v(269)
  and u15 (pstrb_nxt[3], HWRITE, n4[3]);  // ../RTL/cmsdk_ahb_to_apb.v(135)
  or u16 (n4[2], n6[3], n8);  // ../RTL/cmsdk_ahb_to_apb.v(135)
  and u17 (pstrb_nxt[2], HWRITE, n4[2]);  // ../RTL/cmsdk_ahb_to_apb.v(135)
  or u18 (n4[1], n6[1], n7);  // ../RTL/cmsdk_ahb_to_apb.v(135)
  and u19 (pstrb_nxt[1], HWRITE, n4[1]);  // ../RTL/cmsdk_ahb_to_apb.v(135)
  or u20 (n2, state_reg[1], state_reg[2]);  // ../RTL/cmsdk_ahb_to_apb.v(301)
  not u21 (n22[0], PCLKEN);  // ../RTL/cmsdk_ahb_to_apb.v(192)
  buf u22 (PADDR[14], addr_reg[12]);  // ../RTL/cmsdk_ahb_to_apb.v(269)
  not u23 (n31, HRESETn);  // ../RTL/cmsdk_ahb_to_apb.v(140)
  AL_MUX u24 (
    .i0(wr_reg),
    .i1(HWRITE),
    .sel(apb_select),
    .o(n11));  // ../RTL/cmsdk_ahb_to_apb.v(153)
  and u25 (n14, apb_select, HWRITE);  // ../RTL/cmsdk_ahb_to_apb.v(158)
  and u26 (sample_wdata_set, n14, reg_wdata_cfg);  // ../RTL/cmsdk_ahb_to_apb.v(158)
  and u27 (sample_wdata_clr, sample_wdata_reg, PCLKEN);  // ../RTL/cmsdk_ahb_to_apb.v(159)
  buf u28 (PADDR[13], addr_reg[11]);  // ../RTL/cmsdk_ahb_to_apb.v(269)
  buf u29 (PADDR[9], addr_reg[7]);  // ../RTL/cmsdk_ahb_to_apb.v(269)
  buf u3 (PADDR[15], addr_reg[13]);  // ../RTL/cmsdk_ahb_to_apb.v(269)
  or u30 (n15, sample_wdata_set, sample_wdata_clr);  // ../RTL/cmsdk_ahb_to_apb.v(165)
  AL_MUX u31 (
    .i0(sample_wdata_reg),
    .i1(sample_wdata_set),
    .sel(n15),
    .o(n16));  // ../RTL/cmsdk_ahb_to_apb.v(166)
  and u32 (n17, PCLKEN, apb_select);  // ../RTL/cmsdk_ahb_to_apb.v(179)
  and u33 (n18, reg_wdata_cfg, HWRITE);  // ../RTL/cmsdk_ahb_to_apb.v(179)
  not u34 (n19, n18);  // ../RTL/cmsdk_ahb_to_apb.v(179)
  and u35 (n20, n17, n19);  // ../RTL/cmsdk_ahb_to_apb.v(179)
  buf u36 (PADDR[11], addr_reg[9]);  // ../RTL/cmsdk_ahb_to_apb.v(269)
  and u37 (n23, PREADY, PSLVERR);  // ../RTL/cmsdk_ahb_to_apb.v(205)
  and u38 (n24, n23, PCLKEN);  // ../RTL/cmsdk_ahb_to_apb.v(205)
  not u39 (n25, PSLVERR);  // ../RTL/cmsdk_ahb_to_apb.v(208)
  buf u4 (reg_rdata_cfg, 1'b1);  // ../RTL/cmsdk_ahb_to_apb.v(116)
  and u40 (n26, PREADY, n25);  // ../RTL/cmsdk_ahb_to_apb.v(208)
  and u41 (n27, n26, PCLKEN);  // ../RTL/cmsdk_ahb_to_apb.v(208)
  buf u42 (PADDR[8], addr_reg[6]);  // ../RTL/cmsdk_ahb_to_apb.v(269)
  buf u43 (PADDR[7], addr_reg[5]);  // ../RTL/cmsdk_ahb_to_apb.v(269)
  buf u44 (PADDR[6], addr_reg[4]);  // ../RTL/cmsdk_ahb_to_apb.v(269)
  buf u45 (PADDR[5], addr_reg[3]);  // ../RTL/cmsdk_ahb_to_apb.v(269)
  buf u46 (PADDR[4], addr_reg[2]);  // ../RTL/cmsdk_ahb_to_apb.v(269)
  buf u47 (PADDR[3], addr_reg[1]);  // ../RTL/cmsdk_ahb_to_apb.v(269)
  buf u48 (PADDR[2], addr_reg[0]);  // ../RTL/cmsdk_ahb_to_apb.v(269)
  buf u49 (PADDR[1], 1'b0);  // ../RTL/cmsdk_ahb_to_apb.v(269)
  buf u5 (reg_wdata_cfg, 1'b0);  // ../RTL/cmsdk_ahb_to_apb.v(117)
  buf u50 (PPROT[2], pprot_reg[1]);  // ../RTL/cmsdk_ahb_to_apb.v(275)
  buf u51 (PPROT[1], 1'b0);  // ../RTL/cmsdk_ahb_to_apb.v(275)
  buf u52 (PADDR[12], addr_reg[10]);  // ../RTL/cmsdk_ahb_to_apb.v(269)
  buf u53 (PSTRB[3], pstrb_reg[3]);  // ../RTL/cmsdk_ahb_to_apb.v(276)
  or u54 (n4[0], n6[1], n3);  // ../RTL/cmsdk_ahb_to_apb.v(135)
  buf u55 (PSTRB[2], pstrb_reg[2]);  // ../RTL/cmsdk_ahb_to_apb.v(276)
  and u56 (n32, sample_wdata_reg, reg_wdata_cfg);  // ../RTL/cmsdk_ahb_to_apb.v(262)
  and u57 (n33, n32, PCLKEN);  // ../RTL/cmsdk_ahb_to_apb.v(262)
  and u58 (n34, apb_tran_end, reg_rdata_cfg);  // ../RTL/cmsdk_ahb_to_apb.v(264)
  and u59 (n35, n34, PCLKEN);  // ../RTL/cmsdk_ahb_to_apb.v(264)
  and u6 (n0, HSEL, HTRANS[1]);  // ../RTL/cmsdk_ahb_to_apb.v(120)
  or u60 (n6[1], HSIZE[1], n5[1]);  // ../RTL/cmsdk_ahb_to_apb.v(135)
  and u61 (pstrb_nxt[0], HWRITE, n4[0]);  // ../RTL/cmsdk_ahb_to_apb.v(135)
  buf u62 (PWRITE, wr_reg);  // ../RTL/cmsdk_ahb_to_apb.v(270)
  buf u63 (PSTRB[1], pstrb_reg[1]);  // ../RTL/cmsdk_ahb_to_apb.v(276)
  or u64 (PSEL, n38, PENABLE);  // ../RTL/cmsdk_ahb_to_apb.v(273)
  and u65 (n5[3], HSIZE[0], HADDR[1]);  // ../RTL/cmsdk_ahb_to_apb.v(135)
  buf u66 (PADDR[0], 1'b0);  // ../RTL/cmsdk_ahb_to_apb.v(269)
  buf u67 (PPROT[0], pprot_reg[0]);  // ../RTL/cmsdk_ahb_to_apb.v(275)
  not u68 (n39, reg_rdata_cfg);  // ../RTL/cmsdk_ahb_to_apb.v(289)
  and u69 (n40, n39, PREADY);  // ../RTL/cmsdk_ahb_to_apb.v(289)
  and u7 (apb_select, n0, HREADY);  // ../RTL/cmsdk_ahb_to_apb.v(120)
  or u70 (n45, state_reg[0], n2);  // ../RTL/cmsdk_ahb_to_apb.v(301)
  and u71 (n41, n40, n25);  // ../RTL/cmsdk_ahb_to_apb.v(289)
  and u72 (n42, n41, PCLKEN);  // ../RTL/cmsdk_ahb_to_apb.v(289)
  or u73 (HRESP, n43, n44);  // ../RTL/cmsdk_ahb_to_apb.v(299)
  buf u74 (PSTRB[0], pstrb_reg[0]);  // ../RTL/cmsdk_ahb_to_apb.v(276)
  and u75 (n5[1], HSIZE[0], n1);  // ../RTL/cmsdk_ahb_to_apb.v(135)
  or u76 (APBACTIVE, n0, n45);  // ../RTL/cmsdk_ahb_to_apb.v(301)
  and u8 (apb_tran_end, PENABLE, PREADY);  // ../RTL/cmsdk_ahb_to_apb.v(122)
  buf u9 (pprot_nxt[0], HPROT[1]);  // ../RTL/cmsdk_ahb_to_apb.v(124)
  AL_DFF wr_reg_reg (
    .clk(HCLK),
    .d(n11),
    .reset(n31),
    .set(1'b0),
    .q(wr_reg));  // ../RTL/cmsdk_ahb_to_apb.v(153)

endmodule 

module \cmsdk_apb_slave_mux(PORT1_ENABLE=0,PORT2_ENABLE=0,PORT3_ENABLE=0,PORT5_ENABLE=0,PORT6_ENABLE=0,PORT7_ENABLE=0,PORT8_ENABLE=0,PORT9_ENABLE=0,PORT10_ENABLE=0,PORT11_ENABLE=0,PORT12_ENABLE=0,PORT13_ENABLE=0,PORT14_ENABLE=0,PORT15_ENABLE=0)   // ../RTL/cmsdk_apb_slave_mux.v(26)
  (
  DECODE4BIT,
  PRDATA0,
  PRDATA1,
  PRDATA10,
  PRDATA11,
  PRDATA12,
  PRDATA13,
  PRDATA14,
  PRDATA15,
  PRDATA2,
  PRDATA3,
  PRDATA4,
  PRDATA5,
  PRDATA6,
  PRDATA7,
  PRDATA8,
  PRDATA9,
  PREADY0,
  PREADY1,
  PREADY10,
  PREADY11,
  PREADY12,
  PREADY13,
  PREADY14,
  PREADY15,
  PREADY2,
  PREADY3,
  PREADY4,
  PREADY5,
  PREADY6,
  PREADY7,
  PREADY8,
  PREADY9,
  PSEL,
  PSLVERR0,
  PSLVERR1,
  PSLVERR10,
  PSLVERR11,
  PSLVERR12,
  PSLVERR13,
  PSLVERR14,
  PSLVERR15,
  PSLVERR2,
  PSLVERR3,
  PSLVERR4,
  PSLVERR5,
  PSLVERR6,
  PSLVERR7,
  PSLVERR8,
  PSLVERR9,
  PRDATA,
  PREADY,
  PSEL0,
  PSEL1,
  PSEL10,
  PSEL11,
  PSEL12,
  PSEL13,
  PSEL14,
  PSEL15,
  PSEL2,
  PSEL3,
  PSEL4,
  PSEL5,
  PSEL6,
  PSEL7,
  PSEL8,
  PSEL9,
  PSLVERR
  );

  input [3:0] DECODE4BIT;  // ../RTL/cmsdk_apb_slave_mux.v(48)
  input [31:0] PRDATA0;  // ../RTL/cmsdk_apb_slave_mux.v(53)
  input [31:0] PRDATA1;  // ../RTL/cmsdk_apb_slave_mux.v(58)
  input [31:0] PRDATA10;  // ../RTL/cmsdk_apb_slave_mux.v(103)
  input [31:0] PRDATA11;  // ../RTL/cmsdk_apb_slave_mux.v(108)
  input [31:0] PRDATA12;  // ../RTL/cmsdk_apb_slave_mux.v(113)
  input [31:0] PRDATA13;  // ../RTL/cmsdk_apb_slave_mux.v(118)
  input [31:0] PRDATA14;  // ../RTL/cmsdk_apb_slave_mux.v(123)
  input [31:0] PRDATA15;  // ../RTL/cmsdk_apb_slave_mux.v(128)
  input [31:0] PRDATA2;  // ../RTL/cmsdk_apb_slave_mux.v(63)
  input [31:0] PRDATA3;  // ../RTL/cmsdk_apb_slave_mux.v(68)
  input [31:0] PRDATA4;  // ../RTL/cmsdk_apb_slave_mux.v(73)
  input [31:0] PRDATA5;  // ../RTL/cmsdk_apb_slave_mux.v(78)
  input [31:0] PRDATA6;  // ../RTL/cmsdk_apb_slave_mux.v(83)
  input [31:0] PRDATA7;  // ../RTL/cmsdk_apb_slave_mux.v(88)
  input [31:0] PRDATA8;  // ../RTL/cmsdk_apb_slave_mux.v(93)
  input [31:0] PRDATA9;  // ../RTL/cmsdk_apb_slave_mux.v(98)
  input PREADY0;  // ../RTL/cmsdk_apb_slave_mux.v(52)
  input PREADY1;  // ../RTL/cmsdk_apb_slave_mux.v(57)
  input PREADY10;  // ../RTL/cmsdk_apb_slave_mux.v(102)
  input PREADY11;  // ../RTL/cmsdk_apb_slave_mux.v(107)
  input PREADY12;  // ../RTL/cmsdk_apb_slave_mux.v(112)
  input PREADY13;  // ../RTL/cmsdk_apb_slave_mux.v(117)
  input PREADY14;  // ../RTL/cmsdk_apb_slave_mux.v(122)
  input PREADY15;  // ../RTL/cmsdk_apb_slave_mux.v(127)
  input PREADY2;  // ../RTL/cmsdk_apb_slave_mux.v(62)
  input PREADY3;  // ../RTL/cmsdk_apb_slave_mux.v(67)
  input PREADY4;  // ../RTL/cmsdk_apb_slave_mux.v(72)
  input PREADY5;  // ../RTL/cmsdk_apb_slave_mux.v(77)
  input PREADY6;  // ../RTL/cmsdk_apb_slave_mux.v(82)
  input PREADY7;  // ../RTL/cmsdk_apb_slave_mux.v(87)
  input PREADY8;  // ../RTL/cmsdk_apb_slave_mux.v(92)
  input PREADY9;  // ../RTL/cmsdk_apb_slave_mux.v(97)
  input PSEL;  // ../RTL/cmsdk_apb_slave_mux.v(49)
  input PSLVERR0;  // ../RTL/cmsdk_apb_slave_mux.v(54)
  input PSLVERR1;  // ../RTL/cmsdk_apb_slave_mux.v(59)
  input PSLVERR10;  // ../RTL/cmsdk_apb_slave_mux.v(104)
  input PSLVERR11;  // ../RTL/cmsdk_apb_slave_mux.v(109)
  input PSLVERR12;  // ../RTL/cmsdk_apb_slave_mux.v(114)
  input PSLVERR13;  // ../RTL/cmsdk_apb_slave_mux.v(119)
  input PSLVERR14;  // ../RTL/cmsdk_apb_slave_mux.v(124)
  input PSLVERR15;  // ../RTL/cmsdk_apb_slave_mux.v(129)
  input PSLVERR2;  // ../RTL/cmsdk_apb_slave_mux.v(64)
  input PSLVERR3;  // ../RTL/cmsdk_apb_slave_mux.v(69)
  input PSLVERR4;  // ../RTL/cmsdk_apb_slave_mux.v(74)
  input PSLVERR5;  // ../RTL/cmsdk_apb_slave_mux.v(79)
  input PSLVERR6;  // ../RTL/cmsdk_apb_slave_mux.v(84)
  input PSLVERR7;  // ../RTL/cmsdk_apb_slave_mux.v(89)
  input PSLVERR8;  // ../RTL/cmsdk_apb_slave_mux.v(94)
  input PSLVERR9;  // ../RTL/cmsdk_apb_slave_mux.v(99)
  output [31:0] PRDATA;  // ../RTL/cmsdk_apb_slave_mux.v(132)
  output PREADY;  // ../RTL/cmsdk_apb_slave_mux.v(131)
  output PSEL0;  // ../RTL/cmsdk_apb_slave_mux.v(51)
  output PSEL1;  // ../RTL/cmsdk_apb_slave_mux.v(56)
  output PSEL10;  // ../RTL/cmsdk_apb_slave_mux.v(101)
  output PSEL11;  // ../RTL/cmsdk_apb_slave_mux.v(106)
  output PSEL12;  // ../RTL/cmsdk_apb_slave_mux.v(111)
  output PSEL13;  // ../RTL/cmsdk_apb_slave_mux.v(116)
  output PSEL14;  // ../RTL/cmsdk_apb_slave_mux.v(121)
  output PSEL15;  // ../RTL/cmsdk_apb_slave_mux.v(126)
  output PSEL2;  // ../RTL/cmsdk_apb_slave_mux.v(61)
  output PSEL3;  // ../RTL/cmsdk_apb_slave_mux.v(66)
  output PSEL4;  // ../RTL/cmsdk_apb_slave_mux.v(71)
  output PSEL5;  // ../RTL/cmsdk_apb_slave_mux.v(76)
  output PSEL6;  // ../RTL/cmsdk_apb_slave_mux.v(81)
  output PSEL7;  // ../RTL/cmsdk_apb_slave_mux.v(86)
  output PSEL8;  // ../RTL/cmsdk_apb_slave_mux.v(91)
  output PSEL9;  // ../RTL/cmsdk_apb_slave_mux.v(96)
  output PSLVERR;  // ../RTL/cmsdk_apb_slave_mux.v(133)

  parameter PORT0_ENABLE = 1;
  parameter PORT10_ENABLE = 0;
  parameter PORT11_ENABLE = 0;
  parameter PORT12_ENABLE = 0;
  parameter PORT13_ENABLE = 0;
  parameter PORT14_ENABLE = 0;
  parameter PORT15_ENABLE = 0;
  parameter PORT1_ENABLE = 0;
  parameter PORT2_ENABLE = 0;
  parameter PORT3_ENABLE = 0;
  parameter PORT4_ENABLE = 1;
  parameter PORT5_ENABLE = 0;
  parameter PORT6_ENABLE = 0;
  parameter PORT7_ENABLE = 0;
  parameter PORT8_ENABLE = 0;
  parameter PORT9_ENABLE = 0;
  wire [15:0] dec;  // ../RTL/cmsdk_apb_slave_mux.v(148)
  wire [15:0] en;  // ../RTL/cmsdk_apb_slave_mux.v(139)
  wire [31:0] n110;
  wire [31:0] n111;
  wire [31:0] n112;
  wire [31:0] n113;
  wire [31:0] n114;
  wire [31:0] n115;
  wire [31:0] n116;
  wire [31:0] n117;
  wire [31:0] n118;
  wire [31:0] n119;
  wire [31:0] n120;
  wire [31:0] n121;
  wire [31:0] n122;
  wire [31:0] n123;
  wire [31:0] n124;
  wire [31:0] n125;
  wire [31:0] n126;
  wire [31:0] n127;
  wire [31:0] n128;
  wire [31:0] n129;
  wire [31:0] n130;
  wire [31:0] n131;
  wire [31:0] n132;
  wire [31:0] n133;
  wire [31:0] n134;
  wire [31:0] n135;
  wire [31:0] n136;
  wire [31:0] n137;
  wire [31:0] n138;
  wire [31:0] n139;
  wire n0;
  wire n1;
  wire n10;
  wire n100;
  wire n101;
  wire n102;
  wire n103;
  wire n104;
  wire n105;
  wire n106;
  wire n107;
  wire n108;
  wire n109;
  wire n11;
  wire n12;
  wire n13;
  wire n14;
  wire n15;
  wire n16;
  wire n17;
  wire n18;
  wire n19;
  wire n2;
  wire n20;
  wire n21;
  wire n22;
  wire n23;
  wire n24;
  wire n25;
  wire n26;
  wire n27;
  wire n28;
  wire n29;
  wire n3;
  wire n30;
  wire n31;
  wire n32;
  wire n33;
  wire n34;
  wire n35;
  wire n36;
  wire n37;
  wire n38;
  wire n39;
  wire n4;
  wire n40;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n5;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n6;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n65;
  wire n66;
  wire n67;
  wire n68;
  wire n69;
  wire n7;
  wire n70;
  wire n71;
  wire n72;
  wire n73;
  wire n74;
  wire n75;
  wire n76;
  wire n77;
  wire n78;
  wire n79;
  wire n8;
  wire n80;
  wire n81;
  wire n82;
  wire n83;
  wire n84;
  wire n85;
  wire n86;
  wire n87;
  wire n88;
  wire n89;
  wire n9;
  wire n90;
  wire n91;
  wire n92;
  wire n93;
  wire n94;
  wire n95;
  wire n96;
  wire n97;
  wire n98;
  wire n99;

  eq_w4 eq0 (
    .i0(DECODE4BIT),
    .i1(4'b1111),
    .o(dec[15]));  // ../RTL/cmsdk_apb_slave_mux.v(148)
  eq_w4 eq1 (
    .i0(DECODE4BIT),
    .i1(4'b1110),
    .o(dec[14]));  // ../RTL/cmsdk_apb_slave_mux.v(148)
  eq_w4 eq10 (
    .i0(DECODE4BIT),
    .i1(4'b0101),
    .o(dec[5]));  // ../RTL/cmsdk_apb_slave_mux.v(153)
  eq_w4 eq11 (
    .i0(DECODE4BIT),
    .i1(4'b0100),
    .o(dec[4]));  // ../RTL/cmsdk_apb_slave_mux.v(153)
  eq_w4 eq12 (
    .i0(DECODE4BIT),
    .i1(4'b0011),
    .o(dec[3]));  // ../RTL/cmsdk_apb_slave_mux.v(154)
  eq_w4 eq13 (
    .i0(DECODE4BIT),
    .i1(4'b0010),
    .o(dec[2]));  // ../RTL/cmsdk_apb_slave_mux.v(154)
  eq_w4 eq14 (
    .i0(DECODE4BIT),
    .i1(4'b0001),
    .o(dec[1]));  // ../RTL/cmsdk_apb_slave_mux.v(155)
  eq_w4 eq15 (
    .i0(DECODE4BIT),
    .i1(4'b0000),
    .o(dec[0]));  // ../RTL/cmsdk_apb_slave_mux.v(155)
  eq_w4 eq2 (
    .i0(DECODE4BIT),
    .i1(4'b1101),
    .o(dec[13]));  // ../RTL/cmsdk_apb_slave_mux.v(149)
  eq_w4 eq3 (
    .i0(DECODE4BIT),
    .i1(4'b1100),
    .o(dec[12]));  // ../RTL/cmsdk_apb_slave_mux.v(149)
  eq_w4 eq4 (
    .i0(DECODE4BIT),
    .i1(4'b1011),
    .o(dec[11]));  // ../RTL/cmsdk_apb_slave_mux.v(150)
  eq_w4 eq5 (
    .i0(DECODE4BIT),
    .i1(4'b1010),
    .o(dec[10]));  // ../RTL/cmsdk_apb_slave_mux.v(150)
  eq_w4 eq6 (
    .i0(DECODE4BIT),
    .i1(4'b1001),
    .o(dec[9]));  // ../RTL/cmsdk_apb_slave_mux.v(151)
  eq_w4 eq7 (
    .i0(DECODE4BIT),
    .i1(4'b1000),
    .o(dec[8]));  // ../RTL/cmsdk_apb_slave_mux.v(151)
  eq_w4 eq8 (
    .i0(DECODE4BIT),
    .i1(4'b0111),
    .o(dec[7]));  // ../RTL/cmsdk_apb_slave_mux.v(152)
  eq_w4 eq9 (
    .i0(DECODE4BIT),
    .i1(4'b0110),
    .o(dec[6]));  // ../RTL/cmsdk_apb_slave_mux.v(152)
  and u10 (n3, PSEL, dec[3]);  // ../RTL/cmsdk_apb_slave_mux.v(160)
  or u100 (PREADY, n76, n79);  // ../RTL/cmsdk_apb_slave_mux.v(190)
  and u1000 (n115[2], PSEL3, PRDATA3[2]);  // ../RTL/cmsdk_apb_slave_mux.v(212)
  and u1001 (n115[3], PSEL3, PRDATA3[3]);  // ../RTL/cmsdk_apb_slave_mux.v(212)
  and u1002 (n115[4], PSEL3, PRDATA3[4]);  // ../RTL/cmsdk_apb_slave_mux.v(212)
  and u1003 (n115[5], PSEL3, PRDATA3[5]);  // ../RTL/cmsdk_apb_slave_mux.v(212)
  and u1004 (n115[6], PSEL3, PRDATA3[6]);  // ../RTL/cmsdk_apb_slave_mux.v(212)
  and u1005 (n115[7], PSEL3, PRDATA3[7]);  // ../RTL/cmsdk_apb_slave_mux.v(212)
  and u1006 (n115[8], PSEL3, PRDATA3[8]);  // ../RTL/cmsdk_apb_slave_mux.v(212)
  and u1007 (n115[9], PSEL3, PRDATA3[9]);  // ../RTL/cmsdk_apb_slave_mux.v(212)
  and u1008 (n115[10], PSEL3, PRDATA3[10]);  // ../RTL/cmsdk_apb_slave_mux.v(212)
  and u1009 (n115[11], PSEL3, PRDATA3[11]);  // ../RTL/cmsdk_apb_slave_mux.v(212)
  and u101 (n80, PSEL0, PSLVERR0);  // ../RTL/cmsdk_apb_slave_mux.v(192)
  and u1010 (n115[12], PSEL3, PRDATA3[12]);  // ../RTL/cmsdk_apb_slave_mux.v(212)
  and u1011 (n115[13], PSEL3, PRDATA3[13]);  // ../RTL/cmsdk_apb_slave_mux.v(212)
  and u1012 (n115[14], PSEL3, PRDATA3[14]);  // ../RTL/cmsdk_apb_slave_mux.v(212)
  and u1013 (n115[15], PSEL3, PRDATA3[15]);  // ../RTL/cmsdk_apb_slave_mux.v(212)
  and u1014 (n115[16], PSEL3, PRDATA3[16]);  // ../RTL/cmsdk_apb_slave_mux.v(212)
  and u1015 (n115[17], PSEL3, PRDATA3[17]);  // ../RTL/cmsdk_apb_slave_mux.v(212)
  and u1016 (n115[18], PSEL3, PRDATA3[18]);  // ../RTL/cmsdk_apb_slave_mux.v(212)
  and u1017 (n115[19], PSEL3, PRDATA3[19]);  // ../RTL/cmsdk_apb_slave_mux.v(212)
  and u1018 (n115[20], PSEL3, PRDATA3[20]);  // ../RTL/cmsdk_apb_slave_mux.v(212)
  and u1019 (n115[21], PSEL3, PRDATA3[21]);  // ../RTL/cmsdk_apb_slave_mux.v(212)
  and u102 (n81, PSEL1, PSLVERR1);  // ../RTL/cmsdk_apb_slave_mux.v(193)
  and u1020 (n115[22], PSEL3, PRDATA3[22]);  // ../RTL/cmsdk_apb_slave_mux.v(212)
  and u1021 (n115[23], PSEL3, PRDATA3[23]);  // ../RTL/cmsdk_apb_slave_mux.v(212)
  and u1022 (n115[24], PSEL3, PRDATA3[24]);  // ../RTL/cmsdk_apb_slave_mux.v(212)
  and u1023 (n115[25], PSEL3, PRDATA3[25]);  // ../RTL/cmsdk_apb_slave_mux.v(212)
  and u1024 (n115[26], PSEL3, PRDATA3[26]);  // ../RTL/cmsdk_apb_slave_mux.v(212)
  and u1025 (n115[27], PSEL3, PRDATA3[27]);  // ../RTL/cmsdk_apb_slave_mux.v(212)
  and u1026 (n115[28], PSEL3, PRDATA3[28]);  // ../RTL/cmsdk_apb_slave_mux.v(212)
  and u1027 (n115[29], PSEL3, PRDATA3[29]);  // ../RTL/cmsdk_apb_slave_mux.v(212)
  and u1028 (n115[30], PSEL3, PRDATA3[30]);  // ../RTL/cmsdk_apb_slave_mux.v(212)
  and u1029 (n115[31], PSEL3, PRDATA3[31]);  // ../RTL/cmsdk_apb_slave_mux.v(212)
  or u103 (n82, n80, n81);  // ../RTL/cmsdk_apb_slave_mux.v(193)
  or u1030 (n114[1], n112[1], n113[1]);  // ../RTL/cmsdk_apb_slave_mux.v(211)
  or u1031 (n114[2], n112[2], n113[2]);  // ../RTL/cmsdk_apb_slave_mux.v(211)
  or u1032 (n114[3], n112[3], n113[3]);  // ../RTL/cmsdk_apb_slave_mux.v(211)
  or u1033 (n114[4], n112[4], n113[4]);  // ../RTL/cmsdk_apb_slave_mux.v(211)
  or u1034 (n114[5], n112[5], n113[5]);  // ../RTL/cmsdk_apb_slave_mux.v(211)
  or u1035 (n114[6], n112[6], n113[6]);  // ../RTL/cmsdk_apb_slave_mux.v(211)
  or u1036 (n114[7], n112[7], n113[7]);  // ../RTL/cmsdk_apb_slave_mux.v(211)
  or u1037 (n114[8], n112[8], n113[8]);  // ../RTL/cmsdk_apb_slave_mux.v(211)
  or u1038 (n114[9], n112[9], n113[9]);  // ../RTL/cmsdk_apb_slave_mux.v(211)
  or u1039 (n114[10], n112[10], n113[10]);  // ../RTL/cmsdk_apb_slave_mux.v(211)
  and u104 (n83, PSEL2, PSLVERR2);  // ../RTL/cmsdk_apb_slave_mux.v(194)
  or u1040 (n114[11], n112[11], n113[11]);  // ../RTL/cmsdk_apb_slave_mux.v(211)
  or u1041 (n114[12], n112[12], n113[12]);  // ../RTL/cmsdk_apb_slave_mux.v(211)
  or u1042 (n114[13], n112[13], n113[13]);  // ../RTL/cmsdk_apb_slave_mux.v(211)
  or u1043 (n114[14], n112[14], n113[14]);  // ../RTL/cmsdk_apb_slave_mux.v(211)
  or u1044 (n114[15], n112[15], n113[15]);  // ../RTL/cmsdk_apb_slave_mux.v(211)
  or u1045 (n114[16], n112[16], n113[16]);  // ../RTL/cmsdk_apb_slave_mux.v(211)
  or u1046 (n114[17], n112[17], n113[17]);  // ../RTL/cmsdk_apb_slave_mux.v(211)
  or u1047 (n114[18], n112[18], n113[18]);  // ../RTL/cmsdk_apb_slave_mux.v(211)
  or u1048 (n114[19], n112[19], n113[19]);  // ../RTL/cmsdk_apb_slave_mux.v(211)
  or u1049 (n114[20], n112[20], n113[20]);  // ../RTL/cmsdk_apb_slave_mux.v(211)
  or u105 (n84, n82, n83);  // ../RTL/cmsdk_apb_slave_mux.v(194)
  or u1050 (n114[21], n112[21], n113[21]);  // ../RTL/cmsdk_apb_slave_mux.v(211)
  or u1051 (n114[22], n112[22], n113[22]);  // ../RTL/cmsdk_apb_slave_mux.v(211)
  or u1052 (n114[23], n112[23], n113[23]);  // ../RTL/cmsdk_apb_slave_mux.v(211)
  or u1053 (n114[24], n112[24], n113[24]);  // ../RTL/cmsdk_apb_slave_mux.v(211)
  or u1054 (n114[25], n112[25], n113[25]);  // ../RTL/cmsdk_apb_slave_mux.v(211)
  or u1055 (n114[26], n112[26], n113[26]);  // ../RTL/cmsdk_apb_slave_mux.v(211)
  or u1056 (n114[27], n112[27], n113[27]);  // ../RTL/cmsdk_apb_slave_mux.v(211)
  or u1057 (n114[28], n112[28], n113[28]);  // ../RTL/cmsdk_apb_slave_mux.v(211)
  or u1058 (n114[29], n112[29], n113[29]);  // ../RTL/cmsdk_apb_slave_mux.v(211)
  or u1059 (n114[30], n112[30], n113[30]);  // ../RTL/cmsdk_apb_slave_mux.v(211)
  and u106 (n85, PSEL3, PSLVERR3);  // ../RTL/cmsdk_apb_slave_mux.v(195)
  or u1060 (n114[31], n112[31], n113[31]);  // ../RTL/cmsdk_apb_slave_mux.v(211)
  and u1061 (n113[1], PSEL2, PRDATA2[1]);  // ../RTL/cmsdk_apb_slave_mux.v(211)
  and u1062 (n113[2], PSEL2, PRDATA2[2]);  // ../RTL/cmsdk_apb_slave_mux.v(211)
  and u1063 (n113[3], PSEL2, PRDATA2[3]);  // ../RTL/cmsdk_apb_slave_mux.v(211)
  and u1064 (n113[4], PSEL2, PRDATA2[4]);  // ../RTL/cmsdk_apb_slave_mux.v(211)
  and u1065 (n113[5], PSEL2, PRDATA2[5]);  // ../RTL/cmsdk_apb_slave_mux.v(211)
  and u1066 (n113[6], PSEL2, PRDATA2[6]);  // ../RTL/cmsdk_apb_slave_mux.v(211)
  and u1067 (n113[7], PSEL2, PRDATA2[7]);  // ../RTL/cmsdk_apb_slave_mux.v(211)
  and u1068 (n113[8], PSEL2, PRDATA2[8]);  // ../RTL/cmsdk_apb_slave_mux.v(211)
  and u1069 (n113[9], PSEL2, PRDATA2[9]);  // ../RTL/cmsdk_apb_slave_mux.v(211)
  or u107 (n86, n84, n85);  // ../RTL/cmsdk_apb_slave_mux.v(195)
  and u1070 (n113[10], PSEL2, PRDATA2[10]);  // ../RTL/cmsdk_apb_slave_mux.v(211)
  and u1071 (n113[11], PSEL2, PRDATA2[11]);  // ../RTL/cmsdk_apb_slave_mux.v(211)
  and u1072 (n113[12], PSEL2, PRDATA2[12]);  // ../RTL/cmsdk_apb_slave_mux.v(211)
  and u1073 (n113[13], PSEL2, PRDATA2[13]);  // ../RTL/cmsdk_apb_slave_mux.v(211)
  and u1074 (n113[14], PSEL2, PRDATA2[14]);  // ../RTL/cmsdk_apb_slave_mux.v(211)
  and u1075 (n113[15], PSEL2, PRDATA2[15]);  // ../RTL/cmsdk_apb_slave_mux.v(211)
  and u1076 (n113[16], PSEL2, PRDATA2[16]);  // ../RTL/cmsdk_apb_slave_mux.v(211)
  and u1077 (n113[17], PSEL2, PRDATA2[17]);  // ../RTL/cmsdk_apb_slave_mux.v(211)
  and u1078 (n113[18], PSEL2, PRDATA2[18]);  // ../RTL/cmsdk_apb_slave_mux.v(211)
  and u1079 (n113[19], PSEL2, PRDATA2[19]);  // ../RTL/cmsdk_apb_slave_mux.v(211)
  and u108 (n87, PSEL4, PSLVERR4);  // ../RTL/cmsdk_apb_slave_mux.v(196)
  and u1080 (n113[20], PSEL2, PRDATA2[20]);  // ../RTL/cmsdk_apb_slave_mux.v(211)
  and u1081 (n113[21], PSEL2, PRDATA2[21]);  // ../RTL/cmsdk_apb_slave_mux.v(211)
  and u1082 (n113[22], PSEL2, PRDATA2[22]);  // ../RTL/cmsdk_apb_slave_mux.v(211)
  and u1083 (n113[23], PSEL2, PRDATA2[23]);  // ../RTL/cmsdk_apb_slave_mux.v(211)
  and u1084 (n113[24], PSEL2, PRDATA2[24]);  // ../RTL/cmsdk_apb_slave_mux.v(211)
  and u1085 (n113[25], PSEL2, PRDATA2[25]);  // ../RTL/cmsdk_apb_slave_mux.v(211)
  and u1086 (n113[26], PSEL2, PRDATA2[26]);  // ../RTL/cmsdk_apb_slave_mux.v(211)
  and u1087 (n113[27], PSEL2, PRDATA2[27]);  // ../RTL/cmsdk_apb_slave_mux.v(211)
  and u1088 (n113[28], PSEL2, PRDATA2[28]);  // ../RTL/cmsdk_apb_slave_mux.v(211)
  and u1089 (n113[29], PSEL2, PRDATA2[29]);  // ../RTL/cmsdk_apb_slave_mux.v(211)
  or u109 (n88, n86, n87);  // ../RTL/cmsdk_apb_slave_mux.v(196)
  and u1090 (n113[30], PSEL2, PRDATA2[30]);  // ../RTL/cmsdk_apb_slave_mux.v(211)
  and u1091 (n113[31], PSEL2, PRDATA2[31]);  // ../RTL/cmsdk_apb_slave_mux.v(211)
  or u1092 (n112[1], n110[1], n111[1]);  // ../RTL/cmsdk_apb_slave_mux.v(210)
  or u1093 (n112[2], n110[2], n111[2]);  // ../RTL/cmsdk_apb_slave_mux.v(210)
  or u1094 (n112[3], n110[3], n111[3]);  // ../RTL/cmsdk_apb_slave_mux.v(210)
  or u1095 (n112[4], n110[4], n111[4]);  // ../RTL/cmsdk_apb_slave_mux.v(210)
  or u1096 (n112[5], n110[5], n111[5]);  // ../RTL/cmsdk_apb_slave_mux.v(210)
  or u1097 (n112[6], n110[6], n111[6]);  // ../RTL/cmsdk_apb_slave_mux.v(210)
  or u1098 (n112[7], n110[7], n111[7]);  // ../RTL/cmsdk_apb_slave_mux.v(210)
  or u1099 (n112[8], n110[8], n111[8]);  // ../RTL/cmsdk_apb_slave_mux.v(210)
  and u11 (PSEL3, n3, en[3]);  // ../RTL/cmsdk_apb_slave_mux.v(160)
  and u110 (n89, PSEL5, PSLVERR5);  // ../RTL/cmsdk_apb_slave_mux.v(197)
  or u1100 (n112[9], n110[9], n111[9]);  // ../RTL/cmsdk_apb_slave_mux.v(210)
  or u1101 (n112[10], n110[10], n111[10]);  // ../RTL/cmsdk_apb_slave_mux.v(210)
  or u1102 (n112[11], n110[11], n111[11]);  // ../RTL/cmsdk_apb_slave_mux.v(210)
  or u1103 (n112[12], n110[12], n111[12]);  // ../RTL/cmsdk_apb_slave_mux.v(210)
  or u1104 (n112[13], n110[13], n111[13]);  // ../RTL/cmsdk_apb_slave_mux.v(210)
  or u1105 (n112[14], n110[14], n111[14]);  // ../RTL/cmsdk_apb_slave_mux.v(210)
  or u1106 (n112[15], n110[15], n111[15]);  // ../RTL/cmsdk_apb_slave_mux.v(210)
  or u1107 (n112[16], n110[16], n111[16]);  // ../RTL/cmsdk_apb_slave_mux.v(210)
  or u1108 (n112[17], n110[17], n111[17]);  // ../RTL/cmsdk_apb_slave_mux.v(210)
  or u1109 (n112[18], n110[18], n111[18]);  // ../RTL/cmsdk_apb_slave_mux.v(210)
  or u111 (n90, n88, n89);  // ../RTL/cmsdk_apb_slave_mux.v(197)
  or u1110 (n112[19], n110[19], n111[19]);  // ../RTL/cmsdk_apb_slave_mux.v(210)
  or u1111 (n112[20], n110[20], n111[20]);  // ../RTL/cmsdk_apb_slave_mux.v(210)
  or u1112 (n112[21], n110[21], n111[21]);  // ../RTL/cmsdk_apb_slave_mux.v(210)
  or u1113 (n112[22], n110[22], n111[22]);  // ../RTL/cmsdk_apb_slave_mux.v(210)
  or u1114 (n112[23], n110[23], n111[23]);  // ../RTL/cmsdk_apb_slave_mux.v(210)
  or u1115 (n112[24], n110[24], n111[24]);  // ../RTL/cmsdk_apb_slave_mux.v(210)
  or u1116 (n112[25], n110[25], n111[25]);  // ../RTL/cmsdk_apb_slave_mux.v(210)
  or u1117 (n112[26], n110[26], n111[26]);  // ../RTL/cmsdk_apb_slave_mux.v(210)
  or u1118 (n112[27], n110[27], n111[27]);  // ../RTL/cmsdk_apb_slave_mux.v(210)
  or u1119 (n112[28], n110[28], n111[28]);  // ../RTL/cmsdk_apb_slave_mux.v(210)
  and u112 (n91, PSEL6, PSLVERR6);  // ../RTL/cmsdk_apb_slave_mux.v(198)
  or u1120 (n112[29], n110[29], n111[29]);  // ../RTL/cmsdk_apb_slave_mux.v(210)
  or u1121 (n112[30], n110[30], n111[30]);  // ../RTL/cmsdk_apb_slave_mux.v(210)
  or u1122 (n112[31], n110[31], n111[31]);  // ../RTL/cmsdk_apb_slave_mux.v(210)
  buf u1123 (en[1], 1'b0);  // ../RTL/cmsdk_apb_slave_mux.v(139)
  buf u1124 (en[2], 1'b0);  // ../RTL/cmsdk_apb_slave_mux.v(139)
  buf u1125 (en[3], 1'b0);  // ../RTL/cmsdk_apb_slave_mux.v(139)
  buf u1126 (en[4], 1'b1);  // ../RTL/cmsdk_apb_slave_mux.v(139)
  buf u1127 (en[5], 1'b0);  // ../RTL/cmsdk_apb_slave_mux.v(139)
  buf u1128 (en[6], 1'b0);  // ../RTL/cmsdk_apb_slave_mux.v(139)
  buf u1129 (en[7], 1'b0);  // ../RTL/cmsdk_apb_slave_mux.v(139)
  or u113 (n92, n90, n91);  // ../RTL/cmsdk_apb_slave_mux.v(198)
  buf u1130 (en[8], 1'b0);  // ../RTL/cmsdk_apb_slave_mux.v(139)
  buf u1131 (en[9], 1'b0);  // ../RTL/cmsdk_apb_slave_mux.v(139)
  buf u1132 (en[10], 1'b0);  // ../RTL/cmsdk_apb_slave_mux.v(139)
  buf u1133 (en[11], 1'b0);  // ../RTL/cmsdk_apb_slave_mux.v(139)
  buf u1134 (en[12], 1'b0);  // ../RTL/cmsdk_apb_slave_mux.v(139)
  buf u1135 (en[13], 1'b0);  // ../RTL/cmsdk_apb_slave_mux.v(139)
  buf u1136 (en[14], 1'b0);  // ../RTL/cmsdk_apb_slave_mux.v(139)
  buf u1137 (en[15], 1'b0);  // ../RTL/cmsdk_apb_slave_mux.v(139)
  and u114 (n93, PSEL7, PSLVERR7);  // ../RTL/cmsdk_apb_slave_mux.v(199)
  or u115 (n94, n92, n93);  // ../RTL/cmsdk_apb_slave_mux.v(199)
  and u116 (n95, PSEL8, PSLVERR8);  // ../RTL/cmsdk_apb_slave_mux.v(200)
  or u117 (n96, n94, n95);  // ../RTL/cmsdk_apb_slave_mux.v(200)
  and u118 (n97, PSEL9, PSLVERR9);  // ../RTL/cmsdk_apb_slave_mux.v(201)
  or u119 (n98, n96, n97);  // ../RTL/cmsdk_apb_slave_mux.v(201)
  and u12 (n4, PSEL, dec[4]);  // ../RTL/cmsdk_apb_slave_mux.v(161)
  and u120 (n99, PSEL10, PSLVERR10);  // ../RTL/cmsdk_apb_slave_mux.v(202)
  or u121 (n100, n98, n99);  // ../RTL/cmsdk_apb_slave_mux.v(202)
  and u122 (n101, PSEL11, PSLVERR11);  // ../RTL/cmsdk_apb_slave_mux.v(203)
  or u123 (n102, n100, n101);  // ../RTL/cmsdk_apb_slave_mux.v(203)
  and u124 (n103, PSEL12, PSLVERR12);  // ../RTL/cmsdk_apb_slave_mux.v(204)
  or u125 (n104, n102, n103);  // ../RTL/cmsdk_apb_slave_mux.v(204)
  and u126 (n105, PSEL13, PSLVERR13);  // ../RTL/cmsdk_apb_slave_mux.v(205)
  or u127 (n106, n104, n105);  // ../RTL/cmsdk_apb_slave_mux.v(205)
  and u128 (n107, PSEL14, PSLVERR14);  // ../RTL/cmsdk_apb_slave_mux.v(206)
  or u129 (n108, n106, n107);  // ../RTL/cmsdk_apb_slave_mux.v(206)
  and u13 (PSEL4, n4, en[4]);  // ../RTL/cmsdk_apb_slave_mux.v(161)
  and u130 (n109, PSEL15, PSLVERR15);  // ../RTL/cmsdk_apb_slave_mux.v(207)
  or u131 (PSLVERR, n108, n109);  // ../RTL/cmsdk_apb_slave_mux.v(207)
  and u132 (n111[2], PSEL1, PRDATA1[2]);  // ../RTL/cmsdk_apb_slave_mux.v(209)
  and u133 (n111[3], PSEL1, PRDATA1[3]);  // ../RTL/cmsdk_apb_slave_mux.v(209)
  buf u134 (en[0], 1'b1);  // ../RTL/cmsdk_apb_slave_mux.v(139)
  or u135 (n112[0], n110[0], n111[0]);  // ../RTL/cmsdk_apb_slave_mux.v(210)
  and u136 (n113[0], PSEL2, PRDATA2[0]);  // ../RTL/cmsdk_apb_slave_mux.v(211)
  or u137 (n114[0], n112[0], n113[0]);  // ../RTL/cmsdk_apb_slave_mux.v(211)
  and u138 (n115[0], PSEL3, PRDATA3[0]);  // ../RTL/cmsdk_apb_slave_mux.v(212)
  or u139 (n116[0], n114[0], n115[0]);  // ../RTL/cmsdk_apb_slave_mux.v(212)
  and u14 (n5, PSEL, dec[5]);  // ../RTL/cmsdk_apb_slave_mux.v(162)
  and u140 (n117[0], PSEL4, PRDATA4[0]);  // ../RTL/cmsdk_apb_slave_mux.v(213)
  or u141 (n118[0], n116[0], n117[0]);  // ../RTL/cmsdk_apb_slave_mux.v(213)
  and u142 (n119[0], PSEL5, PRDATA5[0]);  // ../RTL/cmsdk_apb_slave_mux.v(214)
  or u143 (n120[0], n118[0], n119[0]);  // ../RTL/cmsdk_apb_slave_mux.v(214)
  and u144 (n121[0], PSEL6, PRDATA6[0]);  // ../RTL/cmsdk_apb_slave_mux.v(215)
  or u145 (n122[0], n120[0], n121[0]);  // ../RTL/cmsdk_apb_slave_mux.v(215)
  and u146 (n123[0], PSEL7, PRDATA7[0]);  // ../RTL/cmsdk_apb_slave_mux.v(216)
  or u147 (n124[0], n122[0], n123[0]);  // ../RTL/cmsdk_apb_slave_mux.v(216)
  and u148 (n125[0], PSEL8, PRDATA8[0]);  // ../RTL/cmsdk_apb_slave_mux.v(217)
  or u149 (n126[0], n124[0], n125[0]);  // ../RTL/cmsdk_apb_slave_mux.v(217)
  and u15 (PSEL5, n5, en[5]);  // ../RTL/cmsdk_apb_slave_mux.v(162)
  and u150 (n127[0], PSEL9, PRDATA9[0]);  // ../RTL/cmsdk_apb_slave_mux.v(218)
  or u151 (n128[0], n126[0], n127[0]);  // ../RTL/cmsdk_apb_slave_mux.v(218)
  and u152 (n129[0], PSEL10, PRDATA10[0]);  // ../RTL/cmsdk_apb_slave_mux.v(219)
  or u153 (n130[0], n128[0], n129[0]);  // ../RTL/cmsdk_apb_slave_mux.v(219)
  and u154 (n131[0], PSEL11, PRDATA11[0]);  // ../RTL/cmsdk_apb_slave_mux.v(220)
  or u155 (n132[0], n130[0], n131[0]);  // ../RTL/cmsdk_apb_slave_mux.v(220)
  and u156 (n133[0], PSEL12, PRDATA12[0]);  // ../RTL/cmsdk_apb_slave_mux.v(221)
  or u157 (n134[0], n132[0], n133[0]);  // ../RTL/cmsdk_apb_slave_mux.v(221)
  and u158 (n135[0], PSEL13, PRDATA13[0]);  // ../RTL/cmsdk_apb_slave_mux.v(222)
  or u159 (n136[0], n134[0], n135[0]);  // ../RTL/cmsdk_apb_slave_mux.v(222)
  and u16 (n6, PSEL, dec[6]);  // ../RTL/cmsdk_apb_slave_mux.v(163)
  and u160 (n137[0], PSEL14, PRDATA14[0]);  // ../RTL/cmsdk_apb_slave_mux.v(223)
  or u161 (n138[0], n136[0], n137[0]);  // ../RTL/cmsdk_apb_slave_mux.v(223)
  and u162 (n139[0], PSEL15, PRDATA15[0]);  // ../RTL/cmsdk_apb_slave_mux.v(224)
  or u163 (PRDATA[0], n138[0], n139[0]);  // ../RTL/cmsdk_apb_slave_mux.v(224)
  and u164 (n111[4], PSEL1, PRDATA1[4]);  // ../RTL/cmsdk_apb_slave_mux.v(209)
  and u165 (n111[5], PSEL1, PRDATA1[5]);  // ../RTL/cmsdk_apb_slave_mux.v(209)
  and u166 (n111[6], PSEL1, PRDATA1[6]);  // ../RTL/cmsdk_apb_slave_mux.v(209)
  and u167 (n111[7], PSEL1, PRDATA1[7]);  // ../RTL/cmsdk_apb_slave_mux.v(209)
  and u168 (n111[8], PSEL1, PRDATA1[8]);  // ../RTL/cmsdk_apb_slave_mux.v(209)
  and u169 (n111[9], PSEL1, PRDATA1[9]);  // ../RTL/cmsdk_apb_slave_mux.v(209)
  and u17 (PSEL6, n6, en[6]);  // ../RTL/cmsdk_apb_slave_mux.v(163)
  and u170 (n111[10], PSEL1, PRDATA1[10]);  // ../RTL/cmsdk_apb_slave_mux.v(209)
  and u171 (n111[11], PSEL1, PRDATA1[11]);  // ../RTL/cmsdk_apb_slave_mux.v(209)
  and u172 (n111[12], PSEL1, PRDATA1[12]);  // ../RTL/cmsdk_apb_slave_mux.v(209)
  and u173 (n111[13], PSEL1, PRDATA1[13]);  // ../RTL/cmsdk_apb_slave_mux.v(209)
  and u174 (n111[14], PSEL1, PRDATA1[14]);  // ../RTL/cmsdk_apb_slave_mux.v(209)
  and u175 (n111[15], PSEL1, PRDATA1[15]);  // ../RTL/cmsdk_apb_slave_mux.v(209)
  and u176 (n111[16], PSEL1, PRDATA1[16]);  // ../RTL/cmsdk_apb_slave_mux.v(209)
  and u177 (n111[17], PSEL1, PRDATA1[17]);  // ../RTL/cmsdk_apb_slave_mux.v(209)
  and u178 (n111[18], PSEL1, PRDATA1[18]);  // ../RTL/cmsdk_apb_slave_mux.v(209)
  and u179 (n111[19], PSEL1, PRDATA1[19]);  // ../RTL/cmsdk_apb_slave_mux.v(209)
  and u18 (n7, PSEL, dec[7]);  // ../RTL/cmsdk_apb_slave_mux.v(164)
  and u180 (n111[20], PSEL1, PRDATA1[20]);  // ../RTL/cmsdk_apb_slave_mux.v(209)
  and u181 (n111[21], PSEL1, PRDATA1[21]);  // ../RTL/cmsdk_apb_slave_mux.v(209)
  and u182 (n111[22], PSEL1, PRDATA1[22]);  // ../RTL/cmsdk_apb_slave_mux.v(209)
  and u183 (n111[23], PSEL1, PRDATA1[23]);  // ../RTL/cmsdk_apb_slave_mux.v(209)
  and u184 (n111[24], PSEL1, PRDATA1[24]);  // ../RTL/cmsdk_apb_slave_mux.v(209)
  and u185 (n111[25], PSEL1, PRDATA1[25]);  // ../RTL/cmsdk_apb_slave_mux.v(209)
  and u186 (n111[26], PSEL1, PRDATA1[26]);  // ../RTL/cmsdk_apb_slave_mux.v(209)
  and u187 (n111[27], PSEL1, PRDATA1[27]);  // ../RTL/cmsdk_apb_slave_mux.v(209)
  and u188 (n111[28], PSEL1, PRDATA1[28]);  // ../RTL/cmsdk_apb_slave_mux.v(209)
  and u189 (n111[29], PSEL1, PRDATA1[29]);  // ../RTL/cmsdk_apb_slave_mux.v(209)
  and u19 (PSEL7, n7, en[7]);  // ../RTL/cmsdk_apb_slave_mux.v(164)
  and u190 (n111[30], PSEL1, PRDATA1[30]);  // ../RTL/cmsdk_apb_slave_mux.v(209)
  and u191 (n111[31], PSEL1, PRDATA1[31]);  // ../RTL/cmsdk_apb_slave_mux.v(209)
  and u192 (n110[0], PSEL0, PRDATA0[0]);  // ../RTL/cmsdk_apb_slave_mux.v(209)
  and u193 (n110[1], PSEL0, PRDATA0[1]);  // ../RTL/cmsdk_apb_slave_mux.v(209)
  and u194 (n110[2], PSEL0, PRDATA0[2]);  // ../RTL/cmsdk_apb_slave_mux.v(209)
  and u195 (n110[3], PSEL0, PRDATA0[3]);  // ../RTL/cmsdk_apb_slave_mux.v(209)
  and u196 (n110[4], PSEL0, PRDATA0[4]);  // ../RTL/cmsdk_apb_slave_mux.v(209)
  and u197 (n110[5], PSEL0, PRDATA0[5]);  // ../RTL/cmsdk_apb_slave_mux.v(209)
  and u198 (n110[6], PSEL0, PRDATA0[6]);  // ../RTL/cmsdk_apb_slave_mux.v(209)
  and u199 (n110[7], PSEL0, PRDATA0[7]);  // ../RTL/cmsdk_apb_slave_mux.v(209)
  and u2 (n111[1], PSEL1, PRDATA1[1]);  // ../RTL/cmsdk_apb_slave_mux.v(209)
  and u20 (n8, PSEL, dec[8]);  // ../RTL/cmsdk_apb_slave_mux.v(165)
  and u200 (n110[8], PSEL0, PRDATA0[8]);  // ../RTL/cmsdk_apb_slave_mux.v(209)
  and u201 (n110[9], PSEL0, PRDATA0[9]);  // ../RTL/cmsdk_apb_slave_mux.v(209)
  and u202 (n110[10], PSEL0, PRDATA0[10]);  // ../RTL/cmsdk_apb_slave_mux.v(209)
  and u203 (n110[11], PSEL0, PRDATA0[11]);  // ../RTL/cmsdk_apb_slave_mux.v(209)
  and u204 (n110[12], PSEL0, PRDATA0[12]);  // ../RTL/cmsdk_apb_slave_mux.v(209)
  and u205 (n110[13], PSEL0, PRDATA0[13]);  // ../RTL/cmsdk_apb_slave_mux.v(209)
  and u206 (n110[14], PSEL0, PRDATA0[14]);  // ../RTL/cmsdk_apb_slave_mux.v(209)
  and u207 (n110[15], PSEL0, PRDATA0[15]);  // ../RTL/cmsdk_apb_slave_mux.v(209)
  and u208 (n110[16], PSEL0, PRDATA0[16]);  // ../RTL/cmsdk_apb_slave_mux.v(209)
  and u209 (n110[17], PSEL0, PRDATA0[17]);  // ../RTL/cmsdk_apb_slave_mux.v(209)
  and u21 (PSEL8, n8, en[8]);  // ../RTL/cmsdk_apb_slave_mux.v(165)
  and u210 (n110[18], PSEL0, PRDATA0[18]);  // ../RTL/cmsdk_apb_slave_mux.v(209)
  and u211 (n110[19], PSEL0, PRDATA0[19]);  // ../RTL/cmsdk_apb_slave_mux.v(209)
  and u212 (n110[20], PSEL0, PRDATA0[20]);  // ../RTL/cmsdk_apb_slave_mux.v(209)
  and u213 (n110[21], PSEL0, PRDATA0[21]);  // ../RTL/cmsdk_apb_slave_mux.v(209)
  and u214 (n110[22], PSEL0, PRDATA0[22]);  // ../RTL/cmsdk_apb_slave_mux.v(209)
  and u215 (n110[23], PSEL0, PRDATA0[23]);  // ../RTL/cmsdk_apb_slave_mux.v(209)
  and u216 (n110[24], PSEL0, PRDATA0[24]);  // ../RTL/cmsdk_apb_slave_mux.v(209)
  and u217 (n110[25], PSEL0, PRDATA0[25]);  // ../RTL/cmsdk_apb_slave_mux.v(209)
  and u218 (n110[26], PSEL0, PRDATA0[26]);  // ../RTL/cmsdk_apb_slave_mux.v(209)
  and u219 (n110[27], PSEL0, PRDATA0[27]);  // ../RTL/cmsdk_apb_slave_mux.v(209)
  and u22 (n9, PSEL, dec[9]);  // ../RTL/cmsdk_apb_slave_mux.v(166)
  and u220 (n110[28], PSEL0, PRDATA0[28]);  // ../RTL/cmsdk_apb_slave_mux.v(209)
  and u221 (n110[29], PSEL0, PRDATA0[29]);  // ../RTL/cmsdk_apb_slave_mux.v(209)
  and u222 (n110[30], PSEL0, PRDATA0[30]);  // ../RTL/cmsdk_apb_slave_mux.v(209)
  and u223 (n110[31], PSEL0, PRDATA0[31]);  // ../RTL/cmsdk_apb_slave_mux.v(209)
  or u224 (PRDATA[1], n138[1], n139[1]);  // ../RTL/cmsdk_apb_slave_mux.v(224)
  or u225 (PRDATA[2], n138[2], n139[2]);  // ../RTL/cmsdk_apb_slave_mux.v(224)
  or u226 (PRDATA[3], n138[3], n139[3]);  // ../RTL/cmsdk_apb_slave_mux.v(224)
  or u227 (PRDATA[4], n138[4], n139[4]);  // ../RTL/cmsdk_apb_slave_mux.v(224)
  or u228 (PRDATA[5], n138[5], n139[5]);  // ../RTL/cmsdk_apb_slave_mux.v(224)
  or u229 (PRDATA[6], n138[6], n139[6]);  // ../RTL/cmsdk_apb_slave_mux.v(224)
  and u23 (PSEL9, n9, en[9]);  // ../RTL/cmsdk_apb_slave_mux.v(166)
  or u230 (PRDATA[7], n138[7], n139[7]);  // ../RTL/cmsdk_apb_slave_mux.v(224)
  or u231 (PRDATA[8], n138[8], n139[8]);  // ../RTL/cmsdk_apb_slave_mux.v(224)
  or u232 (PRDATA[9], n138[9], n139[9]);  // ../RTL/cmsdk_apb_slave_mux.v(224)
  or u233 (PRDATA[10], n138[10], n139[10]);  // ../RTL/cmsdk_apb_slave_mux.v(224)
  or u234 (PRDATA[11], n138[11], n139[11]);  // ../RTL/cmsdk_apb_slave_mux.v(224)
  or u235 (PRDATA[12], n138[12], n139[12]);  // ../RTL/cmsdk_apb_slave_mux.v(224)
  or u236 (PRDATA[13], n138[13], n139[13]);  // ../RTL/cmsdk_apb_slave_mux.v(224)
  or u237 (PRDATA[14], n138[14], n139[14]);  // ../RTL/cmsdk_apb_slave_mux.v(224)
  or u238 (PRDATA[15], n138[15], n139[15]);  // ../RTL/cmsdk_apb_slave_mux.v(224)
  or u239 (PRDATA[16], n138[16], n139[16]);  // ../RTL/cmsdk_apb_slave_mux.v(224)
  and u24 (n10, PSEL, dec[10]);  // ../RTL/cmsdk_apb_slave_mux.v(167)
  or u240 (PRDATA[17], n138[17], n139[17]);  // ../RTL/cmsdk_apb_slave_mux.v(224)
  or u241 (PRDATA[18], n138[18], n139[18]);  // ../RTL/cmsdk_apb_slave_mux.v(224)
  or u242 (PRDATA[19], n138[19], n139[19]);  // ../RTL/cmsdk_apb_slave_mux.v(224)
  or u243 (PRDATA[20], n138[20], n139[20]);  // ../RTL/cmsdk_apb_slave_mux.v(224)
  or u244 (PRDATA[21], n138[21], n139[21]);  // ../RTL/cmsdk_apb_slave_mux.v(224)
  or u245 (PRDATA[22], n138[22], n139[22]);  // ../RTL/cmsdk_apb_slave_mux.v(224)
  or u246 (PRDATA[23], n138[23], n139[23]);  // ../RTL/cmsdk_apb_slave_mux.v(224)
  or u247 (PRDATA[24], n138[24], n139[24]);  // ../RTL/cmsdk_apb_slave_mux.v(224)
  or u248 (PRDATA[25], n138[25], n139[25]);  // ../RTL/cmsdk_apb_slave_mux.v(224)
  or u249 (PRDATA[26], n138[26], n139[26]);  // ../RTL/cmsdk_apb_slave_mux.v(224)
  and u25 (PSEL10, n10, en[10]);  // ../RTL/cmsdk_apb_slave_mux.v(167)
  or u250 (PRDATA[27], n138[27], n139[27]);  // ../RTL/cmsdk_apb_slave_mux.v(224)
  or u251 (PRDATA[28], n138[28], n139[28]);  // ../RTL/cmsdk_apb_slave_mux.v(224)
  or u252 (PRDATA[29], n138[29], n139[29]);  // ../RTL/cmsdk_apb_slave_mux.v(224)
  or u253 (PRDATA[30], n138[30], n139[30]);  // ../RTL/cmsdk_apb_slave_mux.v(224)
  or u254 (PRDATA[31], n138[31], n139[31]);  // ../RTL/cmsdk_apb_slave_mux.v(224)
  and u255 (n139[1], PSEL15, PRDATA15[1]);  // ../RTL/cmsdk_apb_slave_mux.v(224)
  and u256 (n139[2], PSEL15, PRDATA15[2]);  // ../RTL/cmsdk_apb_slave_mux.v(224)
  and u257 (n139[3], PSEL15, PRDATA15[3]);  // ../RTL/cmsdk_apb_slave_mux.v(224)
  and u258 (n139[4], PSEL15, PRDATA15[4]);  // ../RTL/cmsdk_apb_slave_mux.v(224)
  and u259 (n139[5], PSEL15, PRDATA15[5]);  // ../RTL/cmsdk_apb_slave_mux.v(224)
  and u26 (n11, PSEL, dec[11]);  // ../RTL/cmsdk_apb_slave_mux.v(168)
  and u260 (n139[6], PSEL15, PRDATA15[6]);  // ../RTL/cmsdk_apb_slave_mux.v(224)
  and u261 (n139[7], PSEL15, PRDATA15[7]);  // ../RTL/cmsdk_apb_slave_mux.v(224)
  and u262 (n139[8], PSEL15, PRDATA15[8]);  // ../RTL/cmsdk_apb_slave_mux.v(224)
  and u263 (n139[9], PSEL15, PRDATA15[9]);  // ../RTL/cmsdk_apb_slave_mux.v(224)
  and u264 (n139[10], PSEL15, PRDATA15[10]);  // ../RTL/cmsdk_apb_slave_mux.v(224)
  and u265 (n139[11], PSEL15, PRDATA15[11]);  // ../RTL/cmsdk_apb_slave_mux.v(224)
  and u266 (n139[12], PSEL15, PRDATA15[12]);  // ../RTL/cmsdk_apb_slave_mux.v(224)
  and u267 (n139[13], PSEL15, PRDATA15[13]);  // ../RTL/cmsdk_apb_slave_mux.v(224)
  and u268 (n139[14], PSEL15, PRDATA15[14]);  // ../RTL/cmsdk_apb_slave_mux.v(224)
  and u269 (n139[15], PSEL15, PRDATA15[15]);  // ../RTL/cmsdk_apb_slave_mux.v(224)
  and u27 (PSEL11, n11, en[11]);  // ../RTL/cmsdk_apb_slave_mux.v(168)
  and u270 (n139[16], PSEL15, PRDATA15[16]);  // ../RTL/cmsdk_apb_slave_mux.v(224)
  and u271 (n139[17], PSEL15, PRDATA15[17]);  // ../RTL/cmsdk_apb_slave_mux.v(224)
  and u272 (n139[18], PSEL15, PRDATA15[18]);  // ../RTL/cmsdk_apb_slave_mux.v(224)
  and u273 (n139[19], PSEL15, PRDATA15[19]);  // ../RTL/cmsdk_apb_slave_mux.v(224)
  and u274 (n139[20], PSEL15, PRDATA15[20]);  // ../RTL/cmsdk_apb_slave_mux.v(224)
  and u275 (n139[21], PSEL15, PRDATA15[21]);  // ../RTL/cmsdk_apb_slave_mux.v(224)
  and u276 (n139[22], PSEL15, PRDATA15[22]);  // ../RTL/cmsdk_apb_slave_mux.v(224)
  and u277 (n139[23], PSEL15, PRDATA15[23]);  // ../RTL/cmsdk_apb_slave_mux.v(224)
  and u278 (n139[24], PSEL15, PRDATA15[24]);  // ../RTL/cmsdk_apb_slave_mux.v(224)
  and u279 (n139[25], PSEL15, PRDATA15[25]);  // ../RTL/cmsdk_apb_slave_mux.v(224)
  and u28 (n12, PSEL, dec[12]);  // ../RTL/cmsdk_apb_slave_mux.v(169)
  and u280 (n139[26], PSEL15, PRDATA15[26]);  // ../RTL/cmsdk_apb_slave_mux.v(224)
  and u281 (n139[27], PSEL15, PRDATA15[27]);  // ../RTL/cmsdk_apb_slave_mux.v(224)
  and u282 (n139[28], PSEL15, PRDATA15[28]);  // ../RTL/cmsdk_apb_slave_mux.v(224)
  and u283 (n139[29], PSEL15, PRDATA15[29]);  // ../RTL/cmsdk_apb_slave_mux.v(224)
  and u284 (n139[30], PSEL15, PRDATA15[30]);  // ../RTL/cmsdk_apb_slave_mux.v(224)
  and u285 (n139[31], PSEL15, PRDATA15[31]);  // ../RTL/cmsdk_apb_slave_mux.v(224)
  or u286 (n138[1], n136[1], n137[1]);  // ../RTL/cmsdk_apb_slave_mux.v(223)
  or u287 (n138[2], n136[2], n137[2]);  // ../RTL/cmsdk_apb_slave_mux.v(223)
  or u288 (n138[3], n136[3], n137[3]);  // ../RTL/cmsdk_apb_slave_mux.v(223)
  or u289 (n138[4], n136[4], n137[4]);  // ../RTL/cmsdk_apb_slave_mux.v(223)
  and u29 (PSEL12, n12, en[12]);  // ../RTL/cmsdk_apb_slave_mux.v(169)
  or u290 (n138[5], n136[5], n137[5]);  // ../RTL/cmsdk_apb_slave_mux.v(223)
  or u291 (n138[6], n136[6], n137[6]);  // ../RTL/cmsdk_apb_slave_mux.v(223)
  or u292 (n138[7], n136[7], n137[7]);  // ../RTL/cmsdk_apb_slave_mux.v(223)
  or u293 (n138[8], n136[8], n137[8]);  // ../RTL/cmsdk_apb_slave_mux.v(223)
  or u294 (n138[9], n136[9], n137[9]);  // ../RTL/cmsdk_apb_slave_mux.v(223)
  or u295 (n138[10], n136[10], n137[10]);  // ../RTL/cmsdk_apb_slave_mux.v(223)
  or u296 (n138[11], n136[11], n137[11]);  // ../RTL/cmsdk_apb_slave_mux.v(223)
  or u297 (n138[12], n136[12], n137[12]);  // ../RTL/cmsdk_apb_slave_mux.v(223)
  or u298 (n138[13], n136[13], n137[13]);  // ../RTL/cmsdk_apb_slave_mux.v(223)
  or u299 (n138[14], n136[14], n137[14]);  // ../RTL/cmsdk_apb_slave_mux.v(223)
  and u3 (n111[0], PSEL1, PRDATA1[0]);  // ../RTL/cmsdk_apb_slave_mux.v(209)
  and u30 (n13, PSEL, dec[13]);  // ../RTL/cmsdk_apb_slave_mux.v(170)
  or u300 (n138[15], n136[15], n137[15]);  // ../RTL/cmsdk_apb_slave_mux.v(223)
  or u301 (n138[16], n136[16], n137[16]);  // ../RTL/cmsdk_apb_slave_mux.v(223)
  or u302 (n138[17], n136[17], n137[17]);  // ../RTL/cmsdk_apb_slave_mux.v(223)
  or u303 (n138[18], n136[18], n137[18]);  // ../RTL/cmsdk_apb_slave_mux.v(223)
  or u304 (n138[19], n136[19], n137[19]);  // ../RTL/cmsdk_apb_slave_mux.v(223)
  or u305 (n138[20], n136[20], n137[20]);  // ../RTL/cmsdk_apb_slave_mux.v(223)
  or u306 (n138[21], n136[21], n137[21]);  // ../RTL/cmsdk_apb_slave_mux.v(223)
  or u307 (n138[22], n136[22], n137[22]);  // ../RTL/cmsdk_apb_slave_mux.v(223)
  or u308 (n138[23], n136[23], n137[23]);  // ../RTL/cmsdk_apb_slave_mux.v(223)
  or u309 (n138[24], n136[24], n137[24]);  // ../RTL/cmsdk_apb_slave_mux.v(223)
  and u31 (PSEL13, n13, en[13]);  // ../RTL/cmsdk_apb_slave_mux.v(170)
  or u310 (n138[25], n136[25], n137[25]);  // ../RTL/cmsdk_apb_slave_mux.v(223)
  or u311 (n138[26], n136[26], n137[26]);  // ../RTL/cmsdk_apb_slave_mux.v(223)
  or u312 (n138[27], n136[27], n137[27]);  // ../RTL/cmsdk_apb_slave_mux.v(223)
  or u313 (n138[28], n136[28], n137[28]);  // ../RTL/cmsdk_apb_slave_mux.v(223)
  or u314 (n138[29], n136[29], n137[29]);  // ../RTL/cmsdk_apb_slave_mux.v(223)
  or u315 (n138[30], n136[30], n137[30]);  // ../RTL/cmsdk_apb_slave_mux.v(223)
  or u316 (n138[31], n136[31], n137[31]);  // ../RTL/cmsdk_apb_slave_mux.v(223)
  and u317 (n137[1], PSEL14, PRDATA14[1]);  // ../RTL/cmsdk_apb_slave_mux.v(223)
  and u318 (n137[2], PSEL14, PRDATA14[2]);  // ../RTL/cmsdk_apb_slave_mux.v(223)
  and u319 (n137[3], PSEL14, PRDATA14[3]);  // ../RTL/cmsdk_apb_slave_mux.v(223)
  and u32 (n14, PSEL, dec[14]);  // ../RTL/cmsdk_apb_slave_mux.v(171)
  and u320 (n137[4], PSEL14, PRDATA14[4]);  // ../RTL/cmsdk_apb_slave_mux.v(223)
  and u321 (n137[5], PSEL14, PRDATA14[5]);  // ../RTL/cmsdk_apb_slave_mux.v(223)
  and u322 (n137[6], PSEL14, PRDATA14[6]);  // ../RTL/cmsdk_apb_slave_mux.v(223)
  and u323 (n137[7], PSEL14, PRDATA14[7]);  // ../RTL/cmsdk_apb_slave_mux.v(223)
  and u324 (n137[8], PSEL14, PRDATA14[8]);  // ../RTL/cmsdk_apb_slave_mux.v(223)
  and u325 (n137[9], PSEL14, PRDATA14[9]);  // ../RTL/cmsdk_apb_slave_mux.v(223)
  and u326 (n137[10], PSEL14, PRDATA14[10]);  // ../RTL/cmsdk_apb_slave_mux.v(223)
  and u327 (n137[11], PSEL14, PRDATA14[11]);  // ../RTL/cmsdk_apb_slave_mux.v(223)
  and u328 (n137[12], PSEL14, PRDATA14[12]);  // ../RTL/cmsdk_apb_slave_mux.v(223)
  and u329 (n137[13], PSEL14, PRDATA14[13]);  // ../RTL/cmsdk_apb_slave_mux.v(223)
  and u33 (PSEL14, n14, en[14]);  // ../RTL/cmsdk_apb_slave_mux.v(171)
  and u330 (n137[14], PSEL14, PRDATA14[14]);  // ../RTL/cmsdk_apb_slave_mux.v(223)
  and u331 (n137[15], PSEL14, PRDATA14[15]);  // ../RTL/cmsdk_apb_slave_mux.v(223)
  and u332 (n137[16], PSEL14, PRDATA14[16]);  // ../RTL/cmsdk_apb_slave_mux.v(223)
  and u333 (n137[17], PSEL14, PRDATA14[17]);  // ../RTL/cmsdk_apb_slave_mux.v(223)
  and u334 (n137[18], PSEL14, PRDATA14[18]);  // ../RTL/cmsdk_apb_slave_mux.v(223)
  and u335 (n137[19], PSEL14, PRDATA14[19]);  // ../RTL/cmsdk_apb_slave_mux.v(223)
  and u336 (n137[20], PSEL14, PRDATA14[20]);  // ../RTL/cmsdk_apb_slave_mux.v(223)
  and u337 (n137[21], PSEL14, PRDATA14[21]);  // ../RTL/cmsdk_apb_slave_mux.v(223)
  and u338 (n137[22], PSEL14, PRDATA14[22]);  // ../RTL/cmsdk_apb_slave_mux.v(223)
  and u339 (n137[23], PSEL14, PRDATA14[23]);  // ../RTL/cmsdk_apb_slave_mux.v(223)
  and u34 (n15, PSEL, dec[15]);  // ../RTL/cmsdk_apb_slave_mux.v(172)
  and u340 (n137[24], PSEL14, PRDATA14[24]);  // ../RTL/cmsdk_apb_slave_mux.v(223)
  and u341 (n137[25], PSEL14, PRDATA14[25]);  // ../RTL/cmsdk_apb_slave_mux.v(223)
  and u342 (n137[26], PSEL14, PRDATA14[26]);  // ../RTL/cmsdk_apb_slave_mux.v(223)
  and u343 (n137[27], PSEL14, PRDATA14[27]);  // ../RTL/cmsdk_apb_slave_mux.v(223)
  and u344 (n137[28], PSEL14, PRDATA14[28]);  // ../RTL/cmsdk_apb_slave_mux.v(223)
  and u345 (n137[29], PSEL14, PRDATA14[29]);  // ../RTL/cmsdk_apb_slave_mux.v(223)
  and u346 (n137[30], PSEL14, PRDATA14[30]);  // ../RTL/cmsdk_apb_slave_mux.v(223)
  and u347 (n137[31], PSEL14, PRDATA14[31]);  // ../RTL/cmsdk_apb_slave_mux.v(223)
  or u348 (n136[1], n134[1], n135[1]);  // ../RTL/cmsdk_apb_slave_mux.v(222)
  or u349 (n136[2], n134[2], n135[2]);  // ../RTL/cmsdk_apb_slave_mux.v(222)
  and u35 (PSEL15, n15, en[15]);  // ../RTL/cmsdk_apb_slave_mux.v(172)
  or u350 (n136[3], n134[3], n135[3]);  // ../RTL/cmsdk_apb_slave_mux.v(222)
  or u351 (n136[4], n134[4], n135[4]);  // ../RTL/cmsdk_apb_slave_mux.v(222)
  or u352 (n136[5], n134[5], n135[5]);  // ../RTL/cmsdk_apb_slave_mux.v(222)
  or u353 (n136[6], n134[6], n135[6]);  // ../RTL/cmsdk_apb_slave_mux.v(222)
  or u354 (n136[7], n134[7], n135[7]);  // ../RTL/cmsdk_apb_slave_mux.v(222)
  or u355 (n136[8], n134[8], n135[8]);  // ../RTL/cmsdk_apb_slave_mux.v(222)
  or u356 (n136[9], n134[9], n135[9]);  // ../RTL/cmsdk_apb_slave_mux.v(222)
  or u357 (n136[10], n134[10], n135[10]);  // ../RTL/cmsdk_apb_slave_mux.v(222)
  or u358 (n136[11], n134[11], n135[11]);  // ../RTL/cmsdk_apb_slave_mux.v(222)
  or u359 (n136[12], n134[12], n135[12]);  // ../RTL/cmsdk_apb_slave_mux.v(222)
  not u36 (n16, PSEL);  // ../RTL/cmsdk_apb_slave_mux.v(174)
  or u360 (n136[13], n134[13], n135[13]);  // ../RTL/cmsdk_apb_slave_mux.v(222)
  or u361 (n136[14], n134[14], n135[14]);  // ../RTL/cmsdk_apb_slave_mux.v(222)
  or u362 (n136[15], n134[15], n135[15]);  // ../RTL/cmsdk_apb_slave_mux.v(222)
  or u363 (n136[16], n134[16], n135[16]);  // ../RTL/cmsdk_apb_slave_mux.v(222)
  or u364 (n136[17], n134[17], n135[17]);  // ../RTL/cmsdk_apb_slave_mux.v(222)
  or u365 (n136[18], n134[18], n135[18]);  // ../RTL/cmsdk_apb_slave_mux.v(222)
  or u366 (n136[19], n134[19], n135[19]);  // ../RTL/cmsdk_apb_slave_mux.v(222)
  or u367 (n136[20], n134[20], n135[20]);  // ../RTL/cmsdk_apb_slave_mux.v(222)
  or u368 (n136[21], n134[21], n135[21]);  // ../RTL/cmsdk_apb_slave_mux.v(222)
  or u369 (n136[22], n134[22], n135[22]);  // ../RTL/cmsdk_apb_slave_mux.v(222)
  not u37 (n17, en[0]);  // ../RTL/cmsdk_apb_slave_mux.v(175)
  or u370 (n136[23], n134[23], n135[23]);  // ../RTL/cmsdk_apb_slave_mux.v(222)
  or u371 (n136[24], n134[24], n135[24]);  // ../RTL/cmsdk_apb_slave_mux.v(222)
  or u372 (n136[25], n134[25], n135[25]);  // ../RTL/cmsdk_apb_slave_mux.v(222)
  or u373 (n136[26], n134[26], n135[26]);  // ../RTL/cmsdk_apb_slave_mux.v(222)
  or u374 (n136[27], n134[27], n135[27]);  // ../RTL/cmsdk_apb_slave_mux.v(222)
  or u375 (n136[28], n134[28], n135[28]);  // ../RTL/cmsdk_apb_slave_mux.v(222)
  or u376 (n136[29], n134[29], n135[29]);  // ../RTL/cmsdk_apb_slave_mux.v(222)
  or u377 (n136[30], n134[30], n135[30]);  // ../RTL/cmsdk_apb_slave_mux.v(222)
  or u378 (n136[31], n134[31], n135[31]);  // ../RTL/cmsdk_apb_slave_mux.v(222)
  and u379 (n135[1], PSEL13, PRDATA13[1]);  // ../RTL/cmsdk_apb_slave_mux.v(222)
  or u38 (n18, PREADY0, n17);  // ../RTL/cmsdk_apb_slave_mux.v(175)
  and u380 (n135[2], PSEL13, PRDATA13[2]);  // ../RTL/cmsdk_apb_slave_mux.v(222)
  and u381 (n135[3], PSEL13, PRDATA13[3]);  // ../RTL/cmsdk_apb_slave_mux.v(222)
  and u382 (n135[4], PSEL13, PRDATA13[4]);  // ../RTL/cmsdk_apb_slave_mux.v(222)
  and u383 (n135[5], PSEL13, PRDATA13[5]);  // ../RTL/cmsdk_apb_slave_mux.v(222)
  and u384 (n135[6], PSEL13, PRDATA13[6]);  // ../RTL/cmsdk_apb_slave_mux.v(222)
  and u385 (n135[7], PSEL13, PRDATA13[7]);  // ../RTL/cmsdk_apb_slave_mux.v(222)
  and u386 (n135[8], PSEL13, PRDATA13[8]);  // ../RTL/cmsdk_apb_slave_mux.v(222)
  and u387 (n135[9], PSEL13, PRDATA13[9]);  // ../RTL/cmsdk_apb_slave_mux.v(222)
  and u388 (n135[10], PSEL13, PRDATA13[10]);  // ../RTL/cmsdk_apb_slave_mux.v(222)
  and u389 (n135[11], PSEL13, PRDATA13[11]);  // ../RTL/cmsdk_apb_slave_mux.v(222)
  and u39 (n19, dec[0], n18);  // ../RTL/cmsdk_apb_slave_mux.v(175)
  and u390 (n135[12], PSEL13, PRDATA13[12]);  // ../RTL/cmsdk_apb_slave_mux.v(222)
  and u391 (n135[13], PSEL13, PRDATA13[13]);  // ../RTL/cmsdk_apb_slave_mux.v(222)
  and u392 (n135[14], PSEL13, PRDATA13[14]);  // ../RTL/cmsdk_apb_slave_mux.v(222)
  and u393 (n135[15], PSEL13, PRDATA13[15]);  // ../RTL/cmsdk_apb_slave_mux.v(222)
  and u394 (n135[16], PSEL13, PRDATA13[16]);  // ../RTL/cmsdk_apb_slave_mux.v(222)
  and u395 (n135[17], PSEL13, PRDATA13[17]);  // ../RTL/cmsdk_apb_slave_mux.v(222)
  and u396 (n135[18], PSEL13, PRDATA13[18]);  // ../RTL/cmsdk_apb_slave_mux.v(222)
  and u397 (n135[19], PSEL13, PRDATA13[19]);  // ../RTL/cmsdk_apb_slave_mux.v(222)
  and u398 (n135[20], PSEL13, PRDATA13[20]);  // ../RTL/cmsdk_apb_slave_mux.v(222)
  and u399 (n135[21], PSEL13, PRDATA13[21]);  // ../RTL/cmsdk_apb_slave_mux.v(222)
  and u4 (n0, PSEL, dec[0]);  // ../RTL/cmsdk_apb_slave_mux.v(157)
  or u40 (n20, n16, n19);  // ../RTL/cmsdk_apb_slave_mux.v(175)
  and u400 (n135[22], PSEL13, PRDATA13[22]);  // ../RTL/cmsdk_apb_slave_mux.v(222)
  and u401 (n135[23], PSEL13, PRDATA13[23]);  // ../RTL/cmsdk_apb_slave_mux.v(222)
  and u402 (n135[24], PSEL13, PRDATA13[24]);  // ../RTL/cmsdk_apb_slave_mux.v(222)
  and u403 (n135[25], PSEL13, PRDATA13[25]);  // ../RTL/cmsdk_apb_slave_mux.v(222)
  and u404 (n135[26], PSEL13, PRDATA13[26]);  // ../RTL/cmsdk_apb_slave_mux.v(222)
  and u405 (n135[27], PSEL13, PRDATA13[27]);  // ../RTL/cmsdk_apb_slave_mux.v(222)
  and u406 (n135[28], PSEL13, PRDATA13[28]);  // ../RTL/cmsdk_apb_slave_mux.v(222)
  and u407 (n135[29], PSEL13, PRDATA13[29]);  // ../RTL/cmsdk_apb_slave_mux.v(222)
  and u408 (n135[30], PSEL13, PRDATA13[30]);  // ../RTL/cmsdk_apb_slave_mux.v(222)
  and u409 (n135[31], PSEL13, PRDATA13[31]);  // ../RTL/cmsdk_apb_slave_mux.v(222)
  not u41 (n21, en[1]);  // ../RTL/cmsdk_apb_slave_mux.v(176)
  or u410 (n134[1], n132[1], n133[1]);  // ../RTL/cmsdk_apb_slave_mux.v(221)
  or u411 (n134[2], n132[2], n133[2]);  // ../RTL/cmsdk_apb_slave_mux.v(221)
  or u412 (n134[3], n132[3], n133[3]);  // ../RTL/cmsdk_apb_slave_mux.v(221)
  or u413 (n134[4], n132[4], n133[4]);  // ../RTL/cmsdk_apb_slave_mux.v(221)
  or u414 (n134[5], n132[5], n133[5]);  // ../RTL/cmsdk_apb_slave_mux.v(221)
  or u415 (n134[6], n132[6], n133[6]);  // ../RTL/cmsdk_apb_slave_mux.v(221)
  or u416 (n134[7], n132[7], n133[7]);  // ../RTL/cmsdk_apb_slave_mux.v(221)
  or u417 (n134[8], n132[8], n133[8]);  // ../RTL/cmsdk_apb_slave_mux.v(221)
  or u418 (n134[9], n132[9], n133[9]);  // ../RTL/cmsdk_apb_slave_mux.v(221)
  or u419 (n134[10], n132[10], n133[10]);  // ../RTL/cmsdk_apb_slave_mux.v(221)
  or u42 (n22, PREADY1, n21);  // ../RTL/cmsdk_apb_slave_mux.v(176)
  or u420 (n134[11], n132[11], n133[11]);  // ../RTL/cmsdk_apb_slave_mux.v(221)
  or u421 (n134[12], n132[12], n133[12]);  // ../RTL/cmsdk_apb_slave_mux.v(221)
  or u422 (n134[13], n132[13], n133[13]);  // ../RTL/cmsdk_apb_slave_mux.v(221)
  or u423 (n134[14], n132[14], n133[14]);  // ../RTL/cmsdk_apb_slave_mux.v(221)
  or u424 (n134[15], n132[15], n133[15]);  // ../RTL/cmsdk_apb_slave_mux.v(221)
  or u425 (n134[16], n132[16], n133[16]);  // ../RTL/cmsdk_apb_slave_mux.v(221)
  or u426 (n134[17], n132[17], n133[17]);  // ../RTL/cmsdk_apb_slave_mux.v(221)
  or u427 (n134[18], n132[18], n133[18]);  // ../RTL/cmsdk_apb_slave_mux.v(221)
  or u428 (n134[19], n132[19], n133[19]);  // ../RTL/cmsdk_apb_slave_mux.v(221)
  or u429 (n134[20], n132[20], n133[20]);  // ../RTL/cmsdk_apb_slave_mux.v(221)
  and u43 (n23, dec[1], n22);  // ../RTL/cmsdk_apb_slave_mux.v(176)
  or u430 (n134[21], n132[21], n133[21]);  // ../RTL/cmsdk_apb_slave_mux.v(221)
  or u431 (n134[22], n132[22], n133[22]);  // ../RTL/cmsdk_apb_slave_mux.v(221)
  or u432 (n134[23], n132[23], n133[23]);  // ../RTL/cmsdk_apb_slave_mux.v(221)
  or u433 (n134[24], n132[24], n133[24]);  // ../RTL/cmsdk_apb_slave_mux.v(221)
  or u434 (n134[25], n132[25], n133[25]);  // ../RTL/cmsdk_apb_slave_mux.v(221)
  or u435 (n134[26], n132[26], n133[26]);  // ../RTL/cmsdk_apb_slave_mux.v(221)
  or u436 (n134[27], n132[27], n133[27]);  // ../RTL/cmsdk_apb_slave_mux.v(221)
  or u437 (n134[28], n132[28], n133[28]);  // ../RTL/cmsdk_apb_slave_mux.v(221)
  or u438 (n134[29], n132[29], n133[29]);  // ../RTL/cmsdk_apb_slave_mux.v(221)
  or u439 (n134[30], n132[30], n133[30]);  // ../RTL/cmsdk_apb_slave_mux.v(221)
  or u44 (n24, n20, n23);  // ../RTL/cmsdk_apb_slave_mux.v(176)
  or u440 (n134[31], n132[31], n133[31]);  // ../RTL/cmsdk_apb_slave_mux.v(221)
  and u441 (n133[1], PSEL12, PRDATA12[1]);  // ../RTL/cmsdk_apb_slave_mux.v(221)
  and u442 (n133[2], PSEL12, PRDATA12[2]);  // ../RTL/cmsdk_apb_slave_mux.v(221)
  and u443 (n133[3], PSEL12, PRDATA12[3]);  // ../RTL/cmsdk_apb_slave_mux.v(221)
  and u444 (n133[4], PSEL12, PRDATA12[4]);  // ../RTL/cmsdk_apb_slave_mux.v(221)
  and u445 (n133[5], PSEL12, PRDATA12[5]);  // ../RTL/cmsdk_apb_slave_mux.v(221)
  and u446 (n133[6], PSEL12, PRDATA12[6]);  // ../RTL/cmsdk_apb_slave_mux.v(221)
  and u447 (n133[7], PSEL12, PRDATA12[7]);  // ../RTL/cmsdk_apb_slave_mux.v(221)
  and u448 (n133[8], PSEL12, PRDATA12[8]);  // ../RTL/cmsdk_apb_slave_mux.v(221)
  and u449 (n133[9], PSEL12, PRDATA12[9]);  // ../RTL/cmsdk_apb_slave_mux.v(221)
  not u45 (n25, en[2]);  // ../RTL/cmsdk_apb_slave_mux.v(177)
  and u450 (n133[10], PSEL12, PRDATA12[10]);  // ../RTL/cmsdk_apb_slave_mux.v(221)
  and u451 (n133[11], PSEL12, PRDATA12[11]);  // ../RTL/cmsdk_apb_slave_mux.v(221)
  and u452 (n133[12], PSEL12, PRDATA12[12]);  // ../RTL/cmsdk_apb_slave_mux.v(221)
  and u453 (n133[13], PSEL12, PRDATA12[13]);  // ../RTL/cmsdk_apb_slave_mux.v(221)
  and u454 (n133[14], PSEL12, PRDATA12[14]);  // ../RTL/cmsdk_apb_slave_mux.v(221)
  and u455 (n133[15], PSEL12, PRDATA12[15]);  // ../RTL/cmsdk_apb_slave_mux.v(221)
  and u456 (n133[16], PSEL12, PRDATA12[16]);  // ../RTL/cmsdk_apb_slave_mux.v(221)
  and u457 (n133[17], PSEL12, PRDATA12[17]);  // ../RTL/cmsdk_apb_slave_mux.v(221)
  and u458 (n133[18], PSEL12, PRDATA12[18]);  // ../RTL/cmsdk_apb_slave_mux.v(221)
  and u459 (n133[19], PSEL12, PRDATA12[19]);  // ../RTL/cmsdk_apb_slave_mux.v(221)
  or u46 (n26, PREADY2, n25);  // ../RTL/cmsdk_apb_slave_mux.v(177)
  and u460 (n133[20], PSEL12, PRDATA12[20]);  // ../RTL/cmsdk_apb_slave_mux.v(221)
  and u461 (n133[21], PSEL12, PRDATA12[21]);  // ../RTL/cmsdk_apb_slave_mux.v(221)
  and u462 (n133[22], PSEL12, PRDATA12[22]);  // ../RTL/cmsdk_apb_slave_mux.v(221)
  and u463 (n133[23], PSEL12, PRDATA12[23]);  // ../RTL/cmsdk_apb_slave_mux.v(221)
  and u464 (n133[24], PSEL12, PRDATA12[24]);  // ../RTL/cmsdk_apb_slave_mux.v(221)
  and u465 (n133[25], PSEL12, PRDATA12[25]);  // ../RTL/cmsdk_apb_slave_mux.v(221)
  and u466 (n133[26], PSEL12, PRDATA12[26]);  // ../RTL/cmsdk_apb_slave_mux.v(221)
  and u467 (n133[27], PSEL12, PRDATA12[27]);  // ../RTL/cmsdk_apb_slave_mux.v(221)
  and u468 (n133[28], PSEL12, PRDATA12[28]);  // ../RTL/cmsdk_apb_slave_mux.v(221)
  and u469 (n133[29], PSEL12, PRDATA12[29]);  // ../RTL/cmsdk_apb_slave_mux.v(221)
  and u47 (n27, dec[2], n26);  // ../RTL/cmsdk_apb_slave_mux.v(177)
  and u470 (n133[30], PSEL12, PRDATA12[30]);  // ../RTL/cmsdk_apb_slave_mux.v(221)
  and u471 (n133[31], PSEL12, PRDATA12[31]);  // ../RTL/cmsdk_apb_slave_mux.v(221)
  or u472 (n132[1], n130[1], n131[1]);  // ../RTL/cmsdk_apb_slave_mux.v(220)
  or u473 (n132[2], n130[2], n131[2]);  // ../RTL/cmsdk_apb_slave_mux.v(220)
  or u474 (n132[3], n130[3], n131[3]);  // ../RTL/cmsdk_apb_slave_mux.v(220)
  or u475 (n132[4], n130[4], n131[4]);  // ../RTL/cmsdk_apb_slave_mux.v(220)
  or u476 (n132[5], n130[5], n131[5]);  // ../RTL/cmsdk_apb_slave_mux.v(220)
  or u477 (n132[6], n130[6], n131[6]);  // ../RTL/cmsdk_apb_slave_mux.v(220)
  or u478 (n132[7], n130[7], n131[7]);  // ../RTL/cmsdk_apb_slave_mux.v(220)
  or u479 (n132[8], n130[8], n131[8]);  // ../RTL/cmsdk_apb_slave_mux.v(220)
  or u48 (n28, n24, n27);  // ../RTL/cmsdk_apb_slave_mux.v(177)
  or u480 (n132[9], n130[9], n131[9]);  // ../RTL/cmsdk_apb_slave_mux.v(220)
  or u481 (n132[10], n130[10], n131[10]);  // ../RTL/cmsdk_apb_slave_mux.v(220)
  or u482 (n132[11], n130[11], n131[11]);  // ../RTL/cmsdk_apb_slave_mux.v(220)
  or u483 (n132[12], n130[12], n131[12]);  // ../RTL/cmsdk_apb_slave_mux.v(220)
  or u484 (n132[13], n130[13], n131[13]);  // ../RTL/cmsdk_apb_slave_mux.v(220)
  or u485 (n132[14], n130[14], n131[14]);  // ../RTL/cmsdk_apb_slave_mux.v(220)
  or u486 (n132[15], n130[15], n131[15]);  // ../RTL/cmsdk_apb_slave_mux.v(220)
  or u487 (n132[16], n130[16], n131[16]);  // ../RTL/cmsdk_apb_slave_mux.v(220)
  or u488 (n132[17], n130[17], n131[17]);  // ../RTL/cmsdk_apb_slave_mux.v(220)
  or u489 (n132[18], n130[18], n131[18]);  // ../RTL/cmsdk_apb_slave_mux.v(220)
  not u49 (n29, en[3]);  // ../RTL/cmsdk_apb_slave_mux.v(178)
  or u490 (n132[19], n130[19], n131[19]);  // ../RTL/cmsdk_apb_slave_mux.v(220)
  or u491 (n132[20], n130[20], n131[20]);  // ../RTL/cmsdk_apb_slave_mux.v(220)
  or u492 (n132[21], n130[21], n131[21]);  // ../RTL/cmsdk_apb_slave_mux.v(220)
  or u493 (n132[22], n130[22], n131[22]);  // ../RTL/cmsdk_apb_slave_mux.v(220)
  or u494 (n132[23], n130[23], n131[23]);  // ../RTL/cmsdk_apb_slave_mux.v(220)
  or u495 (n132[24], n130[24], n131[24]);  // ../RTL/cmsdk_apb_slave_mux.v(220)
  or u496 (n132[25], n130[25], n131[25]);  // ../RTL/cmsdk_apb_slave_mux.v(220)
  or u497 (n132[26], n130[26], n131[26]);  // ../RTL/cmsdk_apb_slave_mux.v(220)
  or u498 (n132[27], n130[27], n131[27]);  // ../RTL/cmsdk_apb_slave_mux.v(220)
  or u499 (n132[28], n130[28], n131[28]);  // ../RTL/cmsdk_apb_slave_mux.v(220)
  and u5 (PSEL0, n0, en[0]);  // ../RTL/cmsdk_apb_slave_mux.v(157)
  or u50 (n30, PREADY3, n29);  // ../RTL/cmsdk_apb_slave_mux.v(178)
  or u500 (n132[29], n130[29], n131[29]);  // ../RTL/cmsdk_apb_slave_mux.v(220)
  or u501 (n132[30], n130[30], n131[30]);  // ../RTL/cmsdk_apb_slave_mux.v(220)
  or u502 (n132[31], n130[31], n131[31]);  // ../RTL/cmsdk_apb_slave_mux.v(220)
  and u503 (n131[1], PSEL11, PRDATA11[1]);  // ../RTL/cmsdk_apb_slave_mux.v(220)
  and u504 (n131[2], PSEL11, PRDATA11[2]);  // ../RTL/cmsdk_apb_slave_mux.v(220)
  and u505 (n131[3], PSEL11, PRDATA11[3]);  // ../RTL/cmsdk_apb_slave_mux.v(220)
  and u506 (n131[4], PSEL11, PRDATA11[4]);  // ../RTL/cmsdk_apb_slave_mux.v(220)
  and u507 (n131[5], PSEL11, PRDATA11[5]);  // ../RTL/cmsdk_apb_slave_mux.v(220)
  and u508 (n131[6], PSEL11, PRDATA11[6]);  // ../RTL/cmsdk_apb_slave_mux.v(220)
  and u509 (n131[7], PSEL11, PRDATA11[7]);  // ../RTL/cmsdk_apb_slave_mux.v(220)
  and u51 (n31, dec[3], n30);  // ../RTL/cmsdk_apb_slave_mux.v(178)
  and u510 (n131[8], PSEL11, PRDATA11[8]);  // ../RTL/cmsdk_apb_slave_mux.v(220)
  and u511 (n131[9], PSEL11, PRDATA11[9]);  // ../RTL/cmsdk_apb_slave_mux.v(220)
  and u512 (n131[10], PSEL11, PRDATA11[10]);  // ../RTL/cmsdk_apb_slave_mux.v(220)
  and u513 (n131[11], PSEL11, PRDATA11[11]);  // ../RTL/cmsdk_apb_slave_mux.v(220)
  and u514 (n131[12], PSEL11, PRDATA11[12]);  // ../RTL/cmsdk_apb_slave_mux.v(220)
  and u515 (n131[13], PSEL11, PRDATA11[13]);  // ../RTL/cmsdk_apb_slave_mux.v(220)
  and u516 (n131[14], PSEL11, PRDATA11[14]);  // ../RTL/cmsdk_apb_slave_mux.v(220)
  and u517 (n131[15], PSEL11, PRDATA11[15]);  // ../RTL/cmsdk_apb_slave_mux.v(220)
  and u518 (n131[16], PSEL11, PRDATA11[16]);  // ../RTL/cmsdk_apb_slave_mux.v(220)
  and u519 (n131[17], PSEL11, PRDATA11[17]);  // ../RTL/cmsdk_apb_slave_mux.v(220)
  or u52 (n32, n28, n31);  // ../RTL/cmsdk_apb_slave_mux.v(178)
  and u520 (n131[18], PSEL11, PRDATA11[18]);  // ../RTL/cmsdk_apb_slave_mux.v(220)
  and u521 (n131[19], PSEL11, PRDATA11[19]);  // ../RTL/cmsdk_apb_slave_mux.v(220)
  and u522 (n131[20], PSEL11, PRDATA11[20]);  // ../RTL/cmsdk_apb_slave_mux.v(220)
  and u523 (n131[21], PSEL11, PRDATA11[21]);  // ../RTL/cmsdk_apb_slave_mux.v(220)
  and u524 (n131[22], PSEL11, PRDATA11[22]);  // ../RTL/cmsdk_apb_slave_mux.v(220)
  and u525 (n131[23], PSEL11, PRDATA11[23]);  // ../RTL/cmsdk_apb_slave_mux.v(220)
  and u526 (n131[24], PSEL11, PRDATA11[24]);  // ../RTL/cmsdk_apb_slave_mux.v(220)
  and u527 (n131[25], PSEL11, PRDATA11[25]);  // ../RTL/cmsdk_apb_slave_mux.v(220)
  and u528 (n131[26], PSEL11, PRDATA11[26]);  // ../RTL/cmsdk_apb_slave_mux.v(220)
  and u529 (n131[27], PSEL11, PRDATA11[27]);  // ../RTL/cmsdk_apb_slave_mux.v(220)
  not u53 (n33, en[4]);  // ../RTL/cmsdk_apb_slave_mux.v(179)
  and u530 (n131[28], PSEL11, PRDATA11[28]);  // ../RTL/cmsdk_apb_slave_mux.v(220)
  and u531 (n131[29], PSEL11, PRDATA11[29]);  // ../RTL/cmsdk_apb_slave_mux.v(220)
  and u532 (n131[30], PSEL11, PRDATA11[30]);  // ../RTL/cmsdk_apb_slave_mux.v(220)
  and u533 (n131[31], PSEL11, PRDATA11[31]);  // ../RTL/cmsdk_apb_slave_mux.v(220)
  or u534 (n130[1], n128[1], n129[1]);  // ../RTL/cmsdk_apb_slave_mux.v(219)
  or u535 (n130[2], n128[2], n129[2]);  // ../RTL/cmsdk_apb_slave_mux.v(219)
  or u536 (n130[3], n128[3], n129[3]);  // ../RTL/cmsdk_apb_slave_mux.v(219)
  or u537 (n130[4], n128[4], n129[4]);  // ../RTL/cmsdk_apb_slave_mux.v(219)
  or u538 (n130[5], n128[5], n129[5]);  // ../RTL/cmsdk_apb_slave_mux.v(219)
  or u539 (n130[6], n128[6], n129[6]);  // ../RTL/cmsdk_apb_slave_mux.v(219)
  or u54 (n34, PREADY4, n33);  // ../RTL/cmsdk_apb_slave_mux.v(179)
  or u540 (n130[7], n128[7], n129[7]);  // ../RTL/cmsdk_apb_slave_mux.v(219)
  or u541 (n130[8], n128[8], n129[8]);  // ../RTL/cmsdk_apb_slave_mux.v(219)
  or u542 (n130[9], n128[9], n129[9]);  // ../RTL/cmsdk_apb_slave_mux.v(219)
  or u543 (n130[10], n128[10], n129[10]);  // ../RTL/cmsdk_apb_slave_mux.v(219)
  or u544 (n130[11], n128[11], n129[11]);  // ../RTL/cmsdk_apb_slave_mux.v(219)
  or u545 (n130[12], n128[12], n129[12]);  // ../RTL/cmsdk_apb_slave_mux.v(219)
  or u546 (n130[13], n128[13], n129[13]);  // ../RTL/cmsdk_apb_slave_mux.v(219)
  or u547 (n130[14], n128[14], n129[14]);  // ../RTL/cmsdk_apb_slave_mux.v(219)
  or u548 (n130[15], n128[15], n129[15]);  // ../RTL/cmsdk_apb_slave_mux.v(219)
  or u549 (n130[16], n128[16], n129[16]);  // ../RTL/cmsdk_apb_slave_mux.v(219)
  and u55 (n35, dec[4], n34);  // ../RTL/cmsdk_apb_slave_mux.v(179)
  or u550 (n130[17], n128[17], n129[17]);  // ../RTL/cmsdk_apb_slave_mux.v(219)
  or u551 (n130[18], n128[18], n129[18]);  // ../RTL/cmsdk_apb_slave_mux.v(219)
  or u552 (n130[19], n128[19], n129[19]);  // ../RTL/cmsdk_apb_slave_mux.v(219)
  or u553 (n130[20], n128[20], n129[20]);  // ../RTL/cmsdk_apb_slave_mux.v(219)
  or u554 (n130[21], n128[21], n129[21]);  // ../RTL/cmsdk_apb_slave_mux.v(219)
  or u555 (n130[22], n128[22], n129[22]);  // ../RTL/cmsdk_apb_slave_mux.v(219)
  or u556 (n130[23], n128[23], n129[23]);  // ../RTL/cmsdk_apb_slave_mux.v(219)
  or u557 (n130[24], n128[24], n129[24]);  // ../RTL/cmsdk_apb_slave_mux.v(219)
  or u558 (n130[25], n128[25], n129[25]);  // ../RTL/cmsdk_apb_slave_mux.v(219)
  or u559 (n130[26], n128[26], n129[26]);  // ../RTL/cmsdk_apb_slave_mux.v(219)
  or u56 (n36, n32, n35);  // ../RTL/cmsdk_apb_slave_mux.v(179)
  or u560 (n130[27], n128[27], n129[27]);  // ../RTL/cmsdk_apb_slave_mux.v(219)
  or u561 (n130[28], n128[28], n129[28]);  // ../RTL/cmsdk_apb_slave_mux.v(219)
  or u562 (n130[29], n128[29], n129[29]);  // ../RTL/cmsdk_apb_slave_mux.v(219)
  or u563 (n130[30], n128[30], n129[30]);  // ../RTL/cmsdk_apb_slave_mux.v(219)
  or u564 (n130[31], n128[31], n129[31]);  // ../RTL/cmsdk_apb_slave_mux.v(219)
  and u565 (n129[1], PSEL10, PRDATA10[1]);  // ../RTL/cmsdk_apb_slave_mux.v(219)
  and u566 (n129[2], PSEL10, PRDATA10[2]);  // ../RTL/cmsdk_apb_slave_mux.v(219)
  and u567 (n129[3], PSEL10, PRDATA10[3]);  // ../RTL/cmsdk_apb_slave_mux.v(219)
  and u568 (n129[4], PSEL10, PRDATA10[4]);  // ../RTL/cmsdk_apb_slave_mux.v(219)
  and u569 (n129[5], PSEL10, PRDATA10[5]);  // ../RTL/cmsdk_apb_slave_mux.v(219)
  not u57 (n37, en[5]);  // ../RTL/cmsdk_apb_slave_mux.v(180)
  and u570 (n129[6], PSEL10, PRDATA10[6]);  // ../RTL/cmsdk_apb_slave_mux.v(219)
  and u571 (n129[7], PSEL10, PRDATA10[7]);  // ../RTL/cmsdk_apb_slave_mux.v(219)
  and u572 (n129[8], PSEL10, PRDATA10[8]);  // ../RTL/cmsdk_apb_slave_mux.v(219)
  and u573 (n129[9], PSEL10, PRDATA10[9]);  // ../RTL/cmsdk_apb_slave_mux.v(219)
  and u574 (n129[10], PSEL10, PRDATA10[10]);  // ../RTL/cmsdk_apb_slave_mux.v(219)
  and u575 (n129[11], PSEL10, PRDATA10[11]);  // ../RTL/cmsdk_apb_slave_mux.v(219)
  and u576 (n129[12], PSEL10, PRDATA10[12]);  // ../RTL/cmsdk_apb_slave_mux.v(219)
  and u577 (n129[13], PSEL10, PRDATA10[13]);  // ../RTL/cmsdk_apb_slave_mux.v(219)
  and u578 (n129[14], PSEL10, PRDATA10[14]);  // ../RTL/cmsdk_apb_slave_mux.v(219)
  and u579 (n129[15], PSEL10, PRDATA10[15]);  // ../RTL/cmsdk_apb_slave_mux.v(219)
  or u58 (n38, PREADY5, n37);  // ../RTL/cmsdk_apb_slave_mux.v(180)
  and u580 (n129[16], PSEL10, PRDATA10[16]);  // ../RTL/cmsdk_apb_slave_mux.v(219)
  and u581 (n129[17], PSEL10, PRDATA10[17]);  // ../RTL/cmsdk_apb_slave_mux.v(219)
  and u582 (n129[18], PSEL10, PRDATA10[18]);  // ../RTL/cmsdk_apb_slave_mux.v(219)
  and u583 (n129[19], PSEL10, PRDATA10[19]);  // ../RTL/cmsdk_apb_slave_mux.v(219)
  and u584 (n129[20], PSEL10, PRDATA10[20]);  // ../RTL/cmsdk_apb_slave_mux.v(219)
  and u585 (n129[21], PSEL10, PRDATA10[21]);  // ../RTL/cmsdk_apb_slave_mux.v(219)
  and u586 (n129[22], PSEL10, PRDATA10[22]);  // ../RTL/cmsdk_apb_slave_mux.v(219)
  and u587 (n129[23], PSEL10, PRDATA10[23]);  // ../RTL/cmsdk_apb_slave_mux.v(219)
  and u588 (n129[24], PSEL10, PRDATA10[24]);  // ../RTL/cmsdk_apb_slave_mux.v(219)
  and u589 (n129[25], PSEL10, PRDATA10[25]);  // ../RTL/cmsdk_apb_slave_mux.v(219)
  and u59 (n39, dec[5], n38);  // ../RTL/cmsdk_apb_slave_mux.v(180)
  and u590 (n129[26], PSEL10, PRDATA10[26]);  // ../RTL/cmsdk_apb_slave_mux.v(219)
  and u591 (n129[27], PSEL10, PRDATA10[27]);  // ../RTL/cmsdk_apb_slave_mux.v(219)
  and u592 (n129[28], PSEL10, PRDATA10[28]);  // ../RTL/cmsdk_apb_slave_mux.v(219)
  and u593 (n129[29], PSEL10, PRDATA10[29]);  // ../RTL/cmsdk_apb_slave_mux.v(219)
  and u594 (n129[30], PSEL10, PRDATA10[30]);  // ../RTL/cmsdk_apb_slave_mux.v(219)
  and u595 (n129[31], PSEL10, PRDATA10[31]);  // ../RTL/cmsdk_apb_slave_mux.v(219)
  or u596 (n128[1], n126[1], n127[1]);  // ../RTL/cmsdk_apb_slave_mux.v(218)
  or u597 (n128[2], n126[2], n127[2]);  // ../RTL/cmsdk_apb_slave_mux.v(218)
  or u598 (n128[3], n126[3], n127[3]);  // ../RTL/cmsdk_apb_slave_mux.v(218)
  or u599 (n128[4], n126[4], n127[4]);  // ../RTL/cmsdk_apb_slave_mux.v(218)
  and u6 (n1, PSEL, dec[1]);  // ../RTL/cmsdk_apb_slave_mux.v(158)
  or u60 (n40, n36, n39);  // ../RTL/cmsdk_apb_slave_mux.v(180)
  or u600 (n128[5], n126[5], n127[5]);  // ../RTL/cmsdk_apb_slave_mux.v(218)
  or u601 (n128[6], n126[6], n127[6]);  // ../RTL/cmsdk_apb_slave_mux.v(218)
  or u602 (n128[7], n126[7], n127[7]);  // ../RTL/cmsdk_apb_slave_mux.v(218)
  or u603 (n128[8], n126[8], n127[8]);  // ../RTL/cmsdk_apb_slave_mux.v(218)
  or u604 (n128[9], n126[9], n127[9]);  // ../RTL/cmsdk_apb_slave_mux.v(218)
  or u605 (n128[10], n126[10], n127[10]);  // ../RTL/cmsdk_apb_slave_mux.v(218)
  or u606 (n128[11], n126[11], n127[11]);  // ../RTL/cmsdk_apb_slave_mux.v(218)
  or u607 (n128[12], n126[12], n127[12]);  // ../RTL/cmsdk_apb_slave_mux.v(218)
  or u608 (n128[13], n126[13], n127[13]);  // ../RTL/cmsdk_apb_slave_mux.v(218)
  or u609 (n128[14], n126[14], n127[14]);  // ../RTL/cmsdk_apb_slave_mux.v(218)
  not u61 (n41, en[6]);  // ../RTL/cmsdk_apb_slave_mux.v(181)
  or u610 (n128[15], n126[15], n127[15]);  // ../RTL/cmsdk_apb_slave_mux.v(218)
  or u611 (n128[16], n126[16], n127[16]);  // ../RTL/cmsdk_apb_slave_mux.v(218)
  or u612 (n128[17], n126[17], n127[17]);  // ../RTL/cmsdk_apb_slave_mux.v(218)
  or u613 (n128[18], n126[18], n127[18]);  // ../RTL/cmsdk_apb_slave_mux.v(218)
  or u614 (n128[19], n126[19], n127[19]);  // ../RTL/cmsdk_apb_slave_mux.v(218)
  or u615 (n128[20], n126[20], n127[20]);  // ../RTL/cmsdk_apb_slave_mux.v(218)
  or u616 (n128[21], n126[21], n127[21]);  // ../RTL/cmsdk_apb_slave_mux.v(218)
  or u617 (n128[22], n126[22], n127[22]);  // ../RTL/cmsdk_apb_slave_mux.v(218)
  or u618 (n128[23], n126[23], n127[23]);  // ../RTL/cmsdk_apb_slave_mux.v(218)
  or u619 (n128[24], n126[24], n127[24]);  // ../RTL/cmsdk_apb_slave_mux.v(218)
  or u62 (n42, PREADY6, n41);  // ../RTL/cmsdk_apb_slave_mux.v(181)
  or u620 (n128[25], n126[25], n127[25]);  // ../RTL/cmsdk_apb_slave_mux.v(218)
  or u621 (n128[26], n126[26], n127[26]);  // ../RTL/cmsdk_apb_slave_mux.v(218)
  or u622 (n128[27], n126[27], n127[27]);  // ../RTL/cmsdk_apb_slave_mux.v(218)
  or u623 (n128[28], n126[28], n127[28]);  // ../RTL/cmsdk_apb_slave_mux.v(218)
  or u624 (n128[29], n126[29], n127[29]);  // ../RTL/cmsdk_apb_slave_mux.v(218)
  or u625 (n128[30], n126[30], n127[30]);  // ../RTL/cmsdk_apb_slave_mux.v(218)
  or u626 (n128[31], n126[31], n127[31]);  // ../RTL/cmsdk_apb_slave_mux.v(218)
  and u627 (n127[1], PSEL9, PRDATA9[1]);  // ../RTL/cmsdk_apb_slave_mux.v(218)
  and u628 (n127[2], PSEL9, PRDATA9[2]);  // ../RTL/cmsdk_apb_slave_mux.v(218)
  and u629 (n127[3], PSEL9, PRDATA9[3]);  // ../RTL/cmsdk_apb_slave_mux.v(218)
  and u63 (n43, dec[6], n42);  // ../RTL/cmsdk_apb_slave_mux.v(181)
  and u630 (n127[4], PSEL9, PRDATA9[4]);  // ../RTL/cmsdk_apb_slave_mux.v(218)
  and u631 (n127[5], PSEL9, PRDATA9[5]);  // ../RTL/cmsdk_apb_slave_mux.v(218)
  and u632 (n127[6], PSEL9, PRDATA9[6]);  // ../RTL/cmsdk_apb_slave_mux.v(218)
  and u633 (n127[7], PSEL9, PRDATA9[7]);  // ../RTL/cmsdk_apb_slave_mux.v(218)
  and u634 (n127[8], PSEL9, PRDATA9[8]);  // ../RTL/cmsdk_apb_slave_mux.v(218)
  and u635 (n127[9], PSEL9, PRDATA9[9]);  // ../RTL/cmsdk_apb_slave_mux.v(218)
  and u636 (n127[10], PSEL9, PRDATA9[10]);  // ../RTL/cmsdk_apb_slave_mux.v(218)
  and u637 (n127[11], PSEL9, PRDATA9[11]);  // ../RTL/cmsdk_apb_slave_mux.v(218)
  and u638 (n127[12], PSEL9, PRDATA9[12]);  // ../RTL/cmsdk_apb_slave_mux.v(218)
  and u639 (n127[13], PSEL9, PRDATA9[13]);  // ../RTL/cmsdk_apb_slave_mux.v(218)
  or u64 (n44, n40, n43);  // ../RTL/cmsdk_apb_slave_mux.v(181)
  and u640 (n127[14], PSEL9, PRDATA9[14]);  // ../RTL/cmsdk_apb_slave_mux.v(218)
  and u641 (n127[15], PSEL9, PRDATA9[15]);  // ../RTL/cmsdk_apb_slave_mux.v(218)
  and u642 (n127[16], PSEL9, PRDATA9[16]);  // ../RTL/cmsdk_apb_slave_mux.v(218)
  and u643 (n127[17], PSEL9, PRDATA9[17]);  // ../RTL/cmsdk_apb_slave_mux.v(218)
  and u644 (n127[18], PSEL9, PRDATA9[18]);  // ../RTL/cmsdk_apb_slave_mux.v(218)
  and u645 (n127[19], PSEL9, PRDATA9[19]);  // ../RTL/cmsdk_apb_slave_mux.v(218)
  and u646 (n127[20], PSEL9, PRDATA9[20]);  // ../RTL/cmsdk_apb_slave_mux.v(218)
  and u647 (n127[21], PSEL9, PRDATA9[21]);  // ../RTL/cmsdk_apb_slave_mux.v(218)
  and u648 (n127[22], PSEL9, PRDATA9[22]);  // ../RTL/cmsdk_apb_slave_mux.v(218)
  and u649 (n127[23], PSEL9, PRDATA9[23]);  // ../RTL/cmsdk_apb_slave_mux.v(218)
  not u65 (n45, en[7]);  // ../RTL/cmsdk_apb_slave_mux.v(182)
  and u650 (n127[24], PSEL9, PRDATA9[24]);  // ../RTL/cmsdk_apb_slave_mux.v(218)
  and u651 (n127[25], PSEL9, PRDATA9[25]);  // ../RTL/cmsdk_apb_slave_mux.v(218)
  and u652 (n127[26], PSEL9, PRDATA9[26]);  // ../RTL/cmsdk_apb_slave_mux.v(218)
  and u653 (n127[27], PSEL9, PRDATA9[27]);  // ../RTL/cmsdk_apb_slave_mux.v(218)
  and u654 (n127[28], PSEL9, PRDATA9[28]);  // ../RTL/cmsdk_apb_slave_mux.v(218)
  and u655 (n127[29], PSEL9, PRDATA9[29]);  // ../RTL/cmsdk_apb_slave_mux.v(218)
  and u656 (n127[30], PSEL9, PRDATA9[30]);  // ../RTL/cmsdk_apb_slave_mux.v(218)
  and u657 (n127[31], PSEL9, PRDATA9[31]);  // ../RTL/cmsdk_apb_slave_mux.v(218)
  or u658 (n126[1], n124[1], n125[1]);  // ../RTL/cmsdk_apb_slave_mux.v(217)
  or u659 (n126[2], n124[2], n125[2]);  // ../RTL/cmsdk_apb_slave_mux.v(217)
  or u66 (n46, PREADY7, n45);  // ../RTL/cmsdk_apb_slave_mux.v(182)
  or u660 (n126[3], n124[3], n125[3]);  // ../RTL/cmsdk_apb_slave_mux.v(217)
  or u661 (n126[4], n124[4], n125[4]);  // ../RTL/cmsdk_apb_slave_mux.v(217)
  or u662 (n126[5], n124[5], n125[5]);  // ../RTL/cmsdk_apb_slave_mux.v(217)
  or u663 (n126[6], n124[6], n125[6]);  // ../RTL/cmsdk_apb_slave_mux.v(217)
  or u664 (n126[7], n124[7], n125[7]);  // ../RTL/cmsdk_apb_slave_mux.v(217)
  or u665 (n126[8], n124[8], n125[8]);  // ../RTL/cmsdk_apb_slave_mux.v(217)
  or u666 (n126[9], n124[9], n125[9]);  // ../RTL/cmsdk_apb_slave_mux.v(217)
  or u667 (n126[10], n124[10], n125[10]);  // ../RTL/cmsdk_apb_slave_mux.v(217)
  or u668 (n126[11], n124[11], n125[11]);  // ../RTL/cmsdk_apb_slave_mux.v(217)
  or u669 (n126[12], n124[12], n125[12]);  // ../RTL/cmsdk_apb_slave_mux.v(217)
  and u67 (n47, dec[7], n46);  // ../RTL/cmsdk_apb_slave_mux.v(182)
  or u670 (n126[13], n124[13], n125[13]);  // ../RTL/cmsdk_apb_slave_mux.v(217)
  or u671 (n126[14], n124[14], n125[14]);  // ../RTL/cmsdk_apb_slave_mux.v(217)
  or u672 (n126[15], n124[15], n125[15]);  // ../RTL/cmsdk_apb_slave_mux.v(217)
  or u673 (n126[16], n124[16], n125[16]);  // ../RTL/cmsdk_apb_slave_mux.v(217)
  or u674 (n126[17], n124[17], n125[17]);  // ../RTL/cmsdk_apb_slave_mux.v(217)
  or u675 (n126[18], n124[18], n125[18]);  // ../RTL/cmsdk_apb_slave_mux.v(217)
  or u676 (n126[19], n124[19], n125[19]);  // ../RTL/cmsdk_apb_slave_mux.v(217)
  or u677 (n126[20], n124[20], n125[20]);  // ../RTL/cmsdk_apb_slave_mux.v(217)
  or u678 (n126[21], n124[21], n125[21]);  // ../RTL/cmsdk_apb_slave_mux.v(217)
  or u679 (n126[22], n124[22], n125[22]);  // ../RTL/cmsdk_apb_slave_mux.v(217)
  or u68 (n48, n44, n47);  // ../RTL/cmsdk_apb_slave_mux.v(182)
  or u680 (n126[23], n124[23], n125[23]);  // ../RTL/cmsdk_apb_slave_mux.v(217)
  or u681 (n126[24], n124[24], n125[24]);  // ../RTL/cmsdk_apb_slave_mux.v(217)
  or u682 (n126[25], n124[25], n125[25]);  // ../RTL/cmsdk_apb_slave_mux.v(217)
  or u683 (n126[26], n124[26], n125[26]);  // ../RTL/cmsdk_apb_slave_mux.v(217)
  or u684 (n126[27], n124[27], n125[27]);  // ../RTL/cmsdk_apb_slave_mux.v(217)
  or u685 (n126[28], n124[28], n125[28]);  // ../RTL/cmsdk_apb_slave_mux.v(217)
  or u686 (n126[29], n124[29], n125[29]);  // ../RTL/cmsdk_apb_slave_mux.v(217)
  or u687 (n126[30], n124[30], n125[30]);  // ../RTL/cmsdk_apb_slave_mux.v(217)
  or u688 (n126[31], n124[31], n125[31]);  // ../RTL/cmsdk_apb_slave_mux.v(217)
  and u689 (n125[1], PSEL8, PRDATA8[1]);  // ../RTL/cmsdk_apb_slave_mux.v(217)
  not u69 (n49, en[8]);  // ../RTL/cmsdk_apb_slave_mux.v(183)
  and u690 (n125[2], PSEL8, PRDATA8[2]);  // ../RTL/cmsdk_apb_slave_mux.v(217)
  and u691 (n125[3], PSEL8, PRDATA8[3]);  // ../RTL/cmsdk_apb_slave_mux.v(217)
  and u692 (n125[4], PSEL8, PRDATA8[4]);  // ../RTL/cmsdk_apb_slave_mux.v(217)
  and u693 (n125[5], PSEL8, PRDATA8[5]);  // ../RTL/cmsdk_apb_slave_mux.v(217)
  and u694 (n125[6], PSEL8, PRDATA8[6]);  // ../RTL/cmsdk_apb_slave_mux.v(217)
  and u695 (n125[7], PSEL8, PRDATA8[7]);  // ../RTL/cmsdk_apb_slave_mux.v(217)
  and u696 (n125[8], PSEL8, PRDATA8[8]);  // ../RTL/cmsdk_apb_slave_mux.v(217)
  and u697 (n125[9], PSEL8, PRDATA8[9]);  // ../RTL/cmsdk_apb_slave_mux.v(217)
  and u698 (n125[10], PSEL8, PRDATA8[10]);  // ../RTL/cmsdk_apb_slave_mux.v(217)
  and u699 (n125[11], PSEL8, PRDATA8[11]);  // ../RTL/cmsdk_apb_slave_mux.v(217)
  and u7 (PSEL1, n1, en[1]);  // ../RTL/cmsdk_apb_slave_mux.v(158)
  or u70 (n50, PREADY8, n49);  // ../RTL/cmsdk_apb_slave_mux.v(183)
  and u700 (n125[12], PSEL8, PRDATA8[12]);  // ../RTL/cmsdk_apb_slave_mux.v(217)
  and u701 (n125[13], PSEL8, PRDATA8[13]);  // ../RTL/cmsdk_apb_slave_mux.v(217)
  and u702 (n125[14], PSEL8, PRDATA8[14]);  // ../RTL/cmsdk_apb_slave_mux.v(217)
  and u703 (n125[15], PSEL8, PRDATA8[15]);  // ../RTL/cmsdk_apb_slave_mux.v(217)
  and u704 (n125[16], PSEL8, PRDATA8[16]);  // ../RTL/cmsdk_apb_slave_mux.v(217)
  and u705 (n125[17], PSEL8, PRDATA8[17]);  // ../RTL/cmsdk_apb_slave_mux.v(217)
  and u706 (n125[18], PSEL8, PRDATA8[18]);  // ../RTL/cmsdk_apb_slave_mux.v(217)
  and u707 (n125[19], PSEL8, PRDATA8[19]);  // ../RTL/cmsdk_apb_slave_mux.v(217)
  and u708 (n125[20], PSEL8, PRDATA8[20]);  // ../RTL/cmsdk_apb_slave_mux.v(217)
  and u709 (n125[21], PSEL8, PRDATA8[21]);  // ../RTL/cmsdk_apb_slave_mux.v(217)
  and u71 (n51, dec[8], n50);  // ../RTL/cmsdk_apb_slave_mux.v(183)
  and u710 (n125[22], PSEL8, PRDATA8[22]);  // ../RTL/cmsdk_apb_slave_mux.v(217)
  and u711 (n125[23], PSEL8, PRDATA8[23]);  // ../RTL/cmsdk_apb_slave_mux.v(217)
  and u712 (n125[24], PSEL8, PRDATA8[24]);  // ../RTL/cmsdk_apb_slave_mux.v(217)
  and u713 (n125[25], PSEL8, PRDATA8[25]);  // ../RTL/cmsdk_apb_slave_mux.v(217)
  and u714 (n125[26], PSEL8, PRDATA8[26]);  // ../RTL/cmsdk_apb_slave_mux.v(217)
  and u715 (n125[27], PSEL8, PRDATA8[27]);  // ../RTL/cmsdk_apb_slave_mux.v(217)
  and u716 (n125[28], PSEL8, PRDATA8[28]);  // ../RTL/cmsdk_apb_slave_mux.v(217)
  and u717 (n125[29], PSEL8, PRDATA8[29]);  // ../RTL/cmsdk_apb_slave_mux.v(217)
  and u718 (n125[30], PSEL8, PRDATA8[30]);  // ../RTL/cmsdk_apb_slave_mux.v(217)
  and u719 (n125[31], PSEL8, PRDATA8[31]);  // ../RTL/cmsdk_apb_slave_mux.v(217)
  or u72 (n52, n48, n51);  // ../RTL/cmsdk_apb_slave_mux.v(183)
  or u720 (n124[1], n122[1], n123[1]);  // ../RTL/cmsdk_apb_slave_mux.v(216)
  or u721 (n124[2], n122[2], n123[2]);  // ../RTL/cmsdk_apb_slave_mux.v(216)
  or u722 (n124[3], n122[3], n123[3]);  // ../RTL/cmsdk_apb_slave_mux.v(216)
  or u723 (n124[4], n122[4], n123[4]);  // ../RTL/cmsdk_apb_slave_mux.v(216)
  or u724 (n124[5], n122[5], n123[5]);  // ../RTL/cmsdk_apb_slave_mux.v(216)
  or u725 (n124[6], n122[6], n123[6]);  // ../RTL/cmsdk_apb_slave_mux.v(216)
  or u726 (n124[7], n122[7], n123[7]);  // ../RTL/cmsdk_apb_slave_mux.v(216)
  or u727 (n124[8], n122[8], n123[8]);  // ../RTL/cmsdk_apb_slave_mux.v(216)
  or u728 (n124[9], n122[9], n123[9]);  // ../RTL/cmsdk_apb_slave_mux.v(216)
  or u729 (n124[10], n122[10], n123[10]);  // ../RTL/cmsdk_apb_slave_mux.v(216)
  not u73 (n53, en[9]);  // ../RTL/cmsdk_apb_slave_mux.v(184)
  or u730 (n124[11], n122[11], n123[11]);  // ../RTL/cmsdk_apb_slave_mux.v(216)
  or u731 (n124[12], n122[12], n123[12]);  // ../RTL/cmsdk_apb_slave_mux.v(216)
  or u732 (n124[13], n122[13], n123[13]);  // ../RTL/cmsdk_apb_slave_mux.v(216)
  or u733 (n124[14], n122[14], n123[14]);  // ../RTL/cmsdk_apb_slave_mux.v(216)
  or u734 (n124[15], n122[15], n123[15]);  // ../RTL/cmsdk_apb_slave_mux.v(216)
  or u735 (n124[16], n122[16], n123[16]);  // ../RTL/cmsdk_apb_slave_mux.v(216)
  or u736 (n124[17], n122[17], n123[17]);  // ../RTL/cmsdk_apb_slave_mux.v(216)
  or u737 (n124[18], n122[18], n123[18]);  // ../RTL/cmsdk_apb_slave_mux.v(216)
  or u738 (n124[19], n122[19], n123[19]);  // ../RTL/cmsdk_apb_slave_mux.v(216)
  or u739 (n124[20], n122[20], n123[20]);  // ../RTL/cmsdk_apb_slave_mux.v(216)
  or u74 (n54, PREADY9, n53);  // ../RTL/cmsdk_apb_slave_mux.v(184)
  or u740 (n124[21], n122[21], n123[21]);  // ../RTL/cmsdk_apb_slave_mux.v(216)
  or u741 (n124[22], n122[22], n123[22]);  // ../RTL/cmsdk_apb_slave_mux.v(216)
  or u742 (n124[23], n122[23], n123[23]);  // ../RTL/cmsdk_apb_slave_mux.v(216)
  or u743 (n124[24], n122[24], n123[24]);  // ../RTL/cmsdk_apb_slave_mux.v(216)
  or u744 (n124[25], n122[25], n123[25]);  // ../RTL/cmsdk_apb_slave_mux.v(216)
  or u745 (n124[26], n122[26], n123[26]);  // ../RTL/cmsdk_apb_slave_mux.v(216)
  or u746 (n124[27], n122[27], n123[27]);  // ../RTL/cmsdk_apb_slave_mux.v(216)
  or u747 (n124[28], n122[28], n123[28]);  // ../RTL/cmsdk_apb_slave_mux.v(216)
  or u748 (n124[29], n122[29], n123[29]);  // ../RTL/cmsdk_apb_slave_mux.v(216)
  or u749 (n124[30], n122[30], n123[30]);  // ../RTL/cmsdk_apb_slave_mux.v(216)
  and u75 (n55, dec[9], n54);  // ../RTL/cmsdk_apb_slave_mux.v(184)
  or u750 (n124[31], n122[31], n123[31]);  // ../RTL/cmsdk_apb_slave_mux.v(216)
  and u751 (n123[1], PSEL7, PRDATA7[1]);  // ../RTL/cmsdk_apb_slave_mux.v(216)
  and u752 (n123[2], PSEL7, PRDATA7[2]);  // ../RTL/cmsdk_apb_slave_mux.v(216)
  and u753 (n123[3], PSEL7, PRDATA7[3]);  // ../RTL/cmsdk_apb_slave_mux.v(216)
  and u754 (n123[4], PSEL7, PRDATA7[4]);  // ../RTL/cmsdk_apb_slave_mux.v(216)
  and u755 (n123[5], PSEL7, PRDATA7[5]);  // ../RTL/cmsdk_apb_slave_mux.v(216)
  and u756 (n123[6], PSEL7, PRDATA7[6]);  // ../RTL/cmsdk_apb_slave_mux.v(216)
  and u757 (n123[7], PSEL7, PRDATA7[7]);  // ../RTL/cmsdk_apb_slave_mux.v(216)
  and u758 (n123[8], PSEL7, PRDATA7[8]);  // ../RTL/cmsdk_apb_slave_mux.v(216)
  and u759 (n123[9], PSEL7, PRDATA7[9]);  // ../RTL/cmsdk_apb_slave_mux.v(216)
  or u76 (n56, n52, n55);  // ../RTL/cmsdk_apb_slave_mux.v(184)
  and u760 (n123[10], PSEL7, PRDATA7[10]);  // ../RTL/cmsdk_apb_slave_mux.v(216)
  and u761 (n123[11], PSEL7, PRDATA7[11]);  // ../RTL/cmsdk_apb_slave_mux.v(216)
  and u762 (n123[12], PSEL7, PRDATA7[12]);  // ../RTL/cmsdk_apb_slave_mux.v(216)
  and u763 (n123[13], PSEL7, PRDATA7[13]);  // ../RTL/cmsdk_apb_slave_mux.v(216)
  and u764 (n123[14], PSEL7, PRDATA7[14]);  // ../RTL/cmsdk_apb_slave_mux.v(216)
  and u765 (n123[15], PSEL7, PRDATA7[15]);  // ../RTL/cmsdk_apb_slave_mux.v(216)
  and u766 (n123[16], PSEL7, PRDATA7[16]);  // ../RTL/cmsdk_apb_slave_mux.v(216)
  and u767 (n123[17], PSEL7, PRDATA7[17]);  // ../RTL/cmsdk_apb_slave_mux.v(216)
  and u768 (n123[18], PSEL7, PRDATA7[18]);  // ../RTL/cmsdk_apb_slave_mux.v(216)
  and u769 (n123[19], PSEL7, PRDATA7[19]);  // ../RTL/cmsdk_apb_slave_mux.v(216)
  not u77 (n57, en[10]);  // ../RTL/cmsdk_apb_slave_mux.v(185)
  and u770 (n123[20], PSEL7, PRDATA7[20]);  // ../RTL/cmsdk_apb_slave_mux.v(216)
  and u771 (n123[21], PSEL7, PRDATA7[21]);  // ../RTL/cmsdk_apb_slave_mux.v(216)
  and u772 (n123[22], PSEL7, PRDATA7[22]);  // ../RTL/cmsdk_apb_slave_mux.v(216)
  and u773 (n123[23], PSEL7, PRDATA7[23]);  // ../RTL/cmsdk_apb_slave_mux.v(216)
  and u774 (n123[24], PSEL7, PRDATA7[24]);  // ../RTL/cmsdk_apb_slave_mux.v(216)
  and u775 (n123[25], PSEL7, PRDATA7[25]);  // ../RTL/cmsdk_apb_slave_mux.v(216)
  and u776 (n123[26], PSEL7, PRDATA7[26]);  // ../RTL/cmsdk_apb_slave_mux.v(216)
  and u777 (n123[27], PSEL7, PRDATA7[27]);  // ../RTL/cmsdk_apb_slave_mux.v(216)
  and u778 (n123[28], PSEL7, PRDATA7[28]);  // ../RTL/cmsdk_apb_slave_mux.v(216)
  and u779 (n123[29], PSEL7, PRDATA7[29]);  // ../RTL/cmsdk_apb_slave_mux.v(216)
  or u78 (n58, PREADY10, n57);  // ../RTL/cmsdk_apb_slave_mux.v(185)
  and u780 (n123[30], PSEL7, PRDATA7[30]);  // ../RTL/cmsdk_apb_slave_mux.v(216)
  and u781 (n123[31], PSEL7, PRDATA7[31]);  // ../RTL/cmsdk_apb_slave_mux.v(216)
  or u782 (n122[1], n120[1], n121[1]);  // ../RTL/cmsdk_apb_slave_mux.v(215)
  or u783 (n122[2], n120[2], n121[2]);  // ../RTL/cmsdk_apb_slave_mux.v(215)
  or u784 (n122[3], n120[3], n121[3]);  // ../RTL/cmsdk_apb_slave_mux.v(215)
  or u785 (n122[4], n120[4], n121[4]);  // ../RTL/cmsdk_apb_slave_mux.v(215)
  or u786 (n122[5], n120[5], n121[5]);  // ../RTL/cmsdk_apb_slave_mux.v(215)
  or u787 (n122[6], n120[6], n121[6]);  // ../RTL/cmsdk_apb_slave_mux.v(215)
  or u788 (n122[7], n120[7], n121[7]);  // ../RTL/cmsdk_apb_slave_mux.v(215)
  or u789 (n122[8], n120[8], n121[8]);  // ../RTL/cmsdk_apb_slave_mux.v(215)
  and u79 (n59, dec[10], n58);  // ../RTL/cmsdk_apb_slave_mux.v(185)
  or u790 (n122[9], n120[9], n121[9]);  // ../RTL/cmsdk_apb_slave_mux.v(215)
  or u791 (n122[10], n120[10], n121[10]);  // ../RTL/cmsdk_apb_slave_mux.v(215)
  or u792 (n122[11], n120[11], n121[11]);  // ../RTL/cmsdk_apb_slave_mux.v(215)
  or u793 (n122[12], n120[12], n121[12]);  // ../RTL/cmsdk_apb_slave_mux.v(215)
  or u794 (n122[13], n120[13], n121[13]);  // ../RTL/cmsdk_apb_slave_mux.v(215)
  or u795 (n122[14], n120[14], n121[14]);  // ../RTL/cmsdk_apb_slave_mux.v(215)
  or u796 (n122[15], n120[15], n121[15]);  // ../RTL/cmsdk_apb_slave_mux.v(215)
  or u797 (n122[16], n120[16], n121[16]);  // ../RTL/cmsdk_apb_slave_mux.v(215)
  or u798 (n122[17], n120[17], n121[17]);  // ../RTL/cmsdk_apb_slave_mux.v(215)
  or u799 (n122[18], n120[18], n121[18]);  // ../RTL/cmsdk_apb_slave_mux.v(215)
  and u8 (n2, PSEL, dec[2]);  // ../RTL/cmsdk_apb_slave_mux.v(159)
  or u80 (n60, n56, n59);  // ../RTL/cmsdk_apb_slave_mux.v(185)
  or u800 (n122[19], n120[19], n121[19]);  // ../RTL/cmsdk_apb_slave_mux.v(215)
  or u801 (n122[20], n120[20], n121[20]);  // ../RTL/cmsdk_apb_slave_mux.v(215)
  or u802 (n122[21], n120[21], n121[21]);  // ../RTL/cmsdk_apb_slave_mux.v(215)
  or u803 (n122[22], n120[22], n121[22]);  // ../RTL/cmsdk_apb_slave_mux.v(215)
  or u804 (n122[23], n120[23], n121[23]);  // ../RTL/cmsdk_apb_slave_mux.v(215)
  or u805 (n122[24], n120[24], n121[24]);  // ../RTL/cmsdk_apb_slave_mux.v(215)
  or u806 (n122[25], n120[25], n121[25]);  // ../RTL/cmsdk_apb_slave_mux.v(215)
  or u807 (n122[26], n120[26], n121[26]);  // ../RTL/cmsdk_apb_slave_mux.v(215)
  or u808 (n122[27], n120[27], n121[27]);  // ../RTL/cmsdk_apb_slave_mux.v(215)
  or u809 (n122[28], n120[28], n121[28]);  // ../RTL/cmsdk_apb_slave_mux.v(215)
  not u81 (n61, en[11]);  // ../RTL/cmsdk_apb_slave_mux.v(186)
  or u810 (n122[29], n120[29], n121[29]);  // ../RTL/cmsdk_apb_slave_mux.v(215)
  or u811 (n122[30], n120[30], n121[30]);  // ../RTL/cmsdk_apb_slave_mux.v(215)
  or u812 (n122[31], n120[31], n121[31]);  // ../RTL/cmsdk_apb_slave_mux.v(215)
  and u813 (n121[1], PSEL6, PRDATA6[1]);  // ../RTL/cmsdk_apb_slave_mux.v(215)
  and u814 (n121[2], PSEL6, PRDATA6[2]);  // ../RTL/cmsdk_apb_slave_mux.v(215)
  and u815 (n121[3], PSEL6, PRDATA6[3]);  // ../RTL/cmsdk_apb_slave_mux.v(215)
  and u816 (n121[4], PSEL6, PRDATA6[4]);  // ../RTL/cmsdk_apb_slave_mux.v(215)
  and u817 (n121[5], PSEL6, PRDATA6[5]);  // ../RTL/cmsdk_apb_slave_mux.v(215)
  and u818 (n121[6], PSEL6, PRDATA6[6]);  // ../RTL/cmsdk_apb_slave_mux.v(215)
  and u819 (n121[7], PSEL6, PRDATA6[7]);  // ../RTL/cmsdk_apb_slave_mux.v(215)
  or u82 (n62, PREADY11, n61);  // ../RTL/cmsdk_apb_slave_mux.v(186)
  and u820 (n121[8], PSEL6, PRDATA6[8]);  // ../RTL/cmsdk_apb_slave_mux.v(215)
  and u821 (n121[9], PSEL6, PRDATA6[9]);  // ../RTL/cmsdk_apb_slave_mux.v(215)
  and u822 (n121[10], PSEL6, PRDATA6[10]);  // ../RTL/cmsdk_apb_slave_mux.v(215)
  and u823 (n121[11], PSEL6, PRDATA6[11]);  // ../RTL/cmsdk_apb_slave_mux.v(215)
  and u824 (n121[12], PSEL6, PRDATA6[12]);  // ../RTL/cmsdk_apb_slave_mux.v(215)
  and u825 (n121[13], PSEL6, PRDATA6[13]);  // ../RTL/cmsdk_apb_slave_mux.v(215)
  and u826 (n121[14], PSEL6, PRDATA6[14]);  // ../RTL/cmsdk_apb_slave_mux.v(215)
  and u827 (n121[15], PSEL6, PRDATA6[15]);  // ../RTL/cmsdk_apb_slave_mux.v(215)
  and u828 (n121[16], PSEL6, PRDATA6[16]);  // ../RTL/cmsdk_apb_slave_mux.v(215)
  and u829 (n121[17], PSEL6, PRDATA6[17]);  // ../RTL/cmsdk_apb_slave_mux.v(215)
  and u83 (n63, dec[11], n62);  // ../RTL/cmsdk_apb_slave_mux.v(186)
  and u830 (n121[18], PSEL6, PRDATA6[18]);  // ../RTL/cmsdk_apb_slave_mux.v(215)
  and u831 (n121[19], PSEL6, PRDATA6[19]);  // ../RTL/cmsdk_apb_slave_mux.v(215)
  and u832 (n121[20], PSEL6, PRDATA6[20]);  // ../RTL/cmsdk_apb_slave_mux.v(215)
  and u833 (n121[21], PSEL6, PRDATA6[21]);  // ../RTL/cmsdk_apb_slave_mux.v(215)
  and u834 (n121[22], PSEL6, PRDATA6[22]);  // ../RTL/cmsdk_apb_slave_mux.v(215)
  and u835 (n121[23], PSEL6, PRDATA6[23]);  // ../RTL/cmsdk_apb_slave_mux.v(215)
  and u836 (n121[24], PSEL6, PRDATA6[24]);  // ../RTL/cmsdk_apb_slave_mux.v(215)
  and u837 (n121[25], PSEL6, PRDATA6[25]);  // ../RTL/cmsdk_apb_slave_mux.v(215)
  and u838 (n121[26], PSEL6, PRDATA6[26]);  // ../RTL/cmsdk_apb_slave_mux.v(215)
  and u839 (n121[27], PSEL6, PRDATA6[27]);  // ../RTL/cmsdk_apb_slave_mux.v(215)
  or u84 (n64, n60, n63);  // ../RTL/cmsdk_apb_slave_mux.v(186)
  and u840 (n121[28], PSEL6, PRDATA6[28]);  // ../RTL/cmsdk_apb_slave_mux.v(215)
  and u841 (n121[29], PSEL6, PRDATA6[29]);  // ../RTL/cmsdk_apb_slave_mux.v(215)
  and u842 (n121[30], PSEL6, PRDATA6[30]);  // ../RTL/cmsdk_apb_slave_mux.v(215)
  and u843 (n121[31], PSEL6, PRDATA6[31]);  // ../RTL/cmsdk_apb_slave_mux.v(215)
  or u844 (n120[1], n118[1], n119[1]);  // ../RTL/cmsdk_apb_slave_mux.v(214)
  or u845 (n120[2], n118[2], n119[2]);  // ../RTL/cmsdk_apb_slave_mux.v(214)
  or u846 (n120[3], n118[3], n119[3]);  // ../RTL/cmsdk_apb_slave_mux.v(214)
  or u847 (n120[4], n118[4], n119[4]);  // ../RTL/cmsdk_apb_slave_mux.v(214)
  or u848 (n120[5], n118[5], n119[5]);  // ../RTL/cmsdk_apb_slave_mux.v(214)
  or u849 (n120[6], n118[6], n119[6]);  // ../RTL/cmsdk_apb_slave_mux.v(214)
  not u85 (n65, en[12]);  // ../RTL/cmsdk_apb_slave_mux.v(187)
  or u850 (n120[7], n118[7], n119[7]);  // ../RTL/cmsdk_apb_slave_mux.v(214)
  or u851 (n120[8], n118[8], n119[8]);  // ../RTL/cmsdk_apb_slave_mux.v(214)
  or u852 (n120[9], n118[9], n119[9]);  // ../RTL/cmsdk_apb_slave_mux.v(214)
  or u853 (n120[10], n118[10], n119[10]);  // ../RTL/cmsdk_apb_slave_mux.v(214)
  or u854 (n120[11], n118[11], n119[11]);  // ../RTL/cmsdk_apb_slave_mux.v(214)
  or u855 (n120[12], n118[12], n119[12]);  // ../RTL/cmsdk_apb_slave_mux.v(214)
  or u856 (n120[13], n118[13], n119[13]);  // ../RTL/cmsdk_apb_slave_mux.v(214)
  or u857 (n120[14], n118[14], n119[14]);  // ../RTL/cmsdk_apb_slave_mux.v(214)
  or u858 (n120[15], n118[15], n119[15]);  // ../RTL/cmsdk_apb_slave_mux.v(214)
  or u859 (n120[16], n118[16], n119[16]);  // ../RTL/cmsdk_apb_slave_mux.v(214)
  or u86 (n66, PREADY12, n65);  // ../RTL/cmsdk_apb_slave_mux.v(187)
  or u860 (n120[17], n118[17], n119[17]);  // ../RTL/cmsdk_apb_slave_mux.v(214)
  or u861 (n120[18], n118[18], n119[18]);  // ../RTL/cmsdk_apb_slave_mux.v(214)
  or u862 (n120[19], n118[19], n119[19]);  // ../RTL/cmsdk_apb_slave_mux.v(214)
  or u863 (n120[20], n118[20], n119[20]);  // ../RTL/cmsdk_apb_slave_mux.v(214)
  or u864 (n120[21], n118[21], n119[21]);  // ../RTL/cmsdk_apb_slave_mux.v(214)
  or u865 (n120[22], n118[22], n119[22]);  // ../RTL/cmsdk_apb_slave_mux.v(214)
  or u866 (n120[23], n118[23], n119[23]);  // ../RTL/cmsdk_apb_slave_mux.v(214)
  or u867 (n120[24], n118[24], n119[24]);  // ../RTL/cmsdk_apb_slave_mux.v(214)
  or u868 (n120[25], n118[25], n119[25]);  // ../RTL/cmsdk_apb_slave_mux.v(214)
  or u869 (n120[26], n118[26], n119[26]);  // ../RTL/cmsdk_apb_slave_mux.v(214)
  and u87 (n67, dec[12], n66);  // ../RTL/cmsdk_apb_slave_mux.v(187)
  or u870 (n120[27], n118[27], n119[27]);  // ../RTL/cmsdk_apb_slave_mux.v(214)
  or u871 (n120[28], n118[28], n119[28]);  // ../RTL/cmsdk_apb_slave_mux.v(214)
  or u872 (n120[29], n118[29], n119[29]);  // ../RTL/cmsdk_apb_slave_mux.v(214)
  or u873 (n120[30], n118[30], n119[30]);  // ../RTL/cmsdk_apb_slave_mux.v(214)
  or u874 (n120[31], n118[31], n119[31]);  // ../RTL/cmsdk_apb_slave_mux.v(214)
  and u875 (n119[1], PSEL5, PRDATA5[1]);  // ../RTL/cmsdk_apb_slave_mux.v(214)
  and u876 (n119[2], PSEL5, PRDATA5[2]);  // ../RTL/cmsdk_apb_slave_mux.v(214)
  and u877 (n119[3], PSEL5, PRDATA5[3]);  // ../RTL/cmsdk_apb_slave_mux.v(214)
  and u878 (n119[4], PSEL5, PRDATA5[4]);  // ../RTL/cmsdk_apb_slave_mux.v(214)
  and u879 (n119[5], PSEL5, PRDATA5[5]);  // ../RTL/cmsdk_apb_slave_mux.v(214)
  or u88 (n68, n64, n67);  // ../RTL/cmsdk_apb_slave_mux.v(187)
  and u880 (n119[6], PSEL5, PRDATA5[6]);  // ../RTL/cmsdk_apb_slave_mux.v(214)
  and u881 (n119[7], PSEL5, PRDATA5[7]);  // ../RTL/cmsdk_apb_slave_mux.v(214)
  and u882 (n119[8], PSEL5, PRDATA5[8]);  // ../RTL/cmsdk_apb_slave_mux.v(214)
  and u883 (n119[9], PSEL5, PRDATA5[9]);  // ../RTL/cmsdk_apb_slave_mux.v(214)
  and u884 (n119[10], PSEL5, PRDATA5[10]);  // ../RTL/cmsdk_apb_slave_mux.v(214)
  and u885 (n119[11], PSEL5, PRDATA5[11]);  // ../RTL/cmsdk_apb_slave_mux.v(214)
  and u886 (n119[12], PSEL5, PRDATA5[12]);  // ../RTL/cmsdk_apb_slave_mux.v(214)
  and u887 (n119[13], PSEL5, PRDATA5[13]);  // ../RTL/cmsdk_apb_slave_mux.v(214)
  and u888 (n119[14], PSEL5, PRDATA5[14]);  // ../RTL/cmsdk_apb_slave_mux.v(214)
  and u889 (n119[15], PSEL5, PRDATA5[15]);  // ../RTL/cmsdk_apb_slave_mux.v(214)
  not u89 (n69, en[13]);  // ../RTL/cmsdk_apb_slave_mux.v(188)
  and u890 (n119[16], PSEL5, PRDATA5[16]);  // ../RTL/cmsdk_apb_slave_mux.v(214)
  and u891 (n119[17], PSEL5, PRDATA5[17]);  // ../RTL/cmsdk_apb_slave_mux.v(214)
  and u892 (n119[18], PSEL5, PRDATA5[18]);  // ../RTL/cmsdk_apb_slave_mux.v(214)
  and u893 (n119[19], PSEL5, PRDATA5[19]);  // ../RTL/cmsdk_apb_slave_mux.v(214)
  and u894 (n119[20], PSEL5, PRDATA5[20]);  // ../RTL/cmsdk_apb_slave_mux.v(214)
  and u895 (n119[21], PSEL5, PRDATA5[21]);  // ../RTL/cmsdk_apb_slave_mux.v(214)
  and u896 (n119[22], PSEL5, PRDATA5[22]);  // ../RTL/cmsdk_apb_slave_mux.v(214)
  and u897 (n119[23], PSEL5, PRDATA5[23]);  // ../RTL/cmsdk_apb_slave_mux.v(214)
  and u898 (n119[24], PSEL5, PRDATA5[24]);  // ../RTL/cmsdk_apb_slave_mux.v(214)
  and u899 (n119[25], PSEL5, PRDATA5[25]);  // ../RTL/cmsdk_apb_slave_mux.v(214)
  and u9 (PSEL2, n2, en[2]);  // ../RTL/cmsdk_apb_slave_mux.v(159)
  or u90 (n70, PREADY13, n69);  // ../RTL/cmsdk_apb_slave_mux.v(188)
  and u900 (n119[26], PSEL5, PRDATA5[26]);  // ../RTL/cmsdk_apb_slave_mux.v(214)
  and u901 (n119[27], PSEL5, PRDATA5[27]);  // ../RTL/cmsdk_apb_slave_mux.v(214)
  and u902 (n119[28], PSEL5, PRDATA5[28]);  // ../RTL/cmsdk_apb_slave_mux.v(214)
  and u903 (n119[29], PSEL5, PRDATA5[29]);  // ../RTL/cmsdk_apb_slave_mux.v(214)
  and u904 (n119[30], PSEL5, PRDATA5[30]);  // ../RTL/cmsdk_apb_slave_mux.v(214)
  and u905 (n119[31], PSEL5, PRDATA5[31]);  // ../RTL/cmsdk_apb_slave_mux.v(214)
  or u906 (n118[1], n116[1], n117[1]);  // ../RTL/cmsdk_apb_slave_mux.v(213)
  or u907 (n118[2], n116[2], n117[2]);  // ../RTL/cmsdk_apb_slave_mux.v(213)
  or u908 (n118[3], n116[3], n117[3]);  // ../RTL/cmsdk_apb_slave_mux.v(213)
  or u909 (n118[4], n116[4], n117[4]);  // ../RTL/cmsdk_apb_slave_mux.v(213)
  and u91 (n71, dec[13], n70);  // ../RTL/cmsdk_apb_slave_mux.v(188)
  or u910 (n118[5], n116[5], n117[5]);  // ../RTL/cmsdk_apb_slave_mux.v(213)
  or u911 (n118[6], n116[6], n117[6]);  // ../RTL/cmsdk_apb_slave_mux.v(213)
  or u912 (n118[7], n116[7], n117[7]);  // ../RTL/cmsdk_apb_slave_mux.v(213)
  or u913 (n118[8], n116[8], n117[8]);  // ../RTL/cmsdk_apb_slave_mux.v(213)
  or u914 (n118[9], n116[9], n117[9]);  // ../RTL/cmsdk_apb_slave_mux.v(213)
  or u915 (n118[10], n116[10], n117[10]);  // ../RTL/cmsdk_apb_slave_mux.v(213)
  or u916 (n118[11], n116[11], n117[11]);  // ../RTL/cmsdk_apb_slave_mux.v(213)
  or u917 (n118[12], n116[12], n117[12]);  // ../RTL/cmsdk_apb_slave_mux.v(213)
  or u918 (n118[13], n116[13], n117[13]);  // ../RTL/cmsdk_apb_slave_mux.v(213)
  or u919 (n118[14], n116[14], n117[14]);  // ../RTL/cmsdk_apb_slave_mux.v(213)
  or u92 (n72, n68, n71);  // ../RTL/cmsdk_apb_slave_mux.v(188)
  or u920 (n118[15], n116[15], n117[15]);  // ../RTL/cmsdk_apb_slave_mux.v(213)
  or u921 (n118[16], n116[16], n117[16]);  // ../RTL/cmsdk_apb_slave_mux.v(213)
  or u922 (n118[17], n116[17], n117[17]);  // ../RTL/cmsdk_apb_slave_mux.v(213)
  or u923 (n118[18], n116[18], n117[18]);  // ../RTL/cmsdk_apb_slave_mux.v(213)
  or u924 (n118[19], n116[19], n117[19]);  // ../RTL/cmsdk_apb_slave_mux.v(213)
  or u925 (n118[20], n116[20], n117[20]);  // ../RTL/cmsdk_apb_slave_mux.v(213)
  or u926 (n118[21], n116[21], n117[21]);  // ../RTL/cmsdk_apb_slave_mux.v(213)
  or u927 (n118[22], n116[22], n117[22]);  // ../RTL/cmsdk_apb_slave_mux.v(213)
  or u928 (n118[23], n116[23], n117[23]);  // ../RTL/cmsdk_apb_slave_mux.v(213)
  or u929 (n118[24], n116[24], n117[24]);  // ../RTL/cmsdk_apb_slave_mux.v(213)
  not u93 (n73, en[14]);  // ../RTL/cmsdk_apb_slave_mux.v(189)
  or u930 (n118[25], n116[25], n117[25]);  // ../RTL/cmsdk_apb_slave_mux.v(213)
  or u931 (n118[26], n116[26], n117[26]);  // ../RTL/cmsdk_apb_slave_mux.v(213)
  or u932 (n118[27], n116[27], n117[27]);  // ../RTL/cmsdk_apb_slave_mux.v(213)
  or u933 (n118[28], n116[28], n117[28]);  // ../RTL/cmsdk_apb_slave_mux.v(213)
  or u934 (n118[29], n116[29], n117[29]);  // ../RTL/cmsdk_apb_slave_mux.v(213)
  or u935 (n118[30], n116[30], n117[30]);  // ../RTL/cmsdk_apb_slave_mux.v(213)
  or u936 (n118[31], n116[31], n117[31]);  // ../RTL/cmsdk_apb_slave_mux.v(213)
  and u937 (n117[1], PSEL4, PRDATA4[1]);  // ../RTL/cmsdk_apb_slave_mux.v(213)
  and u938 (n117[2], PSEL4, PRDATA4[2]);  // ../RTL/cmsdk_apb_slave_mux.v(213)
  and u939 (n117[3], PSEL4, PRDATA4[3]);  // ../RTL/cmsdk_apb_slave_mux.v(213)
  or u94 (n74, PREADY14, n73);  // ../RTL/cmsdk_apb_slave_mux.v(189)
  and u940 (n117[4], PSEL4, PRDATA4[4]);  // ../RTL/cmsdk_apb_slave_mux.v(213)
  and u941 (n117[5], PSEL4, PRDATA4[5]);  // ../RTL/cmsdk_apb_slave_mux.v(213)
  and u942 (n117[6], PSEL4, PRDATA4[6]);  // ../RTL/cmsdk_apb_slave_mux.v(213)
  and u943 (n117[7], PSEL4, PRDATA4[7]);  // ../RTL/cmsdk_apb_slave_mux.v(213)
  and u944 (n117[8], PSEL4, PRDATA4[8]);  // ../RTL/cmsdk_apb_slave_mux.v(213)
  and u945 (n117[9], PSEL4, PRDATA4[9]);  // ../RTL/cmsdk_apb_slave_mux.v(213)
  and u946 (n117[10], PSEL4, PRDATA4[10]);  // ../RTL/cmsdk_apb_slave_mux.v(213)
  and u947 (n117[11], PSEL4, PRDATA4[11]);  // ../RTL/cmsdk_apb_slave_mux.v(213)
  and u948 (n117[12], PSEL4, PRDATA4[12]);  // ../RTL/cmsdk_apb_slave_mux.v(213)
  and u949 (n117[13], PSEL4, PRDATA4[13]);  // ../RTL/cmsdk_apb_slave_mux.v(213)
  and u95 (n75, dec[14], n74);  // ../RTL/cmsdk_apb_slave_mux.v(189)
  and u950 (n117[14], PSEL4, PRDATA4[14]);  // ../RTL/cmsdk_apb_slave_mux.v(213)
  and u951 (n117[15], PSEL4, PRDATA4[15]);  // ../RTL/cmsdk_apb_slave_mux.v(213)
  and u952 (n117[16], PSEL4, PRDATA4[16]);  // ../RTL/cmsdk_apb_slave_mux.v(213)
  and u953 (n117[17], PSEL4, PRDATA4[17]);  // ../RTL/cmsdk_apb_slave_mux.v(213)
  and u954 (n117[18], PSEL4, PRDATA4[18]);  // ../RTL/cmsdk_apb_slave_mux.v(213)
  and u955 (n117[19], PSEL4, PRDATA4[19]);  // ../RTL/cmsdk_apb_slave_mux.v(213)
  and u956 (n117[20], PSEL4, PRDATA4[20]);  // ../RTL/cmsdk_apb_slave_mux.v(213)
  and u957 (n117[21], PSEL4, PRDATA4[21]);  // ../RTL/cmsdk_apb_slave_mux.v(213)
  and u958 (n117[22], PSEL4, PRDATA4[22]);  // ../RTL/cmsdk_apb_slave_mux.v(213)
  and u959 (n117[23], PSEL4, PRDATA4[23]);  // ../RTL/cmsdk_apb_slave_mux.v(213)
  or u96 (n76, n72, n75);  // ../RTL/cmsdk_apb_slave_mux.v(189)
  and u960 (n117[24], PSEL4, PRDATA4[24]);  // ../RTL/cmsdk_apb_slave_mux.v(213)
  and u961 (n117[25], PSEL4, PRDATA4[25]);  // ../RTL/cmsdk_apb_slave_mux.v(213)
  and u962 (n117[26], PSEL4, PRDATA4[26]);  // ../RTL/cmsdk_apb_slave_mux.v(213)
  and u963 (n117[27], PSEL4, PRDATA4[27]);  // ../RTL/cmsdk_apb_slave_mux.v(213)
  and u964 (n117[28], PSEL4, PRDATA4[28]);  // ../RTL/cmsdk_apb_slave_mux.v(213)
  and u965 (n117[29], PSEL4, PRDATA4[29]);  // ../RTL/cmsdk_apb_slave_mux.v(213)
  and u966 (n117[30], PSEL4, PRDATA4[30]);  // ../RTL/cmsdk_apb_slave_mux.v(213)
  and u967 (n117[31], PSEL4, PRDATA4[31]);  // ../RTL/cmsdk_apb_slave_mux.v(213)
  or u968 (n116[1], n114[1], n115[1]);  // ../RTL/cmsdk_apb_slave_mux.v(212)
  or u969 (n116[2], n114[2], n115[2]);  // ../RTL/cmsdk_apb_slave_mux.v(212)
  not u97 (n77, en[15]);  // ../RTL/cmsdk_apb_slave_mux.v(190)
  or u970 (n116[3], n114[3], n115[3]);  // ../RTL/cmsdk_apb_slave_mux.v(212)
  or u971 (n116[4], n114[4], n115[4]);  // ../RTL/cmsdk_apb_slave_mux.v(212)
  or u972 (n116[5], n114[5], n115[5]);  // ../RTL/cmsdk_apb_slave_mux.v(212)
  or u973 (n116[6], n114[6], n115[6]);  // ../RTL/cmsdk_apb_slave_mux.v(212)
  or u974 (n116[7], n114[7], n115[7]);  // ../RTL/cmsdk_apb_slave_mux.v(212)
  or u975 (n116[8], n114[8], n115[8]);  // ../RTL/cmsdk_apb_slave_mux.v(212)
  or u976 (n116[9], n114[9], n115[9]);  // ../RTL/cmsdk_apb_slave_mux.v(212)
  or u977 (n116[10], n114[10], n115[10]);  // ../RTL/cmsdk_apb_slave_mux.v(212)
  or u978 (n116[11], n114[11], n115[11]);  // ../RTL/cmsdk_apb_slave_mux.v(212)
  or u979 (n116[12], n114[12], n115[12]);  // ../RTL/cmsdk_apb_slave_mux.v(212)
  or u98 (n78, PREADY15, n77);  // ../RTL/cmsdk_apb_slave_mux.v(190)
  or u980 (n116[13], n114[13], n115[13]);  // ../RTL/cmsdk_apb_slave_mux.v(212)
  or u981 (n116[14], n114[14], n115[14]);  // ../RTL/cmsdk_apb_slave_mux.v(212)
  or u982 (n116[15], n114[15], n115[15]);  // ../RTL/cmsdk_apb_slave_mux.v(212)
  or u983 (n116[16], n114[16], n115[16]);  // ../RTL/cmsdk_apb_slave_mux.v(212)
  or u984 (n116[17], n114[17], n115[17]);  // ../RTL/cmsdk_apb_slave_mux.v(212)
  or u985 (n116[18], n114[18], n115[18]);  // ../RTL/cmsdk_apb_slave_mux.v(212)
  or u986 (n116[19], n114[19], n115[19]);  // ../RTL/cmsdk_apb_slave_mux.v(212)
  or u987 (n116[20], n114[20], n115[20]);  // ../RTL/cmsdk_apb_slave_mux.v(212)
  or u988 (n116[21], n114[21], n115[21]);  // ../RTL/cmsdk_apb_slave_mux.v(212)
  or u989 (n116[22], n114[22], n115[22]);  // ../RTL/cmsdk_apb_slave_mux.v(212)
  and u99 (n79, dec[15], n78);  // ../RTL/cmsdk_apb_slave_mux.v(190)
  or u990 (n116[23], n114[23], n115[23]);  // ../RTL/cmsdk_apb_slave_mux.v(212)
  or u991 (n116[24], n114[24], n115[24]);  // ../RTL/cmsdk_apb_slave_mux.v(212)
  or u992 (n116[25], n114[25], n115[25]);  // ../RTL/cmsdk_apb_slave_mux.v(212)
  or u993 (n116[26], n114[26], n115[26]);  // ../RTL/cmsdk_apb_slave_mux.v(212)
  or u994 (n116[27], n114[27], n115[27]);  // ../RTL/cmsdk_apb_slave_mux.v(212)
  or u995 (n116[28], n114[28], n115[28]);  // ../RTL/cmsdk_apb_slave_mux.v(212)
  or u996 (n116[29], n114[29], n115[29]);  // ../RTL/cmsdk_apb_slave_mux.v(212)
  or u997 (n116[30], n114[30], n115[30]);  // ../RTL/cmsdk_apb_slave_mux.v(212)
  or u998 (n116[31], n114[31], n115[31]);  // ../RTL/cmsdk_apb_slave_mux.v(212)
  and u999 (n115[1], PSEL3, PRDATA3[1]);  // ../RTL/cmsdk_apb_slave_mux.v(212)

endmodule 

module eq_w18
  (
  i0,
  i1,
  o
  );

  input [17:0] i0;
  input [17:0] i1;
  output o;



endmodule 

module binary_mux_s1_w18
  (
  i0,
  i1,
  sel,
  o
  );

  input [17:0] i0;
  input [17:0] i1;
  input sel;
  output [17:0] o;



endmodule 

module reg_ar_as_w18
  (
  clk,
  d,
  en,
  reset,
  set,
  q
  );

  input clk;
  input [17:0] d;
  input en;
  input [17:0] reset;
  input [17:0] set;
  output [17:0] q;



endmodule 

module add_pu18_mu18_o18
  (
  i0,
  i1,
  o
  );

  input [17:0] i0;
  input [17:0] i1;
  output [17:0] o;



endmodule 

module eq_w10
  (
  i0,
  i1,
  o
  );

  input [9:0] i0;
  input [9:0] i1;
  output o;



endmodule 

module eq_w7
  (
  i0,
  i1,
  o
  );

  input [6:0] i0;
  input [6:0] i1;
  output o;



endmodule 

module eq_w6
  (
  i0,
  i1,
  o
  );

  input [5:0] i0;
  input [5:0] i1;
  output o;



endmodule 

module binary_mux_s1_w4
  (
  i0,
  i1,
  sel,
  o
  );

  input [3:0] i0;
  input [3:0] i1;
  input sel;
  output [3:0] o;



endmodule 

module binary_mux_s1_w3
  (
  i0,
  i1,
  sel,
  o
  );

  input [2:0] i0;
  input [2:0] i1;
  input sel;
  output [2:0] o;



endmodule 

module binary_mux_s3_w32
  (
  i0,
  i1,
  i2,
  i3,
  i4,
  i5,
  i6,
  i7,
  sel,
  o
  );

  input [31:0] i0;
  input [31:0] i1;
  input [31:0] i2;
  input [31:0] i3;
  input [31:0] i4;
  input [31:0] i5;
  input [31:0] i6;
  input [31:0] i7;
  input [2:0] sel;
  output [31:0] o;



endmodule 

module binary_mux_s4_w32
  (
  i0,
  i1,
  i10,
  i11,
  i12,
  i13,
  i14,
  i15,
  i2,
  i3,
  i4,
  i5,
  i6,
  i7,
  i8,
  i9,
  sel,
  o
  );

  input [31:0] i0;
  input [31:0] i1;
  input [31:0] i10;
  input [31:0] i11;
  input [31:0] i12;
  input [31:0] i13;
  input [31:0] i14;
  input [31:0] i15;
  input [31:0] i2;
  input [31:0] i3;
  input [31:0] i4;
  input [31:0] i5;
  input [31:0] i6;
  input [31:0] i7;
  input [31:0] i8;
  input [31:0] i9;
  input [3:0] sel;
  output [31:0] o;



endmodule 

module reg_ar_as_w4
  (
  clk,
  d,
  en,
  reset,
  set,
  q
  );

  input clk;
  input [3:0] d;
  input en;
  input [3:0] reset;
  input [3:0] set;
  output [3:0] q;



endmodule 

module cortexm0ds_logic  // ../RTL/cortexm0ds_logic.v(27)
  (
  CDBGPWRUPACK,
  DBGRESETn,
  DBGRESTART,
  DCLK,
  ECOREVNUM,
  EDBGRQ,
  FCLK,
  HCLK,
  HRDATA,
  HREADY,
  HRESETn,
  HRESP,
  IRQ,
  IRQLATENCY,
  NMI,
  PORESETn,
  RSTBYPASS,
  RXEV,
  SCLK,
  SE,
  SLEEPHOLDREQn,
  STCALIB,
  STCLKEN,
  SWCLKTCK,
  SWDITMS,
  TDI,
  WICENREQ,
  nTRST,
  CDBGPWRUPREQ,
  CODEHINTDE,
  CODENSEQ,
  DBGRESTARTED,
  GATEHCLK,
  HADDR,
  HALTED,
  HBURST,
  HMASTER,
  HMASTLOCK,
  HPROT,
  HSIZE,
  HTRANS,
  HWDATA,
  HWRITE,
  LOCKUP,
  SLEEPDEEP,
  SLEEPHOLDACKn,
  SLEEPING,
  SPECHTRANS,
  SWDO,
  SWDOEN,
  SYSRESETREQ,
  TDO,
  TXEV,
  WAKEUP,
  WICENACK,
  WICSENSE,
  nTDOEN,
  vis_apsr_o,
  vis_control_o,
  vis_ipsr_o,
  vis_msp_o,
  vis_pc_o,
  vis_primask_o,
  vis_psp_o,
  vis_r0_o,
  vis_r10_o,
  vis_r11_o,
  vis_r12_o,
  vis_r14_o,
  vis_r1_o,
  vis_r2_o,
  vis_r3_o,
  vis_r4_o,
  vis_r5_o,
  vis_r6_o,
  vis_r7_o,
  vis_r8_o,
  vis_r9_o,
  vis_tbit_o
  );

  input CDBGPWRUPACK;  // ../RTL/cortexm0ds_logic.v(92)
  input DBGRESETn;  // ../RTL/cortexm0ds_logic.v(77)
  input DBGRESTART;  // ../RTL/cortexm0ds_logic.v(85)
  input DCLK;  // ../RTL/cortexm0ds_logic.v(75)
  input [27:0] ECOREVNUM;  // ../RTL/cortexm0ds_logic.v(51)
  input EDBGRQ;  // ../RTL/cortexm0ds_logic.v(86)
  input FCLK;  // ../RTL/cortexm0ds_logic.v(72)
  input HCLK;  // ../RTL/cortexm0ds_logic.v(74)
  input [31:0] HRDATA;  // ../RTL/cortexm0ds_logic.v(46)
  input HREADY;  // ../RTL/cortexm0ds_logic.v(81)
  input HRESETn;  // ../RTL/cortexm0ds_logic.v(78)
  input HRESP;  // ../RTL/cortexm0ds_logic.v(82)
  input [31:0] IRQ;  // ../RTL/cortexm0ds_logic.v(48)
  input [7:0] IRQLATENCY;  // ../RTL/cortexm0ds_logic.v(50)
  input NMI;  // ../RTL/cortexm0ds_logic.v(87)
  input PORESETn;  // ../RTL/cortexm0ds_logic.v(76)
  input RSTBYPASS;  // ../RTL/cortexm0ds_logic.v(94)
  input RXEV;  // ../RTL/cortexm0ds_logic.v(88)
  input SCLK;  // ../RTL/cortexm0ds_logic.v(73)
  input SE;  // ../RTL/cortexm0ds_logic.v(93)
  input SLEEPHOLDREQn;  // ../RTL/cortexm0ds_logic.v(90)
  input [25:0] STCALIB;  // ../RTL/cortexm0ds_logic.v(49)
  input STCLKEN;  // ../RTL/cortexm0ds_logic.v(89)
  input SWCLKTCK;  // ../RTL/cortexm0ds_logic.v(79)
  input SWDITMS;  // ../RTL/cortexm0ds_logic.v(83)
  input TDI;  // ../RTL/cortexm0ds_logic.v(84)
  input WICENREQ;  // ../RTL/cortexm0ds_logic.v(91)
  input nTRST;  // ../RTL/cortexm0ds_logic.v(80)
  output CDBGPWRUPREQ;  // ../RTL/cortexm0ds_logic.v(115)
  output [2:0] CODEHINTDE;  // ../RTL/cortexm0ds_logic.v(47)
  output CODENSEQ;  // ../RTL/cortexm0ds_logic.v(98)
  output DBGRESTARTED;  // ../RTL/cortexm0ds_logic.v(104)
  output GATEHCLK;  // ../RTL/cortexm0ds_logic.v(109)
  output [31:0] HADDR;  // ../RTL/cortexm0ds_logic.v(40)
  output HALTED;  // ../RTL/cortexm0ds_logic.v(105)
  output [2:0] HBURST;  // ../RTL/cortexm0ds_logic.v(41)
  output HMASTER;  // ../RTL/cortexm0ds_logic.v(97)
  output HMASTLOCK;  // ../RTL/cortexm0ds_logic.v(95)
  output [3:0] HPROT;  // ../RTL/cortexm0ds_logic.v(42)
  output [2:0] HSIZE;  // ../RTL/cortexm0ds_logic.v(43)
  output [1:0] HTRANS;  // ../RTL/cortexm0ds_logic.v(44)
  output [31:0] HWDATA;  // ../RTL/cortexm0ds_logic.v(45)
  output HWRITE;  // ../RTL/cortexm0ds_logic.v(96)
  output LOCKUP;  // ../RTL/cortexm0ds_logic.v(107)
  output SLEEPDEEP;  // ../RTL/cortexm0ds_logic.v(111)
  output SLEEPHOLDACKn;  // ../RTL/cortexm0ds_logic.v(113)
  output SLEEPING;  // ../RTL/cortexm0ds_logic.v(110)
  output SPECHTRANS;  // ../RTL/cortexm0ds_logic.v(99)
  output SWDO;  // ../RTL/cortexm0ds_logic.v(100)
  output SWDOEN;  // ../RTL/cortexm0ds_logic.v(101)
  output SYSRESETREQ;  // ../RTL/cortexm0ds_logic.v(108)
  output TDO;  // ../RTL/cortexm0ds_logic.v(102)
  output TXEV;  // ../RTL/cortexm0ds_logic.v(106)
  output WAKEUP;  // ../RTL/cortexm0ds_logic.v(112)
  output WICENACK;  // ../RTL/cortexm0ds_logic.v(114)
  output [33:0] WICSENSE;  // ../RTL/cortexm0ds_logic.v(52)
  output nTDOEN;  // ../RTL/cortexm0ds_logic.v(103)
  output [3:0] vis_apsr_o;  // ../RTL/cortexm0ds_logic.v(70)
  output vis_control_o;  // ../RTL/cortexm0ds_logic.v(117)
  output [5:0] vis_ipsr_o;  // ../RTL/cortexm0ds_logic.v(71)
  output [29:0] vis_msp_o;  // ../RTL/cortexm0ds_logic.v(67)
  output [30:0] vis_pc_o;  // ../RTL/cortexm0ds_logic.v(69)
  output vis_primask_o;  // ../RTL/cortexm0ds_logic.v(118)
  output [29:0] vis_psp_o;  // ../RTL/cortexm0ds_logic.v(68)
  output [31:0] vis_r0_o;  // ../RTL/cortexm0ds_logic.v(53)
  output [31:0] vis_r10_o;  // ../RTL/cortexm0ds_logic.v(63)
  output [31:0] vis_r11_o;  // ../RTL/cortexm0ds_logic.v(64)
  output [31:0] vis_r12_o;  // ../RTL/cortexm0ds_logic.v(65)
  output [31:0] vis_r14_o;  // ../RTL/cortexm0ds_logic.v(66)
  output [31:0] vis_r1_o;  // ../RTL/cortexm0ds_logic.v(54)
  output [31:0] vis_r2_o;  // ../RTL/cortexm0ds_logic.v(55)
  output [31:0] vis_r3_o;  // ../RTL/cortexm0ds_logic.v(56)
  output [31:0] vis_r4_o;  // ../RTL/cortexm0ds_logic.v(57)
  output [31:0] vis_r5_o;  // ../RTL/cortexm0ds_logic.v(58)
  output [31:0] vis_r6_o;  // ../RTL/cortexm0ds_logic.v(59)
  output [31:0] vis_r7_o;  // ../RTL/cortexm0ds_logic.v(60)
  output [31:0] vis_r8_o;  // ../RTL/cortexm0ds_logic.v(61)
  output [31:0] vis_r9_o;  // ../RTL/cortexm0ds_logic.v(62)
  output vis_tbit_o;  // ../RTL/cortexm0ds_logic.v(116)

  wire [31:0] Affpw6;  // ../RTL/cortexm0ds_logic.v(1529)
  wire [28:27] Akgpw6;  // ../RTL/cortexm0ds_logic.v(1553)
  wire [2:1] Aphpw6;  // ../RTL/cortexm0ds_logic.v(1580)
  wire [4:0] Aygpw6;  // ../RTL/cortexm0ds_logic.v(1562)
  wire [1:0] B3gpw6;  // ../RTL/cortexm0ds_logic.v(1543)
  wire [23:0] Bagpw6;  // ../RTL/cortexm0ds_logic.v(1547)
  wire [3:0] Cjhpw6;  // ../RTL/cortexm0ds_logic.v(1576)
  wire [7:0] Cyfpw6;  // ../RTL/cortexm0ds_logic.v(1540)
  wire [15:0] D7fpw6;  // ../RTL/cortexm0ds_logic.v(1524)
  wire [4:0] Dhgpw6;  // ../RTL/cortexm0ds_logic.v(1551)
  wire [31:2] E1hpw6;  // ../RTL/cortexm0ds_logic.v(1564)
  wire [31:0] Eafpw6;  // ../RTL/cortexm0ds_logic.v(1526)
  wire [28:27] Engpw6;  // ../RTL/cortexm0ds_logic.v(1555)
  wire [31:0] Fkfpw6;  // ../RTL/cortexm0ds_logic.v(1532)
  wire [4:0] G4hpw6;  // ../RTL/cortexm0ds_logic.v(1566)
  wire [9:0] Gmhpw6;  // ../RTL/cortexm0ds_logic.v(1578)
  wire [28:2] Gqgpw6;  // ../RTL/cortexm0ds_logic.v(1557)
  wire [28:2] Gtgpw6;  // ../RTL/cortexm0ds_logic.v(1559)
  wire [3:0] H2fpw6;  // ../RTL/cortexm0ds_logic.v(1521)
  wire [1:0] H8gpw6;  // ../RTL/cortexm0ds_logic.v(1546)
  wire [16:0] Hrfpw6;  // ../RTL/cortexm0ds_logic.v(1536)
  wire [30:0] Iahpw6;  // ../RTL/cortexm0ds_logic.v(1570)
  wire [31:0] Idfpw6;  // ../RTL/cortexm0ds_logic.v(1528)
  wire [5:0] Ighpw6;  // ../RTL/cortexm0ds_logic.v(1574)
  wire [1:0] Iwfpw6;  // ../RTL/cortexm0ds_logic.v(1539)
  wire [4:0] Jfgpw6;  // ../RTL/cortexm0ds_logic.v(1550)
  wire [31:4] Jshpw6;  // ../RTL/cortexm0ds_logic.v(1582)
  wire [31:2] K7hpw6;  // ../RTL/cortexm0ds_logic.v(1568)
  wire [1:0] L1gpw6;  // ../RTL/cortexm0ds_logic.v(1542)
  wire [23:0] L6gpw6;  // ../RTL/cortexm0ds_logic.v(1545)
  wire [28:27] Ligpw6;  // ../RTL/cortexm0ds_logic.v(1552)
  wire [2:0] Lwgpw6;  // ../RTL/cortexm0ds_logic.v(1561)
  wire [3:0] Mdhpw6;  // ../RTL/cortexm0ds_logic.v(1572)
  wire [31:0] Mifpw6;  // ../RTL/cortexm0ds_logic.v(1531)
  wire [30:2] N5fpw6;  // ../RTL/cortexm0ds_logic.v(1523)
  wire [31:0] Ntkbx6;  // ../RTL/cortexm0ds_logic.v(1719)
  wire [31:0] Nvkbx6;  // ../RTL/cortexm0ds_logic.v(1720)
  wire [33:0] Nxkbx6;  // ../RTL/cortexm0ds_logic.v(1721)
  wire [31:0] Odgpw6;  // ../RTL/cortexm0ds_logic.v(1549)
  wire [33:0] Ozkbx6;  // ../RTL/cortexm0ds_logic.v(1722)
  wire [1:0] Pkhpw6;  // ../RTL/cortexm0ds_logic.v(1577)
  wire [28:27] Plgpw6;  // ../RTL/cortexm0ds_logic.v(1554)
  wire [16:0] Ppfpw6;  // ../RTL/cortexm0ds_logic.v(1535)
  wire [1:0] Pzgpw6;  // ../RTL/cortexm0ds_logic.v(1563)
  wire [30:0] Qbfpw6;  // ../RTL/cortexm0ds_logic.v(1527)
  wire [2:0] R2hpw6;  // ../RTL/cortexm0ds_logic.v(1565)
  wire [63:0] R4gpw6;  // ../RTL/cortexm0ds_logic.v(1544)
  wire [11:0] S8fpw6;  // ../RTL/cortexm0ds_logic.v(1525)
  wire [31:0] Shhpw6;  // ../RTL/cortexm0ds_logic.v(1575)
  wire [1:0] Sqhpw6;  // ../RTL/cortexm0ds_logic.v(1581)
  wire [1:0] Sufpw6;  // ../RTL/cortexm0ds_logic.v(1538)
  wire [31:0] Tgfpw6;  // ../RTL/cortexm0ds_logic.v(1530)
  wire [3:0] Tnhpw6;  // ../RTL/cortexm0ds_logic.v(1579)
  wire [28:2] Togpw6;  // ../RTL/cortexm0ds_logic.v(1556)
  wire [28:2] Trgpw6;  // ../RTL/cortexm0ds_logic.v(1558)
  wire [13:0] Tugpw6;  // ../RTL/cortexm0ds_logic.v(1560)
  wire [23:0] Tzfpw6;  // ../RTL/cortexm0ds_logic.v(1541)
  wire [31:0] Uthpw6;  // ../RTL/cortexm0ds_logic.v(1583)
  wire [1:0] V5hpw6;  // ../RTL/cortexm0ds_logic.v(1567)
  wire [31:0] Vbgpw6;  // ../RTL/cortexm0ds_logic.v(1548)
  wire [7:0] Vnfpw6;  // ../RTL/cortexm0ds_logic.v(1534)
  wire [33:0] Vrkbx6;  // ../RTL/cortexm0ds_logic.v(1718)
  wire [3:0] X3fpw6;  // ../RTL/cortexm0ds_logic.v(1522)
  wire [6:0] X8hpw6;  // ../RTL/cortexm0ds_logic.v(1569)
  wire [8:1] Xlfpw6;  // ../RTL/cortexm0ds_logic.v(1533)
  wire [30:26] Zbhpw6;  // ../RTL/cortexm0ds_logic.v(1571)
  wire [6:0] Zehpw6;  // ../RTL/cortexm0ds_logic.v(1573)
  wire [30:0] Zsfpw6;  // ../RTL/cortexm0ds_logic.v(1537)
  wire [1:0] n101;
  wire [31:0] n111;
  wire [31:0] n112;
  wire [23:0] n114;
  wire [12:0] n1272;
  wire [7:0] n2661;
  wire [31:0] n4277;
  wire [1:0] n5200;
  wire [1:0] n5488;
  wire [1:0] n5968;
  wire [6:0] n7;
  wire A00iu6;  // ../RTL/cortexm0ds_logic.v(303)
  wire A00pw6;  // ../RTL/cortexm0ds_logic.v(1328)
  wire A06ju6;  // ../RTL/cortexm0ds_logic.v(865)
  wire A07iu6;  // ../RTL/cortexm0ds_logic.v(397)
  wire A07pw6;  // ../RTL/cortexm0ds_logic.v(1421)
  wire A08ow6;  // ../RTL/cortexm0ds_logic.v(953)
  wire A0eiu6;  // ../RTL/cortexm0ds_logic.v(491)
  wire A0epw6;  // ../RTL/cortexm0ds_logic.v(1515)
  wire A0fow6;  // ../RTL/cortexm0ds_logic.v(1047)
  wire A0liu6;  // ../RTL/cortexm0ds_logic.v(584)
  wire A0mow6;  // ../RTL/cortexm0ds_logic.v(1141)
  wire A0siu6;  // ../RTL/cortexm0ds_logic.v(678)
  wire A0thu6;  // ../RTL/cortexm0ds_logic.v(210)
  wire A0tow6;  // ../RTL/cortexm0ds_logic.v(1234)
  wire A0ziu6;  // ../RTL/cortexm0ds_logic.v(771)
  wire A15ju6;  // ../RTL/cortexm0ds_logic.v(852)
  wire A16iu6;  // ../RTL/cortexm0ds_logic.v(384)
  wire A16pw6;  // ../RTL/cortexm0ds_logic.v(1408)
  wire A17ow6;  // ../RTL/cortexm0ds_logic.v(940)
  wire A1diu6;  // ../RTL/cortexm0ds_logic.v(478)
  wire A1dpw6;  // ../RTL/cortexm0ds_logic.v(1502)
  wire A1eow6;  // ../RTL/cortexm0ds_logic.v(1034)
  wire A1kiu6;  // ../RTL/cortexm0ds_logic.v(571)
  wire A1low6;  // ../RTL/cortexm0ds_logic.v(1128)
  wire A1qax6;  // ../RTL/cortexm0ds_logic.v(1661)
  wire A1riu6;  // ../RTL/cortexm0ds_logic.v(665)
  wire A1shu6;  // ../RTL/cortexm0ds_logic.v(197)
  wire A1sow6;  // ../RTL/cortexm0ds_logic.v(1221)
  wire A1yiu6;  // ../RTL/cortexm0ds_logic.v(758)
  wire A1zhu6;  // ../RTL/cortexm0ds_logic.v(290)
  wire A1zow6;  // ../RTL/cortexm0ds_logic.v(1315)
  wire A24ju6;  // ../RTL/cortexm0ds_logic.v(839)
  wire A25iu6;  // ../RTL/cortexm0ds_logic.v(371)
  wire A25pw6;  // ../RTL/cortexm0ds_logic.v(1395)
  wire A2ciu6;  // ../RTL/cortexm0ds_logic.v(465)
  wire A2cpw6;  // ../RTL/cortexm0ds_logic.v(1489)
  wire A2dow6;  // ../RTL/cortexm0ds_logic.v(1021)
  wire A2jiu6;  // ../RTL/cortexm0ds_logic.v(558)
  wire A2kow6;  // ../RTL/cortexm0ds_logic.v(1115)
  wire A2lhu6;  // ../RTL/cortexm0ds_logic.v(138)
  wire A2nhu6;  // ../RTL/cortexm0ds_logic.v(144)
  wire A2qiu6;  // ../RTL/cortexm0ds_logic.v(652)
  wire A2rhu6;  // ../RTL/cortexm0ds_logic.v(184)
  wire A2row6;  // ../RTL/cortexm0ds_logic.v(1208)
  wire A2spw6;  // ../RTL/cortexm0ds_logic.v(1602)
  wire A2xiu6;  // ../RTL/cortexm0ds_logic.v(745)
  wire A2yhu6;  // ../RTL/cortexm0ds_logic.v(277)
  wire A2yow6;  // ../RTL/cortexm0ds_logic.v(1302)
  wire A32qw6;  // ../RTL/cortexm0ds_logic.v(1621)
  wire A33ju6;  // ../RTL/cortexm0ds_logic.v(826)
  wire A34iu6;  // ../RTL/cortexm0ds_logic.v(358)
  wire A34pw6;  // ../RTL/cortexm0ds_logic.v(1382)
  wire A3aju6;  // ../RTL/cortexm0ds_logic.v(920)
  wire A3biu6;  // ../RTL/cortexm0ds_logic.v(452)
  wire A3bpw6;  // ../RTL/cortexm0ds_logic.v(1476)
  wire A3cow6;  // ../RTL/cortexm0ds_logic.v(1008)
  wire A3iiu6;  // ../RTL/cortexm0ds_logic.v(545)
  wire A3ipw6;  // ../RTL/cortexm0ds_logic.v(1584)
  wire A3jow6;  // ../RTL/cortexm0ds_logic.v(1102)
  wire A3piu6;  // ../RTL/cortexm0ds_logic.v(639)
  wire A3qax6;  // ../RTL/cortexm0ds_logic.v(1661)
  wire A3qhu6;  // ../RTL/cortexm0ds_logic.v(171)
  wire A3qow6;  // ../RTL/cortexm0ds_logic.v(1195)
  wire A3wiu6;  // ../RTL/cortexm0ds_logic.v(732)
  wire A3xhu6;  // ../RTL/cortexm0ds_logic.v(264)
  wire A3xow6;  // ../RTL/cortexm0ds_logic.v(1289)
  wire A42ju6;  // ../RTL/cortexm0ds_logic.v(813)
  wire A43pw6;  // ../RTL/cortexm0ds_logic.v(1369)
  wire A49ju6;  // ../RTL/cortexm0ds_logic.v(907)
  wire A4aiu6;  // ../RTL/cortexm0ds_logic.v(439)
  wire A4apw6;  // ../RTL/cortexm0ds_logic.v(1463)
  wire A4bow6;  // ../RTL/cortexm0ds_logic.v(995)
  wire A4hiu6;  // ../RTL/cortexm0ds_logic.v(532)
  wire A4iow6;  // ../RTL/cortexm0ds_logic.v(1089)
  wire A4khu6;  // ../RTL/cortexm0ds_logic.v(135)
  wire A4oiu6;  // ../RTL/cortexm0ds_logic.v(626)
  wire A4phu6;  // ../RTL/cortexm0ds_logic.v(158)
  wire A4pow6;  // ../RTL/cortexm0ds_logic.v(1182)
  wire A4viu6;  // ../RTL/cortexm0ds_logic.v(719)
  wire A4whu6;  // ../RTL/cortexm0ds_logic.v(251)
  wire A4wow6;  // ../RTL/cortexm0ds_logic.v(1276)
  wire A51ju6;  // ../RTL/cortexm0ds_logic.v(800)
  wire A52iu6;  // ../RTL/cortexm0ds_logic.v(332)
  wire A52pw6;  // ../RTL/cortexm0ds_logic.v(1356)
  wire A58ju6;  // ../RTL/cortexm0ds_logic.v(894)
  wire A59iu6;  // ../RTL/cortexm0ds_logic.v(426)
  wire A59pw6;  // ../RTL/cortexm0ds_logic.v(1450)
  wire A5aow6;  // ../RTL/cortexm0ds_logic.v(982)
  wire A5giu6;  // ../RTL/cortexm0ds_logic.v(519)
  wire A5how6;  // ../RTL/cortexm0ds_logic.v(1076)
  wire A5ipw6;  // ../RTL/cortexm0ds_logic.v(1584)
  wire A5niu6;  // ../RTL/cortexm0ds_logic.v(613)
  wire A5oow6;  // ../RTL/cortexm0ds_logic.v(1169)
  wire A5qax6;  // ../RTL/cortexm0ds_logic.v(1662)
  wire A5uiu6;  // ../RTL/cortexm0ds_logic.v(706)
  wire A5vhu6;  // ../RTL/cortexm0ds_logic.v(238)
  wire A5vow6;  // ../RTL/cortexm0ds_logic.v(1263)
  wire A60ju6;  // ../RTL/cortexm0ds_logic.v(787)
  wire A61iu6;  // ../RTL/cortexm0ds_logic.v(319)
  wire A61pw6;  // ../RTL/cortexm0ds_logic.v(1343)
  wire A67ju6;  // ../RTL/cortexm0ds_logic.v(881)
  wire A68iu6;  // ../RTL/cortexm0ds_logic.v(413)
  wire A68pw6;  // ../RTL/cortexm0ds_logic.v(1437)
  wire A69ow6;  // ../RTL/cortexm0ds_logic.v(969)
  wire A6cbx6;  // ../RTL/cortexm0ds_logic.v(1701)
  wire A6fiu6;  // ../RTL/cortexm0ds_logic.v(506)
  wire A6gow6;  // ../RTL/cortexm0ds_logic.v(1063)
  wire A6jhu6;  // ../RTL/cortexm0ds_logic.v(133)
  wire A6miu6;  // ../RTL/cortexm0ds_logic.v(600)
  wire A6now6;  // ../RTL/cortexm0ds_logic.v(1156)
  wire A6tiu6;  // ../RTL/cortexm0ds_logic.v(693)
  wire A6uhu6;  // ../RTL/cortexm0ds_logic.v(225)
  wire A6uow6;  // ../RTL/cortexm0ds_logic.v(1250)
  wire A70iu6;  // ../RTL/cortexm0ds_logic.v(306)
  wire A70pw6;  // ../RTL/cortexm0ds_logic.v(1330)
  wire A76ju6;  // ../RTL/cortexm0ds_logic.v(868)
  wire A77iu6;  // ../RTL/cortexm0ds_logic.v(400)
  wire A77pw6;  // ../RTL/cortexm0ds_logic.v(1424)
  wire A78ow6;  // ../RTL/cortexm0ds_logic.v(956)
  wire A7eiu6;  // ../RTL/cortexm0ds_logic.v(493)
  wire A7fow6;  // ../RTL/cortexm0ds_logic.v(1050)
  wire A7liu6;  // ../RTL/cortexm0ds_logic.v(587)
  wire A7mow6;  // ../RTL/cortexm0ds_logic.v(1143)
  wire A7siu6;  // ../RTL/cortexm0ds_logic.v(680)
  wire A7thu6;  // ../RTL/cortexm0ds_logic.v(212)
  wire A7tow6;  // ../RTL/cortexm0ds_logic.v(1237)
  wire A7ziu6;  // ../RTL/cortexm0ds_logic.v(774)
  wire A7zpw6;  // ../RTL/cortexm0ds_logic.v(1615)
  wire A85ju6;  // ../RTL/cortexm0ds_logic.v(855)
  wire A86iu6;  // ../RTL/cortexm0ds_logic.v(387)
  wire A86pw6;  // ../RTL/cortexm0ds_logic.v(1411)
  wire A87ow6;  // ../RTL/cortexm0ds_logic.v(943)
  wire A8diu6;  // ../RTL/cortexm0ds_logic.v(480)
  wire A8dpw6;  // ../RTL/cortexm0ds_logic.v(1505)
  wire A8eow6;  // ../RTL/cortexm0ds_logic.v(1037)
  wire A8ihu6;  // ../RTL/cortexm0ds_logic.v(130)
  wire A8kiu6;  // ../RTL/cortexm0ds_logic.v(574)
  wire A8low6;  // ../RTL/cortexm0ds_logic.v(1130)
  wire A8riu6;  // ../RTL/cortexm0ds_logic.v(667)
  wire A8shu6;  // ../RTL/cortexm0ds_logic.v(199)
  wire A8sow6;  // ../RTL/cortexm0ds_logic.v(1224)
  wire A8yiu6;  // ../RTL/cortexm0ds_logic.v(761)
  wire A8zhu6;  // ../RTL/cortexm0ds_logic.v(293)
  wire A8zow6;  // ../RTL/cortexm0ds_logic.v(1317)
  wire A94ju6;  // ../RTL/cortexm0ds_logic.v(842)
  wire A95iu6;  // ../RTL/cortexm0ds_logic.v(374)
  wire A95pw6;  // ../RTL/cortexm0ds_logic.v(1398)
  wire A96ow6;  // ../RTL/cortexm0ds_logic.v(930)
  wire A9ciu6;  // ../RTL/cortexm0ds_logic.v(467)
  wire A9cpw6;  // ../RTL/cortexm0ds_logic.v(1492)
  wire A9dow6;  // ../RTL/cortexm0ds_logic.v(1024)
  wire A9jiu6;  // ../RTL/cortexm0ds_logic.v(561)
  wire A9kow6;  // ../RTL/cortexm0ds_logic.v(1117)
  wire A9qiu6;  // ../RTL/cortexm0ds_logic.v(654)
  wire A9rhu6;  // ../RTL/cortexm0ds_logic.v(186)
  wire A9row6;  // ../RTL/cortexm0ds_logic.v(1211)
  wire A9xiu6;  // ../RTL/cortexm0ds_logic.v(748)
  wire A9yhu6;  // ../RTL/cortexm0ds_logic.v(280)
  wire A9yow6;  // ../RTL/cortexm0ds_logic.v(1304)
  wire Aa2bx6;  // ../RTL/cortexm0ds_logic.v(1683)
  wire Aa3ju6;  // ../RTL/cortexm0ds_logic.v(829)
  wire Aa4iu6;  // ../RTL/cortexm0ds_logic.v(361)
  wire Aa4pw6;  // ../RTL/cortexm0ds_logic.v(1385)
  wire Aaaju6;  // ../RTL/cortexm0ds_logic.v(922)
  wire Aabiu6;  // ../RTL/cortexm0ds_logic.v(454)
  wire Aabpw6;  // ../RTL/cortexm0ds_logic.v(1479)
  wire Aacow6;  // ../RTL/cortexm0ds_logic.v(1011)
  wire Aaiiu6;  // ../RTL/cortexm0ds_logic.v(548)
  wire Aajow6;  // ../RTL/cortexm0ds_logic.v(1104)
  wire Aapiu6;  // ../RTL/cortexm0ds_logic.v(641)
  wire Aaqhu6;  // ../RTL/cortexm0ds_logic.v(173)
  wire Aaqow6;  // ../RTL/cortexm0ds_logic.v(1198)
  wire Aawiu6;  // ../RTL/cortexm0ds_logic.v(735)
  wire Aaxhu6;  // ../RTL/cortexm0ds_logic.v(267)
  wire Aaxow6;  // ../RTL/cortexm0ds_logic.v(1291)
  wire Ab2ju6;  // ../RTL/cortexm0ds_logic.v(816)
  wire Ab3iu6;  // ../RTL/cortexm0ds_logic.v(348)
  wire Ab3pw6;  // ../RTL/cortexm0ds_logic.v(1372)
  wire Ab9ax6;  // ../RTL/cortexm0ds_logic.v(1630)
  wire Ab9ju6;  // ../RTL/cortexm0ds_logic.v(909)
  wire Abaiu6;  // ../RTL/cortexm0ds_logic.v(441)
  wire Abapw6;  // ../RTL/cortexm0ds_logic.v(1466)
  wire Abbow6;  // ../RTL/cortexm0ds_logic.v(998)
  wire Abfhu6;  // ../RTL/cortexm0ds_logic.v(124)
  wire Abhiu6;  // ../RTL/cortexm0ds_logic.v(535)
  wire Abiow6;  // ../RTL/cortexm0ds_logic.v(1091)
  wire Aboiu6;  // ../RTL/cortexm0ds_logic.v(628)
  wire Abphu6;  // ../RTL/cortexm0ds_logic.v(160)
  wire Abpow6;  // ../RTL/cortexm0ds_logic.v(1185)
  wire Abviu6;  // ../RTL/cortexm0ds_logic.v(722)
  wire Abwhu6;  // ../RTL/cortexm0ds_logic.v(254)
  wire Abwow6;  // ../RTL/cortexm0ds_logic.v(1278)
  wire Ac1ju6;  // ../RTL/cortexm0ds_logic.v(803)
  wire Ac2iu6;  // ../RTL/cortexm0ds_logic.v(335)
  wire Ac2pw6;  // ../RTL/cortexm0ds_logic.v(1359)
  wire Ac8ju6;  // ../RTL/cortexm0ds_logic.v(896)
  wire Ac9iu6;  // ../RTL/cortexm0ds_logic.v(428)
  wire Ac9pw6;  // ../RTL/cortexm0ds_logic.v(1453)
  wire Acaow6;  // ../RTL/cortexm0ds_logic.v(985)
  wire Acebx6;  // ../RTL/cortexm0ds_logic.v(1705)
  wire Acgiu6;  // ../RTL/cortexm0ds_logic.v(522)
  wire Achow6;  // ../RTL/cortexm0ds_logic.v(1078)
  wire Acniu6;  // ../RTL/cortexm0ds_logic.v(615)
  wire Acohu6;  // ../RTL/cortexm0ds_logic.v(147)
  wire Acoow6;  // ../RTL/cortexm0ds_logic.v(1172)
  wire Acuax6;  // ../RTL/cortexm0ds_logic.v(1669)
  wire Acuiu6;  // ../RTL/cortexm0ds_logic.v(709)
  wire Acvhu6;  // ../RTL/cortexm0ds_logic.v(241)
  wire Acvow6;  // ../RTL/cortexm0ds_logic.v(1265)
  wire Ad0ju6;  // ../RTL/cortexm0ds_logic.v(790)
  wire Ad1iu6;  // ../RTL/cortexm0ds_logic.v(322)
  wire Ad1pw6;  // ../RTL/cortexm0ds_logic.v(1346)
  wire Ad7ax6;  // ../RTL/cortexm0ds_logic.v(1626)
  wire Ad7ju6;  // ../RTL/cortexm0ds_logic.v(883)
  wire Ad8iu6;  // ../RTL/cortexm0ds_logic.v(415)
  wire Ad8pw6;  // ../RTL/cortexm0ds_logic.v(1440)
  wire Ad9ow6;  // ../RTL/cortexm0ds_logic.v(972)
  wire Adfiu6;  // ../RTL/cortexm0ds_logic.v(509)
  wire Adgow6;  // ../RTL/cortexm0ds_logic.v(1065)
  wire Admiu6;  // ../RTL/cortexm0ds_logic.v(602)
  wire Adnow6;  // ../RTL/cortexm0ds_logic.v(1159)
  wire Adtiu6;  // ../RTL/cortexm0ds_logic.v(696)
  wire Aduhu6;  // ../RTL/cortexm0ds_logic.v(228)
  wire Aduow6;  // ../RTL/cortexm0ds_logic.v(1252)
  wire Ae0iu6;  // ../RTL/cortexm0ds_logic.v(309)
  wire Ae0pw6;  // ../RTL/cortexm0ds_logic.v(1333)
  wire Ae6ju6;  // ../RTL/cortexm0ds_logic.v(870)
  wire Ae7iu6;  // ../RTL/cortexm0ds_logic.v(402)
  wire Ae7pw6;  // ../RTL/cortexm0ds_logic.v(1427)
  wire Ae8ow6;  // ../RTL/cortexm0ds_logic.v(959)
  wire Aeeiu6;  // ../RTL/cortexm0ds_logic.v(496)
  wire Aefow6;  // ../RTL/cortexm0ds_logic.v(1052)
  wire Aeliu6;  // ../RTL/cortexm0ds_logic.v(589)
  wire Aemow6;  // ../RTL/cortexm0ds_logic.v(1146)
  wire Aesiu6;  // ../RTL/cortexm0ds_logic.v(683)
  wire Aethu6;  // ../RTL/cortexm0ds_logic.v(215)
  wire Aetow6;  // ../RTL/cortexm0ds_logic.v(1239)
  wire Aeziu6;  // ../RTL/cortexm0ds_logic.v(777)
  wire Af5ju6;  // ../RTL/cortexm0ds_logic.v(857)
  wire Af6iu6;  // ../RTL/cortexm0ds_logic.v(389)
  wire Af6pw6;  // ../RTL/cortexm0ds_logic.v(1414)
  wire Af7ow6;  // ../RTL/cortexm0ds_logic.v(946)
  wire Afdiu6;  // ../RTL/cortexm0ds_logic.v(483)
  wire Afdpw6;  // ../RTL/cortexm0ds_logic.v(1507)
  wire Afeow6;  // ../RTL/cortexm0ds_logic.v(1039)
  wire Afkiu6;  // ../RTL/cortexm0ds_logic.v(576)
  wire Aflow6;  // ../RTL/cortexm0ds_logic.v(1133)
  wire Afriu6;  // ../RTL/cortexm0ds_logic.v(670)
  wire Afshu6;  // ../RTL/cortexm0ds_logic.v(202)
  wire Afsow6;  // ../RTL/cortexm0ds_logic.v(1226)
  wire Afyiu6;  // ../RTL/cortexm0ds_logic.v(764)
  wire Afzhu6;  // ../RTL/cortexm0ds_logic.v(296)
  wire Afzow6;  // ../RTL/cortexm0ds_logic.v(1320)
  wire Ag4ju6;  // ../RTL/cortexm0ds_logic.v(844)
  wire Ag5iu6;  // ../RTL/cortexm0ds_logic.v(376)
  wire Ag5pw6;  // ../RTL/cortexm0ds_logic.v(1401)
  wire Ag6ow6;  // ../RTL/cortexm0ds_logic.v(933)
  wire Agciu6;  // ../RTL/cortexm0ds_logic.v(470)
  wire Agcpw6;  // ../RTL/cortexm0ds_logic.v(1494)
  wire Agdow6;  // ../RTL/cortexm0ds_logic.v(1026)
  wire Aghhu6;  // ../RTL/cortexm0ds_logic.v(128)
  wire Agjiu6;  // ../RTL/cortexm0ds_logic.v(563)
  wire Agkow6;  // ../RTL/cortexm0ds_logic.v(1120)
  wire Agqiu6;  // ../RTL/cortexm0ds_logic.v(657)
  wire Agrhu6;  // ../RTL/cortexm0ds_logic.v(189)
  wire Agrow6;  // ../RTL/cortexm0ds_logic.v(1213)
  wire Agxiu6;  // ../RTL/cortexm0ds_logic.v(751)
  wire Agyhu6;  // ../RTL/cortexm0ds_logic.v(283)
  wire Agyow6;  // ../RTL/cortexm0ds_logic.v(1307)
  wire Ah3ju6;  // ../RTL/cortexm0ds_logic.v(831)
  wire Ah4iu6;  // ../RTL/cortexm0ds_logic.v(363)
  wire Ah4pw6;  // ../RTL/cortexm0ds_logic.v(1388)
  wire Ahaju6;  // ../RTL/cortexm0ds_logic.v(925)
  wire Ahbiu6;  // ../RTL/cortexm0ds_logic.v(457)
  wire Ahbpw6;  // ../RTL/cortexm0ds_logic.v(1481)
  wire Ahcow6;  // ../RTL/cortexm0ds_logic.v(1013)
  wire Ahdax6;  // ../RTL/cortexm0ds_logic.v(1638)
  wire Ahdbx6;  // ../RTL/cortexm0ds_logic.v(1704)
  wire Ahghu6;  // ../RTL/cortexm0ds_logic.v(126)
  wire Ahiiu6;  // ../RTL/cortexm0ds_logic.v(550)
  wire Ahjow6;  // ../RTL/cortexm0ds_logic.v(1107)
  wire Ahlpw6;  // ../RTL/cortexm0ds_logic.v(1590)
  wire Ahpiu6;  // ../RTL/cortexm0ds_logic.v(644)
  wire Ahqhu6;  // ../RTL/cortexm0ds_logic.v(176)
  wire Ahqow6;  // ../RTL/cortexm0ds_logic.v(1200)
  wire Ahwiu6;  // ../RTL/cortexm0ds_logic.v(738)
  wire Ahxhu6;  // ../RTL/cortexm0ds_logic.v(270)
  wire Ahxow6;  // ../RTL/cortexm0ds_logic.v(1294)
  wire Ai2ju6;  // ../RTL/cortexm0ds_logic.v(818)
  wire Ai3iu6;  // ../RTL/cortexm0ds_logic.v(350)
  wire Ai3pw6;  // ../RTL/cortexm0ds_logic.v(1375)
  wire Ai9ju6;  // ../RTL/cortexm0ds_logic.v(912)
  wire Aiaiu6;  // ../RTL/cortexm0ds_logic.v(444)
  wire Aiapw6;  // ../RTL/cortexm0ds_logic.v(1468)
  wire Aibow6;  // ../RTL/cortexm0ds_logic.v(1000)
  wire Aihiu6;  // ../RTL/cortexm0ds_logic.v(537)
  wire Aiiow6;  // ../RTL/cortexm0ds_logic.v(1094)
  wire Aioiu6;  // ../RTL/cortexm0ds_logic.v(631)
  wire Aiphu6;  // ../RTL/cortexm0ds_logic.v(163)
  wire Aipow6;  // ../RTL/cortexm0ds_logic.v(1187)
  wire Aiviu6;  // ../RTL/cortexm0ds_logic.v(725)
  wire Aiwhu6;  // ../RTL/cortexm0ds_logic.v(257)
  wire Aiwow6;  // ../RTL/cortexm0ds_logic.v(1281)
  wire Aj1ju6;  // ../RTL/cortexm0ds_logic.v(805)
  wire Aj2iu6;  // ../RTL/cortexm0ds_logic.v(337)
  wire Aj2pw6;  // ../RTL/cortexm0ds_logic.v(1362)
  wire Aj8ju6;  // ../RTL/cortexm0ds_logic.v(899)
  wire Aj9iu6;  // ../RTL/cortexm0ds_logic.v(431)
  wire Aj9pw6;  // ../RTL/cortexm0ds_logic.v(1455)
  wire Ajaow6;  // ../RTL/cortexm0ds_logic.v(987)
  wire Ajgiu6;  // ../RTL/cortexm0ds_logic.v(524)
  wire Ajhow6;  // ../RTL/cortexm0ds_logic.v(1081)
  wire Ajniu6;  // ../RTL/cortexm0ds_logic.v(618)
  wire Ajohu6;  // ../RTL/cortexm0ds_logic.v(150)
  wire Ajoow6;  // ../RTL/cortexm0ds_logic.v(1174)
  wire Ajuiu6;  // ../RTL/cortexm0ds_logic.v(712)
  wire Ajvhu6;  // ../RTL/cortexm0ds_logic.v(244)
  wire Ajvow6;  // ../RTL/cortexm0ds_logic.v(1268)
  wire Ak0ju6;  // ../RTL/cortexm0ds_logic.v(792)
  wire Ak1iu6;  // ../RTL/cortexm0ds_logic.v(324)
  wire Ak1pw6;  // ../RTL/cortexm0ds_logic.v(1349)
  wire Ak7ju6;  // ../RTL/cortexm0ds_logic.v(886)
  wire Ak8iu6;  // ../RTL/cortexm0ds_logic.v(418)
  wire Ak8pw6;  // ../RTL/cortexm0ds_logic.v(1442)
  wire Ak9ow6;  // ../RTL/cortexm0ds_logic.v(974)
  wire Akfiu6;  // ../RTL/cortexm0ds_logic.v(511)
  wire Akgow6;  // ../RTL/cortexm0ds_logic.v(1068)
  wire Akmiu6;  // ../RTL/cortexm0ds_logic.v(605)
  wire Aknow6;  // ../RTL/cortexm0ds_logic.v(1161)
  wire Aktiu6;  // ../RTL/cortexm0ds_logic.v(699)
  wire Akuhu6;  // ../RTL/cortexm0ds_logic.v(231)
  wire Akuow6;  // ../RTL/cortexm0ds_logic.v(1255)
  wire Al0iu6;  // ../RTL/cortexm0ds_logic.v(311)
  wire Al0pw6;  // ../RTL/cortexm0ds_logic.v(1336)
  wire Al6ju6;  // ../RTL/cortexm0ds_logic.v(873)
  wire Al7iu6;  // ../RTL/cortexm0ds_logic.v(405)
  wire Al7pw6;  // ../RTL/cortexm0ds_logic.v(1429)
  wire Al8ow6;  // ../RTL/cortexm0ds_logic.v(961)
  wire Aleiu6;  // ../RTL/cortexm0ds_logic.v(498)
  wire Alfow6;  // ../RTL/cortexm0ds_logic.v(1055)
  wire Alhhu6;  // ../RTL/cortexm0ds_logic.v(129)
  wire Alkhu6;  // ../RTL/cortexm0ds_logic.v(137)
  wire Alliu6;  // ../RTL/cortexm0ds_logic.v(592)
  wire Almow6;  // ../RTL/cortexm0ds_logic.v(1148)
  wire Alsiu6;  // ../RTL/cortexm0ds_logic.v(686)
  wire Althu6;  // ../RTL/cortexm0ds_logic.v(218)
  wire Altow6;  // ../RTL/cortexm0ds_logic.v(1242)
  wire Alziu6;  // ../RTL/cortexm0ds_logic.v(779)
  wire Am5ju6;  // ../RTL/cortexm0ds_logic.v(860)
  wire Am6iu6;  // ../RTL/cortexm0ds_logic.v(392)
  wire Am6pw6;  // ../RTL/cortexm0ds_logic.v(1416)
  wire Am7ow6;  // ../RTL/cortexm0ds_logic.v(948)
  wire Amdiu6;  // ../RTL/cortexm0ds_logic.v(485)
  wire Amdpw6;  // ../RTL/cortexm0ds_logic.v(1510)
  wire Ameow6;  // ../RTL/cortexm0ds_logic.v(1042)
  wire Amkiu6;  // ../RTL/cortexm0ds_logic.v(579)
  wire Amlow6;  // ../RTL/cortexm0ds_logic.v(1135)
  wire Amriu6;  // ../RTL/cortexm0ds_logic.v(673)
  wire Amshu6;  // ../RTL/cortexm0ds_logic.v(205)
  wire Amsow6;  // ../RTL/cortexm0ds_logic.v(1229)
  wire Amupw6;  // ../RTL/cortexm0ds_logic.v(1607)
  wire Amyiu6;  // ../RTL/cortexm0ds_logic.v(766)
  wire Amzhu6;  // ../RTL/cortexm0ds_logic.v(298)
  wire Amzow6;  // ../RTL/cortexm0ds_logic.v(1323)
  wire An4ju6;  // ../RTL/cortexm0ds_logic.v(847)
  wire An5iu6;  // ../RTL/cortexm0ds_logic.v(379)
  wire An5pw6;  // ../RTL/cortexm0ds_logic.v(1403)
  wire An6ow6;  // ../RTL/cortexm0ds_logic.v(935)
  wire Anciu6;  // ../RTL/cortexm0ds_logic.v(472)
  wire Ancpw6;  // ../RTL/cortexm0ds_logic.v(1497)
  wire Andow6;  // ../RTL/cortexm0ds_logic.v(1029)
  wire Aniax6;  // ../RTL/cortexm0ds_logic.v(1648)
  wire Anjhu6;  // ../RTL/cortexm0ds_logic.v(134)
  wire Anjiu6;  // ../RTL/cortexm0ds_logic.v(566)
  wire Ankow6;  // ../RTL/cortexm0ds_logic.v(1122)
  wire Anqiu6;  // ../RTL/cortexm0ds_logic.v(660)
  wire Anrhu6;  // ../RTL/cortexm0ds_logic.v(192)
  wire Anrow6;  // ../RTL/cortexm0ds_logic.v(1216)
  wire Anxiu6;  // ../RTL/cortexm0ds_logic.v(753)
  wire Anyhu6;  // ../RTL/cortexm0ds_logic.v(285)
  wire Anyow6;  // ../RTL/cortexm0ds_logic.v(1310)
  wire Ao3ju6;  // ../RTL/cortexm0ds_logic.v(834)
  wire Ao4iu6;  // ../RTL/cortexm0ds_logic.v(366)
  wire Ao4pw6;  // ../RTL/cortexm0ds_logic.v(1390)
  wire Aoaju6;  // ../RTL/cortexm0ds_logic.v(927)
  wire Aobiu6;  // ../RTL/cortexm0ds_logic.v(459)
  wire Aobpw6;  // ../RTL/cortexm0ds_logic.v(1484)
  wire Aocow6;  // ../RTL/cortexm0ds_logic.v(1016)
  wire Aoeax6;  // ../RTL/cortexm0ds_logic.v(1640)
  wire Aoiiu6;  // ../RTL/cortexm0ds_logic.v(553)
  wire Aojow6;  // ../RTL/cortexm0ds_logic.v(1109)
  wire Aopiu6;  // ../RTL/cortexm0ds_logic.v(647)
  wire Aoqhu6;  // ../RTL/cortexm0ds_logic.v(179)
  wire Aoqow6;  // ../RTL/cortexm0ds_logic.v(1203)
  wire Aowiu6;  // ../RTL/cortexm0ds_logic.v(740)
  wire Aoxhu6;  // ../RTL/cortexm0ds_logic.v(272)
  wire Aoxow6;  // ../RTL/cortexm0ds_logic.v(1297)
  wire Ap2ju6;  // ../RTL/cortexm0ds_logic.v(821)
  wire Ap3iu6;  // ../RTL/cortexm0ds_logic.v(353)
  wire Ap3pw6;  // ../RTL/cortexm0ds_logic.v(1377)
  wire Ap9ju6;  // ../RTL/cortexm0ds_logic.v(914)
  wire Apaiu6;  // ../RTL/cortexm0ds_logic.v(446)
  wire Apapw6;  // ../RTL/cortexm0ds_logic.v(1471)
  wire Apbow6;  // ../RTL/cortexm0ds_logic.v(1003)
  wire Apcax6;  // ../RTL/cortexm0ds_logic.v(1636)
  wire Aphiu6;  // ../RTL/cortexm0ds_logic.v(540)
  wire Apihu6;  // ../RTL/cortexm0ds_logic.v(132)
  wire Apiow6;  // ../RTL/cortexm0ds_logic.v(1096)
  wire Apoiu6;  // ../RTL/cortexm0ds_logic.v(634)
  wire Apphu6;  // ../RTL/cortexm0ds_logic.v(166)
  wire Appow6;  // ../RTL/cortexm0ds_logic.v(1190)
  wire Apviu6;  // ../RTL/cortexm0ds_logic.v(727)
  wire Apwhu6;  // ../RTL/cortexm0ds_logic.v(259)
  wire Apwow6;  // ../RTL/cortexm0ds_logic.v(1284)
  wire Aq1ju6;  // ../RTL/cortexm0ds_logic.v(808)
  wire Aq2iu6;  // ../RTL/cortexm0ds_logic.v(340)
  wire Aq2pw6;  // ../RTL/cortexm0ds_logic.v(1364)
  wire Aq8ju6;  // ../RTL/cortexm0ds_logic.v(901)
  wire Aq9iu6;  // ../RTL/cortexm0ds_logic.v(433)
  wire Aq9pw6;  // ../RTL/cortexm0ds_logic.v(1458)
  wire Aqaow6;  // ../RTL/cortexm0ds_logic.v(990)
  wire Aqgiu6;  // ../RTL/cortexm0ds_logic.v(527)
  wire Aqhow6;  // ../RTL/cortexm0ds_logic.v(1083)
  wire Aqlax6;  // ../RTL/cortexm0ds_logic.v(1654)
  wire Aqniu6;  // ../RTL/cortexm0ds_logic.v(621)
  wire Aqohu6;  // ../RTL/cortexm0ds_logic.v(153)
  wire Aqoow6;  // ../RTL/cortexm0ds_logic.v(1177)
  wire Aquiu6;  // ../RTL/cortexm0ds_logic.v(714)
  wire Aqvhu6;  // ../RTL/cortexm0ds_logic.v(246)
  wire Aqvow6;  // ../RTL/cortexm0ds_logic.v(1271)
  wire Ar0ju6;  // ../RTL/cortexm0ds_logic.v(795)
  wire Ar1bx6;  // ../RTL/cortexm0ds_logic.v(1682)
  wire Ar1iu6;  // ../RTL/cortexm0ds_logic.v(327)
  wire Ar1pw6;  // ../RTL/cortexm0ds_logic.v(1351)
  wire Ar7ju6;  // ../RTL/cortexm0ds_logic.v(888)
  wire Ar8iu6;  // ../RTL/cortexm0ds_logic.v(420)
  wire Ar8pw6;  // ../RTL/cortexm0ds_logic.v(1445)
  wire Ar9ow6;  // ../RTL/cortexm0ds_logic.v(977)
  wire Arehu6;  // ../RTL/cortexm0ds_logic.v(122)
  wire Arfiu6;  // ../RTL/cortexm0ds_logic.v(514)
  wire Argow6;  // ../RTL/cortexm0ds_logic.v(1070)
  wire Armiu6;  // ../RTL/cortexm0ds_logic.v(608)
  wire Arnow6;  // ../RTL/cortexm0ds_logic.v(1164)
  wire Arnpw6;  // ../RTL/cortexm0ds_logic.v(1595)
  wire Artiu6;  // ../RTL/cortexm0ds_logic.v(701)
  wire Aruhu6;  // ../RTL/cortexm0ds_logic.v(233)
  wire Aruow6;  // ../RTL/cortexm0ds_logic.v(1258)
  wire As0iu6;  // ../RTL/cortexm0ds_logic.v(314)
  wire As0pw6;  // ../RTL/cortexm0ds_logic.v(1338)
  wire As6ju6;  // ../RTL/cortexm0ds_logic.v(875)
  wire As7iu6;  // ../RTL/cortexm0ds_logic.v(407)
  wire As7pw6;  // ../RTL/cortexm0ds_logic.v(1432)
  wire As8ow6;  // ../RTL/cortexm0ds_logic.v(964)
  wire Aseiu6;  // ../RTL/cortexm0ds_logic.v(501)
  wire Asfow6;  // ../RTL/cortexm0ds_logic.v(1057)
  wire Asliu6;  // ../RTL/cortexm0ds_logic.v(595)
  wire Asmow6;  // ../RTL/cortexm0ds_logic.v(1151)
  wire Assiu6;  // ../RTL/cortexm0ds_logic.v(688)
  wire Asthu6;  // ../RTL/cortexm0ds_logic.v(220)
  wire Astow6;  // ../RTL/cortexm0ds_logic.v(1245)
  wire Asupw6;  // ../RTL/cortexm0ds_logic.v(1607)
  wire Asziu6;  // ../RTL/cortexm0ds_logic.v(782)
  wire At2bx6;  // ../RTL/cortexm0ds_logic.v(1684)
  wire At5ju6;  // ../RTL/cortexm0ds_logic.v(862)
  wire At6iu6;  // ../RTL/cortexm0ds_logic.v(394)
  wire At6pw6;  // ../RTL/cortexm0ds_logic.v(1419)
  wire At7ow6;  // ../RTL/cortexm0ds_logic.v(951)
  wire Atdiu6;  // ../RTL/cortexm0ds_logic.v(488)
  wire Atdpw6;  // ../RTL/cortexm0ds_logic.v(1512)
  wire Ateow6;  // ../RTL/cortexm0ds_logic.v(1044)
  wire Atkiu6;  // ../RTL/cortexm0ds_logic.v(582)
  wire Atlow6;  // ../RTL/cortexm0ds_logic.v(1138)
  wire Atriu6;  // ../RTL/cortexm0ds_logic.v(675)
  wire Atshu6;  // ../RTL/cortexm0ds_logic.v(207)
  wire Atsow6;  // ../RTL/cortexm0ds_logic.v(1232)
  wire Atyiu6;  // ../RTL/cortexm0ds_logic.v(769)
  wire Atzhu6;  // ../RTL/cortexm0ds_logic.v(301)
  wire Atzow6;  // ../RTL/cortexm0ds_logic.v(1325)
  wire Au4ju6;  // ../RTL/cortexm0ds_logic.v(849)
  wire Au5iu6;  // ../RTL/cortexm0ds_logic.v(381)
  wire Au5pw6;  // ../RTL/cortexm0ds_logic.v(1406)
  wire Au6ow6;  // ../RTL/cortexm0ds_logic.v(938)
  wire Auciu6;  // ../RTL/cortexm0ds_logic.v(475)
  wire Aucpw6;  // ../RTL/cortexm0ds_logic.v(1499)
  wire Audow6;  // ../RTL/cortexm0ds_logic.v(1031)
  wire Aujiu6;  // ../RTL/cortexm0ds_logic.v(569)
  wire Aujpw6;  // ../RTL/cortexm0ds_logic.v(1587)
  wire Aukow6;  // ../RTL/cortexm0ds_logic.v(1125)
  wire Auqiu6;  // ../RTL/cortexm0ds_logic.v(662)
  wire Aurhu6;  // ../RTL/cortexm0ds_logic.v(194)
  wire Aurow6;  // ../RTL/cortexm0ds_logic.v(1219)
  wire Aurpw6;  // ../RTL/cortexm0ds_logic.v(1602)
  wire Auxiu6;  // ../RTL/cortexm0ds_logic.v(756)
  wire Auyax6;  // ../RTL/cortexm0ds_logic.v(1677)
  wire Auyhu6;  // ../RTL/cortexm0ds_logic.v(288)
  wire Auyow6;  // ../RTL/cortexm0ds_logic.v(1312)
  wire Av3ju6;  // ../RTL/cortexm0ds_logic.v(836)
  wire Av4iu6;  // ../RTL/cortexm0ds_logic.v(368)
  wire Av4pw6;  // ../RTL/cortexm0ds_logic.v(1393)
  wire Avbiu6;  // ../RTL/cortexm0ds_logic.v(462)
  wire Avbpw6;  // ../RTL/cortexm0ds_logic.v(1486)
  wire Avcow6;  // ../RTL/cortexm0ds_logic.v(1018)
  wire Aviiu6;  // ../RTL/cortexm0ds_logic.v(556)
  wire Avjow6;  // ../RTL/cortexm0ds_logic.v(1112)
  wire Avmhu6;  // ../RTL/cortexm0ds_logic.v(143)
  wire Avpiu6;  // ../RTL/cortexm0ds_logic.v(649)
  wire Avqhu6;  // ../RTL/cortexm0ds_logic.v(181)
  wire Avqow6;  // ../RTL/cortexm0ds_logic.v(1206)
  wire Avwiu6;  // ../RTL/cortexm0ds_logic.v(743)
  wire Avxhu6;  // ../RTL/cortexm0ds_logic.v(275)
  wire Avxow6;  // ../RTL/cortexm0ds_logic.v(1299)
  wire Avzax6;  // ../RTL/cortexm0ds_logic.v(1679)
  wire Aw2ju6;  // ../RTL/cortexm0ds_logic.v(823)
  wire Aw3iu6;  // ../RTL/cortexm0ds_logic.v(355)
  wire Aw3pw6;  // ../RTL/cortexm0ds_logic.v(1380)
  wire Aw4bx6;  // ../RTL/cortexm0ds_logic.v(1688)
  wire Aw9ju6;  // ../RTL/cortexm0ds_logic.v(917)
  wire Awaiu6;  // ../RTL/cortexm0ds_logic.v(449)
  wire Awapw6;  // ../RTL/cortexm0ds_logic.v(1473)
  wire Awbow6;  // ../RTL/cortexm0ds_logic.v(1005)
  wire Awhiu6;  // ../RTL/cortexm0ds_logic.v(543)
  wire Awiow6;  // ../RTL/cortexm0ds_logic.v(1099)
  wire Awoiu6;  // ../RTL/cortexm0ds_logic.v(636)
  wire Awphu6;  // ../RTL/cortexm0ds_logic.v(168)
  wire Awpow6;  // ../RTL/cortexm0ds_logic.v(1193)
  wire Awupw6;  // ../RTL/cortexm0ds_logic.v(1608)
  wire Awviu6;  // ../RTL/cortexm0ds_logic.v(730)
  wire Awwhu6;  // ../RTL/cortexm0ds_logic.v(262)
  wire Awwow6;  // ../RTL/cortexm0ds_logic.v(1286)
  wire Ax1ju6;  // ../RTL/cortexm0ds_logic.v(810)
  wire Ax2iu6;  // ../RTL/cortexm0ds_logic.v(342)
  wire Ax2pw6;  // ../RTL/cortexm0ds_logic.v(1367)
  wire Ax8ju6;  // ../RTL/cortexm0ds_logic.v(904)
  wire Ax9iu6;  // ../RTL/cortexm0ds_logic.v(436)
  wire Ax9pw6;  // ../RTL/cortexm0ds_logic.v(1460)
  wire Axaow6;  // ../RTL/cortexm0ds_logic.v(992)
  wire Axgiu6;  // ../RTL/cortexm0ds_logic.v(530)
  wire Axhow6;  // ../RTL/cortexm0ds_logic.v(1086)
  wire Axniu6;  // ../RTL/cortexm0ds_logic.v(623)
  wire Axohu6;  // ../RTL/cortexm0ds_logic.v(155)
  wire Axoow6;  // ../RTL/cortexm0ds_logic.v(1180)
  wire Axuiu6;  // ../RTL/cortexm0ds_logic.v(717)
  wire Axvhu6;  // ../RTL/cortexm0ds_logic.v(249)
  wire Axvow6;  // ../RTL/cortexm0ds_logic.v(1273)
  wire Ay0ju6;  // ../RTL/cortexm0ds_logic.v(797)
  wire Ay1iu6;  // ../RTL/cortexm0ds_logic.v(329)
  wire Ay1pw6;  // ../RTL/cortexm0ds_logic.v(1354)
  wire Ay7ju6;  // ../RTL/cortexm0ds_logic.v(891)
  wire Ay8iu6;  // ../RTL/cortexm0ds_logic.v(423)
  wire Ay8pw6;  // ../RTL/cortexm0ds_logic.v(1447)
  wire Ay9ow6;  // ../RTL/cortexm0ds_logic.v(979)
  wire Ayfiu6;  // ../RTL/cortexm0ds_logic.v(517)
  wire Aygow6;  // ../RTL/cortexm0ds_logic.v(1073)
  wire Aylhu6;  // ../RTL/cortexm0ds_logic.v(141)
  wire Aymiu6;  // ../RTL/cortexm0ds_logic.v(610)
  wire Aynow6;  // ../RTL/cortexm0ds_logic.v(1167)
  wire Aytiu6;  // ../RTL/cortexm0ds_logic.v(704)
  wire Ayuhu6;  // ../RTL/cortexm0ds_logic.v(236)
  wire Ayuow6;  // ../RTL/cortexm0ds_logic.v(1260)
  wire Az0iu6;  // ../RTL/cortexm0ds_logic.v(316)
  wire Az0pw6;  // ../RTL/cortexm0ds_logic.v(1341)
  wire Az3bx6;  // ../RTL/cortexm0ds_logic.v(1686)
  wire Az6ju6;  // ../RTL/cortexm0ds_logic.v(878)
  wire Az7iu6;  // ../RTL/cortexm0ds_logic.v(410)
  wire Az7pw6;  // ../RTL/cortexm0ds_logic.v(1434)
  wire Az8ow6;  // ../RTL/cortexm0ds_logic.v(966)
  wire Azeiu6;  // ../RTL/cortexm0ds_logic.v(504)
  wire Azfow6;  // ../RTL/cortexm0ds_logic.v(1060)
  wire Azliu6;  // ../RTL/cortexm0ds_logic.v(597)
  wire Azmow6;  // ../RTL/cortexm0ds_logic.v(1154)
  wire Azpax6;  // ../RTL/cortexm0ds_logic.v(1661)
  wire Azsiu6;  // ../RTL/cortexm0ds_logic.v(691)
  wire Azthu6;  // ../RTL/cortexm0ds_logic.v(223)
  wire Aztow6;  // ../RTL/cortexm0ds_logic.v(1247)
  wire Azziu6;  // ../RTL/cortexm0ds_logic.v(784)
  wire B03ju6;  // ../RTL/cortexm0ds_logic.v(825)
  wire B04iu6;  // ../RTL/cortexm0ds_logic.v(357)
  wire B04pw6;  // ../RTL/cortexm0ds_logic.v(1381)
  wire B0aju6;  // ../RTL/cortexm0ds_logic.v(918)
  wire B0biu6;  // ../RTL/cortexm0ds_logic.v(450)
  wire B0bpw6;  // ../RTL/cortexm0ds_logic.v(1475)
  wire B0cow6;  // ../RTL/cortexm0ds_logic.v(1007)
  wire B0iiu6;  // ../RTL/cortexm0ds_logic.v(544)
  wire B0jow6;  // ../RTL/cortexm0ds_logic.v(1100)
  wire B0piu6;  // ../RTL/cortexm0ds_logic.v(638)
  wire B0qhu6;  // ../RTL/cortexm0ds_logic.v(170)
  wire B0qow6;  // ../RTL/cortexm0ds_logic.v(1194)
  wire B0spw6;  // ../RTL/cortexm0ds_logic.v(1602)
  wire B0wiu6;  // ../RTL/cortexm0ds_logic.v(731)
  wire B0xhu6;  // ../RTL/cortexm0ds_logic.v(263)
  wire B0xow6;  // ../RTL/cortexm0ds_logic.v(1288)
  wire B12ju6;  // ../RTL/cortexm0ds_logic.v(812)
  wire B13iu6;  // ../RTL/cortexm0ds_logic.v(344)
  wire B13pw6;  // ../RTL/cortexm0ds_logic.v(1368)
  wire B19ju6;  // ../RTL/cortexm0ds_logic.v(905)
  wire B1aiu6;  // ../RTL/cortexm0ds_logic.v(437)
  wire B1apw6;  // ../RTL/cortexm0ds_logic.v(1462)
  wire B1bow6;  // ../RTL/cortexm0ds_logic.v(994)
  wire B1hiu6;  // ../RTL/cortexm0ds_logic.v(531)
  wire B1iow6;  // ../RTL/cortexm0ds_logic.v(1087)
  wire B1oiu6;  // ../RTL/cortexm0ds_logic.v(625)
  wire B1phu6;  // ../RTL/cortexm0ds_logic.v(157)
  wire B1pow6;  // ../RTL/cortexm0ds_logic.v(1181)
  wire B1viu6;  // ../RTL/cortexm0ds_logic.v(718)
  wire B1whu6;  // ../RTL/cortexm0ds_logic.v(250)
  wire B1wow6;  // ../RTL/cortexm0ds_logic.v(1275)
  wire B21ju6;  // ../RTL/cortexm0ds_logic.v(799)
  wire B22iu6;  // ../RTL/cortexm0ds_logic.v(331)
  wire B22pw6;  // ../RTL/cortexm0ds_logic.v(1355)
  wire B28ju6;  // ../RTL/cortexm0ds_logic.v(892)
  wire B29iu6;  // ../RTL/cortexm0ds_logic.v(424)
  wire B29pw6;  // ../RTL/cortexm0ds_logic.v(1449)
  wire B2aow6;  // ../RTL/cortexm0ds_logic.v(981)
  wire B2giu6;  // ../RTL/cortexm0ds_logic.v(518)
  wire B2how6;  // ../RTL/cortexm0ds_logic.v(1074)
  wire B2niu6;  // ../RTL/cortexm0ds_logic.v(612)
  wire B2oow6;  // ../RTL/cortexm0ds_logic.v(1168)
  wire B2uiu6;  // ../RTL/cortexm0ds_logic.v(705)
  wire B2vhu6;  // ../RTL/cortexm0ds_logic.v(237)
  wire B2vow6;  // ../RTL/cortexm0ds_logic.v(1262)
  wire B30ju6;  // ../RTL/cortexm0ds_logic.v(786)
  wire B31iu6;  // ../RTL/cortexm0ds_logic.v(318)
  wire B31pw6;  // ../RTL/cortexm0ds_logic.v(1342)
  wire B37ju6;  // ../RTL/cortexm0ds_logic.v(879)
  wire B38iu6;  // ../RTL/cortexm0ds_logic.v(411)
  wire B38pw6;  // ../RTL/cortexm0ds_logic.v(1436)
  wire B39ow6;  // ../RTL/cortexm0ds_logic.v(968)
  wire B3fiu6;  // ../RTL/cortexm0ds_logic.v(505)
  wire B3gbx6;  // ../RTL/cortexm0ds_logic.v(1708)
  wire B3gow6;  // ../RTL/cortexm0ds_logic.v(1061)
  wire B3miu6;  // ../RTL/cortexm0ds_logic.v(599)
  wire B3now6;  // ../RTL/cortexm0ds_logic.v(1155)
  wire B3tiu6;  // ../RTL/cortexm0ds_logic.v(692)
  wire B3uhu6;  // ../RTL/cortexm0ds_logic.v(224)
  wire B3uow6;  // ../RTL/cortexm0ds_logic.v(1249)
  wire B40iu6;  // ../RTL/cortexm0ds_logic.v(305)
  wire B40pw6;  // ../RTL/cortexm0ds_logic.v(1329)
  wire B46ju6;  // ../RTL/cortexm0ds_logic.v(866)
  wire B47iu6;  // ../RTL/cortexm0ds_logic.v(398)
  wire B47pw6;  // ../RTL/cortexm0ds_logic.v(1423)
  wire B48ow6;  // ../RTL/cortexm0ds_logic.v(955)
  wire B4eiu6;  // ../RTL/cortexm0ds_logic.v(492)
  wire B4epw6;  // ../RTL/cortexm0ds_logic.v(1516)
  wire B4fow6;  // ../RTL/cortexm0ds_logic.v(1048)
  wire B4liu6;  // ../RTL/cortexm0ds_logic.v(586)
  wire B4mow6;  // ../RTL/cortexm0ds_logic.v(1142)
  wire B4siu6;  // ../RTL/cortexm0ds_logic.v(679)
  wire B4thu6;  // ../RTL/cortexm0ds_logic.v(211)
  wire B4tow6;  // ../RTL/cortexm0ds_logic.v(1236)
  wire B4uax6;  // ../RTL/cortexm0ds_logic.v(1669)
  wire B4ziu6;  // ../RTL/cortexm0ds_logic.v(773)
  wire B55ju6;  // ../RTL/cortexm0ds_logic.v(853)
  wire B56iu6;  // ../RTL/cortexm0ds_logic.v(385)
  wire B56pw6;  // ../RTL/cortexm0ds_logic.v(1410)
  wire B57ow6;  // ../RTL/cortexm0ds_logic.v(942)
  wire B5diu6;  // ../RTL/cortexm0ds_logic.v(479)
  wire B5dpw6;  // ../RTL/cortexm0ds_logic.v(1503)
  wire B5eow6;  // ../RTL/cortexm0ds_logic.v(1035)
  wire B5kiu6;  // ../RTL/cortexm0ds_logic.v(573)
  wire B5low6;  // ../RTL/cortexm0ds_logic.v(1129)
  wire B5riu6;  // ../RTL/cortexm0ds_logic.v(666)
  wire B5shu6;  // ../RTL/cortexm0ds_logic.v(198)
  wire B5sow6;  // ../RTL/cortexm0ds_logic.v(1223)
  wire B5yiu6;  // ../RTL/cortexm0ds_logic.v(760)
  wire B5zhu6;  // ../RTL/cortexm0ds_logic.v(292)
  wire B5zow6;  // ../RTL/cortexm0ds_logic.v(1316)
  wire B5zpw6;  // ../RTL/cortexm0ds_logic.v(1615)
  wire B64ju6;  // ../RTL/cortexm0ds_logic.v(840)
  wire B65iu6;  // ../RTL/cortexm0ds_logic.v(372)
  wire B65pw6;  // ../RTL/cortexm0ds_logic.v(1397)
  wire B6ciu6;  // ../RTL/cortexm0ds_logic.v(466)
  wire B6cpw6;  // ../RTL/cortexm0ds_logic.v(1490)
  wire B6dow6;  // ../RTL/cortexm0ds_logic.v(1022)
  wire B6jiu6;  // ../RTL/cortexm0ds_logic.v(560)
  wire B6kow6;  // ../RTL/cortexm0ds_logic.v(1116)
  wire B6qiu6;  // ../RTL/cortexm0ds_logic.v(653)
  wire B6rhu6;  // ../RTL/cortexm0ds_logic.v(185)
  wire B6row6;  // ../RTL/cortexm0ds_logic.v(1210)
  wire B6uax6;  // ../RTL/cortexm0ds_logic.v(1669)
  wire B6xiu6;  // ../RTL/cortexm0ds_logic.v(747)
  wire B6yhu6;  // ../RTL/cortexm0ds_logic.v(279)
  wire B6yow6;  // ../RTL/cortexm0ds_logic.v(1303)
  wire B73ju6;  // ../RTL/cortexm0ds_logic.v(827)
  wire B74iu6;  // ../RTL/cortexm0ds_logic.v(359)
  wire B74pw6;  // ../RTL/cortexm0ds_logic.v(1384)
  wire B79bx6;  // ../RTL/cortexm0ds_logic.v(1696)
  wire B7aju6;  // ../RTL/cortexm0ds_logic.v(921)
  wire B7biu6;  // ../RTL/cortexm0ds_logic.v(453)
  wire B7bpw6;  // ../RTL/cortexm0ds_logic.v(1477)
  wire B7cow6;  // ../RTL/cortexm0ds_logic.v(1009)
  wire B7iiu6;  // ../RTL/cortexm0ds_logic.v(547)
  wire B7jow6;  // ../RTL/cortexm0ds_logic.v(1103)
  wire B7lpw6;  // ../RTL/cortexm0ds_logic.v(1590)
  wire B7nhu6;  // ../RTL/cortexm0ds_logic.v(144)
  wire B7piu6;  // ../RTL/cortexm0ds_logic.v(640)
  wire B7qhu6;  // ../RTL/cortexm0ds_logic.v(172)
  wire B7qow6;  // ../RTL/cortexm0ds_logic.v(1197)
  wire B7wiu6;  // ../RTL/cortexm0ds_logic.v(734)
  wire B7xhu6;  // ../RTL/cortexm0ds_logic.v(266)
  wire B7xow6;  // ../RTL/cortexm0ds_logic.v(1290)
  wire B82ju6;  // ../RTL/cortexm0ds_logic.v(814)
  wire B83iu6;  // ../RTL/cortexm0ds_logic.v(346)
  wire B83pw6;  // ../RTL/cortexm0ds_logic.v(1371)
  wire B89ju6;  // ../RTL/cortexm0ds_logic.v(908)
  wire B8aiu6;  // ../RTL/cortexm0ds_logic.v(440)
  wire B8apw6;  // ../RTL/cortexm0ds_logic.v(1464)
  wire B8bow6;  // ../RTL/cortexm0ds_logic.v(996)
  wire B8hiu6;  // ../RTL/cortexm0ds_logic.v(534)
  wire B8iow6;  // ../RTL/cortexm0ds_logic.v(1090)
  wire B8oiu6;  // ../RTL/cortexm0ds_logic.v(627)
  wire B8phu6;  // ../RTL/cortexm0ds_logic.v(159)
  wire B8pow6;  // ../RTL/cortexm0ds_logic.v(1184)
  wire B8uax6;  // ../RTL/cortexm0ds_logic.v(1669)
  wire B8viu6;  // ../RTL/cortexm0ds_logic.v(721)
  wire B8whu6;  // ../RTL/cortexm0ds_logic.v(253)
  wire B8wow6;  // ../RTL/cortexm0ds_logic.v(1277)
  wire B91ju6;  // ../RTL/cortexm0ds_logic.v(801)
  wire B92iu6;  // ../RTL/cortexm0ds_logic.v(333)
  wire B92pw6;  // ../RTL/cortexm0ds_logic.v(1358)
  wire B98ju6;  // ../RTL/cortexm0ds_logic.v(895)
  wire B99iu6;  // ../RTL/cortexm0ds_logic.v(427)
  wire B99pw6;  // ../RTL/cortexm0ds_logic.v(1451)
  wire B9aow6;  // ../RTL/cortexm0ds_logic.v(983)
  wire B9eax6;  // ../RTL/cortexm0ds_logic.v(1639)
  wire B9giu6;  // ../RTL/cortexm0ds_logic.v(521)
  wire B9how6;  // ../RTL/cortexm0ds_logic.v(1077)
  wire B9jbx6;  // ../RTL/cortexm0ds_logic.v(1714)
  wire B9niu6;  // ../RTL/cortexm0ds_logic.v(614)
  wire B9oow6;  // ../RTL/cortexm0ds_logic.v(1171)
  wire B9uiu6;  // ../RTL/cortexm0ds_logic.v(708)
  wire B9vhu6;  // ../RTL/cortexm0ds_logic.v(240)
  wire B9vow6;  // ../RTL/cortexm0ds_logic.v(1264)
  wire Ba0ju6;  // ../RTL/cortexm0ds_logic.v(788)
  wire Ba1iu6;  // ../RTL/cortexm0ds_logic.v(320)
  wire Ba1pw6;  // ../RTL/cortexm0ds_logic.v(1345)
  wire Ba7ju6;  // ../RTL/cortexm0ds_logic.v(882)
  wire Ba8iu6;  // ../RTL/cortexm0ds_logic.v(414)
  wire Ba8pw6;  // ../RTL/cortexm0ds_logic.v(1438)
  wire Ba9ow6;  // ../RTL/cortexm0ds_logic.v(970)
  wire Bafiu6;  // ../RTL/cortexm0ds_logic.v(508)
  wire Bagow6;  // ../RTL/cortexm0ds_logic.v(1064)
  wire Bamiu6;  // ../RTL/cortexm0ds_logic.v(601)
  wire Banow6;  // ../RTL/cortexm0ds_logic.v(1158)
  wire Batiu6;  // ../RTL/cortexm0ds_logic.v(695)
  wire Bauax6;  // ../RTL/cortexm0ds_logic.v(1669)
  wire Bauhu6;  // ../RTL/cortexm0ds_logic.v(227)
  wire Bauow6;  // ../RTL/cortexm0ds_logic.v(1251)
  wire Bb0iu6;  // ../RTL/cortexm0ds_logic.v(307)
  wire Bb0pw6;  // ../RTL/cortexm0ds_logic.v(1332)
  wire Bb6ju6;  // ../RTL/cortexm0ds_logic.v(869)
  wire Bb7iu6;  // ../RTL/cortexm0ds_logic.v(401)
  wire Bb7pw6;  // ../RTL/cortexm0ds_logic.v(1425)
  wire Bb8ow6;  // ../RTL/cortexm0ds_logic.v(957)
  wire Bbeiu6;  // ../RTL/cortexm0ds_logic.v(495)
  wire Bbfow6;  // ../RTL/cortexm0ds_logic.v(1051)
  wire Bbjpw6;  // ../RTL/cortexm0ds_logic.v(1586)
  wire Bbliu6;  // ../RTL/cortexm0ds_logic.v(588)
  wire Bbmow6;  // ../RTL/cortexm0ds_logic.v(1145)
  wire Bbsiu6;  // ../RTL/cortexm0ds_logic.v(682)
  wire Bbthu6;  // ../RTL/cortexm0ds_logic.v(214)
  wire Bbtow6;  // ../RTL/cortexm0ds_logic.v(1238)
  wire Bbziu6;  // ../RTL/cortexm0ds_logic.v(775)
  wire Bc3bx6;  // ../RTL/cortexm0ds_logic.v(1685)
  wire Bc5ju6;  // ../RTL/cortexm0ds_logic.v(856)
  wire Bc6iu6;  // ../RTL/cortexm0ds_logic.v(388)
  wire Bc6pw6;  // ../RTL/cortexm0ds_logic.v(1412)
  wire Bc7ow6;  // ../RTL/cortexm0ds_logic.v(944)
  wire Bcabx6;  // ../RTL/cortexm0ds_logic.v(1698)
  wire Bccax6;  // ../RTL/cortexm0ds_logic.v(1636)
  wire Bcdbx6;  // ../RTL/cortexm0ds_logic.v(1703)
  wire Bcdiu6;  // ../RTL/cortexm0ds_logic.v(482)
  wire Bcdpw6;  // ../RTL/cortexm0ds_logic.v(1506)
  wire Bceow6;  // ../RTL/cortexm0ds_logic.v(1038)
  wire Bcgax6;  // ../RTL/cortexm0ds_logic.v(1643)
  wire Bciax6;  // ../RTL/cortexm0ds_logic.v(1647)
  wire Bckiu6;  // ../RTL/cortexm0ds_logic.v(575)
  wire Bclow6;  // ../RTL/cortexm0ds_logic.v(1132)
  wire Bclpw6;  // ../RTL/cortexm0ds_logic.v(1590)
  wire Bcriu6;  // ../RTL/cortexm0ds_logic.v(669)
  wire Bcshu6;  // ../RTL/cortexm0ds_logic.v(201)
  wire Bcsow6;  // ../RTL/cortexm0ds_logic.v(1225)
  wire Bcyiu6;  // ../RTL/cortexm0ds_logic.v(762)
  wire Bczhu6;  // ../RTL/cortexm0ds_logic.v(294)
  wire Bczow6;  // ../RTL/cortexm0ds_logic.v(1319)
  wire Bd4ju6;  // ../RTL/cortexm0ds_logic.v(843)
  wire Bd5iu6;  // ../RTL/cortexm0ds_logic.v(375)
  wire Bd5pw6;  // ../RTL/cortexm0ds_logic.v(1399)
  wire Bd6ow6;  // ../RTL/cortexm0ds_logic.v(931)
  wire Bdciu6;  // ../RTL/cortexm0ds_logic.v(469)
  wire Bdcpw6;  // ../RTL/cortexm0ds_logic.v(1493)
  wire Bddow6;  // ../RTL/cortexm0ds_logic.v(1025)
  wire Bdjiu6;  // ../RTL/cortexm0ds_logic.v(562)
  wire Bdjpw6;  // ../RTL/cortexm0ds_logic.v(1586)
  wire Bdkow6;  // ../RTL/cortexm0ds_logic.v(1119)
  wire Bdqiu6;  // ../RTL/cortexm0ds_logic.v(656)
  wire Bdrhu6;  // ../RTL/cortexm0ds_logic.v(188)
  wire Bdrow6;  // ../RTL/cortexm0ds_logic.v(1212)
  wire Bdxiu6;  // ../RTL/cortexm0ds_logic.v(749)
  wire Bdyhu6;  // ../RTL/cortexm0ds_logic.v(281)
  wire Bdyow6;  // ../RTL/cortexm0ds_logic.v(1306)
  wire Be3ju6;  // ../RTL/cortexm0ds_logic.v(830)
  wire Be4iu6;  // ../RTL/cortexm0ds_logic.v(362)
  wire Be4pw6;  // ../RTL/cortexm0ds_logic.v(1386)
  wire Beaju6;  // ../RTL/cortexm0ds_logic.v(924)
  wire Bebiu6;  // ../RTL/cortexm0ds_logic.v(456)
  wire Bebpw6;  // ../RTL/cortexm0ds_logic.v(1480)
  wire Becow6;  // ../RTL/cortexm0ds_logic.v(1012)
  wire Beiiu6;  // ../RTL/cortexm0ds_logic.v(549)
  wire Bejow6;  // ../RTL/cortexm0ds_logic.v(1106)
  wire Bepiu6;  // ../RTL/cortexm0ds_logic.v(643)
  wire Beqhu6;  // ../RTL/cortexm0ds_logic.v(175)
  wire Beqow6;  // ../RTL/cortexm0ds_logic.v(1199)
  wire Bewiu6;  // ../RTL/cortexm0ds_logic.v(736)
  wire Bexhu6;  // ../RTL/cortexm0ds_logic.v(268)
  wire Bexow6;  // ../RTL/cortexm0ds_logic.v(1293)
  wire Bf2ju6;  // ../RTL/cortexm0ds_logic.v(817)
  wire Bf3iu6;  // ../RTL/cortexm0ds_logic.v(349)
  wire Bf3pw6;  // ../RTL/cortexm0ds_logic.v(1373)
  wire Bf3qw6;  // ../RTL/cortexm0ds_logic.v(1623)
  wire Bf9ju6;  // ../RTL/cortexm0ds_logic.v(911)
  wire Bfaiu6;  // ../RTL/cortexm0ds_logic.v(443)
  wire Bfapw6;  // ../RTL/cortexm0ds_logic.v(1467)
  wire Bfbow6;  // ../RTL/cortexm0ds_logic.v(999)
  wire Bfhiu6;  // ../RTL/cortexm0ds_logic.v(536)
  wire Bfiow6;  // ../RTL/cortexm0ds_logic.v(1093)
  wire Bfjpw6;  // ../RTL/cortexm0ds_logic.v(1586)
  wire Bfoiu6;  // ../RTL/cortexm0ds_logic.v(630)
  wire Bfphu6;  // ../RTL/cortexm0ds_logic.v(162)
  wire Bfpow6;  // ../RTL/cortexm0ds_logic.v(1186)
  wire Bfviu6;  // ../RTL/cortexm0ds_logic.v(723)
  wire Bfwhu6;  // ../RTL/cortexm0ds_logic.v(255)
  wire Bfwow6;  // ../RTL/cortexm0ds_logic.v(1280)
  wire Bg1ju6;  // ../RTL/cortexm0ds_logic.v(804)
  wire Bg2iu6;  // ../RTL/cortexm0ds_logic.v(336)
  wire Bg2pw6;  // ../RTL/cortexm0ds_logic.v(1360)
  wire Bg8ju6;  // ../RTL/cortexm0ds_logic.v(898)
  wire Bg9iu6;  // ../RTL/cortexm0ds_logic.v(430)
  wire Bg9pw6;  // ../RTL/cortexm0ds_logic.v(1454)
  wire Bgaow6;  // ../RTL/cortexm0ds_logic.v(986)
  wire Bggiu6;  // ../RTL/cortexm0ds_logic.v(523)
  wire Bghow6;  // ../RTL/cortexm0ds_logic.v(1080)
  wire Bgniu6;  // ../RTL/cortexm0ds_logic.v(617)
  wire Bgohu6;  // ../RTL/cortexm0ds_logic.v(149)
  wire Bgoow6;  // ../RTL/cortexm0ds_logic.v(1173)
  wire Bguiu6;  // ../RTL/cortexm0ds_logic.v(710)
  wire Bgvhu6;  // ../RTL/cortexm0ds_logic.v(242)
  wire Bgvow6;  // ../RTL/cortexm0ds_logic.v(1267)
  wire Bh0ju6;  // ../RTL/cortexm0ds_logic.v(791)
  wire Bh1iu6;  // ../RTL/cortexm0ds_logic.v(323)
  wire Bh1pw6;  // ../RTL/cortexm0ds_logic.v(1347)
  wire Bh7ju6;  // ../RTL/cortexm0ds_logic.v(885)
  wire Bh8iu6;  // ../RTL/cortexm0ds_logic.v(417)
  wire Bh8pw6;  // ../RTL/cortexm0ds_logic.v(1441)
  wire Bh9ow6;  // ../RTL/cortexm0ds_logic.v(973)
  wire Bhfiu6;  // ../RTL/cortexm0ds_logic.v(510)
  wire Bhgow6;  // ../RTL/cortexm0ds_logic.v(1067)
  wire Bhmhu6;  // ../RTL/cortexm0ds_logic.v(142)
  wire Bhmiu6;  // ../RTL/cortexm0ds_logic.v(604)
  wire Bhnow6;  // ../RTL/cortexm0ds_logic.v(1160)
  wire Bhtiu6;  // ../RTL/cortexm0ds_logic.v(697)
  wire Bhuhu6;  // ../RTL/cortexm0ds_logic.v(229)
  wire Bhuow6;  // ../RTL/cortexm0ds_logic.v(1254)
  wire Bi0iu6;  // ../RTL/cortexm0ds_logic.v(310)
  wire Bi0pw6;  // ../RTL/cortexm0ds_logic.v(1334)
  wire Bi6ju6;  // ../RTL/cortexm0ds_logic.v(872)
  wire Bi7iu6;  // ../RTL/cortexm0ds_logic.v(404)
  wire Bi7pw6;  // ../RTL/cortexm0ds_logic.v(1428)
  wire Bi8ow6;  // ../RTL/cortexm0ds_logic.v(960)
  wire Biaax6;  // ../RTL/cortexm0ds_logic.v(1632)
  wire Bieiu6;  // ../RTL/cortexm0ds_logic.v(497)
  wire Bifow6;  // ../RTL/cortexm0ds_logic.v(1054)
  wire Biliu6;  // ../RTL/cortexm0ds_logic.v(591)
  wire Bimow6;  // ../RTL/cortexm0ds_logic.v(1147)
  wire Bisiu6;  // ../RTL/cortexm0ds_logic.v(684)
  wire Bithu6;  // ../RTL/cortexm0ds_logic.v(216)
  wire Bitow6;  // ../RTL/cortexm0ds_logic.v(1241)
  wire Biziu6;  // ../RTL/cortexm0ds_logic.v(778)
  wire Bj5ju6;  // ../RTL/cortexm0ds_logic.v(859)
  wire Bj6iu6;  // ../RTL/cortexm0ds_logic.v(391)
  wire Bj6pw6;  // ../RTL/cortexm0ds_logic.v(1415)
  wire Bj7ow6;  // ../RTL/cortexm0ds_logic.v(947)
  wire Bjdiu6;  // ../RTL/cortexm0ds_logic.v(484)
  wire Bjdpw6;  // ../RTL/cortexm0ds_logic.v(1509)
  wire Bjeow6;  // ../RTL/cortexm0ds_logic.v(1041)
  wire Bjkiu6;  // ../RTL/cortexm0ds_logic.v(578)
  wire Bjlow6;  // ../RTL/cortexm0ds_logic.v(1134)
  wire Bjriu6;  // ../RTL/cortexm0ds_logic.v(671)
  wire Bjshu6;  // ../RTL/cortexm0ds_logic.v(203)
  wire Bjsow6;  // ../RTL/cortexm0ds_logic.v(1228)
  wire Bjyiu6;  // ../RTL/cortexm0ds_logic.v(765)
  wire Bjzhu6;  // ../RTL/cortexm0ds_logic.v(297)
  wire Bjzow6;  // ../RTL/cortexm0ds_logic.v(1321)
  wire Bk4ju6;  // ../RTL/cortexm0ds_logic.v(846)
  wire Bk5iu6;  // ../RTL/cortexm0ds_logic.v(378)
  wire Bk5pw6;  // ../RTL/cortexm0ds_logic.v(1402)
  wire Bk6ow6;  // ../RTL/cortexm0ds_logic.v(934)
  wire Bk7ax6;  // ../RTL/cortexm0ds_logic.v(1627)
  wire Bkciu6;  // ../RTL/cortexm0ds_logic.v(471)
  wire Bkcpw6;  // ../RTL/cortexm0ds_logic.v(1496)
  wire Bkdow6;  // ../RTL/cortexm0ds_logic.v(1028)
  wire Bkjiu6;  // ../RTL/cortexm0ds_logic.v(565)
  wire Bkkow6;  // ../RTL/cortexm0ds_logic.v(1121)
  wire Bklhu6;  // ../RTL/cortexm0ds_logic.v(139)
  wire Bkqiu6;  // ../RTL/cortexm0ds_logic.v(658)
  wire Bkrhu6;  // ../RTL/cortexm0ds_logic.v(190)
  wire Bkrow6;  // ../RTL/cortexm0ds_logic.v(1215)
  wire Bkxiu6;  // ../RTL/cortexm0ds_logic.v(752)
  wire Bkyhu6;  // ../RTL/cortexm0ds_logic.v(284)
  wire Bkyow6;  // ../RTL/cortexm0ds_logic.v(1308)
  wire Bl3ju6;  // ../RTL/cortexm0ds_logic.v(833)
  wire Bl4iu6;  // ../RTL/cortexm0ds_logic.v(365)
  wire Bl4pw6;  // ../RTL/cortexm0ds_logic.v(1389)
  wire Blaju6;  // ../RTL/cortexm0ds_logic.v(926)
  wire Blbiu6;  // ../RTL/cortexm0ds_logic.v(458)
  wire Blbpw6;  // ../RTL/cortexm0ds_logic.v(1483)
  wire Blcow6;  // ../RTL/cortexm0ds_logic.v(1015)
  wire Bliiu6;  // ../RTL/cortexm0ds_logic.v(552)
  wire Bljow6;  // ../RTL/cortexm0ds_logic.v(1108)
  wire Blpiu6;  // ../RTL/cortexm0ds_logic.v(645)
  wire Blqhu6;  // ../RTL/cortexm0ds_logic.v(177)
  wire Blqow6;  // ../RTL/cortexm0ds_logic.v(1202)
  wire Blwiu6;  // ../RTL/cortexm0ds_logic.v(739)
  wire Blxhu6;  // ../RTL/cortexm0ds_logic.v(271)
  wire Blxow6;  // ../RTL/cortexm0ds_logic.v(1295)
  wire Bm2ju6;  // ../RTL/cortexm0ds_logic.v(820)
  wire Bm3iu6;  // ../RTL/cortexm0ds_logic.v(352)
  wire Bm3pw6;  // ../RTL/cortexm0ds_logic.v(1376)
  wire Bm9ju6;  // ../RTL/cortexm0ds_logic.v(913)
  wire Bmaiu6;  // ../RTL/cortexm0ds_logic.v(445)
  wire Bmapw6;  // ../RTL/cortexm0ds_logic.v(1470)
  wire Bmbow6;  // ../RTL/cortexm0ds_logic.v(1002)
  wire Bmhiu6;  // ../RTL/cortexm0ds_logic.v(539)
  wire Bmiow6;  // ../RTL/cortexm0ds_logic.v(1095)
  wire Bmoiu6;  // ../RTL/cortexm0ds_logic.v(632)
  wire Bmphu6;  // ../RTL/cortexm0ds_logic.v(164)
  wire Bmpow6;  // ../RTL/cortexm0ds_logic.v(1189)
  wire Bmviu6;  // ../RTL/cortexm0ds_logic.v(726)
  wire Bmwhu6;  // ../RTL/cortexm0ds_logic.v(258)
  wire Bmwow6;  // ../RTL/cortexm0ds_logic.v(1282)
  wire Bn1ju6;  // ../RTL/cortexm0ds_logic.v(807)
  wire Bn2iu6;  // ../RTL/cortexm0ds_logic.v(339)
  wire Bn2pw6;  // ../RTL/cortexm0ds_logic.v(1363)
  wire Bn8ju6;  // ../RTL/cortexm0ds_logic.v(900)
  wire Bn9iu6;  // ../RTL/cortexm0ds_logic.v(432)
  wire Bn9pw6;  // ../RTL/cortexm0ds_logic.v(1457)
  wire Bnaow6;  // ../RTL/cortexm0ds_logic.v(989)
  wire Bngax6;  // ../RTL/cortexm0ds_logic.v(1644)
  wire Bngiu6;  // ../RTL/cortexm0ds_logic.v(526)
  wire Bnhow6;  // ../RTL/cortexm0ds_logic.v(1082)
  wire Bnniu6;  // ../RTL/cortexm0ds_logic.v(619)
  wire Bnohu6;  // ../RTL/cortexm0ds_logic.v(151)
  wire Bnoow6;  // ../RTL/cortexm0ds_logic.v(1176)
  wire Bnuiu6;  // ../RTL/cortexm0ds_logic.v(713)
  wire Bnvhu6;  // ../RTL/cortexm0ds_logic.v(245)
  wire Bnvow6;  // ../RTL/cortexm0ds_logic.v(1269)
  wire Bo0ju6;  // ../RTL/cortexm0ds_logic.v(794)
  wire Bo1iu6;  // ../RTL/cortexm0ds_logic.v(326)
  wire Bo1pw6;  // ../RTL/cortexm0ds_logic.v(1350)
  wire Bo7ju6;  // ../RTL/cortexm0ds_logic.v(887)
  wire Bo8iu6;  // ../RTL/cortexm0ds_logic.v(419)
  wire Bo8pw6;  // ../RTL/cortexm0ds_logic.v(1444)
  wire Bo9ow6;  // ../RTL/cortexm0ds_logic.v(976)
  wire Bofiu6;  // ../RTL/cortexm0ds_logic.v(513)
  wire Bogow6;  // ../RTL/cortexm0ds_logic.v(1069)
  wire Bolax6;  // ../RTL/cortexm0ds_logic.v(1653)
  wire Bomiu6;  // ../RTL/cortexm0ds_logic.v(606)
  wire Bonow6;  // ../RTL/cortexm0ds_logic.v(1163)
  wire Botiu6;  // ../RTL/cortexm0ds_logic.v(700)
  wire Bouhu6;  // ../RTL/cortexm0ds_logic.v(232)
  wire Bouow6;  // ../RTL/cortexm0ds_logic.v(1256)
  wire Bp0iu6;  // ../RTL/cortexm0ds_logic.v(313)
  wire Bp0pw6;  // ../RTL/cortexm0ds_logic.v(1337)
  wire Bp2qw6;  // ../RTL/cortexm0ds_logic.v(1622)
  wire Bp6ju6;  // ../RTL/cortexm0ds_logic.v(874)
  wire Bp7iu6;  // ../RTL/cortexm0ds_logic.v(406)
  wire Bp7pw6;  // ../RTL/cortexm0ds_logic.v(1431)
  wire Bp8ow6;  // ../RTL/cortexm0ds_logic.v(963)
  wire Bpeiu6;  // ../RTL/cortexm0ds_logic.v(500)
  wire Bpfow6;  // ../RTL/cortexm0ds_logic.v(1056)
  wire Bpliu6;  // ../RTL/cortexm0ds_logic.v(593)
  wire Bpmow6;  // ../RTL/cortexm0ds_logic.v(1150)
  wire Bpsiu6;  // ../RTL/cortexm0ds_logic.v(687)
  wire Bpthu6;  // ../RTL/cortexm0ds_logic.v(219)
  wire Bptow6;  // ../RTL/cortexm0ds_logic.v(1243)
  wire Bpziu6;  // ../RTL/cortexm0ds_logic.v(781)
  wire Bq5ju6;  // ../RTL/cortexm0ds_logic.v(861)
  wire Bq6iu6;  // ../RTL/cortexm0ds_logic.v(393)
  wire Bq6pw6;  // ../RTL/cortexm0ds_logic.v(1418)
  wire Bq7ow6;  // ../RTL/cortexm0ds_logic.v(950)
  wire Bq9ax6;  // ../RTL/cortexm0ds_logic.v(1631)
  wire Bqdiu6;  // ../RTL/cortexm0ds_logic.v(487)
  wire Bqdpw6;  // ../RTL/cortexm0ds_logic.v(1511)
  wire Bqeow6;  // ../RTL/cortexm0ds_logic.v(1043)
  wire Bqkiu6;  // ../RTL/cortexm0ds_logic.v(580)
  wire Bqlow6;  // ../RTL/cortexm0ds_logic.v(1137)
  wire Bqriu6;  // ../RTL/cortexm0ds_logic.v(674)
  wire Bqshu6;  // ../RTL/cortexm0ds_logic.v(206)
  wire Bqsow6;  // ../RTL/cortexm0ds_logic.v(1230)
  wire Bqyiu6;  // ../RTL/cortexm0ds_logic.v(768)
  wire Bqzhu6;  // ../RTL/cortexm0ds_logic.v(300)
  wire Bqzow6;  // ../RTL/cortexm0ds_logic.v(1324)
  wire Br4ju6;  // ../RTL/cortexm0ds_logic.v(848)
  wire Br5iu6;  // ../RTL/cortexm0ds_logic.v(380)
  wire Br5pw6;  // ../RTL/cortexm0ds_logic.v(1405)
  wire Br6ow6;  // ../RTL/cortexm0ds_logic.v(937)
  wire Brciu6;  // ../RTL/cortexm0ds_logic.v(474)
  wire Brcpw6;  // ../RTL/cortexm0ds_logic.v(1498)
  wire Brdow6;  // ../RTL/cortexm0ds_logic.v(1030)
  wire Brjiu6;  // ../RTL/cortexm0ds_logic.v(567)
  wire Brkow6;  // ../RTL/cortexm0ds_logic.v(1124)
  wire Brqiu6;  // ../RTL/cortexm0ds_logic.v(661)
  wire Brrhu6;  // ../RTL/cortexm0ds_logic.v(193)
  wire Brrow6;  // ../RTL/cortexm0ds_logic.v(1217)
  wire Brxiu6;  // ../RTL/cortexm0ds_logic.v(755)
  wire Bryhu6;  // ../RTL/cortexm0ds_logic.v(287)
  wire Bryow6;  // ../RTL/cortexm0ds_logic.v(1311)
  wire Bs3ju6;  // ../RTL/cortexm0ds_logic.v(835)
  wire Bs4iu6;  // ../RTL/cortexm0ds_logic.v(367)
  wire Bs4pw6;  // ../RTL/cortexm0ds_logic.v(1392)
  wire Bsaju6;  // ../RTL/cortexm0ds_logic.v(929)
  wire Bsbiu6;  // ../RTL/cortexm0ds_logic.v(461)
  wire Bsbpw6;  // ../RTL/cortexm0ds_logic.v(1485)
  wire Bscow6;  // ../RTL/cortexm0ds_logic.v(1017)
  wire Bsiiu6;  // ../RTL/cortexm0ds_logic.v(554)
  wire Bsjow6;  // ../RTL/cortexm0ds_logic.v(1111)
  wire Bspiu6;  // ../RTL/cortexm0ds_logic.v(648)
  wire Bsqhu6;  // ../RTL/cortexm0ds_logic.v(180)
  wire Bsqow6;  // ../RTL/cortexm0ds_logic.v(1204)
  wire Bsrpw6;  // ../RTL/cortexm0ds_logic.v(1602)
  wire Bswiu6;  // ../RTL/cortexm0ds_logic.v(742)
  wire Bsxhu6;  // ../RTL/cortexm0ds_logic.v(274)
  wire Bsxow6;  // ../RTL/cortexm0ds_logic.v(1298)
  wire Bt2ju6;  // ../RTL/cortexm0ds_logic.v(822)
  wire Bt2qw6;  // ../RTL/cortexm0ds_logic.v(1622)
  wire Bt3iu6;  // ../RTL/cortexm0ds_logic.v(354)
  wire Bt3pw6;  // ../RTL/cortexm0ds_logic.v(1379)
  wire Bt9ju6;  // ../RTL/cortexm0ds_logic.v(916)
  wire Btaiu6;  // ../RTL/cortexm0ds_logic.v(448)
  wire Btapw6;  // ../RTL/cortexm0ds_logic.v(1472)
  wire Btbbx6;  // ../RTL/cortexm0ds_logic.v(1700)
  wire Btbow6;  // ../RTL/cortexm0ds_logic.v(1004)
  wire Bthiu6;  // ../RTL/cortexm0ds_logic.v(541)
  wire Btiow6;  // ../RTL/cortexm0ds_logic.v(1098)
  wire Btoiu6;  // ../RTL/cortexm0ds_logic.v(635)
  wire Btphu6;  // ../RTL/cortexm0ds_logic.v(167)
  wire Btpow6;  // ../RTL/cortexm0ds_logic.v(1191)
  wire Btviu6;  // ../RTL/cortexm0ds_logic.v(729)
  wire Btwhu6;  // ../RTL/cortexm0ds_logic.v(261)
  wire Btwow6;  // ../RTL/cortexm0ds_logic.v(1285)
  wire Bu1ju6;  // ../RTL/cortexm0ds_logic.v(809)
  wire Bu2iu6;  // ../RTL/cortexm0ds_logic.v(341)
  wire Bu2pw6;  // ../RTL/cortexm0ds_logic.v(1366)
  wire Bu6bx6;  // ../RTL/cortexm0ds_logic.v(1691)
  wire Bu8ju6;  // ../RTL/cortexm0ds_logic.v(903)
  wire Bu9iu6;  // ../RTL/cortexm0ds_logic.v(435)
  wire Bu9pw6;  // ../RTL/cortexm0ds_logic.v(1459)
  wire Buabx6;  // ../RTL/cortexm0ds_logic.v(1699)
  wire Buaow6;  // ../RTL/cortexm0ds_logic.v(991)
  wire Bugiu6;  // ../RTL/cortexm0ds_logic.v(528)
  wire Buhow6;  // ../RTL/cortexm0ds_logic.v(1085)
  wire Buniu6;  // ../RTL/cortexm0ds_logic.v(622)
  wire Buohu6;  // ../RTL/cortexm0ds_logic.v(154)
  wire Buoow6;  // ../RTL/cortexm0ds_logic.v(1178)
  wire Buuiu6;  // ../RTL/cortexm0ds_logic.v(716)
  wire Buvhu6;  // ../RTL/cortexm0ds_logic.v(248)
  wire Buvow6;  // ../RTL/cortexm0ds_logic.v(1272)
  wire Bv0ju6;  // ../RTL/cortexm0ds_logic.v(796)
  wire Bv1iu6;  // ../RTL/cortexm0ds_logic.v(328)
  wire Bv1pw6;  // ../RTL/cortexm0ds_logic.v(1353)
  wire Bv7ju6;  // ../RTL/cortexm0ds_logic.v(890)
  wire Bv8iu6;  // ../RTL/cortexm0ds_logic.v(422)
  wire Bv8pw6;  // ../RTL/cortexm0ds_logic.v(1446)
  wire Bv9ow6;  // ../RTL/cortexm0ds_logic.v(978)
  wire Bvaax6;  // ../RTL/cortexm0ds_logic.v(1633)
  wire Bvfbx6;  // ../RTL/cortexm0ds_logic.v(1708)
  wire Bvfiu6;  // ../RTL/cortexm0ds_logic.v(515)
  wire Bvgow6;  // ../RTL/cortexm0ds_logic.v(1072)
  wire Bvmiu6;  // ../RTL/cortexm0ds_logic.v(609)
  wire Bvnow6;  // ../RTL/cortexm0ds_logic.v(1165)
  wire Bvtiu6;  // ../RTL/cortexm0ds_logic.v(703)
  wire Bvuhu6;  // ../RTL/cortexm0ds_logic.v(235)
  wire Bvuow6;  // ../RTL/cortexm0ds_logic.v(1259)
  wire Bw0iu6;  // ../RTL/cortexm0ds_logic.v(315)
  wire Bw0pw6;  // ../RTL/cortexm0ds_logic.v(1340)
  wire Bw6ju6;  // ../RTL/cortexm0ds_logic.v(877)
  wire Bw7iu6;  // ../RTL/cortexm0ds_logic.v(409)
  wire Bw7pw6;  // ../RTL/cortexm0ds_logic.v(1433)
  wire Bw8ow6;  // ../RTL/cortexm0ds_logic.v(965)
  wire Bwdax6;  // ../RTL/cortexm0ds_logic.v(1639)
  wire Bweiu6;  // ../RTL/cortexm0ds_logic.v(502)
  wire Bwfow6;  // ../RTL/cortexm0ds_logic.v(1059)
  wire Bwliu6;  // ../RTL/cortexm0ds_logic.v(596)
  wire Bwmow6;  // ../RTL/cortexm0ds_logic.v(1152)
  wire Bwsiu6;  // ../RTL/cortexm0ds_logic.v(690)
  wire Bwthu6;  // ../RTL/cortexm0ds_logic.v(222)
  wire Bwtow6;  // ../RTL/cortexm0ds_logic.v(1246)
  wire Bwziu6;  // ../RTL/cortexm0ds_logic.v(783)
  wire Bx2qw6;  // ../RTL/cortexm0ds_logic.v(1622)
  wire Bx5ju6;  // ../RTL/cortexm0ds_logic.v(864)
  wire Bx6iu6;  // ../RTL/cortexm0ds_logic.v(396)
  wire Bx6pw6;  // ../RTL/cortexm0ds_logic.v(1420)
  wire Bx7ow6;  // ../RTL/cortexm0ds_logic.v(952)
  wire Bxbax6;  // ../RTL/cortexm0ds_logic.v(1635)
  wire Bxdiu6;  // ../RTL/cortexm0ds_logic.v(489)
  wire Bxdpw6;  // ../RTL/cortexm0ds_logic.v(1514)
  wire Bxeow6;  // ../RTL/cortexm0ds_logic.v(1046)
  wire Bxghu6;  // ../RTL/cortexm0ds_logic.v(127)
  wire Bxkiu6;  // ../RTL/cortexm0ds_logic.v(583)
  wire Bxlow6;  // ../RTL/cortexm0ds_logic.v(1139)
  wire Bxpax6;  // ../RTL/cortexm0ds_logic.v(1661)
  wire Bxriu6;  // ../RTL/cortexm0ds_logic.v(677)
  wire Bxshu6;  // ../RTL/cortexm0ds_logic.v(209)
  wire Bxsow6;  // ../RTL/cortexm0ds_logic.v(1233)
  wire Bxyiu6;  // ../RTL/cortexm0ds_logic.v(770)
  wire Bxzhu6;  // ../RTL/cortexm0ds_logic.v(302)
  wire Bxzow6;  // ../RTL/cortexm0ds_logic.v(1327)
  wire By4ju6;  // ../RTL/cortexm0ds_logic.v(851)
  wire By5iu6;  // ../RTL/cortexm0ds_logic.v(383)
  wire By5pw6;  // ../RTL/cortexm0ds_logic.v(1407)
  wire By6ow6;  // ../RTL/cortexm0ds_logic.v(939)
  wire Byciu6;  // ../RTL/cortexm0ds_logic.v(476)
  wire Bycpw6;  // ../RTL/cortexm0ds_logic.v(1501)
  wire Bydow6;  // ../RTL/cortexm0ds_logic.v(1033)
  wire Byjiu6;  // ../RTL/cortexm0ds_logic.v(570)
  wire Bykow6;  // ../RTL/cortexm0ds_logic.v(1126)
  wire Byqiu6;  // ../RTL/cortexm0ds_logic.v(664)
  wire Byrhu6;  // ../RTL/cortexm0ds_logic.v(196)
  wire Byrow6;  // ../RTL/cortexm0ds_logic.v(1220)
  wire Byxiu6;  // ../RTL/cortexm0ds_logic.v(757)
  wire Byyhu6;  // ../RTL/cortexm0ds_logic.v(289)
  wire Byyow6;  // ../RTL/cortexm0ds_logic.v(1314)
  wire Bz3ju6;  // ../RTL/cortexm0ds_logic.v(838)
  wire Bz4iu6;  // ../RTL/cortexm0ds_logic.v(370)
  wire Bz4pw6;  // ../RTL/cortexm0ds_logic.v(1394)
  wire Bzbiu6;  // ../RTL/cortexm0ds_logic.v(463)
  wire Bzbpw6;  // ../RTL/cortexm0ds_logic.v(1488)
  wire Bzcow6;  // ../RTL/cortexm0ds_logic.v(1020)
  wire Bziiu6;  // ../RTL/cortexm0ds_logic.v(557)
  wire Bzjow6;  // ../RTL/cortexm0ds_logic.v(1113)
  wire Bzpiu6;  // ../RTL/cortexm0ds_logic.v(651)
  wire Bzqhu6;  // ../RTL/cortexm0ds_logic.v(183)
  wire Bzqow6;  // ../RTL/cortexm0ds_logic.v(1207)
  wire Bzwiu6;  // ../RTL/cortexm0ds_logic.v(744)
  wire Bzxhu6;  // ../RTL/cortexm0ds_logic.v(276)
  wire Bzxow6;  // ../RTL/cortexm0ds_logic.v(1301)
  wire C00ju6;  // ../RTL/cortexm0ds_logic.v(785)
  wire C01iu6;  // ../RTL/cortexm0ds_logic.v(317)
  wire C01pw6;  // ../RTL/cortexm0ds_logic.v(1341)
  wire C07bx6;  // ../RTL/cortexm0ds_logic.v(1692)
  wire C07ju6;  // ../RTL/cortexm0ds_logic.v(878)
  wire C08iu6;  // ../RTL/cortexm0ds_logic.v(410)
  wire C08pw6;  // ../RTL/cortexm0ds_logic.v(1435)
  wire C09ow6;  // ../RTL/cortexm0ds_logic.v(967)
  wire C0ehu6;  // ../RTL/cortexm0ds_logic.v(121)
  wire C0fiu6;  // ../RTL/cortexm0ds_logic.v(504)
  wire C0gow6;  // ../RTL/cortexm0ds_logic.v(1060)
  wire C0khu6;  // ../RTL/cortexm0ds_logic.v(135)
  wire C0miu6;  // ../RTL/cortexm0ds_logic.v(598)
  wire C0now6;  // ../RTL/cortexm0ds_logic.v(1154)
  wire C0tiu6;  // ../RTL/cortexm0ds_logic.v(691)
  wire C0uhu6;  // ../RTL/cortexm0ds_logic.v(223)
  wire C0uow6;  // ../RTL/cortexm0ds_logic.v(1248)
  wire C10bx6;  // ../RTL/cortexm0ds_logic.v(1679)
  wire C10iu6;  // ../RTL/cortexm0ds_logic.v(304)
  wire C10pw6;  // ../RTL/cortexm0ds_logic.v(1328)
  wire C14bx6;  // ../RTL/cortexm0ds_logic.v(1686)
  wire C16ju6;  // ../RTL/cortexm0ds_logic.v(865)
  wire C17iu6;  // ../RTL/cortexm0ds_logic.v(397)
  wire C17pw6;  // ../RTL/cortexm0ds_logic.v(1422)
  wire C18ow6;  // ../RTL/cortexm0ds_logic.v(954)
  wire C1eiu6;  // ../RTL/cortexm0ds_logic.v(491)
  wire C1epw6;  // ../RTL/cortexm0ds_logic.v(1515)
  wire C1fax6;  // ../RTL/cortexm0ds_logic.v(1641)
  wire C1fow6;  // ../RTL/cortexm0ds_logic.v(1047)
  wire C1liu6;  // ../RTL/cortexm0ds_logic.v(585)
  wire C1mow6;  // ../RTL/cortexm0ds_logic.v(1141)
  wire C1siu6;  // ../RTL/cortexm0ds_logic.v(678)
  wire C1thu6;  // ../RTL/cortexm0ds_logic.v(210)
  wire C1tow6;  // ../RTL/cortexm0ds_logic.v(1235)
  wire C1wpw6;  // ../RTL/cortexm0ds_logic.v(1610)
  wire C1ziu6;  // ../RTL/cortexm0ds_logic.v(772)
  wire C25ju6;  // ../RTL/cortexm0ds_logic.v(852)
  wire C26iu6;  // ../RTL/cortexm0ds_logic.v(384)
  wire C26pw6;  // ../RTL/cortexm0ds_logic.v(1409)
  wire C27bx6;  // ../RTL/cortexm0ds_logic.v(1692)
  wire C27ow6;  // ../RTL/cortexm0ds_logic.v(941)
  wire C2diu6;  // ../RTL/cortexm0ds_logic.v(478)
  wire C2dpw6;  // ../RTL/cortexm0ds_logic.v(1502)
  wire C2eow6;  // ../RTL/cortexm0ds_logic.v(1034)
  wire C2jhu6;  // ../RTL/cortexm0ds_logic.v(133)
  wire C2kiu6;  // ../RTL/cortexm0ds_logic.v(572)
  wire C2low6;  // ../RTL/cortexm0ds_logic.v(1128)
  wire C2riu6;  // ../RTL/cortexm0ds_logic.v(665)
  wire C2shu6;  // ../RTL/cortexm0ds_logic.v(197)
  wire C2sow6;  // ../RTL/cortexm0ds_logic.v(1222)
  wire C2uax6;  // ../RTL/cortexm0ds_logic.v(1669)
  wire C2yiu6;  // ../RTL/cortexm0ds_logic.v(759)
  wire C2ypw6;  // ../RTL/cortexm0ds_logic.v(1613)
  wire C2zhu6;  // ../RTL/cortexm0ds_logic.v(291)
  wire C2zow6;  // ../RTL/cortexm0ds_logic.v(1315)
  wire C30bx6;  // ../RTL/cortexm0ds_logic.v(1679)
  wire C34ju6;  // ../RTL/cortexm0ds_logic.v(839)
  wire C35iu6;  // ../RTL/cortexm0ds_logic.v(371)
  wire C35pw6;  // ../RTL/cortexm0ds_logic.v(1396)
  wire C37ax6;  // ../RTL/cortexm0ds_logic.v(1626)
  wire C3ciu6;  // ../RTL/cortexm0ds_logic.v(465)
  wire C3cpw6;  // ../RTL/cortexm0ds_logic.v(1489)
  wire C3dow6;  // ../RTL/cortexm0ds_logic.v(1021)
  wire C3jiu6;  // ../RTL/cortexm0ds_logic.v(559)
  wire C3kow6;  // ../RTL/cortexm0ds_logic.v(1115)
  wire C3mhu6;  // ../RTL/cortexm0ds_logic.v(141)
  wire C3qiu6;  // ../RTL/cortexm0ds_logic.v(652)
  wire C3rhu6;  // ../RTL/cortexm0ds_logic.v(184)
  wire C3row6;  // ../RTL/cortexm0ds_logic.v(1209)
  wire C3wpw6;  // ../RTL/cortexm0ds_logic.v(1610)
  wire C3xiu6;  // ../RTL/cortexm0ds_logic.v(746)
  wire C3yhu6;  // ../RTL/cortexm0ds_logic.v(278)
  wire C3yow6;  // ../RTL/cortexm0ds_logic.v(1302)
  wire C3zpw6;  // ../RTL/cortexm0ds_logic.v(1615)
  wire C43ju6;  // ../RTL/cortexm0ds_logic.v(826)
  wire C44iu6;  // ../RTL/cortexm0ds_logic.v(358)
  wire C44pw6;  // ../RTL/cortexm0ds_logic.v(1383)
  wire C47bx6;  // ../RTL/cortexm0ds_logic.v(1692)
  wire C4aju6;  // ../RTL/cortexm0ds_logic.v(920)
  wire C4biu6;  // ../RTL/cortexm0ds_logic.v(452)
  wire C4bpw6;  // ../RTL/cortexm0ds_logic.v(1476)
  wire C4cow6;  // ../RTL/cortexm0ds_logic.v(1008)
  wire C4dax6;  // ../RTL/cortexm0ds_logic.v(1637)
  wire C4ihu6;  // ../RTL/cortexm0ds_logic.v(130)
  wire C4iiu6;  // ../RTL/cortexm0ds_logic.v(546)
  wire C4jow6;  // ../RTL/cortexm0ds_logic.v(1102)
  wire C4piu6;  // ../RTL/cortexm0ds_logic.v(639)
  wire C4qhu6;  // ../RTL/cortexm0ds_logic.v(171)
  wire C4qow6;  // ../RTL/cortexm0ds_logic.v(1196)
  wire C4wiu6;  // ../RTL/cortexm0ds_logic.v(733)
  wire C4xhu6;  // ../RTL/cortexm0ds_logic.v(265)
  wire C4xow6;  // ../RTL/cortexm0ds_logic.v(1289)
  wire C50bx6;  // ../RTL/cortexm0ds_logic.v(1680)
  wire C52ju6;  // ../RTL/cortexm0ds_logic.v(813)
  wire C53iu6;  // ../RTL/cortexm0ds_logic.v(345)
  wire C53pw6;  // ../RTL/cortexm0ds_logic.v(1370)
  wire C59ju6;  // ../RTL/cortexm0ds_logic.v(907)
  wire C5aiu6;  // ../RTL/cortexm0ds_logic.v(439)
  wire C5apw6;  // ../RTL/cortexm0ds_logic.v(1463)
  wire C5bow6;  // ../RTL/cortexm0ds_logic.v(995)
  wire C5gbx6;  // ../RTL/cortexm0ds_logic.v(1708)
  wire C5hiu6;  // ../RTL/cortexm0ds_logic.v(533)
  wire C5iow6;  // ../RTL/cortexm0ds_logic.v(1089)
  wire C5oiu6;  // ../RTL/cortexm0ds_logic.v(626)
  wire C5phu6;  // ../RTL/cortexm0ds_logic.v(158)
  wire C5pow6;  // ../RTL/cortexm0ds_logic.v(1183)
  wire C5viu6;  // ../RTL/cortexm0ds_logic.v(720)
  wire C5whu6;  // ../RTL/cortexm0ds_logic.v(252)
  wire C5wow6;  // ../RTL/cortexm0ds_logic.v(1276)
  wire C5wpw6;  // ../RTL/cortexm0ds_logic.v(1610)
  wire C61ju6;  // ../RTL/cortexm0ds_logic.v(800)
  wire C62iu6;  // ../RTL/cortexm0ds_logic.v(332)
  wire C62pw6;  // ../RTL/cortexm0ds_logic.v(1357)
  wire C67bx6;  // ../RTL/cortexm0ds_logic.v(1692)
  wire C68ju6;  // ../RTL/cortexm0ds_logic.v(894)
  wire C69iu6;  // ../RTL/cortexm0ds_logic.v(426)
  wire C69pw6;  // ../RTL/cortexm0ds_logic.v(1450)
  wire C6aow6;  // ../RTL/cortexm0ds_logic.v(982)
  wire C6giu6;  // ../RTL/cortexm0ds_logic.v(520)
  wire C6how6;  // ../RTL/cortexm0ds_logic.v(1076)
  wire C6niu6;  // ../RTL/cortexm0ds_logic.v(613)
  wire C6oow6;  // ../RTL/cortexm0ds_logic.v(1170)
  wire C6uiu6;  // ../RTL/cortexm0ds_logic.v(707)
  wire C6vhu6;  // ../RTL/cortexm0ds_logic.v(239)
  wire C6vow6;  // ../RTL/cortexm0ds_logic.v(1263)
  wire C70ju6;  // ../RTL/cortexm0ds_logic.v(787)
  wire C71iu6;  // ../RTL/cortexm0ds_logic.v(319)
  wire C71pw6;  // ../RTL/cortexm0ds_logic.v(1344)
  wire C72qw6;  // ../RTL/cortexm0ds_logic.v(1621)
  wire C77ju6;  // ../RTL/cortexm0ds_logic.v(881)
  wire C78iu6;  // ../RTL/cortexm0ds_logic.v(413)
  wire C78pw6;  // ../RTL/cortexm0ds_logic.v(1437)
  wire C79ow6;  // ../RTL/cortexm0ds_logic.v(969)
  wire C7fiu6;  // ../RTL/cortexm0ds_logic.v(507)
  wire C7gow6;  // ../RTL/cortexm0ds_logic.v(1063)
  wire C7miu6;  // ../RTL/cortexm0ds_logic.v(600)
  wire C7now6;  // ../RTL/cortexm0ds_logic.v(1157)
  wire C7tiu6;  // ../RTL/cortexm0ds_logic.v(694)
  wire C7uhu6;  // ../RTL/cortexm0ds_logic.v(226)
  wire C7uow6;  // ../RTL/cortexm0ds_logic.v(1250)
  wire C7wpw6;  // ../RTL/cortexm0ds_logic.v(1610)
  wire C80iu6;  // ../RTL/cortexm0ds_logic.v(306)
  wire C80pw6;  // ../RTL/cortexm0ds_logic.v(1331)
  wire C86ju6;  // ../RTL/cortexm0ds_logic.v(868)
  wire C87bx6;  // ../RTL/cortexm0ds_logic.v(1692)
  wire C87iu6;  // ../RTL/cortexm0ds_logic.v(400)
  wire C87pw6;  // ../RTL/cortexm0ds_logic.v(1424)
  wire C88ow6;  // ../RTL/cortexm0ds_logic.v(956)
  wire C8eiu6;  // ../RTL/cortexm0ds_logic.v(494)
  wire C8fow6;  // ../RTL/cortexm0ds_logic.v(1050)
  wire C8liu6;  // ../RTL/cortexm0ds_logic.v(587)
  wire C8mow6;  // ../RTL/cortexm0ds_logic.v(1144)
  wire C8siu6;  // ../RTL/cortexm0ds_logic.v(681)
  wire C8thu6;  // ../RTL/cortexm0ds_logic.v(213)
  wire C8tow6;  // ../RTL/cortexm0ds_logic.v(1237)
  wire C8ziu6;  // ../RTL/cortexm0ds_logic.v(774)
  wire C95ju6;  // ../RTL/cortexm0ds_logic.v(855)
  wire C96iu6;  // ../RTL/cortexm0ds_logic.v(387)
  wire C96pw6;  // ../RTL/cortexm0ds_logic.v(1411)
  wire C97ow6;  // ../RTL/cortexm0ds_logic.v(943)
  wire C9diu6;  // ../RTL/cortexm0ds_logic.v(481)
  wire C9dpw6;  // ../RTL/cortexm0ds_logic.v(1505)
  wire C9eow6;  // ../RTL/cortexm0ds_logic.v(1037)
  wire C9kiu6;  // ../RTL/cortexm0ds_logic.v(574)
  wire C9low6;  // ../RTL/cortexm0ds_logic.v(1131)
  wire C9riu6;  // ../RTL/cortexm0ds_logic.v(668)
  wire C9shu6;  // ../RTL/cortexm0ds_logic.v(200)
  wire C9sow6;  // ../RTL/cortexm0ds_logic.v(1224)
  wire C9wpw6;  // ../RTL/cortexm0ds_logic.v(1610)
  wire C9yiu6;  // ../RTL/cortexm0ds_logic.v(761)
  wire C9zhu6;  // ../RTL/cortexm0ds_logic.v(293)
  wire C9zow6;  // ../RTL/cortexm0ds_logic.v(1318)
  wire Ca1bx6;  // ../RTL/cortexm0ds_logic.v(1682)
  wire Ca4ju6;  // ../RTL/cortexm0ds_logic.v(842)
  wire Ca5iu6;  // ../RTL/cortexm0ds_logic.v(374)
  wire Ca5pw6;  // ../RTL/cortexm0ds_logic.v(1398)
  wire Ca6ow6;  // ../RTL/cortexm0ds_logic.v(930)
  wire Ca7bx6;  // ../RTL/cortexm0ds_logic.v(1692)
  wire Caciu6;  // ../RTL/cortexm0ds_logic.v(468)
  wire Cacpw6;  // ../RTL/cortexm0ds_logic.v(1492)
  wire Cadow6;  // ../RTL/cortexm0ds_logic.v(1024)
  wire Caehu6;  // ../RTL/cortexm0ds_logic.v(121)
  wire Cajiu6;  // ../RTL/cortexm0ds_logic.v(561)
  wire Cakow6;  // ../RTL/cortexm0ds_logic.v(1118)
  wire Caqiu6;  // ../RTL/cortexm0ds_logic.v(655)
  wire Carhu6;  // ../RTL/cortexm0ds_logic.v(187)
  wire Carow6;  // ../RTL/cortexm0ds_logic.v(1211)
  wire Caxiu6;  // ../RTL/cortexm0ds_logic.v(748)
  wire Cayhu6;  // ../RTL/cortexm0ds_logic.v(280)
  wire Cayow6;  // ../RTL/cortexm0ds_logic.v(1305)
  wire Cb3ju6;  // ../RTL/cortexm0ds_logic.v(829)
  wire Cb4iu6;  // ../RTL/cortexm0ds_logic.v(361)
  wire Cb4pw6;  // ../RTL/cortexm0ds_logic.v(1385)
  wire Cbaju6;  // ../RTL/cortexm0ds_logic.v(923)
  wire Cbbiu6;  // ../RTL/cortexm0ds_logic.v(455)
  wire Cbbpw6;  // ../RTL/cortexm0ds_logic.v(1479)
  wire Cbcow6;  // ../RTL/cortexm0ds_logic.v(1011)
  wire Cbiiu6;  // ../RTL/cortexm0ds_logic.v(548)
  wire Cbjow6;  // ../RTL/cortexm0ds_logic.v(1105)
  wire Cbpiu6;  // ../RTL/cortexm0ds_logic.v(642)
  wire Cbqhu6;  // ../RTL/cortexm0ds_logic.v(174)
  wire Cbqow6;  // ../RTL/cortexm0ds_logic.v(1198)
  wire Cbwiu6;  // ../RTL/cortexm0ds_logic.v(735)
  wire Cbwpw6;  // ../RTL/cortexm0ds_logic.v(1610)
  wire Cbxhu6;  // ../RTL/cortexm0ds_logic.v(267)
  wire Cbxow6;  // ../RTL/cortexm0ds_logic.v(1292)
  wire Cc2bx6;  // ../RTL/cortexm0ds_logic.v(1683)
  wire Cc2ju6;  // ../RTL/cortexm0ds_logic.v(816)
  wire Cc3iu6;  // ../RTL/cortexm0ds_logic.v(348)
  wire Cc3pw6;  // ../RTL/cortexm0ds_logic.v(1372)
  wire Cc7bx6;  // ../RTL/cortexm0ds_logic.v(1692)
  wire Cc9ju6;  // ../RTL/cortexm0ds_logic.v(910)
  wire Ccaiu6;  // ../RTL/cortexm0ds_logic.v(442)
  wire Ccapw6;  // ../RTL/cortexm0ds_logic.v(1466)
  wire Ccbow6;  // ../RTL/cortexm0ds_logic.v(998)
  wire Cccbx6;  // ../RTL/cortexm0ds_logic.v(1701)
  wire Cchax6;  // ../RTL/cortexm0ds_logic.v(1645)
  wire Cchiu6;  // ../RTL/cortexm0ds_logic.v(535)
  wire Cciow6;  // ../RTL/cortexm0ds_logic.v(1092)
  wire Ccoiu6;  // ../RTL/cortexm0ds_logic.v(629)
  wire Ccphu6;  // ../RTL/cortexm0ds_logic.v(161)
  wire Ccpow6;  // ../RTL/cortexm0ds_logic.v(1185)
  wire Ccviu6;  // ../RTL/cortexm0ds_logic.v(722)
  wire Ccwhu6;  // ../RTL/cortexm0ds_logic.v(254)
  wire Ccwow6;  // ../RTL/cortexm0ds_logic.v(1279)
  wire Cd1ju6;  // ../RTL/cortexm0ds_logic.v(803)
  wire Cd2iu6;  // ../RTL/cortexm0ds_logic.v(335)
  wire Cd2pw6;  // ../RTL/cortexm0ds_logic.v(1359)
  wire Cd8ju6;  // ../RTL/cortexm0ds_logic.v(897)
  wire Cd9iu6;  // ../RTL/cortexm0ds_logic.v(429)
  wire Cd9pw6;  // ../RTL/cortexm0ds_logic.v(1453)
  wire Cdaow6;  // ../RTL/cortexm0ds_logic.v(985)
  wire Cdgiu6;  // ../RTL/cortexm0ds_logic.v(522)
  wire Cdhow6;  // ../RTL/cortexm0ds_logic.v(1079)
  wire Cdniu6;  // ../RTL/cortexm0ds_logic.v(616)
  wire Cdohu6;  // ../RTL/cortexm0ds_logic.v(148)
  wire Cdoow6;  // ../RTL/cortexm0ds_logic.v(1172)
  wire Cduiu6;  // ../RTL/cortexm0ds_logic.v(709)
  wire Cdvhu6;  // ../RTL/cortexm0ds_logic.v(241)
  wire Cdvow6;  // ../RTL/cortexm0ds_logic.v(1266)
  wire Cdwpw6;  // ../RTL/cortexm0ds_logic.v(1610)
  wire Ce0ju6;  // ../RTL/cortexm0ds_logic.v(790)
  wire Ce1iu6;  // ../RTL/cortexm0ds_logic.v(322)
  wire Ce1pw6;  // ../RTL/cortexm0ds_logic.v(1346)
  wire Ce7bx6;  // ../RTL/cortexm0ds_logic.v(1692)
  wire Ce7ju6;  // ../RTL/cortexm0ds_logic.v(884)
  wire Ce8iu6;  // ../RTL/cortexm0ds_logic.v(416)
  wire Ce8pw6;  // ../RTL/cortexm0ds_logic.v(1440)
  wire Ce9ow6;  // ../RTL/cortexm0ds_logic.v(972)
  wire Ceabx6;  // ../RTL/cortexm0ds_logic.v(1698)
  wire Cefhu6;  // ../RTL/cortexm0ds_logic.v(124)
  wire Cefiu6;  // ../RTL/cortexm0ds_logic.v(509)
  wire Cegow6;  // ../RTL/cortexm0ds_logic.v(1066)
  wire Cemiu6;  // ../RTL/cortexm0ds_logic.v(603)
  wire Cenow6;  // ../RTL/cortexm0ds_logic.v(1159)
  wire Cetiu6;  // ../RTL/cortexm0ds_logic.v(696)
  wire Ceuhu6;  // ../RTL/cortexm0ds_logic.v(228)
  wire Ceuow6;  // ../RTL/cortexm0ds_logic.v(1253)
  wire Cf0iu6;  // ../RTL/cortexm0ds_logic.v(309)
  wire Cf0pw6;  // ../RTL/cortexm0ds_logic.v(1333)
  wire Cf6ju6;  // ../RTL/cortexm0ds_logic.v(871)
  wire Cf7iu6;  // ../RTL/cortexm0ds_logic.v(403)
  wire Cf7pw6;  // ../RTL/cortexm0ds_logic.v(1427)
  wire Cf8ow6;  // ../RTL/cortexm0ds_logic.v(959)
  wire Cfeiu6;  // ../RTL/cortexm0ds_logic.v(496)
  wire Cffow6;  // ../RTL/cortexm0ds_logic.v(1053)
  wire Cfliu6;  // ../RTL/cortexm0ds_logic.v(590)
  wire Cfmow6;  // ../RTL/cortexm0ds_logic.v(1146)
  wire Cfsiu6;  // ../RTL/cortexm0ds_logic.v(683)
  wire Cfthu6;  // ../RTL/cortexm0ds_logic.v(215)
  wire Cftow6;  // ../RTL/cortexm0ds_logic.v(1240)
  wire Cfvpw6;  // ../RTL/cortexm0ds_logic.v(1609)
  wire Cfwpw6;  // ../RTL/cortexm0ds_logic.v(1610)
  wire Cfziu6;  // ../RTL/cortexm0ds_logic.v(777)
  wire Cg5ju6;  // ../RTL/cortexm0ds_logic.v(858)
  wire Cg6iu6;  // ../RTL/cortexm0ds_logic.v(390)
  wire Cg6pw6;  // ../RTL/cortexm0ds_logic.v(1414)
  wire Cg7bx6;  // ../RTL/cortexm0ds_logic.v(1692)
  wire Cg7ow6;  // ../RTL/cortexm0ds_logic.v(946)
  wire Cgdiu6;  // ../RTL/cortexm0ds_logic.v(483)
  wire Cgdpw6;  // ../RTL/cortexm0ds_logic.v(1508)
  wire Cgeow6;  // ../RTL/cortexm0ds_logic.v(1040)
  wire Cgkiu6;  // ../RTL/cortexm0ds_logic.v(577)
  wire Cglax6;  // ../RTL/cortexm0ds_logic.v(1653)
  wire Cglow6;  // ../RTL/cortexm0ds_logic.v(1133)
  wire Cgriu6;  // ../RTL/cortexm0ds_logic.v(670)
  wire Cgshu6;  // ../RTL/cortexm0ds_logic.v(202)
  wire Cgsow6;  // ../RTL/cortexm0ds_logic.v(1227)
  wire Cgyiu6;  // ../RTL/cortexm0ds_logic.v(764)
  wire Cgzhu6;  // ../RTL/cortexm0ds_logic.v(296)
  wire Cgzow6;  // ../RTL/cortexm0ds_logic.v(1320)
  wire Ch4ju6;  // ../RTL/cortexm0ds_logic.v(845)
  wire Ch5iu6;  // ../RTL/cortexm0ds_logic.v(377)
  wire Ch5pw6;  // ../RTL/cortexm0ds_logic.v(1401)
  wire Ch6ow6;  // ../RTL/cortexm0ds_logic.v(933)
  wire Chciu6;  // ../RTL/cortexm0ds_logic.v(470)
  wire Chcpw6;  // ../RTL/cortexm0ds_logic.v(1495)
  wire Chdow6;  // ../RTL/cortexm0ds_logic.v(1027)
  wire Chjiu6;  // ../RTL/cortexm0ds_logic.v(564)
  wire Chkhu6;  // ../RTL/cortexm0ds_logic.v(136)
  wire Chkow6;  // ../RTL/cortexm0ds_logic.v(1120)
  wire Chqiu6;  // ../RTL/cortexm0ds_logic.v(657)
  wire Chrhu6;  // ../RTL/cortexm0ds_logic.v(189)
  wire Chrow6;  // ../RTL/cortexm0ds_logic.v(1214)
  wire Chwpw6;  // ../RTL/cortexm0ds_logic.v(1610)
  wire Chxiu6;  // ../RTL/cortexm0ds_logic.v(751)
  wire Chyhu6;  // ../RTL/cortexm0ds_logic.v(283)
  wire Chyow6;  // ../RTL/cortexm0ds_logic.v(1307)
  wire Ci3ju6;  // ../RTL/cortexm0ds_logic.v(832)
  wire Ci4iu6;  // ../RTL/cortexm0ds_logic.v(364)
  wire Ci4pw6;  // ../RTL/cortexm0ds_logic.v(1388)
  wire Ci7bx6;  // ../RTL/cortexm0ds_logic.v(1692)
  wire Ciaju6;  // ../RTL/cortexm0ds_logic.v(925)
  wire Cibiu6;  // ../RTL/cortexm0ds_logic.v(457)
  wire Cibpw6;  // ../RTL/cortexm0ds_logic.v(1482)
  wire Cicow6;  // ../RTL/cortexm0ds_logic.v(1014)
  wire Ciiiu6;  // ../RTL/cortexm0ds_logic.v(551)
  wire Cijow6;  // ../RTL/cortexm0ds_logic.v(1107)
  wire Cilax6;  // ../RTL/cortexm0ds_logic.v(1653)
  wire Cipiu6;  // ../RTL/cortexm0ds_logic.v(644)
  wire Ciqhu6;  // ../RTL/cortexm0ds_logic.v(176)
  wire Ciqow6;  // ../RTL/cortexm0ds_logic.v(1201)
  wire Ciwiu6;  // ../RTL/cortexm0ds_logic.v(738)
  wire Cixhu6;  // ../RTL/cortexm0ds_logic.v(270)
  wire Cixow6;  // ../RTL/cortexm0ds_logic.v(1294)
  wire Cj2ju6;  // ../RTL/cortexm0ds_logic.v(819)
  wire Cj3iu6;  // ../RTL/cortexm0ds_logic.v(351)
  wire Cj3pw6;  // ../RTL/cortexm0ds_logic.v(1375)
  wire Cj9ju6;  // ../RTL/cortexm0ds_logic.v(912)
  wire Cjaiu6;  // ../RTL/cortexm0ds_logic.v(444)
  wire Cjapw6;  // ../RTL/cortexm0ds_logic.v(1469)
  wire Cjbow6;  // ../RTL/cortexm0ds_logic.v(1001)
  wire Cjhiu6;  // ../RTL/cortexm0ds_logic.v(538)
  wire Cjiow6;  // ../RTL/cortexm0ds_logic.v(1094)
  wire Cjjhu6;  // ../RTL/cortexm0ds_logic.v(134)
  wire Cjoiu6;  // ../RTL/cortexm0ds_logic.v(631)
  wire Cjphu6;  // ../RTL/cortexm0ds_logic.v(163)
  wire Cjpow6;  // ../RTL/cortexm0ds_logic.v(1188)
  wire Cjqpw6;  // ../RTL/cortexm0ds_logic.v(1600)
  wire Cjviu6;  // ../RTL/cortexm0ds_logic.v(725)
  wire Cjwhu6;  // ../RTL/cortexm0ds_logic.v(257)
  wire Cjwow6;  // ../RTL/cortexm0ds_logic.v(1281)
  wire Cjwpw6;  // ../RTL/cortexm0ds_logic.v(1611)
  wire Ck1ju6;  // ../RTL/cortexm0ds_logic.v(806)
  wire Ck2iu6;  // ../RTL/cortexm0ds_logic.v(338)
  wire Ck2pw6;  // ../RTL/cortexm0ds_logic.v(1362)
  wire Ck7bx6;  // ../RTL/cortexm0ds_logic.v(1693)
  wire Ck8ju6;  // ../RTL/cortexm0ds_logic.v(899)
  wire Ck9iu6;  // ../RTL/cortexm0ds_logic.v(431)
  wire Ck9pw6;  // ../RTL/cortexm0ds_logic.v(1456)
  wire Ckaow6;  // ../RTL/cortexm0ds_logic.v(988)
  wire Ckgiu6;  // ../RTL/cortexm0ds_logic.v(525)
  wire Ckhow6;  // ../RTL/cortexm0ds_logic.v(1081)
  wire Cklax6;  // ../RTL/cortexm0ds_logic.v(1653)
  wire Ckniu6;  // ../RTL/cortexm0ds_logic.v(618)
  wire Ckohu6;  // ../RTL/cortexm0ds_logic.v(150)
  wire Ckoow6;  // ../RTL/cortexm0ds_logic.v(1175)
  wire Ckuiu6;  // ../RTL/cortexm0ds_logic.v(712)
  wire Ckvhu6;  // ../RTL/cortexm0ds_logic.v(244)
  wire Ckvow6;  // ../RTL/cortexm0ds_logic.v(1268)
  wire Cl0ju6;  // ../RTL/cortexm0ds_logic.v(793)
  wire Cl1iu6;  // ../RTL/cortexm0ds_logic.v(325)
  wire Cl1pw6;  // ../RTL/cortexm0ds_logic.v(1349)
  wire Cl7ju6;  // ../RTL/cortexm0ds_logic.v(886)
  wire Cl8iu6;  // ../RTL/cortexm0ds_logic.v(418)
  wire Cl8pw6;  // ../RTL/cortexm0ds_logic.v(1443)
  wire Cl9ow6;  // ../RTL/cortexm0ds_logic.v(975)
  wire Clfiu6;  // ../RTL/cortexm0ds_logic.v(512)
  wire Clgow6;  // ../RTL/cortexm0ds_logic.v(1068)
  wire Clihu6;  // ../RTL/cortexm0ds_logic.v(131)
  wire Clmiu6;  // ../RTL/cortexm0ds_logic.v(605)
  wire Clnow6;  // ../RTL/cortexm0ds_logic.v(1162)
  wire Cltiu6;  // ../RTL/cortexm0ds_logic.v(699)
  wire Cluhu6;  // ../RTL/cortexm0ds_logic.v(231)
  wire Cluow6;  // ../RTL/cortexm0ds_logic.v(1255)
  wire Cm0iu6;  // ../RTL/cortexm0ds_logic.v(312)
  wire Cm0pw6;  // ../RTL/cortexm0ds_logic.v(1336)
  wire Cm6ju6;  // ../RTL/cortexm0ds_logic.v(873)
  wire Cm7bx6;  // ../RTL/cortexm0ds_logic.v(1693)
  wire Cm7iu6;  // ../RTL/cortexm0ds_logic.v(405)
  wire Cm7pw6;  // ../RTL/cortexm0ds_logic.v(1430)
  wire Cm8ow6;  // ../RTL/cortexm0ds_logic.v(962)
  wire Cmeiu6;  // ../RTL/cortexm0ds_logic.v(499)
  wire Cmfow6;  // ../RTL/cortexm0ds_logic.v(1055)
  wire Cmlax6;  // ../RTL/cortexm0ds_logic.v(1653)
  wire Cmliu6;  // ../RTL/cortexm0ds_logic.v(592)
  wire Cmmow6;  // ../RTL/cortexm0ds_logic.v(1149)
  wire Cmsiu6;  // ../RTL/cortexm0ds_logic.v(686)
  wire Cmthu6;  // ../RTL/cortexm0ds_logic.v(218)
  wire Cmtow6;  // ../RTL/cortexm0ds_logic.v(1242)
  wire Cmziu6;  // ../RTL/cortexm0ds_logic.v(780)
  wire Cn5ju6;  // ../RTL/cortexm0ds_logic.v(860)
  wire Cn6iu6;  // ../RTL/cortexm0ds_logic.v(392)
  wire Cn6pw6;  // ../RTL/cortexm0ds_logic.v(1417)
  wire Cn7ow6;  // ../RTL/cortexm0ds_logic.v(949)
  wire Cncbx6;  // ../RTL/cortexm0ds_logic.v(1702)
  wire Cndbx6;  // ../RTL/cortexm0ds_logic.v(1704)
  wire Cndiu6;  // ../RTL/cortexm0ds_logic.v(486)
  wire Cndpw6;  // ../RTL/cortexm0ds_logic.v(1510)
  wire Cneow6;  // ../RTL/cortexm0ds_logic.v(1042)
  wire Cnkiu6;  // ../RTL/cortexm0ds_logic.v(579)
  wire Cnlow6;  // ../RTL/cortexm0ds_logic.v(1136)
  wire Cnriu6;  // ../RTL/cortexm0ds_logic.v(673)
  wire Cnshu6;  // ../RTL/cortexm0ds_logic.v(205)
  wire Cnsow6;  // ../RTL/cortexm0ds_logic.v(1229)
  wire Cnyiu6;  // ../RTL/cortexm0ds_logic.v(767)
  wire Cnzhu6;  // ../RTL/cortexm0ds_logic.v(299)
  wire Cnzow6;  // ../RTL/cortexm0ds_logic.v(1323)
  wire Co4ju6;  // ../RTL/cortexm0ds_logic.v(847)
  wire Co5iu6;  // ../RTL/cortexm0ds_logic.v(379)
  wire Co5pw6;  // ../RTL/cortexm0ds_logic.v(1404)
  wire Co6ow6;  // ../RTL/cortexm0ds_logic.v(936)
  wire Co7bx6;  // ../RTL/cortexm0ds_logic.v(1693)
  wire Cociu6;  // ../RTL/cortexm0ds_logic.v(473)
  wire Cocpw6;  // ../RTL/cortexm0ds_logic.v(1497)
  wire Codow6;  // ../RTL/cortexm0ds_logic.v(1029)
  wire Cojiu6;  // ../RTL/cortexm0ds_logic.v(566)
  wire Cokbx6;  // ../RTL/cortexm0ds_logic.v(1717)
  wire Cokow6;  // ../RTL/cortexm0ds_logic.v(1123)
  wire Coqiu6;  // ../RTL/cortexm0ds_logic.v(660)
  wire Corhu6;  // ../RTL/cortexm0ds_logic.v(192)
  wire Corow6;  // ../RTL/cortexm0ds_logic.v(1216)
  wire Coupw6;  // ../RTL/cortexm0ds_logic.v(1607)
  wire Coxiu6;  // ../RTL/cortexm0ds_logic.v(754)
  wire Coyhu6;  // ../RTL/cortexm0ds_logic.v(286)
  wire Coyow6;  // ../RTL/cortexm0ds_logic.v(1310)
  wire Cp3ju6;  // ../RTL/cortexm0ds_logic.v(834)
  wire Cp4iu6;  // ../RTL/cortexm0ds_logic.v(366)
  wire Cp4pw6;  // ../RTL/cortexm0ds_logic.v(1391)
  wire Cpaju6;  // ../RTL/cortexm0ds_logic.v(928)
  wire Cpbiu6;  // ../RTL/cortexm0ds_logic.v(460)
  wire Cpbpw6;  // ../RTL/cortexm0ds_logic.v(1484)
  wire Cpcow6;  // ../RTL/cortexm0ds_logic.v(1016)
  wire Cpiiu6;  // ../RTL/cortexm0ds_logic.v(553)
  wire Cpjow6;  // ../RTL/cortexm0ds_logic.v(1110)
  wire Cppiu6;  // ../RTL/cortexm0ds_logic.v(647)
  wire Cpqhu6;  // ../RTL/cortexm0ds_logic.v(179)
  wire Cpqow6;  // ../RTL/cortexm0ds_logic.v(1203)
  wire Cpwiu6;  // ../RTL/cortexm0ds_logic.v(741)
  wire Cpxhu6;  // ../RTL/cortexm0ds_logic.v(273)
  wire Cpxow6;  // ../RTL/cortexm0ds_logic.v(1297)
  wire Cq2ju6;  // ../RTL/cortexm0ds_logic.v(821)
  wire Cq3iu6;  // ../RTL/cortexm0ds_logic.v(353)
  wire Cq3pw6;  // ../RTL/cortexm0ds_logic.v(1378)
  wire Cq3qw6;  // ../RTL/cortexm0ds_logic.v(1624)
  wire Cq7bx6;  // ../RTL/cortexm0ds_logic.v(1693)
  wire Cq9ju6;  // ../RTL/cortexm0ds_logic.v(915)
  wire Cqapw6;  // ../RTL/cortexm0ds_logic.v(1471)
  wire Cqbow6;  // ../RTL/cortexm0ds_logic.v(1003)
  wire Cqhiu6;  // ../RTL/cortexm0ds_logic.v(540)
  wire Cqiow6;  // ../RTL/cortexm0ds_logic.v(1097)
  wire Cqoiu6;  // ../RTL/cortexm0ds_logic.v(634)
  wire Cqphu6;  // ../RTL/cortexm0ds_logic.v(166)
  wire Cqpow6;  // ../RTL/cortexm0ds_logic.v(1190)
  wire Cqrpw6;  // ../RTL/cortexm0ds_logic.v(1602)
  wire Cqviu6;  // ../RTL/cortexm0ds_logic.v(728)
  wire Cqwhu6;  // ../RTL/cortexm0ds_logic.v(260)
  wire Cqwow6;  // ../RTL/cortexm0ds_logic.v(1284)
  wire Cr1ju6;  // ../RTL/cortexm0ds_logic.v(808)
  wire Cr2iu6;  // ../RTL/cortexm0ds_logic.v(340)
  wire Cr2pw6;  // ../RTL/cortexm0ds_logic.v(1365)
  wire Cr8ju6;  // ../RTL/cortexm0ds_logic.v(902)
  wire Cr9iu6;  // ../RTL/cortexm0ds_logic.v(434)
  wire Cr9pw6;  // ../RTL/cortexm0ds_logic.v(1458)
  wire Craow6;  // ../RTL/cortexm0ds_logic.v(990)
  wire Crgiu6;  // ../RTL/cortexm0ds_logic.v(527)
  wire Crhow6;  // ../RTL/cortexm0ds_logic.v(1084)
  wire Crniu6;  // ../RTL/cortexm0ds_logic.v(621)
  wire Crohu6;  // ../RTL/cortexm0ds_logic.v(153)
  wire Croow6;  // ../RTL/cortexm0ds_logic.v(1177)
  wire Cruiu6;  // ../RTL/cortexm0ds_logic.v(715)
  wire Crvhu6;  // ../RTL/cortexm0ds_logic.v(247)
  wire Crvow6;  // ../RTL/cortexm0ds_logic.v(1271)
  wire Cs0ju6;  // ../RTL/cortexm0ds_logic.v(795)
  wire Cs1iu6;  // ../RTL/cortexm0ds_logic.v(327)
  wire Cs1pw6;  // ../RTL/cortexm0ds_logic.v(1352)
  wire Cs6bx6;  // ../RTL/cortexm0ds_logic.v(1691)
  wire Cs7ju6;  // ../RTL/cortexm0ds_logic.v(889)
  wire Cs8iu6;  // ../RTL/cortexm0ds_logic.v(421)
  wire Cs8pw6;  // ../RTL/cortexm0ds_logic.v(1445)
  wire Cs9ow6;  // ../RTL/cortexm0ds_logic.v(977)
  wire Csfiu6;  // ../RTL/cortexm0ds_logic.v(514)
  wire Csgow6;  // ../RTL/cortexm0ds_logic.v(1071)
  wire Csmiu6;  // ../RTL/cortexm0ds_logic.v(608)
  wire Csnow6;  // ../RTL/cortexm0ds_logic.v(1164)
  wire Cstiu6;  // ../RTL/cortexm0ds_logic.v(702)
  wire Csuhu6;  // ../RTL/cortexm0ds_logic.v(234)
  wire Csuow6;  // ../RTL/cortexm0ds_logic.v(1258)
  wire Ct0iu6;  // ../RTL/cortexm0ds_logic.v(314)
  wire Ct0pw6;  // ../RTL/cortexm0ds_logic.v(1339)
  wire Ct6ju6;  // ../RTL/cortexm0ds_logic.v(876)
  wire Ct7iu6;  // ../RTL/cortexm0ds_logic.v(408)
  wire Ct7pw6;  // ../RTL/cortexm0ds_logic.v(1432)
  wire Ct8ow6;  // ../RTL/cortexm0ds_logic.v(964)
  wire Cteiu6;  // ../RTL/cortexm0ds_logic.v(501)
  wire Ctfow6;  // ../RTL/cortexm0ds_logic.v(1058)
  wire Ctliu6;  // ../RTL/cortexm0ds_logic.v(595)
  wire Ctmow6;  // ../RTL/cortexm0ds_logic.v(1151)
  wire Ctsiu6;  // ../RTL/cortexm0ds_logic.v(689)
  wire Ctthu6;  // ../RTL/cortexm0ds_logic.v(221)
  wire Cttow6;  // ../RTL/cortexm0ds_logic.v(1245)
  wire Ctziu6;  // ../RTL/cortexm0ds_logic.v(782)
  wire Cu5ju6;  // ../RTL/cortexm0ds_logic.v(863)
  wire Cu6iu6;  // ../RTL/cortexm0ds_logic.v(395)
  wire Cu6pw6;  // ../RTL/cortexm0ds_logic.v(1419)
  wire Cu7ow6;  // ../RTL/cortexm0ds_logic.v(951)
  wire Cudiu6;  // ../RTL/cortexm0ds_logic.v(488)
  wire Cudpw6;  // ../RTL/cortexm0ds_logic.v(1513)
  wire Cuehu6;  // ../RTL/cortexm0ds_logic.v(123)
  wire Cueow6;  // ../RTL/cortexm0ds_logic.v(1045)
  wire Cukiu6;  // ../RTL/cortexm0ds_logic.v(582)
  wire Culow6;  // ../RTL/cortexm0ds_logic.v(1138)
  wire Curiu6;  // ../RTL/cortexm0ds_logic.v(676)
  wire Cushu6;  // ../RTL/cortexm0ds_logic.v(208)
  wire Cusow6;  // ../RTL/cortexm0ds_logic.v(1232)
  wire Cuyiu6;  // ../RTL/cortexm0ds_logic.v(769)
  wire Cuzhu6;  // ../RTL/cortexm0ds_logic.v(301)
  wire Cuzow6;  // ../RTL/cortexm0ds_logic.v(1326)
  wire Cv4ju6;  // ../RTL/cortexm0ds_logic.v(850)
  wire Cv5iu6;  // ../RTL/cortexm0ds_logic.v(382)
  wire Cv5pw6;  // ../RTL/cortexm0ds_logic.v(1406)
  wire Cv6ow6;  // ../RTL/cortexm0ds_logic.v(938)
  wire Cvciu6;  // ../RTL/cortexm0ds_logic.v(475)
  wire Cvcpw6;  // ../RTL/cortexm0ds_logic.v(1500)
  wire Cvdow6;  // ../RTL/cortexm0ds_logic.v(1032)
  wire Cvjiu6;  // ../RTL/cortexm0ds_logic.v(569)
  wire Cvkow6;  // ../RTL/cortexm0ds_logic.v(1125)
  wire Cvpax6;  // ../RTL/cortexm0ds_logic.v(1661)
  wire Cvqiu6;  // ../RTL/cortexm0ds_logic.v(663)
  wire Cvrhu6;  // ../RTL/cortexm0ds_logic.v(195)
  wire Cvrow6;  // ../RTL/cortexm0ds_logic.v(1219)
  wire Cvxiu6;  // ../RTL/cortexm0ds_logic.v(756)
  wire Cvyhu6;  // ../RTL/cortexm0ds_logic.v(288)
  wire Cvyow6;  // ../RTL/cortexm0ds_logic.v(1313)
  wire Cw3ju6;  // ../RTL/cortexm0ds_logic.v(837)
  wire Cw4iu6;  // ../RTL/cortexm0ds_logic.v(369)
  wire Cw4pw6;  // ../RTL/cortexm0ds_logic.v(1393)
  wire Cwbiu6;  // ../RTL/cortexm0ds_logic.v(462)
  wire Cwbpw6;  // ../RTL/cortexm0ds_logic.v(1487)
  wire Cwcow6;  // ../RTL/cortexm0ds_logic.v(1019)
  wire Cwiiu6;  // ../RTL/cortexm0ds_logic.v(556)
  wire Cwjow6;  // ../RTL/cortexm0ds_logic.v(1112)
  wire Cwpiu6;  // ../RTL/cortexm0ds_logic.v(650)
  wire Cwqhu6;  // ../RTL/cortexm0ds_logic.v(182)
  wire Cwqow6;  // ../RTL/cortexm0ds_logic.v(1206)
  wire Cwwiu6;  // ../RTL/cortexm0ds_logic.v(743)
  wire Cwxhu6;  // ../RTL/cortexm0ds_logic.v(275)
  wire Cwxow6;  // ../RTL/cortexm0ds_logic.v(1300)
  wire Cwyax6;  // ../RTL/cortexm0ds_logic.v(1677)
  wire Cx2ju6;  // ../RTL/cortexm0ds_logic.v(824)
  wire Cx3iu6;  // ../RTL/cortexm0ds_logic.v(356)
  wire Cx3pw6;  // ../RTL/cortexm0ds_logic.v(1380)
  wire Cx9ju6;  // ../RTL/cortexm0ds_logic.v(917)
  wire Cxaiu6;  // ../RTL/cortexm0ds_logic.v(449)
  wire Cxapw6;  // ../RTL/cortexm0ds_logic.v(1474)
  wire Cxbow6;  // ../RTL/cortexm0ds_logic.v(1006)
  wire Cxcbx6;  // ../RTL/cortexm0ds_logic.v(1702)
  wire Cxhiu6;  // ../RTL/cortexm0ds_logic.v(543)
  wire Cxiow6;  // ../RTL/cortexm0ds_logic.v(1099)
  wire Cxoiu6;  // ../RTL/cortexm0ds_logic.v(637)
  wire Cxphu6;  // ../RTL/cortexm0ds_logic.v(169)
  wire Cxpow6;  // ../RTL/cortexm0ds_logic.v(1193)
  wire Cxviu6;  // ../RTL/cortexm0ds_logic.v(730)
  wire Cxwhu6;  // ../RTL/cortexm0ds_logic.v(262)
  wire Cxwow6;  // ../RTL/cortexm0ds_logic.v(1287)
  wire Cxzax6;  // ../RTL/cortexm0ds_logic.v(1679)
  wire Cy1ju6;  // ../RTL/cortexm0ds_logic.v(811)
  wire Cy2iu6;  // ../RTL/cortexm0ds_logic.v(343)
  wire Cy2pw6;  // ../RTL/cortexm0ds_logic.v(1367)
  wire Cy4bx6;  // ../RTL/cortexm0ds_logic.v(1688)
  wire Cy8ju6;  // ../RTL/cortexm0ds_logic.v(904)
  wire Cy9iu6;  // ../RTL/cortexm0ds_logic.v(436)
  wire Cy9pw6;  // ../RTL/cortexm0ds_logic.v(1461)
  wire Cyaow6;  // ../RTL/cortexm0ds_logic.v(993)
  wire Cydbx6;  // ../RTL/cortexm0ds_logic.v(1704)
  wire Cygiu6;  // ../RTL/cortexm0ds_logic.v(530)
  wire Cyhow6;  // ../RTL/cortexm0ds_logic.v(1086)
  wire Cykhu6;  // ../RTL/cortexm0ds_logic.v(138)
  wire Cynhu6;  // ../RTL/cortexm0ds_logic.v(146)
  wire Cyniu6;  // ../RTL/cortexm0ds_logic.v(624)
  wire Cyohu6;  // ../RTL/cortexm0ds_logic.v(156)
  wire Cyoow6;  // ../RTL/cortexm0ds_logic.v(1180)
  wire Cyuiu6;  // ../RTL/cortexm0ds_logic.v(717)
  wire Cyvhu6;  // ../RTL/cortexm0ds_logic.v(249)
  wire Cyvow6;  // ../RTL/cortexm0ds_logic.v(1274)
  wire Cz0ju6;  // ../RTL/cortexm0ds_logic.v(798)
  wire Cz1iu6;  // ../RTL/cortexm0ds_logic.v(330)
  wire Cz1pw6;  // ../RTL/cortexm0ds_logic.v(1354)
  wire Cz7ju6;  // ../RTL/cortexm0ds_logic.v(891)
  wire Cz8iu6;  // ../RTL/cortexm0ds_logic.v(423)
  wire Cz8pw6;  // ../RTL/cortexm0ds_logic.v(1448)
  wire Cz9ow6;  // ../RTL/cortexm0ds_logic.v(980)
  wire Czfiu6;  // ../RTL/cortexm0ds_logic.v(517)
  wire Czgow6;  // ../RTL/cortexm0ds_logic.v(1073)
  wire Czmiu6;  // ../RTL/cortexm0ds_logic.v(611)
  wire Cznow6;  // ../RTL/cortexm0ds_logic.v(1167)
  wire Cztiu6;  // ../RTL/cortexm0ds_logic.v(704)
  wire Czuhu6;  // ../RTL/cortexm0ds_logic.v(236)
  wire Czuow6;  // ../RTL/cortexm0ds_logic.v(1261)
  wire Czzax6;  // ../RTL/cortexm0ds_logic.v(1679)
  wire D04ju6;  // ../RTL/cortexm0ds_logic.v(838)
  wire D05iu6;  // ../RTL/cortexm0ds_logic.v(370)
  wire D05pw6;  // ../RTL/cortexm0ds_logic.v(1395)
  wire D0ciu6;  // ../RTL/cortexm0ds_logic.v(464)
  wire D0cpw6;  // ../RTL/cortexm0ds_logic.v(1488)
  wire D0dow6;  // ../RTL/cortexm0ds_logic.v(1020)
  wire D0jiu6;  // ../RTL/cortexm0ds_logic.v(557)
  wire D0kow6;  // ../RTL/cortexm0ds_logic.v(1114)
  wire D0qiu6;  // ../RTL/cortexm0ds_logic.v(651)
  wire D0rhu6;  // ../RTL/cortexm0ds_logic.v(183)
  wire D0row6;  // ../RTL/cortexm0ds_logic.v(1207)
  wire D0uax6;  // ../RTL/cortexm0ds_logic.v(1669)
  wire D0xiu6;  // ../RTL/cortexm0ds_logic.v(745)
  wire D0yhu6;  // ../RTL/cortexm0ds_logic.v(277)
  wire D0yow6;  // ../RTL/cortexm0ds_logic.v(1301)
  wire D12qw6;  // ../RTL/cortexm0ds_logic.v(1621)
  wire D13ju6;  // ../RTL/cortexm0ds_logic.v(825)
  wire D14iu6;  // ../RTL/cortexm0ds_logic.v(357)
  wire D14pw6;  // ../RTL/cortexm0ds_logic.v(1382)
  wire D1aax6;  // ../RTL/cortexm0ds_logic.v(1631)
  wire D1aju6;  // ../RTL/cortexm0ds_logic.v(919)
  wire D1biu6;  // ../RTL/cortexm0ds_logic.v(451)
  wire D1bpw6;  // ../RTL/cortexm0ds_logic.v(1475)
  wire D1cow6;  // ../RTL/cortexm0ds_logic.v(1007)
  wire D1iiu6;  // ../RTL/cortexm0ds_logic.v(544)
  wire D1jow6;  // ../RTL/cortexm0ds_logic.v(1101)
  wire D1piu6;  // ../RTL/cortexm0ds_logic.v(638)
  wire D1qhu6;  // ../RTL/cortexm0ds_logic.v(170)
  wire D1qow6;  // ../RTL/cortexm0ds_logic.v(1194)
  wire D1wiu6;  // ../RTL/cortexm0ds_logic.v(732)
  wire D1xhu6;  // ../RTL/cortexm0ds_logic.v(264)
  wire D1xow6;  // ../RTL/cortexm0ds_logic.v(1288)
  wire D1zpw6;  // ../RTL/cortexm0ds_logic.v(1615)
  wire D22ju6;  // ../RTL/cortexm0ds_logic.v(812)
  wire D23iu6;  // ../RTL/cortexm0ds_logic.v(344)
  wire D23pw6;  // ../RTL/cortexm0ds_logic.v(1369)
  wire D29ju6;  // ../RTL/cortexm0ds_logic.v(906)
  wire D2aiu6;  // ../RTL/cortexm0ds_logic.v(438)
  wire D2apw6;  // ../RTL/cortexm0ds_logic.v(1462)
  wire D2bow6;  // ../RTL/cortexm0ds_logic.v(994)
  wire D2hiu6;  // ../RTL/cortexm0ds_logic.v(531)
  wire D2iow6;  // ../RTL/cortexm0ds_logic.v(1088)
  wire D2oiu6;  // ../RTL/cortexm0ds_logic.v(625)
  wire D2opw6;  // ../RTL/cortexm0ds_logic.v(1595)
  wire D2phu6;  // ../RTL/cortexm0ds_logic.v(157)
  wire D2pow6;  // ../RTL/cortexm0ds_logic.v(1181)
  wire D2rpw6;  // ../RTL/cortexm0ds_logic.v(1601)
  wire D2viu6;  // ../RTL/cortexm0ds_logic.v(719)
  wire D2whu6;  // ../RTL/cortexm0ds_logic.v(251)
  wire D2wow6;  // ../RTL/cortexm0ds_logic.v(1275)
  wire D31ju6;  // ../RTL/cortexm0ds_logic.v(799)
  wire D32iu6;  // ../RTL/cortexm0ds_logic.v(331)
  wire D32pw6;  // ../RTL/cortexm0ds_logic.v(1356)
  wire D38ju6;  // ../RTL/cortexm0ds_logic.v(893)
  wire D39iu6;  // ../RTL/cortexm0ds_logic.v(425)
  wire D39pw6;  // ../RTL/cortexm0ds_logic.v(1449)
  wire D3aow6;  // ../RTL/cortexm0ds_logic.v(981)
  wire D3giu6;  // ../RTL/cortexm0ds_logic.v(518)
  wire D3how6;  // ../RTL/cortexm0ds_logic.v(1075)
  wire D3niu6;  // ../RTL/cortexm0ds_logic.v(612)
  wire D3oow6;  // ../RTL/cortexm0ds_logic.v(1168)
  wire D3uiu6;  // ../RTL/cortexm0ds_logic.v(706)
  wire D3vhu6;  // ../RTL/cortexm0ds_logic.v(238)
  wire D3vow6;  // ../RTL/cortexm0ds_logic.v(1262)
  wire D40ju6;  // ../RTL/cortexm0ds_logic.v(786)
  wire D41iu6;  // ../RTL/cortexm0ds_logic.v(318)
  wire D41pw6;  // ../RTL/cortexm0ds_logic.v(1343)
  wire D43qw6;  // ../RTL/cortexm0ds_logic.v(1623)
  wire D46bx6;  // ../RTL/cortexm0ds_logic.v(1690)
  wire D47ju6;  // ../RTL/cortexm0ds_logic.v(880)
  wire D48iu6;  // ../RTL/cortexm0ds_logic.v(412)
  wire D48pw6;  // ../RTL/cortexm0ds_logic.v(1436)
  wire D49ow6;  // ../RTL/cortexm0ds_logic.v(968)
  wire D4fiu6;  // ../RTL/cortexm0ds_logic.v(505)
  wire D4gow6;  // ../RTL/cortexm0ds_logic.v(1062)
  wire D4miu6;  // ../RTL/cortexm0ds_logic.v(599)
  wire D4now6;  // ../RTL/cortexm0ds_logic.v(1155)
  wire D4tiu6;  // ../RTL/cortexm0ds_logic.v(693)
  wire D4uhu6;  // ../RTL/cortexm0ds_logic.v(225)
  wire D4uow6;  // ../RTL/cortexm0ds_logic.v(1249)
  wire D50iu6;  // ../RTL/cortexm0ds_logic.v(305)
  wire D50pw6;  // ../RTL/cortexm0ds_logic.v(1330)
  wire D56ju6;  // ../RTL/cortexm0ds_logic.v(867)
  wire D57iu6;  // ../RTL/cortexm0ds_logic.v(399)
  wire D57pw6;  // ../RTL/cortexm0ds_logic.v(1423)
  wire D58ow6;  // ../RTL/cortexm0ds_logic.v(955)
  wire D5eiu6;  // ../RTL/cortexm0ds_logic.v(492)
  wire D5epw6;  // ../RTL/cortexm0ds_logic.v(1517)
  wire D5fow6;  // ../RTL/cortexm0ds_logic.v(1049)
  wire D5liu6;  // ../RTL/cortexm0ds_logic.v(586)
  wire D5mow6;  // ../RTL/cortexm0ds_logic.v(1142)
  wire D5siu6;  // ../RTL/cortexm0ds_logic.v(680)
  wire D5thu6;  // ../RTL/cortexm0ds_logic.v(212)
  wire D5tow6;  // ../RTL/cortexm0ds_logic.v(1236)
  wire D5ziu6;  // ../RTL/cortexm0ds_logic.v(773)
  wire D65ju6;  // ../RTL/cortexm0ds_logic.v(854)
  wire D66bx6;  // ../RTL/cortexm0ds_logic.v(1690)
  wire D66iu6;  // ../RTL/cortexm0ds_logic.v(386)
  wire D66pw6;  // ../RTL/cortexm0ds_logic.v(1410)
  wire D67ow6;  // ../RTL/cortexm0ds_logic.v(942)
  wire D6diu6;  // ../RTL/cortexm0ds_logic.v(479)
  wire D6dpw6;  // ../RTL/cortexm0ds_logic.v(1504)
  wire D6eow6;  // ../RTL/cortexm0ds_logic.v(1036)
  wire D6kiu6;  // ../RTL/cortexm0ds_logic.v(573)
  wire D6low6;  // ../RTL/cortexm0ds_logic.v(1129)
  wire D6riu6;  // ../RTL/cortexm0ds_logic.v(667)
  wire D6shu6;  // ../RTL/cortexm0ds_logic.v(199)
  wire D6sow6;  // ../RTL/cortexm0ds_logic.v(1223)
  wire D6yiu6;  // ../RTL/cortexm0ds_logic.v(760)
  wire D6zhu6;  // ../RTL/cortexm0ds_logic.v(292)
  wire D6zow6;  // ../RTL/cortexm0ds_logic.v(1317)
  wire D70bx6;  // ../RTL/cortexm0ds_logic.v(1680)
  wire D74ju6;  // ../RTL/cortexm0ds_logic.v(841)
  wire D75iu6;  // ../RTL/cortexm0ds_logic.v(373)
  wire D75pw6;  // ../RTL/cortexm0ds_logic.v(1397)
  wire D7ciu6;  // ../RTL/cortexm0ds_logic.v(466)
  wire D7cpw6;  // ../RTL/cortexm0ds_logic.v(1491)
  wire D7dow6;  // ../RTL/cortexm0ds_logic.v(1023)
  wire D7gbx6;  // ../RTL/cortexm0ds_logic.v(1709)
  wire D7jiu6;  // ../RTL/cortexm0ds_logic.v(560)
  wire D7kow6;  // ../RTL/cortexm0ds_logic.v(1116)
  wire D7qiu6;  // ../RTL/cortexm0ds_logic.v(654)
  wire D7rhu6;  // ../RTL/cortexm0ds_logic.v(186)
  wire D7row6;  // ../RTL/cortexm0ds_logic.v(1210)
  wire D7xiu6;  // ../RTL/cortexm0ds_logic.v(747)
  wire D7yhu6;  // ../RTL/cortexm0ds_logic.v(279)
  wire D7yow6;  // ../RTL/cortexm0ds_logic.v(1304)
  wire D83ju6;  // ../RTL/cortexm0ds_logic.v(828)
  wire D84iu6;  // ../RTL/cortexm0ds_logic.v(360)
  wire D84pw6;  // ../RTL/cortexm0ds_logic.v(1384)
  wire D86bx6;  // ../RTL/cortexm0ds_logic.v(1690)
  wire D8aju6;  // ../RTL/cortexm0ds_logic.v(921)
  wire D8biu6;  // ../RTL/cortexm0ds_logic.v(453)
  wire D8bpw6;  // ../RTL/cortexm0ds_logic.v(1478)
  wire D8cow6;  // ../RTL/cortexm0ds_logic.v(1010)
  wire D8hhu6;  // ../RTL/cortexm0ds_logic.v(128)
  wire D8iiu6;  // ../RTL/cortexm0ds_logic.v(547)
  wire D8jow6;  // ../RTL/cortexm0ds_logic.v(1103)
  wire D8piu6;  // ../RTL/cortexm0ds_logic.v(641)
  wire D8qhu6;  // ../RTL/cortexm0ds_logic.v(173)
  wire D8qow6;  // ../RTL/cortexm0ds_logic.v(1197)
  wire D8wiu6;  // ../RTL/cortexm0ds_logic.v(734)
  wire D8xhu6;  // ../RTL/cortexm0ds_logic.v(266)
  wire D8xow6;  // ../RTL/cortexm0ds_logic.v(1291)
  wire D92ju6;  // ../RTL/cortexm0ds_logic.v(815)
  wire D93iu6;  // ../RTL/cortexm0ds_logic.v(347)
  wire D93pw6;  // ../RTL/cortexm0ds_logic.v(1371)
  wire D99ax6;  // ../RTL/cortexm0ds_logic.v(1630)
  wire D99ju6;  // ../RTL/cortexm0ds_logic.v(908)
  wire D9aiu6;  // ../RTL/cortexm0ds_logic.v(440)
  wire D9apw6;  // ../RTL/cortexm0ds_logic.v(1465)
  wire D9bow6;  // ../RTL/cortexm0ds_logic.v(997)
  wire D9hiu6;  // ../RTL/cortexm0ds_logic.v(534)
  wire D9iow6;  // ../RTL/cortexm0ds_logic.v(1090)
  wire D9oiu6;  // ../RTL/cortexm0ds_logic.v(628)
  wire D9phu6;  // ../RTL/cortexm0ds_logic.v(160)
  wire D9pow6;  // ../RTL/cortexm0ds_logic.v(1184)
  wire D9viu6;  // ../RTL/cortexm0ds_logic.v(721)
  wire D9whu6;  // ../RTL/cortexm0ds_logic.v(253)
  wire D9wow6;  // ../RTL/cortexm0ds_logic.v(1278)
  wire Da1ju6;  // ../RTL/cortexm0ds_logic.v(802)
  wire Da2iu6;  // ../RTL/cortexm0ds_logic.v(334)
  wire Da2pw6;  // ../RTL/cortexm0ds_logic.v(1358)
  wire Da6bx6;  // ../RTL/cortexm0ds_logic.v(1690)
  wire Da8ju6;  // ../RTL/cortexm0ds_logic.v(895)
  wire Da9iu6;  // ../RTL/cortexm0ds_logic.v(427)
  wire Da9pw6;  // ../RTL/cortexm0ds_logic.v(1452)
  wire Daaow6;  // ../RTL/cortexm0ds_logic.v(984)
  wire Daebx6;  // ../RTL/cortexm0ds_logic.v(1705)
  wire Dagiu6;  // ../RTL/cortexm0ds_logic.v(521)
  wire Dahow6;  // ../RTL/cortexm0ds_logic.v(1077)
  wire Daiax6;  // ../RTL/cortexm0ds_logic.v(1647)
  wire Daniu6;  // ../RTL/cortexm0ds_logic.v(615)
  wire Daoow6;  // ../RTL/cortexm0ds_logic.v(1171)
  wire Dauiu6;  // ../RTL/cortexm0ds_logic.v(708)
  wire Davhu6;  // ../RTL/cortexm0ds_logic.v(240)
  wire Davow6;  // ../RTL/cortexm0ds_logic.v(1265)
  wire Db0ju6;  // ../RTL/cortexm0ds_logic.v(789)
  wire Db1iu6;  // ../RTL/cortexm0ds_logic.v(321)
  wire Db1pw6;  // ../RTL/cortexm0ds_logic.v(1345)
  wire Db7ju6;  // ../RTL/cortexm0ds_logic.v(882)
  wire Db8iu6;  // ../RTL/cortexm0ds_logic.v(414)
  wire Db8pw6;  // ../RTL/cortexm0ds_logic.v(1439)
  wire Db9ow6;  // ../RTL/cortexm0ds_logic.v(971)
  wire Dbfiu6;  // ../RTL/cortexm0ds_logic.v(508)
  wire Dbgow6;  // ../RTL/cortexm0ds_logic.v(1064)
  wire Dbmiu6;  // ../RTL/cortexm0ds_logic.v(602)
  wire Dbnow6;  // ../RTL/cortexm0ds_logic.v(1158)
  wire Dbtiu6;  // ../RTL/cortexm0ds_logic.v(695)
  wire Dbuhu6;  // ../RTL/cortexm0ds_logic.v(227)
  wire Dbuow6;  // ../RTL/cortexm0ds_logic.v(1252)
  wire Dc0iu6;  // ../RTL/cortexm0ds_logic.v(308)
  wire Dc0pw6;  // ../RTL/cortexm0ds_logic.v(1332)
  wire Dc6bx6;  // ../RTL/cortexm0ds_logic.v(1690)
  wire Dc6ju6;  // ../RTL/cortexm0ds_logic.v(869)
  wire Dc7iu6;  // ../RTL/cortexm0ds_logic.v(401)
  wire Dc7pw6;  // ../RTL/cortexm0ds_logic.v(1426)
  wire Dc8ow6;  // ../RTL/cortexm0ds_logic.v(958)
  wire Dceiu6;  // ../RTL/cortexm0ds_logic.v(495)
  wire Dcfow6;  // ../RTL/cortexm0ds_logic.v(1051)
  wire Dcliu6;  // ../RTL/cortexm0ds_logic.v(589)
  wire Dcmow6;  // ../RTL/cortexm0ds_logic.v(1145)
  wire Dcsiu6;  // ../RTL/cortexm0ds_logic.v(682)
  wire Dcthu6;  // ../RTL/cortexm0ds_logic.v(214)
  wire Dctow6;  // ../RTL/cortexm0ds_logic.v(1239)
  wire Dcziu6;  // ../RTL/cortexm0ds_logic.v(776)
  wire Dd5ju6;  // ../RTL/cortexm0ds_logic.v(856)
  wire Dd6iu6;  // ../RTL/cortexm0ds_logic.v(388)
  wire Dd6pw6;  // ../RTL/cortexm0ds_logic.v(1413)
  wire Dd7ow6;  // ../RTL/cortexm0ds_logic.v(945)
  wire Dddiu6;  // ../RTL/cortexm0ds_logic.v(482)
  wire Dddpw6;  // ../RTL/cortexm0ds_logic.v(1506)
  wire Ddeow6;  // ../RTL/cortexm0ds_logic.v(1038)
  wire Ddkiu6;  // ../RTL/cortexm0ds_logic.v(576)
  wire Ddlow6;  // ../RTL/cortexm0ds_logic.v(1132)
  wire Ddriu6;  // ../RTL/cortexm0ds_logic.v(669)
  wire Ddshu6;  // ../RTL/cortexm0ds_logic.v(201)
  wire Ddsow6;  // ../RTL/cortexm0ds_logic.v(1226)
  wire Ddyiu6;  // ../RTL/cortexm0ds_logic.v(763)
  wire Ddzhu6;  // ../RTL/cortexm0ds_logic.v(295)
  wire Ddzow6;  // ../RTL/cortexm0ds_logic.v(1319)
  wire De4ju6;  // ../RTL/cortexm0ds_logic.v(843)
  wire De5iu6;  // ../RTL/cortexm0ds_logic.v(375)
  wire De5pw6;  // ../RTL/cortexm0ds_logic.v(1400)
  wire De6bx6;  // ../RTL/cortexm0ds_logic.v(1690)
  wire De6ow6;  // ../RTL/cortexm0ds_logic.v(932)
  wire Deciu6;  // ../RTL/cortexm0ds_logic.v(469)
  wire Decpw6;  // ../RTL/cortexm0ds_logic.v(1493)
  wire Dedow6;  // ../RTL/cortexm0ds_logic.v(1025)
  wire Dejiu6;  // ../RTL/cortexm0ds_logic.v(563)
  wire Dekow6;  // ../RTL/cortexm0ds_logic.v(1119)
  wire Delax6;  // ../RTL/cortexm0ds_logic.v(1653)
  wire Deqiu6;  // ../RTL/cortexm0ds_logic.v(656)
  wire Derhu6;  // ../RTL/cortexm0ds_logic.v(188)
  wire Derow6;  // ../RTL/cortexm0ds_logic.v(1213)
  wire Dexiu6;  // ../RTL/cortexm0ds_logic.v(750)
  wire Deyhu6;  // ../RTL/cortexm0ds_logic.v(282)
  wire Deyow6;  // ../RTL/cortexm0ds_logic.v(1306)
  wire Df3ju6;  // ../RTL/cortexm0ds_logic.v(830)
  wire Df4iu6;  // ../RTL/cortexm0ds_logic.v(362)
  wire Df4pw6;  // ../RTL/cortexm0ds_logic.v(1387)
  wire Dfaju6;  // ../RTL/cortexm0ds_logic.v(924)
  wire Dfbax6;  // ../RTL/cortexm0ds_logic.v(1634)
  wire Dfbiu6;  // ../RTL/cortexm0ds_logic.v(456)
  wire Dfbpw6;  // ../RTL/cortexm0ds_logic.v(1480)
  wire Dfcow6;  // ../RTL/cortexm0ds_logic.v(1012)
  wire Dfiiu6;  // ../RTL/cortexm0ds_logic.v(550)
  wire Dfjow6;  // ../RTL/cortexm0ds_logic.v(1106)
  wire Dfpiu6;  // ../RTL/cortexm0ds_logic.v(643)
  wire Dfqhu6;  // ../RTL/cortexm0ds_logic.v(175)
  wire Dfqow6;  // ../RTL/cortexm0ds_logic.v(1200)
  wire Dfwiu6;  // ../RTL/cortexm0ds_logic.v(737)
  wire Dfxhu6;  // ../RTL/cortexm0ds_logic.v(269)
  wire Dfxow6;  // ../RTL/cortexm0ds_logic.v(1293)
  wire Dg2ju6;  // ../RTL/cortexm0ds_logic.v(817)
  wire Dg2qw6;  // ../RTL/cortexm0ds_logic.v(1621)
  wire Dg3iu6;  // ../RTL/cortexm0ds_logic.v(349)
  wire Dg3pw6;  // ../RTL/cortexm0ds_logic.v(1374)
  wire Dg6bx6;  // ../RTL/cortexm0ds_logic.v(1691)
  wire Dg9ju6;  // ../RTL/cortexm0ds_logic.v(911)
  wire Dgaiu6;  // ../RTL/cortexm0ds_logic.v(443)
  wire Dgapw6;  // ../RTL/cortexm0ds_logic.v(1467)
  wire Dgbow6;  // ../RTL/cortexm0ds_logic.v(999)
  wire Dghiu6;  // ../RTL/cortexm0ds_logic.v(537)
  wire Dgiow6;  // ../RTL/cortexm0ds_logic.v(1093)
  wire Dgoiu6;  // ../RTL/cortexm0ds_logic.v(630)
  wire Dgphu6;  // ../RTL/cortexm0ds_logic.v(162)
  wire Dgpow6;  // ../RTL/cortexm0ds_logic.v(1187)
  wire Dgviu6;  // ../RTL/cortexm0ds_logic.v(724)
  wire Dgwhu6;  // ../RTL/cortexm0ds_logic.v(256)
  wire Dgwow6;  // ../RTL/cortexm0ds_logic.v(1280)
  wire Dh1ju6;  // ../RTL/cortexm0ds_logic.v(804)
  wire Dh2iu6;  // ../RTL/cortexm0ds_logic.v(336)
  wire Dh2pw6;  // ../RTL/cortexm0ds_logic.v(1361)
  wire Dh8ju6;  // ../RTL/cortexm0ds_logic.v(898)
  wire Dh9iu6;  // ../RTL/cortexm0ds_logic.v(430)
  wire Dh9pw6;  // ../RTL/cortexm0ds_logic.v(1454)
  wire Dhaow6;  // ../RTL/cortexm0ds_logic.v(986)
  wire Dhfhu6;  // ../RTL/cortexm0ds_logic.v(124)
  wire Dhgiu6;  // ../RTL/cortexm0ds_logic.v(524)
  wire Dhhow6;  // ../RTL/cortexm0ds_logic.v(1080)
  wire Dhniu6;  // ../RTL/cortexm0ds_logic.v(617)
  wire Dhohu6;  // ../RTL/cortexm0ds_logic.v(149)
  wire Dhoow6;  // ../RTL/cortexm0ds_logic.v(1174)
  wire Dhuiu6;  // ../RTL/cortexm0ds_logic.v(711)
  wire Dhvhu6;  // ../RTL/cortexm0ds_logic.v(243)
  wire Dhvow6;  // ../RTL/cortexm0ds_logic.v(1267)
  wire Di0ju6;  // ../RTL/cortexm0ds_logic.v(791)
  wire Di1iu6;  // ../RTL/cortexm0ds_logic.v(323)
  wire Di1pw6;  // ../RTL/cortexm0ds_logic.v(1348)
  wire Di3qw6;  // ../RTL/cortexm0ds_logic.v(1624)
  wire Di6bx6;  // ../RTL/cortexm0ds_logic.v(1691)
  wire Di7ju6;  // ../RTL/cortexm0ds_logic.v(885)
  wire Di8iu6;  // ../RTL/cortexm0ds_logic.v(417)
  wire Di8pw6;  // ../RTL/cortexm0ds_logic.v(1441)
  wire Di9ow6;  // ../RTL/cortexm0ds_logic.v(973)
  wire Difiu6;  // ../RTL/cortexm0ds_logic.v(511)
  wire Digow6;  // ../RTL/cortexm0ds_logic.v(1067)
  wire Dimiu6;  // ../RTL/cortexm0ds_logic.v(604)
  wire Dinow6;  // ../RTL/cortexm0ds_logic.v(1161)
  wire Ditiu6;  // ../RTL/cortexm0ds_logic.v(698)
  wire Diuhu6;  // ../RTL/cortexm0ds_logic.v(230)
  wire Diuow6;  // ../RTL/cortexm0ds_logic.v(1254)
  wire Dj0iu6;  // ../RTL/cortexm0ds_logic.v(310)
  wire Dj0pw6;  // ../RTL/cortexm0ds_logic.v(1335)
  wire Dj6ju6;  // ../RTL/cortexm0ds_logic.v(872)
  wire Dj7iu6;  // ../RTL/cortexm0ds_logic.v(404)
  wire Dj7pw6;  // ../RTL/cortexm0ds_logic.v(1428)
  wire Dj8ow6;  // ../RTL/cortexm0ds_logic.v(960)
  wire Djeiu6;  // ../RTL/cortexm0ds_logic.v(498)
  wire Djfow6;  // ../RTL/cortexm0ds_logic.v(1054)
  wire Djliu6;  // ../RTL/cortexm0ds_logic.v(591)
  wire Djmow6;  // ../RTL/cortexm0ds_logic.v(1148)
  wire Djsiu6;  // ../RTL/cortexm0ds_logic.v(685)
  wire Djthu6;  // ../RTL/cortexm0ds_logic.v(217)
  wire Djtow6;  // ../RTL/cortexm0ds_logic.v(1241)
  wire Djziu6;  // ../RTL/cortexm0ds_logic.v(778)
  wire Dk5ju6;  // ../RTL/cortexm0ds_logic.v(859)
  wire Dk6bx6;  // ../RTL/cortexm0ds_logic.v(1691)
  wire Dk6iu6;  // ../RTL/cortexm0ds_logic.v(391)
  wire Dk6pw6;  // ../RTL/cortexm0ds_logic.v(1415)
  wire Dk7ow6;  // ../RTL/cortexm0ds_logic.v(947)
  wire Dk9bx6;  // ../RTL/cortexm0ds_logic.v(1696)
  wire Dkdiu6;  // ../RTL/cortexm0ds_logic.v(485)
  wire Dkdpw6;  // ../RTL/cortexm0ds_logic.v(1509)
  wire Dkeow6;  // ../RTL/cortexm0ds_logic.v(1041)
  wire Dkfhu6;  // ../RTL/cortexm0ds_logic.v(124)
  wire Dkkiu6;  // ../RTL/cortexm0ds_logic.v(578)
  wire Dklow6;  // ../RTL/cortexm0ds_logic.v(1135)
  wire Dkriu6;  // ../RTL/cortexm0ds_logic.v(672)
  wire Dkshu6;  // ../RTL/cortexm0ds_logic.v(204)
  wire Dksow6;  // ../RTL/cortexm0ds_logic.v(1228)
  wire Dkyiu6;  // ../RTL/cortexm0ds_logic.v(765)
  wire Dkzhu6;  // ../RTL/cortexm0ds_logic.v(297)
  wire Dkzow6;  // ../RTL/cortexm0ds_logic.v(1322)
  wire Dl4ju6;  // ../RTL/cortexm0ds_logic.v(846)
  wire Dl5iu6;  // ../RTL/cortexm0ds_logic.v(378)
  wire Dl5pw6;  // ../RTL/cortexm0ds_logic.v(1402)
  wire Dl6ow6;  // ../RTL/cortexm0ds_logic.v(934)
  wire Dlciu6;  // ../RTL/cortexm0ds_logic.v(472)
  wire Dlcpw6;  // ../RTL/cortexm0ds_logic.v(1496)
  wire Dldow6;  // ../RTL/cortexm0ds_logic.v(1028)
  wire Dljiu6;  // ../RTL/cortexm0ds_logic.v(565)
  wire Dlkow6;  // ../RTL/cortexm0ds_logic.v(1122)
  wire Dlqiu6;  // ../RTL/cortexm0ds_logic.v(659)
  wire Dlrhu6;  // ../RTL/cortexm0ds_logic.v(191)
  wire Dlrow6;  // ../RTL/cortexm0ds_logic.v(1215)
  wire Dlxiu6;  // ../RTL/cortexm0ds_logic.v(752)
  wire Dlyhu6;  // ../RTL/cortexm0ds_logic.v(284)
  wire Dlyow6;  // ../RTL/cortexm0ds_logic.v(1309)
  wire Dm3ju6;  // ../RTL/cortexm0ds_logic.v(833)
  wire Dm4iu6;  // ../RTL/cortexm0ds_logic.v(365)
  wire Dm4pw6;  // ../RTL/cortexm0ds_logic.v(1389)
  wire Dm6bx6;  // ../RTL/cortexm0ds_logic.v(1691)
  wire Dmaju6;  // ../RTL/cortexm0ds_logic.v(927)
  wire Dmbiu6;  // ../RTL/cortexm0ds_logic.v(459)
  wire Dmbpw6;  // ../RTL/cortexm0ds_logic.v(1483)
  wire Dmcow6;  // ../RTL/cortexm0ds_logic.v(1015)
  wire Dmeax6;  // ../RTL/cortexm0ds_logic.v(1640)
  wire Dmiiu6;  // ../RTL/cortexm0ds_logic.v(552)
  wire Dmjow6;  // ../RTL/cortexm0ds_logic.v(1109)
  wire Dmmhu6;  // ../RTL/cortexm0ds_logic.v(142)
  wire Dmpiu6;  // ../RTL/cortexm0ds_logic.v(646)
  wire Dmqhu6;  // ../RTL/cortexm0ds_logic.v(178)
  wire Dmqow6;  // ../RTL/cortexm0ds_logic.v(1202)
  wire Dmwiu6;  // ../RTL/cortexm0ds_logic.v(739)
  wire Dmxhu6;  // ../RTL/cortexm0ds_logic.v(271)
  wire Dmxow6;  // ../RTL/cortexm0ds_logic.v(1296)
  wire Dn2ju6;  // ../RTL/cortexm0ds_logic.v(820)
  wire Dn3iu6;  // ../RTL/cortexm0ds_logic.v(352)
  wire Dn3pw6;  // ../RTL/cortexm0ds_logic.v(1376)
  wire Dn9ju6;  // ../RTL/cortexm0ds_logic.v(914)
  wire Dnaiu6;  // ../RTL/cortexm0ds_logic.v(446)
  wire Dnapw6;  // ../RTL/cortexm0ds_logic.v(1470)
  wire Dnbow6;  // ../RTL/cortexm0ds_logic.v(1002)
  wire Dncax6;  // ../RTL/cortexm0ds_logic.v(1636)
  wire Dnfhu6;  // ../RTL/cortexm0ds_logic.v(124)
  wire Dnhiu6;  // ../RTL/cortexm0ds_logic.v(539)
  wire Dniow6;  // ../RTL/cortexm0ds_logic.v(1096)
  wire Dnoiu6;  // ../RTL/cortexm0ds_logic.v(633)
  wire Dnphu6;  // ../RTL/cortexm0ds_logic.v(165)
  wire Dnpow6;  // ../RTL/cortexm0ds_logic.v(1189)
  wire Dnviu6;  // ../RTL/cortexm0ds_logic.v(726)
  wire Dnwhu6;  // ../RTL/cortexm0ds_logic.v(258)
  wire Dnwow6;  // ../RTL/cortexm0ds_logic.v(1283)
  wire Do1ju6;  // ../RTL/cortexm0ds_logic.v(807)
  wire Do2iu6;  // ../RTL/cortexm0ds_logic.v(339)
  wire Do2pw6;  // ../RTL/cortexm0ds_logic.v(1363)
  wire Do6bx6;  // ../RTL/cortexm0ds_logic.v(1691)
  wire Do8ju6;  // ../RTL/cortexm0ds_logic.v(901)
  wire Do9iu6;  // ../RTL/cortexm0ds_logic.v(433)
  wire Do9pw6;  // ../RTL/cortexm0ds_logic.v(1457)
  wire Doaow6;  // ../RTL/cortexm0ds_logic.v(989)
  wire Dogiu6;  // ../RTL/cortexm0ds_logic.v(526)
  wire Dohow6;  // ../RTL/cortexm0ds_logic.v(1083)
  wire Doniu6;  // ../RTL/cortexm0ds_logic.v(620)
  wire Doohu6;  // ../RTL/cortexm0ds_logic.v(152)
  wire Dooow6;  // ../RTL/cortexm0ds_logic.v(1176)
  wire Dorpw6;  // ../RTL/cortexm0ds_logic.v(1602)
  wire Douiu6;  // ../RTL/cortexm0ds_logic.v(713)
  wire Dovhu6;  // ../RTL/cortexm0ds_logic.v(245)
  wire Dovow6;  // ../RTL/cortexm0ds_logic.v(1270)
  wire Dp0ju6;  // ../RTL/cortexm0ds_logic.v(794)
  wire Dp1iu6;  // ../RTL/cortexm0ds_logic.v(326)
  wire Dp1pw6;  // ../RTL/cortexm0ds_logic.v(1350)
  wire Dp7ju6;  // ../RTL/cortexm0ds_logic.v(888)
  wire Dp8iu6;  // ../RTL/cortexm0ds_logic.v(420)
  wire Dp8pw6;  // ../RTL/cortexm0ds_logic.v(1444)
  wire Dp9ow6;  // ../RTL/cortexm0ds_logic.v(976)
  wire Dpfiu6;  // ../RTL/cortexm0ds_logic.v(513)
  wire Dpgow6;  // ../RTL/cortexm0ds_logic.v(1070)
  wire Dplhu6;  // ../RTL/cortexm0ds_logic.v(140)
  wire Dpmiu6;  // ../RTL/cortexm0ds_logic.v(607)
  wire Dpnow6;  // ../RTL/cortexm0ds_logic.v(1163)
  wire Dptiu6;  // ../RTL/cortexm0ds_logic.v(700)
  wire Dpuhu6;  // ../RTL/cortexm0ds_logic.v(232)
  wire Dpuow6;  // ../RTL/cortexm0ds_logic.v(1257)
  wire Dpwpw6;  // ../RTL/cortexm0ds_logic.v(1611)
  wire Dq0iu6;  // ../RTL/cortexm0ds_logic.v(313)
  wire Dq0pw6;  // ../RTL/cortexm0ds_logic.v(1337)
  wire Dq6bx6;  // ../RTL/cortexm0ds_logic.v(1691)
  wire Dq6ju6;  // ../RTL/cortexm0ds_logic.v(875)
  wire Dq7iu6;  // ../RTL/cortexm0ds_logic.v(407)
  wire Dq7pw6;  // ../RTL/cortexm0ds_logic.v(1431)
  wire Dq8ow6;  // ../RTL/cortexm0ds_logic.v(963)
  wire Dqeiu6;  // ../RTL/cortexm0ds_logic.v(500)
  wire Dqfhu6;  // ../RTL/cortexm0ds_logic.v(125)
  wire Dqfow6;  // ../RTL/cortexm0ds_logic.v(1057)
  wire Dqkbx6;  // ../RTL/cortexm0ds_logic.v(1717)
  wire Dqliu6;  // ../RTL/cortexm0ds_logic.v(594)
  wire Dqmow6;  // ../RTL/cortexm0ds_logic.v(1150)
  wire Dqsiu6;  // ../RTL/cortexm0ds_logic.v(687)
  wire Dqthu6;  // ../RTL/cortexm0ds_logic.v(219)
  wire Dqtow6;  // ../RTL/cortexm0ds_logic.v(1244)
  wire Dqziu6;  // ../RTL/cortexm0ds_logic.v(781)
  wire Dr5ju6;  // ../RTL/cortexm0ds_logic.v(862)
  wire Dr6iu6;  // ../RTL/cortexm0ds_logic.v(394)
  wire Dr6pw6;  // ../RTL/cortexm0ds_logic.v(1418)
  wire Dr7ow6;  // ../RTL/cortexm0ds_logic.v(950)
  wire Drcbx6;  // ../RTL/cortexm0ds_logic.v(1702)
  wire Drdiu6;  // ../RTL/cortexm0ds_logic.v(487)
  wire Drdpw6;  // ../RTL/cortexm0ds_logic.v(1512)
  wire Dreow6;  // ../RTL/cortexm0ds_logic.v(1044)
  wire Drhax6;  // ../RTL/cortexm0ds_logic.v(1646)
  wire Drhhu6;  // ../RTL/cortexm0ds_logic.v(129)
  wire Drkiu6;  // ../RTL/cortexm0ds_logic.v(581)
  wire Drlow6;  // ../RTL/cortexm0ds_logic.v(1137)
  wire Drriu6;  // ../RTL/cortexm0ds_logic.v(674)
  wire Drshu6;  // ../RTL/cortexm0ds_logic.v(206)
  wire Drsow6;  // ../RTL/cortexm0ds_logic.v(1231)
  wire Dryiu6;  // ../RTL/cortexm0ds_logic.v(768)
  wire Drzhu6;  // ../RTL/cortexm0ds_logic.v(300)
  wire Drzow6;  // ../RTL/cortexm0ds_logic.v(1324)
  wire Ds4ju6;  // ../RTL/cortexm0ds_logic.v(849)
  wire Ds5iu6;  // ../RTL/cortexm0ds_logic.v(381)
  wire Ds5pw6;  // ../RTL/cortexm0ds_logic.v(1405)
  wire Ds6ow6;  // ../RTL/cortexm0ds_logic.v(937)
  wire Dsciu6;  // ../RTL/cortexm0ds_logic.v(474)
  wire Dscpw6;  // ../RTL/cortexm0ds_logic.v(1499)
  wire Dsdow6;  // ../RTL/cortexm0ds_logic.v(1031)
  wire Dsjiu6;  // ../RTL/cortexm0ds_logic.v(568)
  wire Dskow6;  // ../RTL/cortexm0ds_logic.v(1124)
  wire Dsqiu6;  // ../RTL/cortexm0ds_logic.v(661)
  wire Dsrhu6;  // ../RTL/cortexm0ds_logic.v(193)
  wire Dsrow6;  // ../RTL/cortexm0ds_logic.v(1218)
  wire Dsxiu6;  // ../RTL/cortexm0ds_logic.v(755)
  wire Dsyhu6;  // ../RTL/cortexm0ds_logic.v(287)
  wire Dsyow6;  // ../RTL/cortexm0ds_logic.v(1311)
  wire Dt1bx6;  // ../RTL/cortexm0ds_logic.v(1682)
  wire Dt3ju6;  // ../RTL/cortexm0ds_logic.v(836)
  wire Dt4iu6;  // ../RTL/cortexm0ds_logic.v(368)
  wire Dt4pw6;  // ../RTL/cortexm0ds_logic.v(1392)
  wire Dtaju6;  // ../RTL/cortexm0ds_logic.v(929)
  wire Dtbiu6;  // ../RTL/cortexm0ds_logic.v(461)
  wire Dtbpw6;  // ../RTL/cortexm0ds_logic.v(1486)
  wire Dtcow6;  // ../RTL/cortexm0ds_logic.v(1018)
  wire Dtiiu6;  // ../RTL/cortexm0ds_logic.v(555)
  wire Dtjow6;  // ../RTL/cortexm0ds_logic.v(1111)
  wire Dtnhu6;  // ../RTL/cortexm0ds_logic.v(145)
  wire Dtpax6;  // ../RTL/cortexm0ds_logic.v(1661)
  wire Dtpiu6;  // ../RTL/cortexm0ds_logic.v(648)
  wire Dtqhu6;  // ../RTL/cortexm0ds_logic.v(180)
  wire Dtqow6;  // ../RTL/cortexm0ds_logic.v(1205)
  wire Dtwiu6;  // ../RTL/cortexm0ds_logic.v(742)
  wire Dtxhu6;  // ../RTL/cortexm0ds_logic.v(274)
  wire Dtxow6;  // ../RTL/cortexm0ds_logic.v(1298)
  wire Du2ju6;  // ../RTL/cortexm0ds_logic.v(823)
  wire Du3iu6;  // ../RTL/cortexm0ds_logic.v(355)
  wire Du3pw6;  // ../RTL/cortexm0ds_logic.v(1379)
  wire Du9ju6;  // ../RTL/cortexm0ds_logic.v(916)
  wire Duaiu6;  // ../RTL/cortexm0ds_logic.v(448)
  wire Duapw6;  // ../RTL/cortexm0ds_logic.v(1473)
  wire Dubow6;  // ../RTL/cortexm0ds_logic.v(1005)
  wire Dugax6;  // ../RTL/cortexm0ds_logic.v(1644)
  wire Duhiu6;  // ../RTL/cortexm0ds_logic.v(542)
  wire Duiow6;  // ../RTL/cortexm0ds_logic.v(1098)
  wire Duoiu6;  // ../RTL/cortexm0ds_logic.v(635)
  wire Duphu6;  // ../RTL/cortexm0ds_logic.v(167)
  wire Dupow6;  // ../RTL/cortexm0ds_logic.v(1192)
  wire Duviu6;  // ../RTL/cortexm0ds_logic.v(729)
  wire Duwhu6;  // ../RTL/cortexm0ds_logic.v(261)
  wire Duwow6;  // ../RTL/cortexm0ds_logic.v(1285)
  wire Dv1ju6;  // ../RTL/cortexm0ds_logic.v(810)
  wire Dv2bx6;  // ../RTL/cortexm0ds_logic.v(1684)
  wire Dv2iu6;  // ../RTL/cortexm0ds_logic.v(342)
  wire Dv2pw6;  // ../RTL/cortexm0ds_logic.v(1366)
  wire Dv8ju6;  // ../RTL/cortexm0ds_logic.v(903)
  wire Dv9iu6;  // ../RTL/cortexm0ds_logic.v(435)
  wire Dv9pw6;  // ../RTL/cortexm0ds_logic.v(1460)
  wire Dvaow6;  // ../RTL/cortexm0ds_logic.v(992)
  wire Dvghu6;  // ../RTL/cortexm0ds_logic.v(127)
  wire Dvgiu6;  // ../RTL/cortexm0ds_logic.v(529)
  wire Dvhow6;  // ../RTL/cortexm0ds_logic.v(1085)
  wire Dvniu6;  // ../RTL/cortexm0ds_logic.v(622)
  wire Dvohu6;  // ../RTL/cortexm0ds_logic.v(154)
  wire Dvoow6;  // ../RTL/cortexm0ds_logic.v(1179)
  wire Dvuiu6;  // ../RTL/cortexm0ds_logic.v(716)
  wire Dvvhu6;  // ../RTL/cortexm0ds_logic.v(248)
  wire Dvvow6;  // ../RTL/cortexm0ds_logic.v(1272)
  wire Dw0ju6;  // ../RTL/cortexm0ds_logic.v(797)
  wire Dw1iu6;  // ../RTL/cortexm0ds_logic.v(329)
  wire Dw1pw6;  // ../RTL/cortexm0ds_logic.v(1353)
  wire Dw7ju6;  // ../RTL/cortexm0ds_logic.v(890)
  wire Dw8iu6;  // ../RTL/cortexm0ds_logic.v(422)
  wire Dw8pw6;  // ../RTL/cortexm0ds_logic.v(1447)
  wire Dw9ow6;  // ../RTL/cortexm0ds_logic.v(979)
  wire Dwfiu6;  // ../RTL/cortexm0ds_logic.v(516)
  wire Dwgow6;  // ../RTL/cortexm0ds_logic.v(1072)
  wire Dwmiu6;  // ../RTL/cortexm0ds_logic.v(609)
  wire Dwnow6;  // ../RTL/cortexm0ds_logic.v(1166)
  wire Dwtiu6;  // ../RTL/cortexm0ds_logic.v(703)
  wire Dwuhu6;  // ../RTL/cortexm0ds_logic.v(235)
  wire Dwuow6;  // ../RTL/cortexm0ds_logic.v(1259)
  wire Dx0iu6;  // ../RTL/cortexm0ds_logic.v(316)
  wire Dx0pw6;  // ../RTL/cortexm0ds_logic.v(1340)
  wire Dx6ju6;  // ../RTL/cortexm0ds_logic.v(877)
  wire Dx7iu6;  // ../RTL/cortexm0ds_logic.v(409)
  wire Dx7pw6;  // ../RTL/cortexm0ds_logic.v(1434)
  wire Dx8ow6;  // ../RTL/cortexm0ds_logic.v(966)
  wire Dxeiu6;  // ../RTL/cortexm0ds_logic.v(503)
  wire Dxfhu6;  // ../RTL/cortexm0ds_logic.v(125)
  wire Dxfow6;  // ../RTL/cortexm0ds_logic.v(1059)
  wire Dxliu6;  // ../RTL/cortexm0ds_logic.v(596)
  wire Dxmow6;  // ../RTL/cortexm0ds_logic.v(1153)
  wire Dxsiu6;  // ../RTL/cortexm0ds_logic.v(690)
  wire Dxthu6;  // ../RTL/cortexm0ds_logic.v(222)
  wire Dxtow6;  // ../RTL/cortexm0ds_logic.v(1246)
  wire Dxvpw6;  // ../RTL/cortexm0ds_logic.v(1609)
  wire Dxziu6;  // ../RTL/cortexm0ds_logic.v(784)
  wire Dy5ju6;  // ../RTL/cortexm0ds_logic.v(864)
  wire Dy6iu6;  // ../RTL/cortexm0ds_logic.v(396)
  wire Dy6pw6;  // ../RTL/cortexm0ds_logic.v(1421)
  wire Dy7ow6;  // ../RTL/cortexm0ds_logic.v(953)
  wire Dydiu6;  // ../RTL/cortexm0ds_logic.v(490)
  wire Dydpw6;  // ../RTL/cortexm0ds_logic.v(1514)
  wire Dyeow6;  // ../RTL/cortexm0ds_logic.v(1046)
  wire Dykiu6;  // ../RTL/cortexm0ds_logic.v(583)
  wire Dylow6;  // ../RTL/cortexm0ds_logic.v(1140)
  wire Dyriu6;  // ../RTL/cortexm0ds_logic.v(677)
  wire Dyshu6;  // ../RTL/cortexm0ds_logic.v(209)
  wire Dysow6;  // ../RTL/cortexm0ds_logic.v(1233)
  wire Dyyiu6;  // ../RTL/cortexm0ds_logic.v(771)
  wire Dyzhu6;  // ../RTL/cortexm0ds_logic.v(303)
  wire Dyzow6;  // ../RTL/cortexm0ds_logic.v(1327)
  wire Dz4ju6;  // ../RTL/cortexm0ds_logic.v(851)
  wire Dz5iu6;  // ../RTL/cortexm0ds_logic.v(383)
  wire Dz5pw6;  // ../RTL/cortexm0ds_logic.v(1408)
  wire Dz6ow6;  // ../RTL/cortexm0ds_logic.v(940)
  wire Dzciu6;  // ../RTL/cortexm0ds_logic.v(477)
  wire Dzcpw6;  // ../RTL/cortexm0ds_logic.v(1501)
  wire Dzdow6;  // ../RTL/cortexm0ds_logic.v(1033)
  wire Dzjiu6;  // ../RTL/cortexm0ds_logic.v(570)
  wire Dzkow6;  // ../RTL/cortexm0ds_logic.v(1127)
  wire Dzqiu6;  // ../RTL/cortexm0ds_logic.v(664)
  wire Dzrhu6;  // ../RTL/cortexm0ds_logic.v(196)
  wire Dzrow6;  // ../RTL/cortexm0ds_logic.v(1220)
  wire Dzvpw6;  // ../RTL/cortexm0ds_logic.v(1610)
  wire Dzxiu6;  // ../RTL/cortexm0ds_logic.v(758)
  wire Dzyhu6;  // ../RTL/cortexm0ds_logic.v(290)
  wire Dzyow6;  // ../RTL/cortexm0ds_logic.v(1314)
  wire E01ju6;  // ../RTL/cortexm0ds_logic.v(798)
  wire E02iu6;  // ../RTL/cortexm0ds_logic.v(330)
  wire E02pw6;  // ../RTL/cortexm0ds_logic.v(1355)
  wire E05bx6;  // ../RTL/cortexm0ds_logic.v(1688)
  wire E08ju6;  // ../RTL/cortexm0ds_logic.v(892)
  wire E09iu6;  // ../RTL/cortexm0ds_logic.v(424)
  wire E09pw6;  // ../RTL/cortexm0ds_logic.v(1448)
  wire E0aow6;  // ../RTL/cortexm0ds_logic.v(980)
  wire E0giu6;  // ../RTL/cortexm0ds_logic.v(517)
  wire E0how6;  // ../RTL/cortexm0ds_logic.v(1074)
  wire E0ihu6;  // ../RTL/cortexm0ds_logic.v(130)
  wire E0niu6;  // ../RTL/cortexm0ds_logic.v(611)
  wire E0oow6;  // ../RTL/cortexm0ds_logic.v(1167)
  wire E0uiu6;  // ../RTL/cortexm0ds_logic.v(705)
  wire E0vhu6;  // ../RTL/cortexm0ds_logic.v(237)
  wire E0vow6;  // ../RTL/cortexm0ds_logic.v(1261)
  wire E10ju6;  // ../RTL/cortexm0ds_logic.v(785)
  wire E11iu6;  // ../RTL/cortexm0ds_logic.v(317)
  wire E11pw6;  // ../RTL/cortexm0ds_logic.v(1342)
  wire E17ju6;  // ../RTL/cortexm0ds_logic.v(879)
  wire E18iu6;  // ../RTL/cortexm0ds_logic.v(411)
  wire E18pw6;  // ../RTL/cortexm0ds_logic.v(1435)
  wire E19ow6;  // ../RTL/cortexm0ds_logic.v(967)
  wire E1fiu6;  // ../RTL/cortexm0ds_logic.v(504)
  wire E1gow6;  // ../RTL/cortexm0ds_logic.v(1061)
  wire E1miu6;  // ../RTL/cortexm0ds_logic.v(598)
  wire E1now6;  // ../RTL/cortexm0ds_logic.v(1154)
  wire E1npw6;  // ../RTL/cortexm0ds_logic.v(1593)
  wire E1tiu6;  // ../RTL/cortexm0ds_logic.v(692)
  wire E1uhu6;  // ../RTL/cortexm0ds_logic.v(224)
  wire E1uow6;  // ../RTL/cortexm0ds_logic.v(1248)
  wire E20iu6;  // ../RTL/cortexm0ds_logic.v(304)
  wire E20pw6;  // ../RTL/cortexm0ds_logic.v(1329)
  wire E26ju6;  // ../RTL/cortexm0ds_logic.v(866)
  wire E27iu6;  // ../RTL/cortexm0ds_logic.v(398)
  wire E27pw6;  // ../RTL/cortexm0ds_logic.v(1422)
  wire E28ow6;  // ../RTL/cortexm0ds_logic.v(954)
  wire E2eiu6;  // ../RTL/cortexm0ds_logic.v(491)
  wire E2epw6;  // ../RTL/cortexm0ds_logic.v(1516)
  wire E2fow6;  // ../RTL/cortexm0ds_logic.v(1048)
  wire E2liu6;  // ../RTL/cortexm0ds_logic.v(585)
  wire E2mow6;  // ../RTL/cortexm0ds_logic.v(1141)
  wire E2siu6;  // ../RTL/cortexm0ds_logic.v(679)
  wire E2thu6;  // ../RTL/cortexm0ds_logic.v(211)
  wire E2tow6;  // ../RTL/cortexm0ds_logic.v(1235)
  wire E2ziu6;  // ../RTL/cortexm0ds_logic.v(772)
  wire E34bx6;  // ../RTL/cortexm0ds_logic.v(1686)
  wire E35ju6;  // ../RTL/cortexm0ds_logic.v(853)
  wire E36iu6;  // ../RTL/cortexm0ds_logic.v(385)
  wire E36pw6;  // ../RTL/cortexm0ds_logic.v(1409)
  wire E37ow6;  // ../RTL/cortexm0ds_logic.v(941)
  wire E3diu6;  // ../RTL/cortexm0ds_logic.v(478)
  wire E3dpw6;  // ../RTL/cortexm0ds_logic.v(1503)
  wire E3eow6;  // ../RTL/cortexm0ds_logic.v(1035)
  wire E3kiu6;  // ../RTL/cortexm0ds_logic.v(572)
  wire E3low6;  // ../RTL/cortexm0ds_logic.v(1128)
  wire E3npw6;  // ../RTL/cortexm0ds_logic.v(1593)
  wire E3riu6;  // ../RTL/cortexm0ds_logic.v(666)
  wire E3shu6;  // ../RTL/cortexm0ds_logic.v(198)
  wire E3sow6;  // ../RTL/cortexm0ds_logic.v(1222)
  wire E3yiu6;  // ../RTL/cortexm0ds_logic.v(759)
  wire E3zhu6;  // ../RTL/cortexm0ds_logic.v(291)
  wire E3zow6;  // ../RTL/cortexm0ds_logic.v(1316)
  wire E44ju6;  // ../RTL/cortexm0ds_logic.v(840)
  wire E45iu6;  // ../RTL/cortexm0ds_logic.v(372)
  wire E45pw6;  // ../RTL/cortexm0ds_logic.v(1396)
  wire E4ciu6;  // ../RTL/cortexm0ds_logic.v(465)
  wire E4cpw6;  // ../RTL/cortexm0ds_logic.v(1490)
  wire E4dow6;  // ../RTL/cortexm0ds_logic.v(1022)
  wire E4jiu6;  // ../RTL/cortexm0ds_logic.v(559)
  wire E4kow6;  // ../RTL/cortexm0ds_logic.v(1115)
  wire E4qiu6;  // ../RTL/cortexm0ds_logic.v(653)
  wire E4rhu6;  // ../RTL/cortexm0ds_logic.v(185)
  wire E4row6;  // ../RTL/cortexm0ds_logic.v(1209)
  wire E4xiu6;  // ../RTL/cortexm0ds_logic.v(746)
  wire E4yhu6;  // ../RTL/cortexm0ds_logic.v(278)
  wire E4yow6;  // ../RTL/cortexm0ds_logic.v(1303)
  wire E53ju6;  // ../RTL/cortexm0ds_logic.v(827)
  wire E54iu6;  // ../RTL/cortexm0ds_logic.v(359)
  wire E54pw6;  // ../RTL/cortexm0ds_logic.v(1383)
  wire E5aju6;  // ../RTL/cortexm0ds_logic.v(920)
  wire E5biu6;  // ../RTL/cortexm0ds_logic.v(452)
  wire E5bpw6;  // ../RTL/cortexm0ds_logic.v(1477)
  wire E5cow6;  // ../RTL/cortexm0ds_logic.v(1009)
  wire E5ehu6;  // ../RTL/cortexm0ds_logic.v(121)
  wire E5hhu6;  // ../RTL/cortexm0ds_logic.v(128)
  wire E5iiu6;  // ../RTL/cortexm0ds_logic.v(546)
  wire E5jow6;  // ../RTL/cortexm0ds_logic.v(1102)
  wire E5npw6;  // ../RTL/cortexm0ds_logic.v(1594)
  wire E5pax6;  // ../RTL/cortexm0ds_logic.v(1660)
  wire E5piu6;  // ../RTL/cortexm0ds_logic.v(640)
  wire E5qhu6;  // ../RTL/cortexm0ds_logic.v(172)
  wire E5qow6;  // ../RTL/cortexm0ds_logic.v(1196)
  wire E5wiu6;  // ../RTL/cortexm0ds_logic.v(733)
  wire E5xhu6;  // ../RTL/cortexm0ds_logic.v(265)
  wire E5xow6;  // ../RTL/cortexm0ds_logic.v(1290)
  wire E62ju6;  // ../RTL/cortexm0ds_logic.v(814)
  wire E63iu6;  // ../RTL/cortexm0ds_logic.v(346)
  wire E63pw6;  // ../RTL/cortexm0ds_logic.v(1370)
  wire E69ju6;  // ../RTL/cortexm0ds_logic.v(907)
  wire E6aiu6;  // ../RTL/cortexm0ds_logic.v(439)
  wire E6apw6;  // ../RTL/cortexm0ds_logic.v(1464)
  wire E6bow6;  // ../RTL/cortexm0ds_logic.v(996)
  wire E6hiu6;  // ../RTL/cortexm0ds_logic.v(533)
  wire E6iax6;  // ../RTL/cortexm0ds_logic.v(1647)
  wire E6iow6;  // ../RTL/cortexm0ds_logic.v(1089)
  wire E6oiu6;  // ../RTL/cortexm0ds_logic.v(627)
  wire E6phu6;  // ../RTL/cortexm0ds_logic.v(159)
  wire E6pow6;  // ../RTL/cortexm0ds_logic.v(1183)
  wire E6viu6;  // ../RTL/cortexm0ds_logic.v(720)
  wire E6whu6;  // ../RTL/cortexm0ds_logic.v(252)
  wire E6wow6;  // ../RTL/cortexm0ds_logic.v(1277)
  wire E71ju6;  // ../RTL/cortexm0ds_logic.v(801)
  wire E72iu6;  // ../RTL/cortexm0ds_logic.v(333)
  wire E72pw6;  // ../RTL/cortexm0ds_logic.v(1357)
  wire E78ju6;  // ../RTL/cortexm0ds_logic.v(894)
  wire E79iu6;  // ../RTL/cortexm0ds_logic.v(426)
  wire E79pw6;  // ../RTL/cortexm0ds_logic.v(1451)
  wire E7aow6;  // ../RTL/cortexm0ds_logic.v(983)
  wire E7giu6;  // ../RTL/cortexm0ds_logic.v(520)
  wire E7how6;  // ../RTL/cortexm0ds_logic.v(1076)
  wire E7niu6;  // ../RTL/cortexm0ds_logic.v(614)
  wire E7npw6;  // ../RTL/cortexm0ds_logic.v(1594)
  wire E7oow6;  // ../RTL/cortexm0ds_logic.v(1170)
  wire E7pax6;  // ../RTL/cortexm0ds_logic.v(1660)
  wire E7uiu6;  // ../RTL/cortexm0ds_logic.v(707)
  wire E7vhu6;  // ../RTL/cortexm0ds_logic.v(239)
  wire E7vow6;  // ../RTL/cortexm0ds_logic.v(1264)
  wire E80ju6;  // ../RTL/cortexm0ds_logic.v(788)
  wire E81iu6;  // ../RTL/cortexm0ds_logic.v(320)
  wire E81pw6;  // ../RTL/cortexm0ds_logic.v(1344)
  wire E87ju6;  // ../RTL/cortexm0ds_logic.v(881)
  wire E88iu6;  // ../RTL/cortexm0ds_logic.v(413)
  wire E88pw6;  // ../RTL/cortexm0ds_logic.v(1438)
  wire E89ow6;  // ../RTL/cortexm0ds_logic.v(970)
  wire E8fiu6;  // ../RTL/cortexm0ds_logic.v(507)
  wire E8gow6;  // ../RTL/cortexm0ds_logic.v(1063)
  wire E8iax6;  // ../RTL/cortexm0ds_logic.v(1647)
  wire E8mhu6;  // ../RTL/cortexm0ds_logic.v(141)
  wire E8miu6;  // ../RTL/cortexm0ds_logic.v(601)
  wire E8now6;  // ../RTL/cortexm0ds_logic.v(1157)
  wire E8tiu6;  // ../RTL/cortexm0ds_logic.v(694)
  wire E8uhu6;  // ../RTL/cortexm0ds_logic.v(226)
  wire E8uow6;  // ../RTL/cortexm0ds_logic.v(1251)
  wire E90bx6;  // ../RTL/cortexm0ds_logic.v(1680)
  wire E90iu6;  // ../RTL/cortexm0ds_logic.v(307)
  wire E90pw6;  // ../RTL/cortexm0ds_logic.v(1331)
  wire E96ju6;  // ../RTL/cortexm0ds_logic.v(868)
  wire E97ax6;  // ../RTL/cortexm0ds_logic.v(1626)
  wire E97iu6;  // ../RTL/cortexm0ds_logic.v(400)
  wire E97pw6;  // ../RTL/cortexm0ds_logic.v(1425)
  wire E98ow6;  // ../RTL/cortexm0ds_logic.v(957)
  wire E9eiu6;  // ../RTL/cortexm0ds_logic.v(494)
  wire E9fow6;  // ../RTL/cortexm0ds_logic.v(1050)
  wire E9liu6;  // ../RTL/cortexm0ds_logic.v(588)
  wire E9mow6;  // ../RTL/cortexm0ds_logic.v(1144)
  wire E9npw6;  // ../RTL/cortexm0ds_logic.v(1594)
  wire E9pax6;  // ../RTL/cortexm0ds_logic.v(1660)
  wire E9siu6;  // ../RTL/cortexm0ds_logic.v(681)
  wire E9thu6;  // ../RTL/cortexm0ds_logic.v(213)
  wire E9tow6;  // ../RTL/cortexm0ds_logic.v(1238)
  wire E9ziu6;  // ../RTL/cortexm0ds_logic.v(775)
  wire Ea5ju6;  // ../RTL/cortexm0ds_logic.v(855)
  wire Ea6iu6;  // ../RTL/cortexm0ds_logic.v(387)
  wire Ea6pw6;  // ../RTL/cortexm0ds_logic.v(1412)
  wire Ea7ow6;  // ../RTL/cortexm0ds_logic.v(944)
  wire Eadiu6;  // ../RTL/cortexm0ds_logic.v(481)
  wire Eadpw6;  // ../RTL/cortexm0ds_logic.v(1505)
  wire Eaeow6;  // ../RTL/cortexm0ds_logic.v(1037)
  wire Eafax6;  // ../RTL/cortexm0ds_logic.v(1641)
  wire Eagax6;  // ../RTL/cortexm0ds_logic.v(1643)
  wire Eakiu6;  // ../RTL/cortexm0ds_logic.v(575)
  wire Ealow6;  // ../RTL/cortexm0ds_logic.v(1131)
  wire Eariu6;  // ../RTL/cortexm0ds_logic.v(668)
  wire Eashu6;  // ../RTL/cortexm0ds_logic.v(200)
  wire Easow6;  // ../RTL/cortexm0ds_logic.v(1225)
  wire Eayiu6;  // ../RTL/cortexm0ds_logic.v(762)
  wire Eazhu6;  // ../RTL/cortexm0ds_logic.v(294)
  wire Eazow6;  // ../RTL/cortexm0ds_logic.v(1318)
  wire Eb4ju6;  // ../RTL/cortexm0ds_logic.v(842)
  wire Eb5iu6;  // ../RTL/cortexm0ds_logic.v(374)
  wire Eb5pw6;  // ../RTL/cortexm0ds_logic.v(1399)
  wire Eb6ow6;  // ../RTL/cortexm0ds_logic.v(931)
  wire Ebciu6;  // ../RTL/cortexm0ds_logic.v(468)
  wire Ebcpw6;  // ../RTL/cortexm0ds_logic.v(1492)
  wire Ebdow6;  // ../RTL/cortexm0ds_logic.v(1024)
  wire Ebjiu6;  // ../RTL/cortexm0ds_logic.v(562)
  wire Ebkow6;  // ../RTL/cortexm0ds_logic.v(1118)
  wire Eblhu6;  // ../RTL/cortexm0ds_logic.v(139)
  wire Ebnpw6;  // ../RTL/cortexm0ds_logic.v(1594)
  wire Ebpax6;  // ../RTL/cortexm0ds_logic.v(1660)
  wire Ebqiu6;  // ../RTL/cortexm0ds_logic.v(655)
  wire Ebrhu6;  // ../RTL/cortexm0ds_logic.v(187)
  wire Ebrow6;  // ../RTL/cortexm0ds_logic.v(1212)
  wire Ebxiu6;  // ../RTL/cortexm0ds_logic.v(749)
  wire Ebyhu6;  // ../RTL/cortexm0ds_logic.v(281)
  wire Ebyow6;  // ../RTL/cortexm0ds_logic.v(1305)
  wire Ec3ju6;  // ../RTL/cortexm0ds_logic.v(829)
  wire Ec4iu6;  // ../RTL/cortexm0ds_logic.v(361)
  wire Ec4pw6;  // ../RTL/cortexm0ds_logic.v(1386)
  wire Ecaju6;  // ../RTL/cortexm0ds_logic.v(923)
  wire Ecbiu6;  // ../RTL/cortexm0ds_logic.v(455)
  wire Ecbpw6;  // ../RTL/cortexm0ds_logic.v(1479)
  wire Eccow6;  // ../RTL/cortexm0ds_logic.v(1011)
  wire Eciiu6;  // ../RTL/cortexm0ds_logic.v(549)
  wire Ecjow6;  // ../RTL/cortexm0ds_logic.v(1105)
  wire Eclax6;  // ../RTL/cortexm0ds_logic.v(1653)
  wire Ecpiu6;  // ../RTL/cortexm0ds_logic.v(642)
  wire Ecqhu6;  // ../RTL/cortexm0ds_logic.v(174)
  wire Ecqow6;  // ../RTL/cortexm0ds_logic.v(1199)
  wire Ectax6;  // ../RTL/cortexm0ds_logic.v(1667)
  wire Ecwiu6;  // ../RTL/cortexm0ds_logic.v(736)
  wire Ecxhu6;  // ../RTL/cortexm0ds_logic.v(268)
  wire Ecxow6;  // ../RTL/cortexm0ds_logic.v(1292)
  wire Ed2ju6;  // ../RTL/cortexm0ds_logic.v(816)
  wire Ed3iu6;  // ../RTL/cortexm0ds_logic.v(348)
  wire Ed3pw6;  // ../RTL/cortexm0ds_logic.v(1373)
  wire Ed9ju6;  // ../RTL/cortexm0ds_logic.v(910)
  wire Edaiu6;  // ../RTL/cortexm0ds_logic.v(442)
  wire Edapw6;  // ../RTL/cortexm0ds_logic.v(1466)
  wire Edbow6;  // ../RTL/cortexm0ds_logic.v(998)
  wire Edehu6;  // ../RTL/cortexm0ds_logic.v(121)
  wire Edhiu6;  // ../RTL/cortexm0ds_logic.v(536)
  wire Ediow6;  // ../RTL/cortexm0ds_logic.v(1092)
  wire Edkhu6;  // ../RTL/cortexm0ds_logic.v(136)
  wire Ednpw6;  // ../RTL/cortexm0ds_logic.v(1594)
  wire Edoiu6;  // ../RTL/cortexm0ds_logic.v(629)
  wire Edpax6;  // ../RTL/cortexm0ds_logic.v(1660)
  wire Edphu6;  // ../RTL/cortexm0ds_logic.v(161)
  wire Edpow6;  // ../RTL/cortexm0ds_logic.v(1186)
  wire Edviu6;  // ../RTL/cortexm0ds_logic.v(723)
  wire Edwhu6;  // ../RTL/cortexm0ds_logic.v(255)
  wire Edwow6;  // ../RTL/cortexm0ds_logic.v(1279)
  wire Ee1ju6;  // ../RTL/cortexm0ds_logic.v(803)
  wire Ee2iu6;  // ../RTL/cortexm0ds_logic.v(335)
  wire Ee2pw6;  // ../RTL/cortexm0ds_logic.v(1360)
  wire Ee3bx6;  // ../RTL/cortexm0ds_logic.v(1685)
  wire Ee8ju6;  // ../RTL/cortexm0ds_logic.v(897)
  wire Ee9iu6;  // ../RTL/cortexm0ds_logic.v(429)
  wire Ee9pw6;  // ../RTL/cortexm0ds_logic.v(1453)
  wire Eeaow6;  // ../RTL/cortexm0ds_logic.v(985)
  wire Eegiu6;  // ../RTL/cortexm0ds_logic.v(523)
  wire Eehow6;  // ../RTL/cortexm0ds_logic.v(1079)
  wire Eeniu6;  // ../RTL/cortexm0ds_logic.v(616)
  wire Eeohu6;  // ../RTL/cortexm0ds_logic.v(148)
  wire Eeoow6;  // ../RTL/cortexm0ds_logic.v(1173)
  wire Eetax6;  // ../RTL/cortexm0ds_logic.v(1667)
  wire Eeuiu6;  // ../RTL/cortexm0ds_logic.v(710)
  wire Eevhu6;  // ../RTL/cortexm0ds_logic.v(242)
  wire Eevow6;  // ../RTL/cortexm0ds_logic.v(1266)
  wire Ef0ju6;  // ../RTL/cortexm0ds_logic.v(790)
  wire Ef1iu6;  // ../RTL/cortexm0ds_logic.v(322)
  wire Ef1pw6;  // ../RTL/cortexm0ds_logic.v(1347)
  wire Ef7ju6;  // ../RTL/cortexm0ds_logic.v(884)
  wire Ef8iu6;  // ../RTL/cortexm0ds_logic.v(416)
  wire Ef8pw6;  // ../RTL/cortexm0ds_logic.v(1440)
  wire Ef9ow6;  // ../RTL/cortexm0ds_logic.v(972)
  wire Efdax6;  // ../RTL/cortexm0ds_logic.v(1638)
  wire Effiu6;  // ../RTL/cortexm0ds_logic.v(510)
  wire Efgow6;  // ../RTL/cortexm0ds_logic.v(1066)
  wire Efjhu6;  // ../RTL/cortexm0ds_logic.v(134)
  wire Efmiu6;  // ../RTL/cortexm0ds_logic.v(603)
  wire Efnow6;  // ../RTL/cortexm0ds_logic.v(1160)
  wire Efnpw6;  // ../RTL/cortexm0ds_logic.v(1594)
  wire Efpax6;  // ../RTL/cortexm0ds_logic.v(1660)
  wire Eftiu6;  // ../RTL/cortexm0ds_logic.v(697)
  wire Efuhu6;  // ../RTL/cortexm0ds_logic.v(229)
  wire Efuow6;  // ../RTL/cortexm0ds_logic.v(1253)
  wire Eg0iu6;  // ../RTL/cortexm0ds_logic.v(309)
  wire Eg0pw6;  // ../RTL/cortexm0ds_logic.v(1334)
  wire Eg6ju6;  // ../RTL/cortexm0ds_logic.v(871)
  wire Eg7iu6;  // ../RTL/cortexm0ds_logic.v(403)
  wire Eg7pw6;  // ../RTL/cortexm0ds_logic.v(1427)
  wire Eg8ow6;  // ../RTL/cortexm0ds_logic.v(959)
  wire Egaax6;  // ../RTL/cortexm0ds_logic.v(1632)
  wire Egeiu6;  // ../RTL/cortexm0ds_logic.v(497)
  wire Egfow6;  // ../RTL/cortexm0ds_logic.v(1053)
  wire Eghbx6;  // ../RTL/cortexm0ds_logic.v(1711)
  wire Egliu6;  // ../RTL/cortexm0ds_logic.v(590)
  wire Egmow6;  // ../RTL/cortexm0ds_logic.v(1147)
  wire Egsiu6;  // ../RTL/cortexm0ds_logic.v(684)
  wire Egtax6;  // ../RTL/cortexm0ds_logic.v(1668)
  wire Egthu6;  // ../RTL/cortexm0ds_logic.v(216)
  wire Egtow6;  // ../RTL/cortexm0ds_logic.v(1240)
  wire Egziu6;  // ../RTL/cortexm0ds_logic.v(777)
  wire Eh5ju6;  // ../RTL/cortexm0ds_logic.v(858)
  wire Eh6iu6;  // ../RTL/cortexm0ds_logic.v(390)
  wire Eh6pw6;  // ../RTL/cortexm0ds_logic.v(1414)
  wire Eh7ow6;  // ../RTL/cortexm0ds_logic.v(946)
  wire Ehdiu6;  // ../RTL/cortexm0ds_logic.v(484)
  wire Ehdpw6;  // ../RTL/cortexm0ds_logic.v(1508)
  wire Eheow6;  // ../RTL/cortexm0ds_logic.v(1040)
  wire Ehihu6;  // ../RTL/cortexm0ds_logic.v(131)
  wire Ehkiu6;  // ../RTL/cortexm0ds_logic.v(577)
  wire Ehlow6;  // ../RTL/cortexm0ds_logic.v(1134)
  wire Ehnpw6;  // ../RTL/cortexm0ds_logic.v(1594)
  wire Ehpax6;  // ../RTL/cortexm0ds_logic.v(1660)
  wire Ehqpw6;  // ../RTL/cortexm0ds_logic.v(1600)
  wire Ehriu6;  // ../RTL/cortexm0ds_logic.v(671)
  wire Ehshu6;  // ../RTL/cortexm0ds_logic.v(203)
  wire Ehsow6;  // ../RTL/cortexm0ds_logic.v(1227)
  wire Ehyiu6;  // ../RTL/cortexm0ds_logic.v(764)
  wire Ehzhu6;  // ../RTL/cortexm0ds_logic.v(296)
  wire Ehzow6;  // ../RTL/cortexm0ds_logic.v(1321)
  wire Ei4ju6;  // ../RTL/cortexm0ds_logic.v(845)
  wire Ei5iu6;  // ../RTL/cortexm0ds_logic.v(377)
  wire Ei5pw6;  // ../RTL/cortexm0ds_logic.v(1401)
  wire Ei6ow6;  // ../RTL/cortexm0ds_logic.v(933)
  wire Eiciu6;  // ../RTL/cortexm0ds_logic.v(471)
  wire Eicpw6;  // ../RTL/cortexm0ds_logic.v(1495)
  wire Eidow6;  // ../RTL/cortexm0ds_logic.v(1027)
  wire Eijiu6;  // ../RTL/cortexm0ds_logic.v(564)
  wire Eikow6;  // ../RTL/cortexm0ds_logic.v(1121)
  wire Eiqiu6;  // ../RTL/cortexm0ds_logic.v(658)
  wire Eirhu6;  // ../RTL/cortexm0ds_logic.v(190)
  wire Eirow6;  // ../RTL/cortexm0ds_logic.v(1214)
  wire Eitax6;  // ../RTL/cortexm0ds_logic.v(1668)
  wire Eixiu6;  // ../RTL/cortexm0ds_logic.v(751)
  wire Eiyhu6;  // ../RTL/cortexm0ds_logic.v(283)
  wire Eiyow6;  // ../RTL/cortexm0ds_logic.v(1308)
  wire Ej3ju6;  // ../RTL/cortexm0ds_logic.v(832)
  wire Ej4iu6;  // ../RTL/cortexm0ds_logic.v(364)
  wire Ej4pw6;  // ../RTL/cortexm0ds_logic.v(1388)
  wire Ejaju6;  // ../RTL/cortexm0ds_logic.v(926)
  wire Ejbiu6;  // ../RTL/cortexm0ds_logic.v(458)
  wire Ejbpw6;  // ../RTL/cortexm0ds_logic.v(1482)
  wire Ejcow6;  // ../RTL/cortexm0ds_logic.v(1014)
  wire Ejiiu6;  // ../RTL/cortexm0ds_logic.v(551)
  wire Ejjow6;  // ../RTL/cortexm0ds_logic.v(1108)
  wire Ejnpw6;  // ../RTL/cortexm0ds_logic.v(1594)
  wire Ejpax6;  // ../RTL/cortexm0ds_logic.v(1660)
  wire Ejpiu6;  // ../RTL/cortexm0ds_logic.v(645)
  wire Ejqhu6;  // ../RTL/cortexm0ds_logic.v(177)
  wire Ejqow6;  // ../RTL/cortexm0ds_logic.v(1201)
  wire Ejwiu6;  // ../RTL/cortexm0ds_logic.v(738)
  wire Ejxhu6;  // ../RTL/cortexm0ds_logic.v(270)
  wire Ejxow6;  // ../RTL/cortexm0ds_logic.v(1295)
  wire Ek2ju6;  // ../RTL/cortexm0ds_logic.v(819)
  wire Ek3iu6;  // ../RTL/cortexm0ds_logic.v(351)
  wire Ek3pw6;  // ../RTL/cortexm0ds_logic.v(1375)
  wire Ek9ju6;  // ../RTL/cortexm0ds_logic.v(913)
  wire Ekaiu6;  // ../RTL/cortexm0ds_logic.v(445)
  wire Ekapw6;  // ../RTL/cortexm0ds_logic.v(1469)
  wire Ekbow6;  // ../RTL/cortexm0ds_logic.v(1001)
  wire Ekhiu6;  // ../RTL/cortexm0ds_logic.v(538)
  wire Ekiow6;  // ../RTL/cortexm0ds_logic.v(1095)
  wire Ekoiu6;  // ../RTL/cortexm0ds_logic.v(632)
  wire Ekphu6;  // ../RTL/cortexm0ds_logic.v(164)
  wire Ekpow6;  // ../RTL/cortexm0ds_logic.v(1188)
  wire Ektax6;  // ../RTL/cortexm0ds_logic.v(1668)
  wire Ekviu6;  // ../RTL/cortexm0ds_logic.v(725)
  wire Ekwhu6;  // ../RTL/cortexm0ds_logic.v(257)
  wire Ekwow6;  // ../RTL/cortexm0ds_logic.v(1282)
  wire El1ju6;  // ../RTL/cortexm0ds_logic.v(806)
  wire El2iu6;  // ../RTL/cortexm0ds_logic.v(338)
  wire El2pw6;  // ../RTL/cortexm0ds_logic.v(1362)
  wire El8ju6;  // ../RTL/cortexm0ds_logic.v(900)
  wire El9iu6;  // ../RTL/cortexm0ds_logic.v(432)
  wire El9pw6;  // ../RTL/cortexm0ds_logic.v(1456)
  wire Elaow6;  // ../RTL/cortexm0ds_logic.v(988)
  wire Elgax6;  // ../RTL/cortexm0ds_logic.v(1644)
  wire Elgiu6;  // ../RTL/cortexm0ds_logic.v(525)
  wire Elhow6;  // ../RTL/cortexm0ds_logic.v(1082)
  wire Eliax6;  // ../RTL/cortexm0ds_logic.v(1648)
  wire Elniu6;  // ../RTL/cortexm0ds_logic.v(619)
  wire Elnpw6;  // ../RTL/cortexm0ds_logic.v(1594)
  wire Elohu6;  // ../RTL/cortexm0ds_logic.v(151)
  wire Eloow6;  // ../RTL/cortexm0ds_logic.v(1175)
  wire Elpax6;  // ../RTL/cortexm0ds_logic.v(1661)
  wire Eluiu6;  // ../RTL/cortexm0ds_logic.v(712)
  wire Elvhu6;  // ../RTL/cortexm0ds_logic.v(244)
  wire Elvow6;  // ../RTL/cortexm0ds_logic.v(1269)
  wire Em0ju6;  // ../RTL/cortexm0ds_logic.v(793)
  wire Em1iu6;  // ../RTL/cortexm0ds_logic.v(325)
  wire Em1pw6;  // ../RTL/cortexm0ds_logic.v(1349)
  wire Em7ju6;  // ../RTL/cortexm0ds_logic.v(887)
  wire Em8iu6;  // ../RTL/cortexm0ds_logic.v(419)
  wire Em8pw6;  // ../RTL/cortexm0ds_logic.v(1443)
  wire Em9ow6;  // ../RTL/cortexm0ds_logic.v(975)
  wire Emfiu6;  // ../RTL/cortexm0ds_logic.v(512)
  wire Emgow6;  // ../RTL/cortexm0ds_logic.v(1069)
  wire Emmiu6;  // ../RTL/cortexm0ds_logic.v(606)
  wire Emnow6;  // ../RTL/cortexm0ds_logic.v(1162)
  wire Emrpw6;  // ../RTL/cortexm0ds_logic.v(1602)
  wire Emtax6;  // ../RTL/cortexm0ds_logic.v(1668)
  wire Emtiu6;  // ../RTL/cortexm0ds_logic.v(699)
  wire Emuhu6;  // ../RTL/cortexm0ds_logic.v(231)
  wire Emuow6;  // ../RTL/cortexm0ds_logic.v(1256)
  wire En0iu6;  // ../RTL/cortexm0ds_logic.v(312)
  wire En0pw6;  // ../RTL/cortexm0ds_logic.v(1336)
  wire En6ju6;  // ../RTL/cortexm0ds_logic.v(874)
  wire En7iu6;  // ../RTL/cortexm0ds_logic.v(406)
  wire En7pw6;  // ../RTL/cortexm0ds_logic.v(1430)
  wire En8ow6;  // ../RTL/cortexm0ds_logic.v(962)
  wire Eneiu6;  // ../RTL/cortexm0ds_logic.v(499)
  wire Enfow6;  // ../RTL/cortexm0ds_logic.v(1056)
  wire Enliu6;  // ../RTL/cortexm0ds_logic.v(593)
  wire Enmow6;  // ../RTL/cortexm0ds_logic.v(1149)
  wire Enpax6;  // ../RTL/cortexm0ds_logic.v(1661)
  wire Ensiu6;  // ../RTL/cortexm0ds_logic.v(686)
  wire Enthu6;  // ../RTL/cortexm0ds_logic.v(218)
  wire Entow6;  // ../RTL/cortexm0ds_logic.v(1243)
  wire Enziu6;  // ../RTL/cortexm0ds_logic.v(780)
  wire Eo5ju6;  // ../RTL/cortexm0ds_logic.v(861)
  wire Eo6iu6;  // ../RTL/cortexm0ds_logic.v(393)
  wire Eo6pw6;  // ../RTL/cortexm0ds_logic.v(1417)
  wire Eo7ow6;  // ../RTL/cortexm0ds_logic.v(949)
  wire Eodiu6;  // ../RTL/cortexm0ds_logic.v(486)
  wire Eodpw6;  // ../RTL/cortexm0ds_logic.v(1511)
  wire Eoeow6;  // ../RTL/cortexm0ds_logic.v(1043)
  wire Eokiu6;  // ../RTL/cortexm0ds_logic.v(580)
  wire Eolow6;  // ../RTL/cortexm0ds_logic.v(1136)
  wire Eoriu6;  // ../RTL/cortexm0ds_logic.v(673)
  wire Eoshu6;  // ../RTL/cortexm0ds_logic.v(205)
  wire Eosow6;  // ../RTL/cortexm0ds_logic.v(1230)
  wire Eotax6;  // ../RTL/cortexm0ds_logic.v(1668)
  wire Eoyiu6;  // ../RTL/cortexm0ds_logic.v(767)
  wire Eozhu6;  // ../RTL/cortexm0ds_logic.v(299)
  wire Eozow6;  // ../RTL/cortexm0ds_logic.v(1323)
  wire Ep4ju6;  // ../RTL/cortexm0ds_logic.v(848)
  wire Ep5iu6;  // ../RTL/cortexm0ds_logic.v(380)
  wire Ep5pw6;  // ../RTL/cortexm0ds_logic.v(1404)
  wire Ep6ow6;  // ../RTL/cortexm0ds_logic.v(936)
  wire Epciu6;  // ../RTL/cortexm0ds_logic.v(473)
  wire Epcpw6;  // ../RTL/cortexm0ds_logic.v(1498)
  wire Epdow6;  // ../RTL/cortexm0ds_logic.v(1030)
  wire Epjiu6;  // ../RTL/cortexm0ds_logic.v(567)
  wire Epkow6;  // ../RTL/cortexm0ds_logic.v(1123)
  wire Eppax6;  // ../RTL/cortexm0ds_logic.v(1661)
  wire Epqiu6;  // ../RTL/cortexm0ds_logic.v(660)
  wire Eprhu6;  // ../RTL/cortexm0ds_logic.v(192)
  wire Eprow6;  // ../RTL/cortexm0ds_logic.v(1217)
  wire Epxiu6;  // ../RTL/cortexm0ds_logic.v(754)
  wire Epyhu6;  // ../RTL/cortexm0ds_logic.v(286)
  wire Epyow6;  // ../RTL/cortexm0ds_logic.v(1310)
  wire Eq3ju6;  // ../RTL/cortexm0ds_logic.v(835)
  wire Eq4iu6;  // ../RTL/cortexm0ds_logic.v(367)
  wire Eq4pw6;  // ../RTL/cortexm0ds_logic.v(1391)
  wire Eqaju6;  // ../RTL/cortexm0ds_logic.v(928)
  wire Eqbiu6;  // ../RTL/cortexm0ds_logic.v(460)
  wire Eqbpw6;  // ../RTL/cortexm0ds_logic.v(1485)
  wire Eqcow6;  // ../RTL/cortexm0ds_logic.v(1017)
  wire Eqiiu6;  // ../RTL/cortexm0ds_logic.v(554)
  wire Eqjow6;  // ../RTL/cortexm0ds_logic.v(1110)
  wire Eqpiu6;  // ../RTL/cortexm0ds_logic.v(647)
  wire Eqqhu6;  // ../RTL/cortexm0ds_logic.v(179)
  wire Eqqow6;  // ../RTL/cortexm0ds_logic.v(1204)
  wire Eqtax6;  // ../RTL/cortexm0ds_logic.v(1668)
  wire Equpw6;  // ../RTL/cortexm0ds_logic.v(1607)
  wire Eqwiu6;  // ../RTL/cortexm0ds_logic.v(741)
  wire Eqxhu6;  // ../RTL/cortexm0ds_logic.v(273)
  wire Eqxow6;  // ../RTL/cortexm0ds_logic.v(1297)
  wire Er2ju6;  // ../RTL/cortexm0ds_logic.v(822)
  wire Er3iu6;  // ../RTL/cortexm0ds_logic.v(354)
  wire Er3pw6;  // ../RTL/cortexm0ds_logic.v(1378)
  wire Er9ju6;  // ../RTL/cortexm0ds_logic.v(915)
  wire Eraiu6;  // ../RTL/cortexm0ds_logic.v(447)
  wire Erapw6;  // ../RTL/cortexm0ds_logic.v(1472)
  wire Erbbx6;  // ../RTL/cortexm0ds_logic.v(1700)
  wire Erbow6;  // ../RTL/cortexm0ds_logic.v(1004)
  wire Erhiu6;  // ../RTL/cortexm0ds_logic.v(541)
  wire Eriow6;  // ../RTL/cortexm0ds_logic.v(1097)
  wire Eroiu6;  // ../RTL/cortexm0ds_logic.v(634)
  wire Erpax6;  // ../RTL/cortexm0ds_logic.v(1661)
  wire Erphu6;  // ../RTL/cortexm0ds_logic.v(166)
  wire Erpow6;  // ../RTL/cortexm0ds_logic.v(1191)
  wire Erviu6;  // ../RTL/cortexm0ds_logic.v(728)
  wire Erwhu6;  // ../RTL/cortexm0ds_logic.v(260)
  wire Erwow6;  // ../RTL/cortexm0ds_logic.v(1284)
  wire Es1ju6;  // ../RTL/cortexm0ds_logic.v(809)
  wire Es2iu6;  // ../RTL/cortexm0ds_logic.v(341)
  wire Es2pw6;  // ../RTL/cortexm0ds_logic.v(1365)
  wire Es8ju6;  // ../RTL/cortexm0ds_logic.v(902)
  wire Es9iu6;  // ../RTL/cortexm0ds_logic.v(434)
  wire Es9pw6;  // ../RTL/cortexm0ds_logic.v(1459)
  wire Esabx6;  // ../RTL/cortexm0ds_logic.v(1698)
  wire Esaow6;  // ../RTL/cortexm0ds_logic.v(991)
  wire Esgiu6;  // ../RTL/cortexm0ds_logic.v(528)
  wire Eshow6;  // ../RTL/cortexm0ds_logic.v(1084)
  wire Esniu6;  // ../RTL/cortexm0ds_logic.v(621)
  wire Esohu6;  // ../RTL/cortexm0ds_logic.v(153)
  wire Esoow6;  // ../RTL/cortexm0ds_logic.v(1178)
  wire Estax6;  // ../RTL/cortexm0ds_logic.v(1668)
  wire Esuiu6;  // ../RTL/cortexm0ds_logic.v(715)
  wire Esvhu6;  // ../RTL/cortexm0ds_logic.v(247)
  wire Esvow6;  // ../RTL/cortexm0ds_logic.v(1271)
  wire Et0ju6;  // ../RTL/cortexm0ds_logic.v(796)
  wire Et1iu6;  // ../RTL/cortexm0ds_logic.v(328)
  wire Et1pw6;  // ../RTL/cortexm0ds_logic.v(1352)
  wire Et7ju6;  // ../RTL/cortexm0ds_logic.v(889)
  wire Et8iu6;  // ../RTL/cortexm0ds_logic.v(421)
  wire Et8pw6;  // ../RTL/cortexm0ds_logic.v(1446)
  wire Et9ow6;  // ../RTL/cortexm0ds_logic.v(978)
  wire Etfbx6;  // ../RTL/cortexm0ds_logic.v(1708)
  wire Etfiu6;  // ../RTL/cortexm0ds_logic.v(515)
  wire Etgow6;  // ../RTL/cortexm0ds_logic.v(1071)
  wire Etmiu6;  // ../RTL/cortexm0ds_logic.v(608)
  wire Etnow6;  // ../RTL/cortexm0ds_logic.v(1165)
  wire Ettiu6;  // ../RTL/cortexm0ds_logic.v(702)
  wire Etuhu6;  // ../RTL/cortexm0ds_logic.v(234)
  wire Etuow6;  // ../RTL/cortexm0ds_logic.v(1258)
  wire Eu0iu6;  // ../RTL/cortexm0ds_logic.v(315)
  wire Eu0pw6;  // ../RTL/cortexm0ds_logic.v(1339)
  wire Eu6ju6;  // ../RTL/cortexm0ds_logic.v(876)
  wire Eu7iu6;  // ../RTL/cortexm0ds_logic.v(408)
  wire Eu7pw6;  // ../RTL/cortexm0ds_logic.v(1433)
  wire Eu8ow6;  // ../RTL/cortexm0ds_logic.v(965)
  wire Eudax6;  // ../RTL/cortexm0ds_logic.v(1639)
  wire Eueiu6;  // ../RTL/cortexm0ds_logic.v(502)
  wire Eufow6;  // ../RTL/cortexm0ds_logic.v(1058)
  wire Eukhu6;  // ../RTL/cortexm0ds_logic.v(137)
  wire Euliu6;  // ../RTL/cortexm0ds_logic.v(595)
  wire Eumow6;  // ../RTL/cortexm0ds_logic.v(1152)
  wire Eusiu6;  // ../RTL/cortexm0ds_logic.v(689)
  wire Eutax6;  // ../RTL/cortexm0ds_logic.v(1668)
  wire Euthu6;  // ../RTL/cortexm0ds_logic.v(221)
  wire Eutow6;  // ../RTL/cortexm0ds_logic.v(1245)
  wire Euziu6;  // ../RTL/cortexm0ds_logic.v(783)
  wire Ev5ju6;  // ../RTL/cortexm0ds_logic.v(863)
  wire Ev6iu6;  // ../RTL/cortexm0ds_logic.v(395)
  wire Ev6pw6;  // ../RTL/cortexm0ds_logic.v(1420)
  wire Ev7ow6;  // ../RTL/cortexm0ds_logic.v(952)
  wire Evbax6;  // ../RTL/cortexm0ds_logic.v(1635)
  wire Evdiu6;  // ../RTL/cortexm0ds_logic.v(489)
  wire Evdpw6;  // ../RTL/cortexm0ds_logic.v(1513)
  wire Eveow6;  // ../RTL/cortexm0ds_logic.v(1045)
  wire Evhpw6;  // ../RTL/cortexm0ds_logic.v(1584)
  wire Evkiu6;  // ../RTL/cortexm0ds_logic.v(582)
  wire Evlow6;  // ../RTL/cortexm0ds_logic.v(1139)
  wire Evriu6;  // ../RTL/cortexm0ds_logic.v(676)
  wire Evshu6;  // ../RTL/cortexm0ds_logic.v(208)
  wire Evsow6;  // ../RTL/cortexm0ds_logic.v(1232)
  wire Evyiu6;  // ../RTL/cortexm0ds_logic.v(770)
  wire Evypw6;  // ../RTL/cortexm0ds_logic.v(1615)
  wire Evzhu6;  // ../RTL/cortexm0ds_logic.v(302)
  wire Evzow6;  // ../RTL/cortexm0ds_logic.v(1326)
  wire Ew4ju6;  // ../RTL/cortexm0ds_logic.v(850)
  wire Ew5iu6;  // ../RTL/cortexm0ds_logic.v(382)
  wire Ew5pw6;  // ../RTL/cortexm0ds_logic.v(1407)
  wire Ew6ow6;  // ../RTL/cortexm0ds_logic.v(939)
  wire Ewciu6;  // ../RTL/cortexm0ds_logic.v(476)
  wire Ewcpw6;  // ../RTL/cortexm0ds_logic.v(1500)
  wire Ewdow6;  // ../RTL/cortexm0ds_logic.v(1032)
  wire Ewjhu6;  // ../RTL/cortexm0ds_logic.v(135)
  wire Ewjiu6;  // ../RTL/cortexm0ds_logic.v(569)
  wire Ewkow6;  // ../RTL/cortexm0ds_logic.v(1126)
  wire Ewqiu6;  // ../RTL/cortexm0ds_logic.v(663)
  wire Ewrhu6;  // ../RTL/cortexm0ds_logic.v(195)
  wire Ewrow6;  // ../RTL/cortexm0ds_logic.v(1219)
  wire Ewtax6;  // ../RTL/cortexm0ds_logic.v(1668)
  wire Ewxiu6;  // ../RTL/cortexm0ds_logic.v(757)
  wire Ewyhu6;  // ../RTL/cortexm0ds_logic.v(289)
  wire Ewyow6;  // ../RTL/cortexm0ds_logic.v(1313)
  wire Ex3ju6;  // ../RTL/cortexm0ds_logic.v(837)
  wire Ex4iu6;  // ../RTL/cortexm0ds_logic.v(369)
  wire Ex4pw6;  // ../RTL/cortexm0ds_logic.v(1394)
  wire Exbiu6;  // ../RTL/cortexm0ds_logic.v(463)
  wire Exbpw6;  // ../RTL/cortexm0ds_logic.v(1487)
  wire Excow6;  // ../RTL/cortexm0ds_logic.v(1019)
  wire Exehu6;  // ../RTL/cortexm0ds_logic.v(123)
  wire Exiiu6;  // ../RTL/cortexm0ds_logic.v(556)
  wire Exjow6;  // ../RTL/cortexm0ds_logic.v(1113)
  wire Expiu6;  // ../RTL/cortexm0ds_logic.v(650)
  wire Exqhu6;  // ../RTL/cortexm0ds_logic.v(182)
  wire Exqow6;  // ../RTL/cortexm0ds_logic.v(1206)
  wire Exwiu6;  // ../RTL/cortexm0ds_logic.v(744)
  wire Exxhu6;  // ../RTL/cortexm0ds_logic.v(276)
  wire Exxow6;  // ../RTL/cortexm0ds_logic.v(1300)
  wire Exypw6;  // ../RTL/cortexm0ds_logic.v(1615)
  wire Ey2ju6;  // ../RTL/cortexm0ds_logic.v(824)
  wire Ey3iu6;  // ../RTL/cortexm0ds_logic.v(356)
  wire Ey3pw6;  // ../RTL/cortexm0ds_logic.v(1381)
  wire Ey9ju6;  // ../RTL/cortexm0ds_logic.v(918)
  wire Eyaiu6;  // ../RTL/cortexm0ds_logic.v(450)
  wire Eyapw6;  // ../RTL/cortexm0ds_logic.v(1474)
  wire Eybow6;  // ../RTL/cortexm0ds_logic.v(1006)
  wire Eyhiu6;  // ../RTL/cortexm0ds_logic.v(543)
  wire Eyihu6;  // ../RTL/cortexm0ds_logic.v(132)
  wire Eyiow6;  // ../RTL/cortexm0ds_logic.v(1100)
  wire Eyoiu6;  // ../RTL/cortexm0ds_logic.v(637)
  wire Eyphu6;  // ../RTL/cortexm0ds_logic.v(169)
  wire Eypow6;  // ../RTL/cortexm0ds_logic.v(1193)
  wire Eytax6;  // ../RTL/cortexm0ds_logic.v(1668)
  wire Eyviu6;  // ../RTL/cortexm0ds_logic.v(731)
  wire Eywhu6;  // ../RTL/cortexm0ds_logic.v(263)
  wire Eywow6;  // ../RTL/cortexm0ds_logic.v(1287)
  wire Eyyax6;  // ../RTL/cortexm0ds_logic.v(1677)
  wire Ez1ju6;  // ../RTL/cortexm0ds_logic.v(811)
  wire Ez1qw6;  // ../RTL/cortexm0ds_logic.v(1621)
  wire Ez2iu6;  // ../RTL/cortexm0ds_logic.v(343)
  wire Ez2pw6;  // ../RTL/cortexm0ds_logic.v(1368)
  wire Ez8ju6;  // ../RTL/cortexm0ds_logic.v(905)
  wire Ez9iu6;  // ../RTL/cortexm0ds_logic.v(437)
  wire Ez9pw6;  // ../RTL/cortexm0ds_logic.v(1461)
  wire Ezaow6;  // ../RTL/cortexm0ds_logic.v(993)
  wire Ezgiu6;  // ../RTL/cortexm0ds_logic.v(530)
  wire Ezhow6;  // ../RTL/cortexm0ds_logic.v(1087)
  wire Ezniu6;  // ../RTL/cortexm0ds_logic.v(624)
  wire Ezohu6;  // ../RTL/cortexm0ds_logic.v(156)
  wire Ezoow6;  // ../RTL/cortexm0ds_logic.v(1180)
  wire Ezuiu6;  // ../RTL/cortexm0ds_logic.v(718)
  wire Ezvhu6;  // ../RTL/cortexm0ds_logic.v(250)
  wire Ezvow6;  // ../RTL/cortexm0ds_logic.v(1274)
  wire Ezypw6;  // ../RTL/cortexm0ds_logic.v(1615)
  wire F05ju6;  // ../RTL/cortexm0ds_logic.v(852)
  wire F06iu6;  // ../RTL/cortexm0ds_logic.v(384)
  wire F06pw6;  // ../RTL/cortexm0ds_logic.v(1408)
  wire F07ow6;  // ../RTL/cortexm0ds_logic.v(940)
  wire F0diu6;  // ../RTL/cortexm0ds_logic.v(477)
  wire F0dpw6;  // ../RTL/cortexm0ds_logic.v(1502)
  wire F0eow6;  // ../RTL/cortexm0ds_logic.v(1034)
  wire F0kiu6;  // ../RTL/cortexm0ds_logic.v(571)
  wire F0low6;  // ../RTL/cortexm0ds_logic.v(1127)
  wire F0riu6;  // ../RTL/cortexm0ds_logic.v(664)
  wire F0shu6;  // ../RTL/cortexm0ds_logic.v(196)
  wire F0sow6;  // ../RTL/cortexm0ds_logic.v(1221)
  wire F0yiu6;  // ../RTL/cortexm0ds_logic.v(758)
  wire F0zhu6;  // ../RTL/cortexm0ds_logic.v(290)
  wire F0zow6;  // ../RTL/cortexm0ds_logic.v(1314)
  wire F14ju6;  // ../RTL/cortexm0ds_logic.v(839)
  wire F15iu6;  // ../RTL/cortexm0ds_logic.v(371)
  wire F15pw6;  // ../RTL/cortexm0ds_logic.v(1395)
  wire F17ax6;  // ../RTL/cortexm0ds_logic.v(1626)
  wire F1ciu6;  // ../RTL/cortexm0ds_logic.v(464)
  wire F1cpw6;  // ../RTL/cortexm0ds_logic.v(1489)
  wire F1dow6;  // ../RTL/cortexm0ds_logic.v(1021)
  wire F1jiu6;  // ../RTL/cortexm0ds_logic.v(558)
  wire F1kow6;  // ../RTL/cortexm0ds_logic.v(1114)
  wire F1pax6;  // ../RTL/cortexm0ds_logic.v(1660)
  wire F1qiu6;  // ../RTL/cortexm0ds_logic.v(651)
  wire F1rhu6;  // ../RTL/cortexm0ds_logic.v(183)
  wire F1row6;  // ../RTL/cortexm0ds_logic.v(1208)
  wire F1xiu6;  // ../RTL/cortexm0ds_logic.v(745)
  wire F1yhu6;  // ../RTL/cortexm0ds_logic.v(277)
  wire F1yow6;  // ../RTL/cortexm0ds_logic.v(1301)
  wire F23ju6;  // ../RTL/cortexm0ds_logic.v(826)
  wire F24iu6;  // ../RTL/cortexm0ds_logic.v(358)
  wire F24pw6;  // ../RTL/cortexm0ds_logic.v(1382)
  wire F26bx6;  // ../RTL/cortexm0ds_logic.v(1690)
  wire F2aju6;  // ../RTL/cortexm0ds_logic.v(919)
  wire F2biu6;  // ../RTL/cortexm0ds_logic.v(451)
  wire F2bpw6;  // ../RTL/cortexm0ds_logic.v(1476)
  wire F2cow6;  // ../RTL/cortexm0ds_logic.v(1008)
  wire F2dax6;  // ../RTL/cortexm0ds_logic.v(1637)
  wire F2iiu6;  // ../RTL/cortexm0ds_logic.v(545)
  wire F2jow6;  // ../RTL/cortexm0ds_logic.v(1101)
  wire F2piu6;  // ../RTL/cortexm0ds_logic.v(638)
  wire F2qhu6;  // ../RTL/cortexm0ds_logic.v(170)
  wire F2qow6;  // ../RTL/cortexm0ds_logic.v(1195)
  wire F2tax6;  // ../RTL/cortexm0ds_logic.v(1667)
  wire F2wiu6;  // ../RTL/cortexm0ds_logic.v(732)
  wire F2xhu6;  // ../RTL/cortexm0ds_logic.v(264)
  wire F2xow6;  // ../RTL/cortexm0ds_logic.v(1288)
  wire F32ju6;  // ../RTL/cortexm0ds_logic.v(813)
  wire F33iu6;  // ../RTL/cortexm0ds_logic.v(345)
  wire F33pw6;  // ../RTL/cortexm0ds_logic.v(1369)
  wire F39ju6;  // ../RTL/cortexm0ds_logic.v(906)
  wire F3aiu6;  // ../RTL/cortexm0ds_logic.v(438)
  wire F3apw6;  // ../RTL/cortexm0ds_logic.v(1463)
  wire F3bow6;  // ../RTL/cortexm0ds_logic.v(995)
  wire F3hiu6;  // ../RTL/cortexm0ds_logic.v(532)
  wire F3iow6;  // ../RTL/cortexm0ds_logic.v(1088)
  wire F3oiu6;  // ../RTL/cortexm0ds_logic.v(625)
  wire F3pax6;  // ../RTL/cortexm0ds_logic.v(1660)
  wire F3phu6;  // ../RTL/cortexm0ds_logic.v(157)
  wire F3pow6;  // ../RTL/cortexm0ds_logic.v(1182)
  wire F3viu6;  // ../RTL/cortexm0ds_logic.v(719)
  wire F3whu6;  // ../RTL/cortexm0ds_logic.v(251)
  wire F3wow6;  // ../RTL/cortexm0ds_logic.v(1275)
  wire F41ju6;  // ../RTL/cortexm0ds_logic.v(800)
  wire F42iu6;  // ../RTL/cortexm0ds_logic.v(332)
  wire F42pw6;  // ../RTL/cortexm0ds_logic.v(1356)
  wire F48ju6;  // ../RTL/cortexm0ds_logic.v(893)
  wire F49iu6;  // ../RTL/cortexm0ds_logic.v(425)
  wire F49pw6;  // ../RTL/cortexm0ds_logic.v(1450)
  wire F4aow6;  // ../RTL/cortexm0ds_logic.v(982)
  wire F4giu6;  // ../RTL/cortexm0ds_logic.v(519)
  wire F4how6;  // ../RTL/cortexm0ds_logic.v(1075)
  wire F4iax6;  // ../RTL/cortexm0ds_logic.v(1647)
  wire F4ibx6;  // ../RTL/cortexm0ds_logic.v(1712)
  wire F4niu6;  // ../RTL/cortexm0ds_logic.v(612)
  wire F4oow6;  // ../RTL/cortexm0ds_logic.v(1169)
  wire F4tax6;  // ../RTL/cortexm0ds_logic.v(1667)
  wire F4uiu6;  // ../RTL/cortexm0ds_logic.v(706)
  wire F4vhu6;  // ../RTL/cortexm0ds_logic.v(238)
  wire F4vow6;  // ../RTL/cortexm0ds_logic.v(1262)
  wire F50ju6;  // ../RTL/cortexm0ds_logic.v(787)
  wire F51iu6;  // ../RTL/cortexm0ds_logic.v(319)
  wire F51pw6;  // ../RTL/cortexm0ds_logic.v(1343)
  wire F57ju6;  // ../RTL/cortexm0ds_logic.v(880)
  wire F58iu6;  // ../RTL/cortexm0ds_logic.v(412)
  wire F58pw6;  // ../RTL/cortexm0ds_logic.v(1437)
  wire F59bx6;  // ../RTL/cortexm0ds_logic.v(1695)
  wire F59ow6;  // ../RTL/cortexm0ds_logic.v(969)
  wire F5fiu6;  // ../RTL/cortexm0ds_logic.v(506)
  wire F5gow6;  // ../RTL/cortexm0ds_logic.v(1062)
  wire F5miu6;  // ../RTL/cortexm0ds_logic.v(599)
  wire F5now6;  // ../RTL/cortexm0ds_logic.v(1156)
  wire F5tiu6;  // ../RTL/cortexm0ds_logic.v(693)
  wire F5uhu6;  // ../RTL/cortexm0ds_logic.v(225)
  wire F5uow6;  // ../RTL/cortexm0ds_logic.v(1249)
  wire F60iu6;  // ../RTL/cortexm0ds_logic.v(306)
  wire F60pw6;  // ../RTL/cortexm0ds_logic.v(1330)
  wire F66ju6;  // ../RTL/cortexm0ds_logic.v(867)
  wire F67iu6;  // ../RTL/cortexm0ds_logic.v(399)
  wire F67pw6;  // ../RTL/cortexm0ds_logic.v(1424)
  wire F68ow6;  // ../RTL/cortexm0ds_logic.v(956)
  wire F6dbx6;  // ../RTL/cortexm0ds_logic.v(1703)
  wire F6eiu6;  // ../RTL/cortexm0ds_logic.v(493)
  wire F6fow6;  // ../RTL/cortexm0ds_logic.v(1049)
  wire F6liu6;  // ../RTL/cortexm0ds_logic.v(586)
  wire F6mow6;  // ../RTL/cortexm0ds_logic.v(1143)
  wire F6siu6;  // ../RTL/cortexm0ds_logic.v(680)
  wire F6tax6;  // ../RTL/cortexm0ds_logic.v(1667)
  wire F6thu6;  // ../RTL/cortexm0ds_logic.v(212)
  wire F6tow6;  // ../RTL/cortexm0ds_logic.v(1236)
  wire F6ziu6;  // ../RTL/cortexm0ds_logic.v(774)
  wire F75ju6;  // ../RTL/cortexm0ds_logic.v(854)
  wire F76iu6;  // ../RTL/cortexm0ds_logic.v(386)
  wire F76pw6;  // ../RTL/cortexm0ds_logic.v(1411)
  wire F77ow6;  // ../RTL/cortexm0ds_logic.v(943)
  wire F7diu6;  // ../RTL/cortexm0ds_logic.v(480)
  wire F7dpw6;  // ../RTL/cortexm0ds_logic.v(1504)
  wire F7eax6;  // ../RTL/cortexm0ds_logic.v(1639)
  wire F7eow6;  // ../RTL/cortexm0ds_logic.v(1036)
  wire F7jbx6;  // ../RTL/cortexm0ds_logic.v(1714)
  wire F7kiu6;  // ../RTL/cortexm0ds_logic.v(573)
  wire F7low6;  // ../RTL/cortexm0ds_logic.v(1130)
  wire F7riu6;  // ../RTL/cortexm0ds_logic.v(667)
  wire F7shu6;  // ../RTL/cortexm0ds_logic.v(199)
  wire F7sow6;  // ../RTL/cortexm0ds_logic.v(1223)
  wire F7yiu6;  // ../RTL/cortexm0ds_logic.v(761)
  wire F7zhu6;  // ../RTL/cortexm0ds_logic.v(293)
  wire F7zow6;  // ../RTL/cortexm0ds_logic.v(1317)
  wire F84ju6;  // ../RTL/cortexm0ds_logic.v(841)
  wire F85iu6;  // ../RTL/cortexm0ds_logic.v(373)
  wire F85pw6;  // ../RTL/cortexm0ds_logic.v(1398)
  wire F86ow6;  // ../RTL/cortexm0ds_logic.v(930)
  wire F8cbx6;  // ../RTL/cortexm0ds_logic.v(1701)
  wire F8ciu6;  // ../RTL/cortexm0ds_logic.v(467)
  wire F8cpw6;  // ../RTL/cortexm0ds_logic.v(1491)
  wire F8dbx6;  // ../RTL/cortexm0ds_logic.v(1703)
  wire F8dow6;  // ../RTL/cortexm0ds_logic.v(1023)
  wire F8jiu6;  // ../RTL/cortexm0ds_logic.v(560)
  wire F8kow6;  // ../RTL/cortexm0ds_logic.v(1117)
  wire F8qiu6;  // ../RTL/cortexm0ds_logic.v(654)
  wire F8rhu6;  // ../RTL/cortexm0ds_logic.v(186)
  wire F8row6;  // ../RTL/cortexm0ds_logic.v(1210)
  wire F8tax6;  // ../RTL/cortexm0ds_logic.v(1667)
  wire F8xiu6;  // ../RTL/cortexm0ds_logic.v(748)
  wire F8yhu6;  // ../RTL/cortexm0ds_logic.v(280)
  wire F8yow6;  // ../RTL/cortexm0ds_logic.v(1304)
  wire F93ju6;  // ../RTL/cortexm0ds_logic.v(828)
  wire F94iu6;  // ../RTL/cortexm0ds_logic.v(360)
  wire F94pw6;  // ../RTL/cortexm0ds_logic.v(1385)
  wire F9aju6;  // ../RTL/cortexm0ds_logic.v(922)
  wire F9biu6;  // ../RTL/cortexm0ds_logic.v(454)
  wire F9bpw6;  // ../RTL/cortexm0ds_logic.v(1478)
  wire F9cow6;  // ../RTL/cortexm0ds_logic.v(1010)
  wire F9gbx6;  // ../RTL/cortexm0ds_logic.v(1709)
  wire F9iiu6;  // ../RTL/cortexm0ds_logic.v(547)
  wire F9jow6;  // ../RTL/cortexm0ds_logic.v(1104)
  wire F9piu6;  // ../RTL/cortexm0ds_logic.v(641)
  wire F9qhu6;  // ../RTL/cortexm0ds_logic.v(173)
  wire F9qow6;  // ../RTL/cortexm0ds_logic.v(1197)
  wire F9vpw6;  // ../RTL/cortexm0ds_logic.v(1608)
  wire F9wiu6;  // ../RTL/cortexm0ds_logic.v(735)
  wire F9xhu6;  // ../RTL/cortexm0ds_logic.v(267)
  wire F9xow6;  // ../RTL/cortexm0ds_logic.v(1291)
  wire Fa2ju6;  // ../RTL/cortexm0ds_logic.v(815)
  wire Fa3iu6;  // ../RTL/cortexm0ds_logic.v(347)
  wire Fa3pw6;  // ../RTL/cortexm0ds_logic.v(1372)
  wire Fa9ju6;  // ../RTL/cortexm0ds_logic.v(909)
  wire Faaiu6;  // ../RTL/cortexm0ds_logic.v(441)
  wire Faapw6;  // ../RTL/cortexm0ds_logic.v(1465)
  wire Fabow6;  // ../RTL/cortexm0ds_logic.v(997)
  wire Facax6;  // ../RTL/cortexm0ds_logic.v(1636)
  wire Facbx6;  // ../RTL/cortexm0ds_logic.v(1701)
  wire Fahax6;  // ../RTL/cortexm0ds_logic.v(1645)
  wire Fahiu6;  // ../RTL/cortexm0ds_logic.v(534)
  wire Faiow6;  // ../RTL/cortexm0ds_logic.v(1091)
  wire Fanhu6;  // ../RTL/cortexm0ds_logic.v(144)
  wire Faoiu6;  // ../RTL/cortexm0ds_logic.v(628)
  wire Faphu6;  // ../RTL/cortexm0ds_logic.v(160)
  wire Fapow6;  // ../RTL/cortexm0ds_logic.v(1184)
  wire Fatax6;  // ../RTL/cortexm0ds_logic.v(1667)
  wire Faviu6;  // ../RTL/cortexm0ds_logic.v(722)
  wire Fawhu6;  // ../RTL/cortexm0ds_logic.v(254)
  wire Fawow6;  // ../RTL/cortexm0ds_logic.v(1278)
  wire Fb0bx6;  // ../RTL/cortexm0ds_logic.v(1680)
  wire Fb1ju6;  // ../RTL/cortexm0ds_logic.v(802)
  wire Fb2iu6;  // ../RTL/cortexm0ds_logic.v(334)
  wire Fb2pw6;  // ../RTL/cortexm0ds_logic.v(1359)
  wire Fb8ju6;  // ../RTL/cortexm0ds_logic.v(896)
  wire Fb9iu6;  // ../RTL/cortexm0ds_logic.v(428)
  wire Fb9pw6;  // ../RTL/cortexm0ds_logic.v(1452)
  wire Fbaow6;  // ../RTL/cortexm0ds_logic.v(984)
  wire Fbgiu6;  // ../RTL/cortexm0ds_logic.v(521)
  wire Fbhow6;  // ../RTL/cortexm0ds_logic.v(1078)
  wire Fbniu6;  // ../RTL/cortexm0ds_logic.v(615)
  wire Fbohu6;  // ../RTL/cortexm0ds_logic.v(147)
  wire Fboow6;  // ../RTL/cortexm0ds_logic.v(1171)
  wire Fbuiu6;  // ../RTL/cortexm0ds_logic.v(709)
  wire Fbvhu6;  // ../RTL/cortexm0ds_logic.v(241)
  wire Fbvow6;  // ../RTL/cortexm0ds_logic.v(1265)
  wire Fc0ju6;  // ../RTL/cortexm0ds_logic.v(789)
  wire Fc1bx6;  // ../RTL/cortexm0ds_logic.v(1682)
  wire Fc1iu6;  // ../RTL/cortexm0ds_logic.v(321)
  wire Fc1pw6;  // ../RTL/cortexm0ds_logic.v(1346)
  wire Fc7ju6;  // ../RTL/cortexm0ds_logic.v(883)
  wire Fc8iu6;  // ../RTL/cortexm0ds_logic.v(415)
  wire Fc8pw6;  // ../RTL/cortexm0ds_logic.v(1439)
  wire Fc9ow6;  // ../RTL/cortexm0ds_logic.v(971)
  wire Fcfiu6;  // ../RTL/cortexm0ds_logic.v(508)
  wire Fcgow6;  // ../RTL/cortexm0ds_logic.v(1065)
  wire Fcmiu6;  // ../RTL/cortexm0ds_logic.v(602)
  wire Fcnow6;  // ../RTL/cortexm0ds_logic.v(1158)
  wire Fctiu6;  // ../RTL/cortexm0ds_logic.v(696)
  wire Fcuhu6;  // ../RTL/cortexm0ds_logic.v(228)
  wire Fcuow6;  // ../RTL/cortexm0ds_logic.v(1252)
  wire Fd0iu6;  // ../RTL/cortexm0ds_logic.v(308)
  wire Fd0pw6;  // ../RTL/cortexm0ds_logic.v(1333)
  wire Fd6ju6;  // ../RTL/cortexm0ds_logic.v(870)
  wire Fd7iu6;  // ../RTL/cortexm0ds_logic.v(402)
  wire Fd7pw6;  // ../RTL/cortexm0ds_logic.v(1426)
  wire Fd8ow6;  // ../RTL/cortexm0ds_logic.v(958)
  wire Fdeiu6;  // ../RTL/cortexm0ds_logic.v(495)
  wire Fdfow6;  // ../RTL/cortexm0ds_logic.v(1052)
  wire Fdliu6;  // ../RTL/cortexm0ds_logic.v(589)
  wire Fdmow6;  // ../RTL/cortexm0ds_logic.v(1145)
  wire Fdsiu6;  // ../RTL/cortexm0ds_logic.v(683)
  wire Fdthu6;  // ../RTL/cortexm0ds_logic.v(215)
  wire Fdtow6;  // ../RTL/cortexm0ds_logic.v(1239)
  wire Fdziu6;  // ../RTL/cortexm0ds_logic.v(776)
  wire Fe2bx6;  // ../RTL/cortexm0ds_logic.v(1683)
  wire Fe5ju6;  // ../RTL/cortexm0ds_logic.v(857)
  wire Fe6iu6;  // ../RTL/cortexm0ds_logic.v(389)
  wire Fe6pw6;  // ../RTL/cortexm0ds_logic.v(1413)
  wire Fe7ow6;  // ../RTL/cortexm0ds_logic.v(945)
  wire Fediu6;  // ../RTL/cortexm0ds_logic.v(482)
  wire Fedpw6;  // ../RTL/cortexm0ds_logic.v(1507)
  wire Feeow6;  // ../RTL/cortexm0ds_logic.v(1039)
  wire Fekiu6;  // ../RTL/cortexm0ds_logic.v(576)
  wire Felow6;  // ../RTL/cortexm0ds_logic.v(1132)
  wire Feriu6;  // ../RTL/cortexm0ds_logic.v(670)
  wire Feshu6;  // ../RTL/cortexm0ds_logic.v(202)
  wire Fesow6;  // ../RTL/cortexm0ds_logic.v(1226)
  wire Feyiu6;  // ../RTL/cortexm0ds_logic.v(763)
  wire Fezhu6;  // ../RTL/cortexm0ds_logic.v(295)
  wire Fezow6;  // ../RTL/cortexm0ds_logic.v(1320)
  wire Ff4ju6;  // ../RTL/cortexm0ds_logic.v(844)
  wire Ff5iu6;  // ../RTL/cortexm0ds_logic.v(376)
  wire Ff5pw6;  // ../RTL/cortexm0ds_logic.v(1400)
  wire Ff6ow6;  // ../RTL/cortexm0ds_logic.v(932)
  wire Ffciu6;  // ../RTL/cortexm0ds_logic.v(469)
  wire Ffcpw6;  // ../RTL/cortexm0ds_logic.v(1494)
  wire Ffdow6;  // ../RTL/cortexm0ds_logic.v(1026)
  wire Ffjiu6;  // ../RTL/cortexm0ds_logic.v(563)
  wire Ffkow6;  // ../RTL/cortexm0ds_logic.v(1119)
  wire Ffqiu6;  // ../RTL/cortexm0ds_logic.v(657)
  wire Ffrhu6;  // ../RTL/cortexm0ds_logic.v(189)
  wire Ffrow6;  // ../RTL/cortexm0ds_logic.v(1213)
  wire Ffxiu6;  // ../RTL/cortexm0ds_logic.v(750)
  wire Ffyhu6;  // ../RTL/cortexm0ds_logic.v(282)
  wire Ffyow6;  // ../RTL/cortexm0ds_logic.v(1307)
  wire Fg3ju6;  // ../RTL/cortexm0ds_logic.v(831)
  wire Fg4iu6;  // ../RTL/cortexm0ds_logic.v(363)
  wire Fg4pw6;  // ../RTL/cortexm0ds_logic.v(1387)
  wire Fgaju6;  // ../RTL/cortexm0ds_logic.v(924)
  wire Fgbiu6;  // ../RTL/cortexm0ds_logic.v(456)
  wire Fgbpw6;  // ../RTL/cortexm0ds_logic.v(1481)
  wire Fgcow6;  // ../RTL/cortexm0ds_logic.v(1013)
  wire Fgiiu6;  // ../RTL/cortexm0ds_logic.v(550)
  wire Fgjow6;  // ../RTL/cortexm0ds_logic.v(1106)
  wire Fgpiu6;  // ../RTL/cortexm0ds_logic.v(644)
  wire Fgqhu6;  // ../RTL/cortexm0ds_logic.v(176)
  wire Fgqow6;  // ../RTL/cortexm0ds_logic.v(1200)
  wire Fgwiu6;  // ../RTL/cortexm0ds_logic.v(737)
  wire Fgxhu6;  // ../RTL/cortexm0ds_logic.v(269)
  wire Fgxow6;  // ../RTL/cortexm0ds_logic.v(1294)
  wire Fh2ju6;  // ../RTL/cortexm0ds_logic.v(818)
  wire Fh3iu6;  // ../RTL/cortexm0ds_logic.v(350)
  wire Fh3pw6;  // ../RTL/cortexm0ds_logic.v(1374)
  wire Fh9ju6;  // ../RTL/cortexm0ds_logic.v(911)
  wire Fhaiu6;  // ../RTL/cortexm0ds_logic.v(443)
  wire Fhapw6;  // ../RTL/cortexm0ds_logic.v(1468)
  wire Fhbow6;  // ../RTL/cortexm0ds_logic.v(1000)
  wire Fhhiu6;  // ../RTL/cortexm0ds_logic.v(537)
  wire Fhiow6;  // ../RTL/cortexm0ds_logic.v(1093)
  wire Fhoiu6;  // ../RTL/cortexm0ds_logic.v(631)
  wire Fhphu6;  // ../RTL/cortexm0ds_logic.v(163)
  wire Fhpow6;  // ../RTL/cortexm0ds_logic.v(1187)
  wire Fhviu6;  // ../RTL/cortexm0ds_logic.v(724)
  wire Fhwhu6;  // ../RTL/cortexm0ds_logic.v(256)
  wire Fhwow6;  // ../RTL/cortexm0ds_logic.v(1281)
  wire Fi1ju6;  // ../RTL/cortexm0ds_logic.v(805)
  wire Fi2iu6;  // ../RTL/cortexm0ds_logic.v(337)
  wire Fi2pw6;  // ../RTL/cortexm0ds_logic.v(1361)
  wire Fi8ju6;  // ../RTL/cortexm0ds_logic.v(898)
  wire Fi9iu6;  // ../RTL/cortexm0ds_logic.v(430)
  wire Fi9pw6;  // ../RTL/cortexm0ds_logic.v(1455)
  wire Fiaow6;  // ../RTL/cortexm0ds_logic.v(987)
  wire Figiu6;  // ../RTL/cortexm0ds_logic.v(524)
  wire Fihow6;  // ../RTL/cortexm0ds_logic.v(1080)
  wire Finiu6;  // ../RTL/cortexm0ds_logic.v(618)
  wire Fiohu6;  // ../RTL/cortexm0ds_logic.v(150)
  wire Fioow6;  // ../RTL/cortexm0ds_logic.v(1174)
  wire Fiuiu6;  // ../RTL/cortexm0ds_logic.v(711)
  wire Fivhu6;  // ../RTL/cortexm0ds_logic.v(243)
  wire Fivow6;  // ../RTL/cortexm0ds_logic.v(1268)
  wire Fj0ju6;  // ../RTL/cortexm0ds_logic.v(792)
  wire Fj1iu6;  // ../RTL/cortexm0ds_logic.v(324)
  wire Fj1pw6;  // ../RTL/cortexm0ds_logic.v(1348)
  wire Fj7ju6;  // ../RTL/cortexm0ds_logic.v(885)
  wire Fj8ax6;  // ../RTL/cortexm0ds_logic.v(1628)
  wire Fj8iu6;  // ../RTL/cortexm0ds_logic.v(417)
  wire Fj8pw6;  // ../RTL/cortexm0ds_logic.v(1442)
  wire Fj9ow6;  // ../RTL/cortexm0ds_logic.v(974)
  wire Fjdbx6;  // ../RTL/cortexm0ds_logic.v(1704)
  wire Fjfiu6;  // ../RTL/cortexm0ds_logic.v(511)
  wire Fjgow6;  // ../RTL/cortexm0ds_logic.v(1067)
  wire Fjmiu6;  // ../RTL/cortexm0ds_logic.v(605)
  wire Fjnow6;  // ../RTL/cortexm0ds_logic.v(1161)
  wire Fjtiu6;  // ../RTL/cortexm0ds_logic.v(698)
  wire Fjuhu6;  // ../RTL/cortexm0ds_logic.v(230)
  wire Fjuow6;  // ../RTL/cortexm0ds_logic.v(1255)
  wire Fk0iu6;  // ../RTL/cortexm0ds_logic.v(311)
  wire Fk0pw6;  // ../RTL/cortexm0ds_logic.v(1335)
  wire Fk6ju6;  // ../RTL/cortexm0ds_logic.v(872)
  wire Fk7iu6;  // ../RTL/cortexm0ds_logic.v(404)
  wire Fk7pw6;  // ../RTL/cortexm0ds_logic.v(1429)
  wire Fk8ow6;  // ../RTL/cortexm0ds_logic.v(961)
  wire Fkeiu6;  // ../RTL/cortexm0ds_logic.v(498)
  wire Fkfow6;  // ../RTL/cortexm0ds_logic.v(1054)
  wire Fkliu6;  // ../RTL/cortexm0ds_logic.v(592)
  wire Fkmow6;  // ../RTL/cortexm0ds_logic.v(1148)
  wire Fkrpw6;  // ../RTL/cortexm0ds_logic.v(1602)
  wire Fksiu6;  // ../RTL/cortexm0ds_logic.v(685)
  wire Fkthu6;  // ../RTL/cortexm0ds_logic.v(217)
  wire Fktow6;  // ../RTL/cortexm0ds_logic.v(1242)
  wire Fkziu6;  // ../RTL/cortexm0ds_logic.v(779)
  wire Fl2qw6;  // ../RTL/cortexm0ds_logic.v(1622)
  wire Fl5ju6;  // ../RTL/cortexm0ds_logic.v(859)
  wire Fl6iu6;  // ../RTL/cortexm0ds_logic.v(391)
  wire Fl6pw6;  // ../RTL/cortexm0ds_logic.v(1416)
  wire Fl7ow6;  // ../RTL/cortexm0ds_logic.v(948)
  wire Fldbx6;  // ../RTL/cortexm0ds_logic.v(1704)
  wire Fldiu6;  // ../RTL/cortexm0ds_logic.v(485)
  wire Fldpw6;  // ../RTL/cortexm0ds_logic.v(1509)
  wire Fleow6;  // ../RTL/cortexm0ds_logic.v(1041)
  wire Flkiu6;  // ../RTL/cortexm0ds_logic.v(579)
  wire Fllow6;  // ../RTL/cortexm0ds_logic.v(1135)
  wire Flriu6;  // ../RTL/cortexm0ds_logic.v(672)
  wire Flshu6;  // ../RTL/cortexm0ds_logic.v(204)
  wire Flsow6;  // ../RTL/cortexm0ds_logic.v(1229)
  wire Flyiu6;  // ../RTL/cortexm0ds_logic.v(766)
  wire Flzhu6;  // ../RTL/cortexm0ds_logic.v(298)
  wire Flzow6;  // ../RTL/cortexm0ds_logic.v(1322)
  wire Fm4ju6;  // ../RTL/cortexm0ds_logic.v(846)
  wire Fm5iu6;  // ../RTL/cortexm0ds_logic.v(378)
  wire Fm5pw6;  // ../RTL/cortexm0ds_logic.v(1403)
  wire Fm6ow6;  // ../RTL/cortexm0ds_logic.v(935)
  wire Fm7ax6;  // ../RTL/cortexm0ds_logic.v(1627)
  wire Fmciu6;  // ../RTL/cortexm0ds_logic.v(472)
  wire Fmcpw6;  // ../RTL/cortexm0ds_logic.v(1496)
  wire Fmdhu6;  // ../RTL/cortexm0ds_logic.v(120)
  wire Fmdow6;  // ../RTL/cortexm0ds_logic.v(1028)
  wire Fmjiu6;  // ../RTL/cortexm0ds_logic.v(566)
  wire Fmkow6;  // ../RTL/cortexm0ds_logic.v(1122)
  wire Fmqiu6;  // ../RTL/cortexm0ds_logic.v(659)
  wire Fmrhu6;  // ../RTL/cortexm0ds_logic.v(191)
  wire Fmrow6;  // ../RTL/cortexm0ds_logic.v(1216)
  wire Fmxiu6;  // ../RTL/cortexm0ds_logic.v(753)
  wire Fmyhu6;  // ../RTL/cortexm0ds_logic.v(285)
  wire Fmyow6;  // ../RTL/cortexm0ds_logic.v(1309)
  wire Fn3ju6;  // ../RTL/cortexm0ds_logic.v(833)
  wire Fn4iu6;  // ../RTL/cortexm0ds_logic.v(365)
  wire Fn4pw6;  // ../RTL/cortexm0ds_logic.v(1390)
  wire Fnaju6;  // ../RTL/cortexm0ds_logic.v(927)
  wire Fnbiu6;  // ../RTL/cortexm0ds_logic.v(459)
  wire Fnbpw6;  // ../RTL/cortexm0ds_logic.v(1483)
  wire Fncow6;  // ../RTL/cortexm0ds_logic.v(1015)
  wire Fniiu6;  // ../RTL/cortexm0ds_logic.v(553)
  wire Fnjow6;  // ../RTL/cortexm0ds_logic.v(1109)
  wire Fnnhu6;  // ../RTL/cortexm0ds_logic.v(145)
  wire Fnnpw6;  // ../RTL/cortexm0ds_logic.v(1594)
  wire Fnpiu6;  // ../RTL/cortexm0ds_logic.v(646)
  wire Fnqhu6;  // ../RTL/cortexm0ds_logic.v(178)
  wire Fnqow6;  // ../RTL/cortexm0ds_logic.v(1203)
  wire Fnwiu6;  // ../RTL/cortexm0ds_logic.v(740)
  wire Fnxhu6;  // ../RTL/cortexm0ds_logic.v(272)
  wire Fnxow6;  // ../RTL/cortexm0ds_logic.v(1296)
  wire Fo2ju6;  // ../RTL/cortexm0ds_logic.v(820)
  wire Fo3iu6;  // ../RTL/cortexm0ds_logic.v(352)
  wire Fo3pw6;  // ../RTL/cortexm0ds_logic.v(1377)
  wire Fo9ax6;  // ../RTL/cortexm0ds_logic.v(1631)
  wire Fo9ju6;  // ../RTL/cortexm0ds_logic.v(914)
  wire Foaiu6;  // ../RTL/cortexm0ds_logic.v(446)
  wire Foapw6;  // ../RTL/cortexm0ds_logic.v(1470)
  wire Fobow6;  // ../RTL/cortexm0ds_logic.v(1002)
  wire Fohiu6;  // ../RTL/cortexm0ds_logic.v(540)
  wire Foiow6;  // ../RTL/cortexm0ds_logic.v(1096)
  wire Fooiu6;  // ../RTL/cortexm0ds_logic.v(633)
  wire Fophu6;  // ../RTL/cortexm0ds_logic.v(165)
  wire Fopow6;  // ../RTL/cortexm0ds_logic.v(1190)
  wire Foviu6;  // ../RTL/cortexm0ds_logic.v(727)
  wire Fowhu6;  // ../RTL/cortexm0ds_logic.v(259)
  wire Fowow6;  // ../RTL/cortexm0ds_logic.v(1283)
  wire Fp1ju6;  // ../RTL/cortexm0ds_logic.v(807)
  wire Fp2iu6;  // ../RTL/cortexm0ds_logic.v(339)
  wire Fp2pw6;  // ../RTL/cortexm0ds_logic.v(1364)
  wire Fp8ju6;  // ../RTL/cortexm0ds_logic.v(901)
  wire Fp9iu6;  // ../RTL/cortexm0ds_logic.v(433)
  wire Fp9pw6;  // ../RTL/cortexm0ds_logic.v(1457)
  wire Fpaow6;  // ../RTL/cortexm0ds_logic.v(989)
  wire Fpgiu6;  // ../RTL/cortexm0ds_logic.v(527)
  wire Fphow6;  // ../RTL/cortexm0ds_logic.v(1083)
  wire Fpniu6;  // ../RTL/cortexm0ds_logic.v(620)
  wire Fpnpw6;  // ../RTL/cortexm0ds_logic.v(1595)
  wire Fpohu6;  // ../RTL/cortexm0ds_logic.v(152)
  wire Fpoow6;  // ../RTL/cortexm0ds_logic.v(1177)
  wire Fpuiu6;  // ../RTL/cortexm0ds_logic.v(714)
  wire Fpvhu6;  // ../RTL/cortexm0ds_logic.v(246)
  wire Fpvow6;  // ../RTL/cortexm0ds_logic.v(1270)
  wire Fq0ju6;  // ../RTL/cortexm0ds_logic.v(794)
  wire Fq1iu6;  // ../RTL/cortexm0ds_logic.v(326)
  wire Fq1pw6;  // ../RTL/cortexm0ds_logic.v(1351)
  wire Fq7ju6;  // ../RTL/cortexm0ds_logic.v(888)
  wire Fq8iu6;  // ../RTL/cortexm0ds_logic.v(420)
  wire Fq8pw6;  // ../RTL/cortexm0ds_logic.v(1444)
  wire Fq9ow6;  // ../RTL/cortexm0ds_logic.v(976)
  wire Fqfiu6;  // ../RTL/cortexm0ds_logic.v(514)
  wire Fqgow6;  // ../RTL/cortexm0ds_logic.v(1070)
  wire Fqmiu6;  // ../RTL/cortexm0ds_logic.v(607)
  wire Fqnow6;  // ../RTL/cortexm0ds_logic.v(1164)
  wire Fqtiu6;  // ../RTL/cortexm0ds_logic.v(701)
  wire Fquhu6;  // ../RTL/cortexm0ds_logic.v(233)
  wire Fquow6;  // ../RTL/cortexm0ds_logic.v(1257)
  wire Fr0iu6;  // ../RTL/cortexm0ds_logic.v(313)
  wire Fr0pw6;  // ../RTL/cortexm0ds_logic.v(1338)
  wire Fr6ju6;  // ../RTL/cortexm0ds_logic.v(875)
  wire Fr7iu6;  // ../RTL/cortexm0ds_logic.v(407)
  wire Fr7pw6;  // ../RTL/cortexm0ds_logic.v(1431)
  wire Fr8ow6;  // ../RTL/cortexm0ds_logic.v(963)
  wire Freiu6;  // ../RTL/cortexm0ds_logic.v(501)
  wire Frfow6;  // ../RTL/cortexm0ds_logic.v(1057)
  wire Frliu6;  // ../RTL/cortexm0ds_logic.v(594)
  wire Frmhu6;  // ../RTL/cortexm0ds_logic.v(143)
  wire Frmow6;  // ../RTL/cortexm0ds_logic.v(1151)
  wire Frsiu6;  // ../RTL/cortexm0ds_logic.v(688)
  wire Frthu6;  // ../RTL/cortexm0ds_logic.v(220)
  wire Frtow6;  // ../RTL/cortexm0ds_logic.v(1244)
  wire Frziu6;  // ../RTL/cortexm0ds_logic.v(781)
  wire Fs5ju6;  // ../RTL/cortexm0ds_logic.v(862)
  wire Fs6iu6;  // ../RTL/cortexm0ds_logic.v(394)
  wire Fs6pw6;  // ../RTL/cortexm0ds_logic.v(1418)
  wire Fs7ow6;  // ../RTL/cortexm0ds_logic.v(950)
  wire Fsdhu6;  // ../RTL/cortexm0ds_logic.v(120)
  wire Fsdiu6;  // ../RTL/cortexm0ds_logic.v(488)
  wire Fsdpw6;  // ../RTL/cortexm0ds_logic.v(1512)
  wire Fseow6;  // ../RTL/cortexm0ds_logic.v(1044)
  wire Fskiu6;  // ../RTL/cortexm0ds_logic.v(581)
  wire Fslow6;  // ../RTL/cortexm0ds_logic.v(1138)
  wire Fsriu6;  // ../RTL/cortexm0ds_logic.v(675)
  wire Fsshu6;  // ../RTL/cortexm0ds_logic.v(207)
  wire Fssow6;  // ../RTL/cortexm0ds_logic.v(1231)
  wire Fsyiu6;  // ../RTL/cortexm0ds_logic.v(768)
  wire Fszhu6;  // ../RTL/cortexm0ds_logic.v(300)
  wire Fszow6;  // ../RTL/cortexm0ds_logic.v(1325)
  wire Ft4ju6;  // ../RTL/cortexm0ds_logic.v(849)
  wire Ft5iu6;  // ../RTL/cortexm0ds_logic.v(381)
  wire Ft5pw6;  // ../RTL/cortexm0ds_logic.v(1405)
  wire Ft6ow6;  // ../RTL/cortexm0ds_logic.v(937)
  wire Ftaax6;  // ../RTL/cortexm0ds_logic.v(1633)
  wire Ftciu6;  // ../RTL/cortexm0ds_logic.v(475)
  wire Ftcpw6;  // ../RTL/cortexm0ds_logic.v(1499)
  wire Ftdow6;  // ../RTL/cortexm0ds_logic.v(1031)
  wire Ftghu6;  // ../RTL/cortexm0ds_logic.v(127)
  wire Ftjiu6;  // ../RTL/cortexm0ds_logic.v(568)
  wire Ftkow6;  // ../RTL/cortexm0ds_logic.v(1125)
  wire Ftqiu6;  // ../RTL/cortexm0ds_logic.v(662)
  wire Ftrhu6;  // ../RTL/cortexm0ds_logic.v(194)
  wire Ftrow6;  // ../RTL/cortexm0ds_logic.v(1218)
  wire Ftxiu6;  // ../RTL/cortexm0ds_logic.v(755)
  wire Ftyhu6;  // ../RTL/cortexm0ds_logic.v(287)
  wire Ftyow6;  // ../RTL/cortexm0ds_logic.v(1312)
  wire Ftypw6;  // ../RTL/cortexm0ds_logic.v(1615)
  wire Fu3ju6;  // ../RTL/cortexm0ds_logic.v(836)
  wire Fu4iu6;  // ../RTL/cortexm0ds_logic.v(368)
  wire Fu4pw6;  // ../RTL/cortexm0ds_logic.v(1392)
  wire Fubiu6;  // ../RTL/cortexm0ds_logic.v(462)
  wire Fubpw6;  // ../RTL/cortexm0ds_logic.v(1486)
  wire Fucow6;  // ../RTL/cortexm0ds_logic.v(1018)
  wire Fuiiu6;  // ../RTL/cortexm0ds_logic.v(555)
  wire Fujow6;  // ../RTL/cortexm0ds_logic.v(1112)
  wire Fulhu6;  // ../RTL/cortexm0ds_logic.v(140)
  wire Fupiu6;  // ../RTL/cortexm0ds_logic.v(649)
  wire Fuqhu6;  // ../RTL/cortexm0ds_logic.v(181)
  wire Fuqow6;  // ../RTL/cortexm0ds_logic.v(1205)
  wire Fuwiu6;  // ../RTL/cortexm0ds_logic.v(742)
  wire Fuxhu6;  // ../RTL/cortexm0ds_logic.v(274)
  wire Fuxow6;  // ../RTL/cortexm0ds_logic.v(1299)
  wire Fv2ju6;  // ../RTL/cortexm0ds_logic.v(823)
  wire Fv3iu6;  // ../RTL/cortexm0ds_logic.v(355)
  wire Fv3pw6;  // ../RTL/cortexm0ds_logic.v(1379)
  wire Fv9ju6;  // ../RTL/cortexm0ds_logic.v(917)
  wire Fvaiu6;  // ../RTL/cortexm0ds_logic.v(449)
  wire Fvapw6;  // ../RTL/cortexm0ds_logic.v(1473)
  wire Fvbow6;  // ../RTL/cortexm0ds_logic.v(1005)
  wire Fvcbx6;  // ../RTL/cortexm0ds_logic.v(1702)
  wire Fvdhu6;  // ../RTL/cortexm0ds_logic.v(120)
  wire Fvhiu6;  // ../RTL/cortexm0ds_logic.v(542)
  wire Fviow6;  // ../RTL/cortexm0ds_logic.v(1099)
  wire Fvoax6;  // ../RTL/cortexm0ds_logic.v(1659)
  wire Fvoiu6;  // ../RTL/cortexm0ds_logic.v(636)
  wire Fvphu6;  // ../RTL/cortexm0ds_logic.v(168)
  wire Fvpow6;  // ../RTL/cortexm0ds_logic.v(1192)
  wire Fvviu6;  // ../RTL/cortexm0ds_logic.v(729)
  wire Fvwhu6;  // ../RTL/cortexm0ds_logic.v(261)
  wire Fvwow6;  // ../RTL/cortexm0ds_logic.v(1286)
  wire Fw1ju6;  // ../RTL/cortexm0ds_logic.v(810)
  wire Fw2iu6;  // ../RTL/cortexm0ds_logic.v(342)
  wire Fw2pw6;  // ../RTL/cortexm0ds_logic.v(1366)
  wire Fw8ju6;  // ../RTL/cortexm0ds_logic.v(904)
  wire Fw9iu6;  // ../RTL/cortexm0ds_logic.v(436)
  wire Fw9pw6;  // ../RTL/cortexm0ds_logic.v(1460)
  wire Fwaow6;  // ../RTL/cortexm0ds_logic.v(992)
  wire Fwgiu6;  // ../RTL/cortexm0ds_logic.v(529)
  wire Fwhow6;  // ../RTL/cortexm0ds_logic.v(1086)
  wire Fwniu6;  // ../RTL/cortexm0ds_logic.v(623)
  wire Fwohu6;  // ../RTL/cortexm0ds_logic.v(155)
  wire Fwoow6;  // ../RTL/cortexm0ds_logic.v(1179)
  wire Fwuiu6;  // ../RTL/cortexm0ds_logic.v(716)
  wire Fwvhu6;  // ../RTL/cortexm0ds_logic.v(248)
  wire Fwvow6;  // ../RTL/cortexm0ds_logic.v(1273)
  wire Fx0ju6;  // ../RTL/cortexm0ds_logic.v(797)
  wire Fx1iu6;  // ../RTL/cortexm0ds_logic.v(329)
  wire Fx1pw6;  // ../RTL/cortexm0ds_logic.v(1353)
  wire Fx1qw6;  // ../RTL/cortexm0ds_logic.v(1620)
  wire Fx7ju6;  // ../RTL/cortexm0ds_logic.v(891)
  wire Fx8iu6;  // ../RTL/cortexm0ds_logic.v(423)
  wire Fx8pw6;  // ../RTL/cortexm0ds_logic.v(1447)
  wire Fx9ow6;  // ../RTL/cortexm0ds_logic.v(979)
  wire Fxfiu6;  // ../RTL/cortexm0ds_logic.v(516)
  wire Fxgow6;  // ../RTL/cortexm0ds_logic.v(1073)
  wire Fxmiu6;  // ../RTL/cortexm0ds_logic.v(610)
  wire Fxnow6;  // ../RTL/cortexm0ds_logic.v(1166)
  wire Fxoax6;  // ../RTL/cortexm0ds_logic.v(1659)
  wire Fxtiu6;  // ../RTL/cortexm0ds_logic.v(703)
  wire Fxuhu6;  // ../RTL/cortexm0ds_logic.v(235)
  wire Fxuow6;  // ../RTL/cortexm0ds_logic.v(1260)
  wire Fy0iu6;  // ../RTL/cortexm0ds_logic.v(316)
  wire Fy0pw6;  // ../RTL/cortexm0ds_logic.v(1340)
  wire Fy6ju6;  // ../RTL/cortexm0ds_logic.v(878)
  wire Fy7iu6;  // ../RTL/cortexm0ds_logic.v(410)
  wire Fy7pw6;  // ../RTL/cortexm0ds_logic.v(1434)
  wire Fy8ow6;  // ../RTL/cortexm0ds_logic.v(966)
  wire Fyeiu6;  // ../RTL/cortexm0ds_logic.v(503)
  wire Fyfow6;  // ../RTL/cortexm0ds_logic.v(1060)
  wire Fyliu6;  // ../RTL/cortexm0ds_logic.v(597)
  wire Fymow6;  // ../RTL/cortexm0ds_logic.v(1153)
  wire Fysiu6;  // ../RTL/cortexm0ds_logic.v(690)
  wire Fythu6;  // ../RTL/cortexm0ds_logic.v(222)
  wire Fytow6;  // ../RTL/cortexm0ds_logic.v(1247)
  wire Fyziu6;  // ../RTL/cortexm0ds_logic.v(784)
  wire Fz5ju6;  // ../RTL/cortexm0ds_logic.v(865)
  wire Fz6iu6;  // ../RTL/cortexm0ds_logic.v(397)
  wire Fz6pw6;  // ../RTL/cortexm0ds_logic.v(1421)
  wire Fz7ow6;  // ../RTL/cortexm0ds_logic.v(953)
  wire Fzdiu6;  // ../RTL/cortexm0ds_logic.v(490)
  wire Fzdpw6;  // ../RTL/cortexm0ds_logic.v(1515)
  wire Fzeow6;  // ../RTL/cortexm0ds_logic.v(1047)
  wire Fzkiu6;  // ../RTL/cortexm0ds_logic.v(584)
  wire Fzlow6;  // ../RTL/cortexm0ds_logic.v(1140)
  wire Fzmpw6;  // ../RTL/cortexm0ds_logic.v(1593)
  wire Fzoax6;  // ../RTL/cortexm0ds_logic.v(1659)
  wire Fzriu6;  // ../RTL/cortexm0ds_logic.v(677)
  wire Fzshu6;  // ../RTL/cortexm0ds_logic.v(209)
  wire Fzsow6;  // ../RTL/cortexm0ds_logic.v(1234)
  wire Fzyiu6;  // ../RTL/cortexm0ds_logic.v(771)
  wire Fzzhu6;  // ../RTL/cortexm0ds_logic.v(303)
  wire Fzzow6;  // ../RTL/cortexm0ds_logic.v(1327)
  wire G02ju6;  // ../RTL/cortexm0ds_logic.v(812)
  wire G03iu6;  // ../RTL/cortexm0ds_logic.v(344)
  wire G03pw6;  // ../RTL/cortexm0ds_logic.v(1368)
  wire G09ju6;  // ../RTL/cortexm0ds_logic.v(905)
  wire G0aiu6;  // ../RTL/cortexm0ds_logic.v(437)
  wire G0apw6;  // ../RTL/cortexm0ds_logic.v(1462)
  wire G0bow6;  // ../RTL/cortexm0ds_logic.v(994)
  wire G0fhu6;  // ../RTL/cortexm0ds_logic.v(123)
  wire G0hiu6;  // ../RTL/cortexm0ds_logic.v(531)
  wire G0iow6;  // ../RTL/cortexm0ds_logic.v(1087)
  wire G0oiu6;  // ../RTL/cortexm0ds_logic.v(624)
  wire G0phu6;  // ../RTL/cortexm0ds_logic.v(156)
  wire G0pow6;  // ../RTL/cortexm0ds_logic.v(1181)
  wire G0tax6;  // ../RTL/cortexm0ds_logic.v(1667)
  wire G0viu6;  // ../RTL/cortexm0ds_logic.v(718)
  wire G0whu6;  // ../RTL/cortexm0ds_logic.v(250)
  wire G0wow6;  // ../RTL/cortexm0ds_logic.v(1274)
  wire G0zax6;  // ../RTL/cortexm0ds_logic.v(1678)
  wire G11ju6;  // ../RTL/cortexm0ds_logic.v(799)
  wire G12iu6;  // ../RTL/cortexm0ds_logic.v(331)
  wire G12pw6;  // ../RTL/cortexm0ds_logic.v(1355)
  wire G18ju6;  // ../RTL/cortexm0ds_logic.v(892)
  wire G19iu6;  // ../RTL/cortexm0ds_logic.v(424)
  wire G19pw6;  // ../RTL/cortexm0ds_logic.v(1449)
  wire G1aow6;  // ../RTL/cortexm0ds_logic.v(981)
  wire G1giu6;  // ../RTL/cortexm0ds_logic.v(518)
  wire G1how6;  // ../RTL/cortexm0ds_logic.v(1074)
  wire G1niu6;  // ../RTL/cortexm0ds_logic.v(611)
  wire G1oow6;  // ../RTL/cortexm0ds_logic.v(1168)
  wire G1uiu6;  // ../RTL/cortexm0ds_logic.v(705)
  wire G1vhu6;  // ../RTL/cortexm0ds_logic.v(237)
  wire G1vow6;  // ../RTL/cortexm0ds_logic.v(1261)
  wire G20ju6;  // ../RTL/cortexm0ds_logic.v(786)
  wire G21iu6;  // ../RTL/cortexm0ds_logic.v(318)
  wire G21pw6;  // ../RTL/cortexm0ds_logic.v(1342)
  wire G25bx6;  // ../RTL/cortexm0ds_logic.v(1688)
  wire G27ju6;  // ../RTL/cortexm0ds_logic.v(879)
  wire G28iu6;  // ../RTL/cortexm0ds_logic.v(411)
  wire G28pw6;  // ../RTL/cortexm0ds_logic.v(1436)
  wire G29ow6;  // ../RTL/cortexm0ds_logic.v(968)
  wire G2fiu6;  // ../RTL/cortexm0ds_logic.v(505)
  wire G2gow6;  // ../RTL/cortexm0ds_logic.v(1061)
  wire G2iax6;  // ../RTL/cortexm0ds_logic.v(1647)
  wire G2miu6;  // ../RTL/cortexm0ds_logic.v(598)
  wire G2now6;  // ../RTL/cortexm0ds_logic.v(1155)
  wire G2ohu6;  // ../RTL/cortexm0ds_logic.v(146)
  wire G2tiu6;  // ../RTL/cortexm0ds_logic.v(692)
  wire G2uhu6;  // ../RTL/cortexm0ds_logic.v(224)
  wire G2uow6;  // ../RTL/cortexm0ds_logic.v(1248)
  wire G30iu6;  // ../RTL/cortexm0ds_logic.v(305)
  wire G30pw6;  // ../RTL/cortexm0ds_logic.v(1329)
  wire G36ju6;  // ../RTL/cortexm0ds_logic.v(866)
  wire G37iu6;  // ../RTL/cortexm0ds_logic.v(398)
  wire G37pw6;  // ../RTL/cortexm0ds_logic.v(1423)
  wire G38ow6;  // ../RTL/cortexm0ds_logic.v(955)
  wire G3eiu6;  // ../RTL/cortexm0ds_logic.v(492)
  wire G3epw6;  // ../RTL/cortexm0ds_logic.v(1516)
  wire G3fow6;  // ../RTL/cortexm0ds_logic.v(1048)
  wire G3liu6;  // ../RTL/cortexm0ds_logic.v(585)
  wire G3mow6;  // ../RTL/cortexm0ds_logic.v(1142)
  wire G3siu6;  // ../RTL/cortexm0ds_logic.v(679)
  wire G3thu6;  // ../RTL/cortexm0ds_logic.v(211)
  wire G3tow6;  // ../RTL/cortexm0ds_logic.v(1235)
  wire G3ziu6;  // ../RTL/cortexm0ds_logic.v(773)
  wire G45ju6;  // ../RTL/cortexm0ds_logic.v(853)
  wire G46iu6;  // ../RTL/cortexm0ds_logic.v(385)
  wire G46pw6;  // ../RTL/cortexm0ds_logic.v(1410)
  wire G47ow6;  // ../RTL/cortexm0ds_logic.v(942)
  wire G4diu6;  // ../RTL/cortexm0ds_logic.v(479)
  wire G4dpw6;  // ../RTL/cortexm0ds_logic.v(1503)
  wire G4eow6;  // ../RTL/cortexm0ds_logic.v(1035)
  wire G4kiu6;  // ../RTL/cortexm0ds_logic.v(572)
  wire G4low6;  // ../RTL/cortexm0ds_logic.v(1129)
  wire G4riu6;  // ../RTL/cortexm0ds_logic.v(666)
  wire G4shu6;  // ../RTL/cortexm0ds_logic.v(198)
  wire G4sow6;  // ../RTL/cortexm0ds_logic.v(1222)
  wire G4yiu6;  // ../RTL/cortexm0ds_logic.v(760)
  wire G4zhu6;  // ../RTL/cortexm0ds_logic.v(292)
  wire G4zow6;  // ../RTL/cortexm0ds_logic.v(1316)
  wire G54bx6;  // ../RTL/cortexm0ds_logic.v(1686)
  wire G54ju6;  // ../RTL/cortexm0ds_logic.v(840)
  wire G55iu6;  // ../RTL/cortexm0ds_logic.v(372)
  wire G55pw6;  // ../RTL/cortexm0ds_logic.v(1397)
  wire G5ciu6;  // ../RTL/cortexm0ds_logic.v(466)
  wire G5cpw6;  // ../RTL/cortexm0ds_logic.v(1490)
  wire G5dow6;  // ../RTL/cortexm0ds_logic.v(1022)
  wire G5jiu6;  // ../RTL/cortexm0ds_logic.v(559)
  wire G5kow6;  // ../RTL/cortexm0ds_logic.v(1116)
  wire G5qiu6;  // ../RTL/cortexm0ds_logic.v(653)
  wire G5rhu6;  // ../RTL/cortexm0ds_logic.v(185)
  wire G5row6;  // ../RTL/cortexm0ds_logic.v(1209)
  wire G5xiu6;  // ../RTL/cortexm0ds_logic.v(747)
  wire G5yhu6;  // ../RTL/cortexm0ds_logic.v(279)
  wire G5yow6;  // ../RTL/cortexm0ds_logic.v(1303)
  wire G63ju6;  // ../RTL/cortexm0ds_logic.v(827)
  wire G64iu6;  // ../RTL/cortexm0ds_logic.v(359)
  wire G64pw6;  // ../RTL/cortexm0ds_logic.v(1384)
  wire G6aju6;  // ../RTL/cortexm0ds_logic.v(921)
  wire G6biu6;  // ../RTL/cortexm0ds_logic.v(453)
  wire G6bpw6;  // ../RTL/cortexm0ds_logic.v(1477)
  wire G6cow6;  // ../RTL/cortexm0ds_logic.v(1009)
  wire G6iiu6;  // ../RTL/cortexm0ds_logic.v(546)
  wire G6jow6;  // ../RTL/cortexm0ds_logic.v(1103)
  wire G6piu6;  // ../RTL/cortexm0ds_logic.v(640)
  wire G6qhu6;  // ../RTL/cortexm0ds_logic.v(172)
  wire G6qow6;  // ../RTL/cortexm0ds_logic.v(1196)
  wire G6wiu6;  // ../RTL/cortexm0ds_logic.v(734)
  wire G6xhu6;  // ../RTL/cortexm0ds_logic.v(266)
  wire G6xow6;  // ../RTL/cortexm0ds_logic.v(1290)
  wire G72ju6;  // ../RTL/cortexm0ds_logic.v(814)
  wire G73iu6;  // ../RTL/cortexm0ds_logic.v(346)
  wire G73pw6;  // ../RTL/cortexm0ds_logic.v(1371)
  wire G79ax6;  // ../RTL/cortexm0ds_logic.v(1630)
  wire G79ju6;  // ../RTL/cortexm0ds_logic.v(908)
  wire G7aiu6;  // ../RTL/cortexm0ds_logic.v(440)
  wire G7apw6;  // ../RTL/cortexm0ds_logic.v(1464)
  wire G7bow6;  // ../RTL/cortexm0ds_logic.v(996)
  wire G7hiu6;  // ../RTL/cortexm0ds_logic.v(533)
  wire G7iow6;  // ../RTL/cortexm0ds_logic.v(1090)
  wire G7lhu6;  // ../RTL/cortexm0ds_logic.v(138)
  wire G7oiu6;  // ../RTL/cortexm0ds_logic.v(627)
  wire G7phu6;  // ../RTL/cortexm0ds_logic.v(159)
  wire G7pow6;  // ../RTL/cortexm0ds_logic.v(1183)
  wire G7viu6;  // ../RTL/cortexm0ds_logic.v(721)
  wire G7whu6;  // ../RTL/cortexm0ds_logic.v(253)
  wire G7wow6;  // ../RTL/cortexm0ds_logic.v(1277)
  wire G81ju6;  // ../RTL/cortexm0ds_logic.v(801)
  wire G82iu6;  // ../RTL/cortexm0ds_logic.v(333)
  wire G82pw6;  // ../RTL/cortexm0ds_logic.v(1358)
  wire G88ju6;  // ../RTL/cortexm0ds_logic.v(895)
  wire G89iu6;  // ../RTL/cortexm0ds_logic.v(427)
  wire G89pw6;  // ../RTL/cortexm0ds_logic.v(1451)
  wire G8aow6;  // ../RTL/cortexm0ds_logic.v(983)
  wire G8ebx6;  // ../RTL/cortexm0ds_logic.v(1705)
  wire G8giu6;  // ../RTL/cortexm0ds_logic.v(520)
  wire G8how6;  // ../RTL/cortexm0ds_logic.v(1077)
  wire G8niu6;  // ../RTL/cortexm0ds_logic.v(614)
  wire G8oow6;  // ../RTL/cortexm0ds_logic.v(1170)
  wire G8uiu6;  // ../RTL/cortexm0ds_logic.v(708)
  wire G8vhu6;  // ../RTL/cortexm0ds_logic.v(240)
  wire G8vow6;  // ../RTL/cortexm0ds_logic.v(1264)
  wire G90ju6;  // ../RTL/cortexm0ds_logic.v(788)
  wire G91iu6;  // ../RTL/cortexm0ds_logic.v(320)
  wire G91pw6;  // ../RTL/cortexm0ds_logic.v(1345)
  wire G97ju6;  // ../RTL/cortexm0ds_logic.v(882)
  wire G98iu6;  // ../RTL/cortexm0ds_logic.v(414)
  wire G98pw6;  // ../RTL/cortexm0ds_logic.v(1438)
  wire G99ow6;  // ../RTL/cortexm0ds_logic.v(970)
  wire G9fiu6;  // ../RTL/cortexm0ds_logic.v(507)
  wire G9gow6;  // ../RTL/cortexm0ds_logic.v(1064)
  wire G9khu6;  // ../RTL/cortexm0ds_logic.v(136)
  wire G9miu6;  // ../RTL/cortexm0ds_logic.v(601)
  wire G9now6;  // ../RTL/cortexm0ds_logic.v(1157)
  wire G9tiu6;  // ../RTL/cortexm0ds_logic.v(695)
  wire G9uhu6;  // ../RTL/cortexm0ds_logic.v(227)
  wire G9uow6;  // ../RTL/cortexm0ds_logic.v(1251)
  wire Ga0iu6;  // ../RTL/cortexm0ds_logic.v(307)
  wire Ga0pw6;  // ../RTL/cortexm0ds_logic.v(1332)
  wire Ga6ju6;  // ../RTL/cortexm0ds_logic.v(869)
  wire Ga7iu6;  // ../RTL/cortexm0ds_logic.v(401)
  wire Ga7pw6;  // ../RTL/cortexm0ds_logic.v(1425)
  wire Ga8ow6;  // ../RTL/cortexm0ds_logic.v(957)
  wire Gaeiu6;  // ../RTL/cortexm0ds_logic.v(494)
  wire Gafow6;  // ../RTL/cortexm0ds_logic.v(1051)
  wire Galiu6;  // ../RTL/cortexm0ds_logic.v(588)
  wire Gamow6;  // ../RTL/cortexm0ds_logic.v(1144)
  wire Gasiu6;  // ../RTL/cortexm0ds_logic.v(682)
  wire Gathu6;  // ../RTL/cortexm0ds_logic.v(214)
  wire Gatow6;  // ../RTL/cortexm0ds_logic.v(1238)
  wire Gaziu6;  // ../RTL/cortexm0ds_logic.v(775)
  wire Gb5ju6;  // ../RTL/cortexm0ds_logic.v(856)
  wire Gb6iu6;  // ../RTL/cortexm0ds_logic.v(388)
  wire Gb6pw6;  // ../RTL/cortexm0ds_logic.v(1412)
  wire Gb7ow6;  // ../RTL/cortexm0ds_logic.v(944)
  wire Gbdiu6;  // ../RTL/cortexm0ds_logic.v(481)
  wire Gbdpw6;  // ../RTL/cortexm0ds_logic.v(1506)
  wire Gbeow6;  // ../RTL/cortexm0ds_logic.v(1038)
  wire Gbjhu6;  // ../RTL/cortexm0ds_logic.v(133)
  wire Gbkiu6;  // ../RTL/cortexm0ds_logic.v(575)
  wire Gblow6;  // ../RTL/cortexm0ds_logic.v(1131)
  wire Gbriu6;  // ../RTL/cortexm0ds_logic.v(669)
  wire Gbshu6;  // ../RTL/cortexm0ds_logic.v(201)
  wire Gbsow6;  // ../RTL/cortexm0ds_logic.v(1225)
  wire Gbvpw6;  // ../RTL/cortexm0ds_logic.v(1608)
  wire Gbyiu6;  // ../RTL/cortexm0ds_logic.v(762)
  wire Gbzhu6;  // ../RTL/cortexm0ds_logic.v(294)
  wire Gbzow6;  // ../RTL/cortexm0ds_logic.v(1319)
  wire Gc1qw6;  // ../RTL/cortexm0ds_logic.v(1619)
  wire Gc4ju6;  // ../RTL/cortexm0ds_logic.v(843)
  wire Gc5iu6;  // ../RTL/cortexm0ds_logic.v(375)
  wire Gc5pw6;  // ../RTL/cortexm0ds_logic.v(1399)
  wire Gc6ow6;  // ../RTL/cortexm0ds_logic.v(931)
  wire Gcciu6;  // ../RTL/cortexm0ds_logic.v(468)
  wire Gccpw6;  // ../RTL/cortexm0ds_logic.v(1493)
  wire Gcdow6;  // ../RTL/cortexm0ds_logic.v(1025)
  wire Gcjiu6;  // ../RTL/cortexm0ds_logic.v(562)
  wire Gckow6;  // ../RTL/cortexm0ds_logic.v(1118)
  wire Gcqiu6;  // ../RTL/cortexm0ds_logic.v(656)
  wire Gcrhu6;  // ../RTL/cortexm0ds_logic.v(188)
  wire Gcrow6;  // ../RTL/cortexm0ds_logic.v(1212)
  wire Gcxiu6;  // ../RTL/cortexm0ds_logic.v(749)
  wire Gcyhu6;  // ../RTL/cortexm0ds_logic.v(281)
  wire Gcyow6;  // ../RTL/cortexm0ds_logic.v(1306)
  wire Gd0bx6;  // ../RTL/cortexm0ds_logic.v(1680)
  wire Gd3ju6;  // ../RTL/cortexm0ds_logic.v(830)
  wire Gd4iu6;  // ../RTL/cortexm0ds_logic.v(362)
  wire Gd4pw6;  // ../RTL/cortexm0ds_logic.v(1386)
  wire Gdaju6;  // ../RTL/cortexm0ds_logic.v(923)
  wire Gdbiu6;  // ../RTL/cortexm0ds_logic.v(455)
  wire Gdbpw6;  // ../RTL/cortexm0ds_logic.v(1480)
  wire Gdcow6;  // ../RTL/cortexm0ds_logic.v(1012)
  wire Gdihu6;  // ../RTL/cortexm0ds_logic.v(131)
  wire Gdiiu6;  // ../RTL/cortexm0ds_logic.v(549)
  wire Gdjow6;  // ../RTL/cortexm0ds_logic.v(1105)
  wire Gdmhu6;  // ../RTL/cortexm0ds_logic.v(142)
  wire Gdpiu6;  // ../RTL/cortexm0ds_logic.v(643)
  wire Gdqhu6;  // ../RTL/cortexm0ds_logic.v(175)
  wire Gdqow6;  // ../RTL/cortexm0ds_logic.v(1199)
  wire Gdwiu6;  // ../RTL/cortexm0ds_logic.v(736)
  wire Gdxhu6;  // ../RTL/cortexm0ds_logic.v(268)
  wire Gdxow6;  // ../RTL/cortexm0ds_logic.v(1293)
  wire Ge2ju6;  // ../RTL/cortexm0ds_logic.v(817)
  wire Ge3iu6;  // ../RTL/cortexm0ds_logic.v(349)
  wire Ge3pw6;  // ../RTL/cortexm0ds_logic.v(1373)
  wire Ge9ju6;  // ../RTL/cortexm0ds_logic.v(910)
  wire Geaiu6;  // ../RTL/cortexm0ds_logic.v(442)
  wire Geapw6;  // ../RTL/cortexm0ds_logic.v(1467)
  wire Gebow6;  // ../RTL/cortexm0ds_logic.v(999)
  wire Gehiu6;  // ../RTL/cortexm0ds_logic.v(536)
  wire Geiow6;  // ../RTL/cortexm0ds_logic.v(1092)
  wire Geoiu6;  // ../RTL/cortexm0ds_logic.v(630)
  wire Gephu6;  // ../RTL/cortexm0ds_logic.v(162)
  wire Gepow6;  // ../RTL/cortexm0ds_logic.v(1186)
  wire Geviu6;  // ../RTL/cortexm0ds_logic.v(723)
  wire Gewhu6;  // ../RTL/cortexm0ds_logic.v(255)
  wire Gewow6;  // ../RTL/cortexm0ds_logic.v(1280)
  wire Gf1ju6;  // ../RTL/cortexm0ds_logic.v(804)
  wire Gf2iu6;  // ../RTL/cortexm0ds_logic.v(336)
  wire Gf2pw6;  // ../RTL/cortexm0ds_logic.v(1360)
  wire Gf8ju6;  // ../RTL/cortexm0ds_logic.v(897)
  wire Gf9iu6;  // ../RTL/cortexm0ds_logic.v(429)
  wire Gf9pw6;  // ../RTL/cortexm0ds_logic.v(1454)
  wire Gfaow6;  // ../RTL/cortexm0ds_logic.v(986)
  wire Gfghu6;  // ../RTL/cortexm0ds_logic.v(126)
  wire Gfgiu6;  // ../RTL/cortexm0ds_logic.v(523)
  wire Gfhow6;  // ../RTL/cortexm0ds_logic.v(1079)
  wire Gfniu6;  // ../RTL/cortexm0ds_logic.v(617)
  wire Gfohu6;  // ../RTL/cortexm0ds_logic.v(149)
  wire Gfoow6;  // ../RTL/cortexm0ds_logic.v(1173)
  wire Gfuiu6;  // ../RTL/cortexm0ds_logic.v(710)
  wire Gfvhu6;  // ../RTL/cortexm0ds_logic.v(242)
  wire Gfvow6;  // ../RTL/cortexm0ds_logic.v(1267)
  wire Gg0ju6;  // ../RTL/cortexm0ds_logic.v(791)
  wire Gg1iu6;  // ../RTL/cortexm0ds_logic.v(323)
  wire Gg1pw6;  // ../RTL/cortexm0ds_logic.v(1347)
  wire Gg7ju6;  // ../RTL/cortexm0ds_logic.v(884)
  wire Gg8iu6;  // ../RTL/cortexm0ds_logic.v(416)
  wire Gg8pw6;  // ../RTL/cortexm0ds_logic.v(1441)
  wire Gg9ow6;  // ../RTL/cortexm0ds_logic.v(973)
  wire Ggabx6;  // ../RTL/cortexm0ds_logic.v(1698)
  wire Ggehu6;  // ../RTL/cortexm0ds_logic.v(122)
  wire Ggfiu6;  // ../RTL/cortexm0ds_logic.v(510)
  wire Gggow6;  // ../RTL/cortexm0ds_logic.v(1066)
  wire Gglhu6;  // ../RTL/cortexm0ds_logic.v(139)
  wire Ggmiu6;  // ../RTL/cortexm0ds_logic.v(604)
  wire Ggnow6;  // ../RTL/cortexm0ds_logic.v(1160)
  wire Ggtiu6;  // ../RTL/cortexm0ds_logic.v(697)
  wire Gguhu6;  // ../RTL/cortexm0ds_logic.v(229)
  wire Gguow6;  // ../RTL/cortexm0ds_logic.v(1254)
  wire Gh0iu6;  // ../RTL/cortexm0ds_logic.v(310)
  wire Gh0pw6;  // ../RTL/cortexm0ds_logic.v(1334)
  wire Gh6ju6;  // ../RTL/cortexm0ds_logic.v(871)
  wire Gh7iu6;  // ../RTL/cortexm0ds_logic.v(403)
  wire Gh7pw6;  // ../RTL/cortexm0ds_logic.v(1428)
  wire Gh8ow6;  // ../RTL/cortexm0ds_logic.v(960)
  wire Gheiu6;  // ../RTL/cortexm0ds_logic.v(497)
  wire Ghfow6;  // ../RTL/cortexm0ds_logic.v(1053)
  wire Ghliu6;  // ../RTL/cortexm0ds_logic.v(591)
  wire Ghmow6;  // ../RTL/cortexm0ds_logic.v(1147)
  wire Ghsiu6;  // ../RTL/cortexm0ds_logic.v(684)
  wire Ghthu6;  // ../RTL/cortexm0ds_logic.v(216)
  wire Ghtow6;  // ../RTL/cortexm0ds_logic.v(1241)
  wire Ghziu6;  // ../RTL/cortexm0ds_logic.v(778)
  wire Gi5ju6;  // ../RTL/cortexm0ds_logic.v(858)
  wire Gi6iu6;  // ../RTL/cortexm0ds_logic.v(390)
  wire Gi6pw6;  // ../RTL/cortexm0ds_logic.v(1415)
  wire Gi7ow6;  // ../RTL/cortexm0ds_logic.v(947)
  wire Gidiu6;  // ../RTL/cortexm0ds_logic.v(484)
  wire Gidpw6;  // ../RTL/cortexm0ds_logic.v(1508)
  wire Gieow6;  // ../RTL/cortexm0ds_logic.v(1040)
  wire Gihbx6;  // ../RTL/cortexm0ds_logic.v(1711)
  wire Gikiu6;  // ../RTL/cortexm0ds_logic.v(578)
  wire Gilow6;  // ../RTL/cortexm0ds_logic.v(1134)
  wire Giriu6;  // ../RTL/cortexm0ds_logic.v(671)
  wire Gishu6;  // ../RTL/cortexm0ds_logic.v(203)
  wire Gisow6;  // ../RTL/cortexm0ds_logic.v(1228)
  wire Giyiu6;  // ../RTL/cortexm0ds_logic.v(765)
  wire Gizhu6;  // ../RTL/cortexm0ds_logic.v(297)
  wire Gizow6;  // ../RTL/cortexm0ds_logic.v(1321)
  wire Gj4ju6;  // ../RTL/cortexm0ds_logic.v(845)
  wire Gj5iu6;  // ../RTL/cortexm0ds_logic.v(377)
  wire Gj5pw6;  // ../RTL/cortexm0ds_logic.v(1402)
  wire Gj6ow6;  // ../RTL/cortexm0ds_logic.v(934)
  wire Gjciu6;  // ../RTL/cortexm0ds_logic.v(471)
  wire Gjcpw6;  // ../RTL/cortexm0ds_logic.v(1495)
  wire Gjdow6;  // ../RTL/cortexm0ds_logic.v(1027)
  wire Gjjiu6;  // ../RTL/cortexm0ds_logic.v(565)
  wire Gjkow6;  // ../RTL/cortexm0ds_logic.v(1121)
  wire Gjqiu6;  // ../RTL/cortexm0ds_logic.v(658)
  wire Gjrhu6;  // ../RTL/cortexm0ds_logic.v(190)
  wire Gjrow6;  // ../RTL/cortexm0ds_logic.v(1215)
  wire Gjxiu6;  // ../RTL/cortexm0ds_logic.v(752)
  wire Gjyhu6;  // ../RTL/cortexm0ds_logic.v(284)
  wire Gjyow6;  // ../RTL/cortexm0ds_logic.v(1308)
  wire Gk3ju6;  // ../RTL/cortexm0ds_logic.v(832)
  wire Gk4iu6;  // ../RTL/cortexm0ds_logic.v(364)
  wire Gk4pw6;  // ../RTL/cortexm0ds_logic.v(1389)
  wire Gkaju6;  // ../RTL/cortexm0ds_logic.v(926)
  wire Gkbiu6;  // ../RTL/cortexm0ds_logic.v(458)
  wire Gkbpw6;  // ../RTL/cortexm0ds_logic.v(1482)
  wire Gkcow6;  // ../RTL/cortexm0ds_logic.v(1014)
  wire Gkeax6;  // ../RTL/cortexm0ds_logic.v(1640)
  wire Gkiiu6;  // ../RTL/cortexm0ds_logic.v(552)
  wire Gkjow6;  // ../RTL/cortexm0ds_logic.v(1108)
  wire Gkpiu6;  // ../RTL/cortexm0ds_logic.v(645)
  wire Gkqhu6;  // ../RTL/cortexm0ds_logic.v(177)
  wire Gkqow6;  // ../RTL/cortexm0ds_logic.v(1202)
  wire Gkwiu6;  // ../RTL/cortexm0ds_logic.v(739)
  wire Gkxhu6;  // ../RTL/cortexm0ds_logic.v(271)
  wire Gkxow6;  // ../RTL/cortexm0ds_logic.v(1295)
  wire Gl1qw6;  // ../RTL/cortexm0ds_logic.v(1620)
  wire Gl2ju6;  // ../RTL/cortexm0ds_logic.v(819)
  wire Gl3iu6;  // ../RTL/cortexm0ds_logic.v(351)
  wire Gl3pw6;  // ../RTL/cortexm0ds_logic.v(1376)
  wire Gl9ju6;  // ../RTL/cortexm0ds_logic.v(913)
  wire Glaiu6;  // ../RTL/cortexm0ds_logic.v(445)
  wire Glapw6;  // ../RTL/cortexm0ds_logic.v(1469)
  wire Glbow6;  // ../RTL/cortexm0ds_logic.v(1001)
  wire Glhiu6;  // ../RTL/cortexm0ds_logic.v(539)
  wire Gliow6;  // ../RTL/cortexm0ds_logic.v(1095)
  wire Gloiu6;  // ../RTL/cortexm0ds_logic.v(632)
  wire Glphu6;  // ../RTL/cortexm0ds_logic.v(164)
  wire Glpow6;  // ../RTL/cortexm0ds_logic.v(1189)
  wire Glviu6;  // ../RTL/cortexm0ds_logic.v(726)
  wire Glwhu6;  // ../RTL/cortexm0ds_logic.v(258)
  wire Glwow6;  // ../RTL/cortexm0ds_logic.v(1282)
  wire Gm1ju6;  // ../RTL/cortexm0ds_logic.v(806)
  wire Gm2iu6;  // ../RTL/cortexm0ds_logic.v(338)
  wire Gm2pw6;  // ../RTL/cortexm0ds_logic.v(1363)
  wire Gm8ju6;  // ../RTL/cortexm0ds_logic.v(900)
  wire Gm9iu6;  // ../RTL/cortexm0ds_logic.v(432)
  wire Gm9pw6;  // ../RTL/cortexm0ds_logic.v(1456)
  wire Gmaow6;  // ../RTL/cortexm0ds_logic.v(988)
  wire Gmgiu6;  // ../RTL/cortexm0ds_logic.v(526)
  wire Gmhow6;  // ../RTL/cortexm0ds_logic.v(1082)
  wire Gmniu6;  // ../RTL/cortexm0ds_logic.v(619)
  wire Gmohu6;  // ../RTL/cortexm0ds_logic.v(151)
  wire Gmoow6;  // ../RTL/cortexm0ds_logic.v(1176)
  wire Gmuiu6;  // ../RTL/cortexm0ds_logic.v(713)
  wire Gmvhu6;  // ../RTL/cortexm0ds_logic.v(245)
  wire Gmvow6;  // ../RTL/cortexm0ds_logic.v(1269)
  wire Gn0ju6;  // ../RTL/cortexm0ds_logic.v(793)
  wire Gn1iu6;  // ../RTL/cortexm0ds_logic.v(325)
  wire Gn1pw6;  // ../RTL/cortexm0ds_logic.v(1350)
  wire Gn7ju6;  // ../RTL/cortexm0ds_logic.v(887)
  wire Gn8iu6;  // ../RTL/cortexm0ds_logic.v(419)
  wire Gn8pw6;  // ../RTL/cortexm0ds_logic.v(1443)
  wire Gn9ow6;  // ../RTL/cortexm0ds_logic.v(975)
  wire Gnfiu6;  // ../RTL/cortexm0ds_logic.v(513)
  wire Gngow6;  // ../RTL/cortexm0ds_logic.v(1069)
  wire Gnmiu6;  // ../RTL/cortexm0ds_logic.v(606)
  wire Gnnow6;  // ../RTL/cortexm0ds_logic.v(1163)
  wire Gnqpw6;  // ../RTL/cortexm0ds_logic.v(1600)
  wire Gntiu6;  // ../RTL/cortexm0ds_logic.v(700)
  wire Gnuhu6;  // ../RTL/cortexm0ds_logic.v(232)
  wire Gnuow6;  // ../RTL/cortexm0ds_logic.v(1256)
  wire Go0iu6;  // ../RTL/cortexm0ds_logic.v(312)
  wire Go0pw6;  // ../RTL/cortexm0ds_logic.v(1337)
  wire Go6ju6;  // ../RTL/cortexm0ds_logic.v(874)
  wire Go7iu6;  // ../RTL/cortexm0ds_logic.v(406)
  wire Go7pw6;  // ../RTL/cortexm0ds_logic.v(1430)
  wire Go8ow6;  // ../RTL/cortexm0ds_logic.v(962)
  wire Goeiu6;  // ../RTL/cortexm0ds_logic.v(500)
  wire Gofow6;  // ../RTL/cortexm0ds_logic.v(1056)
  wire Goliu6;  // ../RTL/cortexm0ds_logic.v(593)
  wire Golpw6;  // ../RTL/cortexm0ds_logic.v(1591)
  wire Gomow6;  // ../RTL/cortexm0ds_logic.v(1150)
  wire Gosiu6;  // ../RTL/cortexm0ds_logic.v(687)
  wire Gothu6;  // ../RTL/cortexm0ds_logic.v(219)
  wire Gotow6;  // ../RTL/cortexm0ds_logic.v(1243)
  wire Goziu6;  // ../RTL/cortexm0ds_logic.v(780)
  wire Gp5ju6;  // ../RTL/cortexm0ds_logic.v(861)
  wire Gp6ax6;  // ../RTL/cortexm0ds_logic.v(1625)
  wire Gp6iu6;  // ../RTL/cortexm0ds_logic.v(393)
  wire Gp6pw6;  // ../RTL/cortexm0ds_logic.v(1417)
  wire Gp7ow6;  // ../RTL/cortexm0ds_logic.v(949)
  wire Gpdiu6;  // ../RTL/cortexm0ds_logic.v(487)
  wire Gpdpw6;  // ../RTL/cortexm0ds_logic.v(1511)
  wire Gpeow6;  // ../RTL/cortexm0ds_logic.v(1043)
  wire Gpkiu6;  // ../RTL/cortexm0ds_logic.v(580)
  wire Gplow6;  // ../RTL/cortexm0ds_logic.v(1137)
  wire Gpqpw6;  // ../RTL/cortexm0ds_logic.v(1600)
  wire Gpriu6;  // ../RTL/cortexm0ds_logic.v(674)
  wire Gpshu6;  // ../RTL/cortexm0ds_logic.v(206)
  wire Gpsow6;  // ../RTL/cortexm0ds_logic.v(1230)
  wire Gpyiu6;  // ../RTL/cortexm0ds_logic.v(767)
  wire Gpzhu6;  // ../RTL/cortexm0ds_logic.v(299)
  wire Gpzow6;  // ../RTL/cortexm0ds_logic.v(1324)
  wire Gq4ju6;  // ../RTL/cortexm0ds_logic.v(848)
  wire Gq5iu6;  // ../RTL/cortexm0ds_logic.v(380)
  wire Gq5pw6;  // ../RTL/cortexm0ds_logic.v(1404)
  wire Gq6ow6;  // ../RTL/cortexm0ds_logic.v(936)
  wire Gqciu6;  // ../RTL/cortexm0ds_logic.v(474)
  wire Gqcpw6;  // ../RTL/cortexm0ds_logic.v(1498)
  wire Gqdow6;  // ../RTL/cortexm0ds_logic.v(1030)
  wire Gqjiu6;  // ../RTL/cortexm0ds_logic.v(567)
  wire Gqkhu6;  // ../RTL/cortexm0ds_logic.v(137)
  wire Gqkow6;  // ../RTL/cortexm0ds_logic.v(1124)
  wire Gqqiu6;  // ../RTL/cortexm0ds_logic.v(661)
  wire Gqrhu6;  // ../RTL/cortexm0ds_logic.v(193)
  wire Gqrow6;  // ../RTL/cortexm0ds_logic.v(1217)
  wire Gqxiu6;  // ../RTL/cortexm0ds_logic.v(754)
  wire Gqyhu6;  // ../RTL/cortexm0ds_logic.v(286)
  wire Gqyow6;  // ../RTL/cortexm0ds_logic.v(1311)
  wire Gr2qw6;  // ../RTL/cortexm0ds_logic.v(1622)
  wire Gr3ju6;  // ../RTL/cortexm0ds_logic.v(835)
  wire Gr4iu6;  // ../RTL/cortexm0ds_logic.v(367)
  wire Gr4pw6;  // ../RTL/cortexm0ds_logic.v(1391)
  wire Gr6ax6;  // ../RTL/cortexm0ds_logic.v(1625)
  wire Graju6;  // ../RTL/cortexm0ds_logic.v(929)
  wire Grbiu6;  // ../RTL/cortexm0ds_logic.v(461)
  wire Grbpw6;  // ../RTL/cortexm0ds_logic.v(1485)
  wire Grcow6;  // ../RTL/cortexm0ds_logic.v(1017)
  wire Griiu6;  // ../RTL/cortexm0ds_logic.v(554)
  wire Grjow6;  // ../RTL/cortexm0ds_logic.v(1111)
  wire Grpiu6;  // ../RTL/cortexm0ds_logic.v(648)
  wire Grqhu6;  // ../RTL/cortexm0ds_logic.v(180)
  wire Grqow6;  // ../RTL/cortexm0ds_logic.v(1204)
  wire Grwiu6;  // ../RTL/cortexm0ds_logic.v(741)
  wire Grxhu6;  // ../RTL/cortexm0ds_logic.v(273)
  wire Grxow6;  // ../RTL/cortexm0ds_logic.v(1298)
  wire Gs2ju6;  // ../RTL/cortexm0ds_logic.v(822)
  wire Gs3iu6;  // ../RTL/cortexm0ds_logic.v(354)
  wire Gs3pw6;  // ../RTL/cortexm0ds_logic.v(1378)
  wire Gs9ju6;  // ../RTL/cortexm0ds_logic.v(916)
  wire Gsaiu6;  // ../RTL/cortexm0ds_logic.v(448)
  wire Gsapw6;  // ../RTL/cortexm0ds_logic.v(1472)
  wire Gsbow6;  // ../RTL/cortexm0ds_logic.v(1004)
  wire Gshiu6;  // ../RTL/cortexm0ds_logic.v(541)
  wire Gsiow6;  // ../RTL/cortexm0ds_logic.v(1098)
  wire Gsjhu6;  // ../RTL/cortexm0ds_logic.v(135)
  wire Gsoiu6;  // ../RTL/cortexm0ds_logic.v(635)
  wire Gsphu6;  // ../RTL/cortexm0ds_logic.v(167)
  wire Gspow6;  // ../RTL/cortexm0ds_logic.v(1191)
  wire Gsviu6;  // ../RTL/cortexm0ds_logic.v(728)
  wire Gswhu6;  // ../RTL/cortexm0ds_logic.v(260)
  wire Gswow6;  // ../RTL/cortexm0ds_logic.v(1285)
  wire Gt1ju6;  // ../RTL/cortexm0ds_logic.v(809)
  wire Gt2iu6;  // ../RTL/cortexm0ds_logic.v(341)
  wire Gt2pw6;  // ../RTL/cortexm0ds_logic.v(1365)
  wire Gt6ax6;  // ../RTL/cortexm0ds_logic.v(1625)
  wire Gt8ju6;  // ../RTL/cortexm0ds_logic.v(903)
  wire Gt9iu6;  // ../RTL/cortexm0ds_logic.v(435)
  wire Gt9pw6;  // ../RTL/cortexm0ds_logic.v(1459)
  wire Gtaow6;  // ../RTL/cortexm0ds_logic.v(991)
  wire Gtgiu6;  // ../RTL/cortexm0ds_logic.v(528)
  wire Gthow6;  // ../RTL/cortexm0ds_logic.v(1085)
  wire Gtniu6;  // ../RTL/cortexm0ds_logic.v(622)
  wire Gtoax6;  // ../RTL/cortexm0ds_logic.v(1659)
  wire Gtohu6;  // ../RTL/cortexm0ds_logic.v(154)
  wire Gtoow6;  // ../RTL/cortexm0ds_logic.v(1178)
  wire Gtuiu6;  // ../RTL/cortexm0ds_logic.v(715)
  wire Gtvhu6;  // ../RTL/cortexm0ds_logic.v(247)
  wire Gtvow6;  // ../RTL/cortexm0ds_logic.v(1272)
  wire Gu0ju6;  // ../RTL/cortexm0ds_logic.v(796)
  wire Gu1iu6;  // ../RTL/cortexm0ds_logic.v(328)
  wire Gu1pw6;  // ../RTL/cortexm0ds_logic.v(1352)
  wire Gu7ju6;  // ../RTL/cortexm0ds_logic.v(890)
  wire Gu8iu6;  // ../RTL/cortexm0ds_logic.v(422)
  wire Gu8pw6;  // ../RTL/cortexm0ds_logic.v(1446)
  wire Gu9ow6;  // ../RTL/cortexm0ds_logic.v(978)
  wire Gufiu6;  // ../RTL/cortexm0ds_logic.v(515)
  wire Gugow6;  // ../RTL/cortexm0ds_logic.v(1072)
  wire Guihu6;  // ../RTL/cortexm0ds_logic.v(132)
  wire Gumiu6;  // ../RTL/cortexm0ds_logic.v(609)
  wire Gunow6;  // ../RTL/cortexm0ds_logic.v(1165)
  wire Gutiu6;  // ../RTL/cortexm0ds_logic.v(702)
  wire Guuhu6;  // ../RTL/cortexm0ds_logic.v(234)
  wire Guuow6;  // ../RTL/cortexm0ds_logic.v(1259)
  wire Gv0iu6;  // ../RTL/cortexm0ds_logic.v(315)
  wire Gv0pw6;  // ../RTL/cortexm0ds_logic.v(1339)
  wire Gv1bx6;  // ../RTL/cortexm0ds_logic.v(1683)
  wire Gv1qw6;  // ../RTL/cortexm0ds_logic.v(1620)
  wire Gv6ax6;  // ../RTL/cortexm0ds_logic.v(1625)
  wire Gv6ju6;  // ../RTL/cortexm0ds_logic.v(877)
  wire Gv7iu6;  // ../RTL/cortexm0ds_logic.v(409)
  wire Gv7pw6;  // ../RTL/cortexm0ds_logic.v(1433)
  wire Gv8ow6;  // ../RTL/cortexm0ds_logic.v(965)
  wire Gveiu6;  // ../RTL/cortexm0ds_logic.v(502)
  wire Gvfow6;  // ../RTL/cortexm0ds_logic.v(1059)
  wire Gvliu6;  // ../RTL/cortexm0ds_logic.v(596)
  wire Gvmow6;  // ../RTL/cortexm0ds_logic.v(1152)
  wire Gvmpw6;  // ../RTL/cortexm0ds_logic.v(1593)
  wire Gvsiu6;  // ../RTL/cortexm0ds_logic.v(689)
  wire Gvthu6;  // ../RTL/cortexm0ds_logic.v(221)
  wire Gvtow6;  // ../RTL/cortexm0ds_logic.v(1246)
  wire Gvziu6;  // ../RTL/cortexm0ds_logic.v(783)
  wire Gw5ju6;  // ../RTL/cortexm0ds_logic.v(864)
  wire Gw6bx6;  // ../RTL/cortexm0ds_logic.v(1691)
  wire Gw6iu6;  // ../RTL/cortexm0ds_logic.v(396)
  wire Gw6pw6;  // ../RTL/cortexm0ds_logic.v(1420)
  wire Gw7ow6;  // ../RTL/cortexm0ds_logic.v(952)
  wire Gwdiu6;  // ../RTL/cortexm0ds_logic.v(489)
  wire Gwdpw6;  // ../RTL/cortexm0ds_logic.v(1514)
  wire Gweow6;  // ../RTL/cortexm0ds_logic.v(1046)
  wire Gwhhu6;  // ../RTL/cortexm0ds_logic.v(129)
  wire Gwkiu6;  // ../RTL/cortexm0ds_logic.v(583)
  wire Gwlow6;  // ../RTL/cortexm0ds_logic.v(1139)
  wire Gwnhu6;  // ../RTL/cortexm0ds_logic.v(146)
  wire Gwriu6;  // ../RTL/cortexm0ds_logic.v(676)
  wire Gwshu6;  // ../RTL/cortexm0ds_logic.v(208)
  wire Gwsow6;  // ../RTL/cortexm0ds_logic.v(1233)
  wire Gwwpw6;  // ../RTL/cortexm0ds_logic.v(1611)
  wire Gwxpw6;  // ../RTL/cortexm0ds_logic.v(1613)
  wire Gwyiu6;  // ../RTL/cortexm0ds_logic.v(770)
  wire Gwzhu6;  // ../RTL/cortexm0ds_logic.v(302)
  wire Gwzow6;  // ../RTL/cortexm0ds_logic.v(1326)
  wire Gx2bx6;  // ../RTL/cortexm0ds_logic.v(1684)
  wire Gx4ju6;  // ../RTL/cortexm0ds_logic.v(851)
  wire Gx5iu6;  // ../RTL/cortexm0ds_logic.v(383)
  wire Gx5pw6;  // ../RTL/cortexm0ds_logic.v(1407)
  wire Gx6ax6;  // ../RTL/cortexm0ds_logic.v(1625)
  wire Gx6ow6;  // ../RTL/cortexm0ds_logic.v(939)
  wire Gxciu6;  // ../RTL/cortexm0ds_logic.v(476)
  wire Gxcpw6;  // ../RTL/cortexm0ds_logic.v(1501)
  wire Gxdow6;  // ../RTL/cortexm0ds_logic.v(1033)
  wire Gxjiu6;  // ../RTL/cortexm0ds_logic.v(570)
  wire Gxkow6;  // ../RTL/cortexm0ds_logic.v(1126)
  wire Gxmpw6;  // ../RTL/cortexm0ds_logic.v(1593)
  wire Gxqiu6;  // ../RTL/cortexm0ds_logic.v(663)
  wire Gxrhu6;  // ../RTL/cortexm0ds_logic.v(195)
  wire Gxrow6;  // ../RTL/cortexm0ds_logic.v(1220)
  wire Gxxiu6;  // ../RTL/cortexm0ds_logic.v(757)
  wire Gxyhu6;  // ../RTL/cortexm0ds_logic.v(289)
  wire Gxyow6;  // ../RTL/cortexm0ds_logic.v(1313)
  wire Gy3ju6;  // ../RTL/cortexm0ds_logic.v(838)
  wire Gy4iu6;  // ../RTL/cortexm0ds_logic.v(370)
  wire Gy4pw6;  // ../RTL/cortexm0ds_logic.v(1394)
  wire Gybiu6;  // ../RTL/cortexm0ds_logic.v(463)
  wire Gybpw6;  // ../RTL/cortexm0ds_logic.v(1488)
  wire Gycow6;  // ../RTL/cortexm0ds_logic.v(1020)
  wire Gyiiu6;  // ../RTL/cortexm0ds_logic.v(557)
  wire Gyjow6;  // ../RTL/cortexm0ds_logic.v(1113)
  wire Gylpw6;  // ../RTL/cortexm0ds_logic.v(1591)
  wire Gypiu6;  // ../RTL/cortexm0ds_logic.v(650)
  wire Gyqhu6;  // ../RTL/cortexm0ds_logic.v(182)
  wire Gyqow6;  // ../RTL/cortexm0ds_logic.v(1207)
  wire Gywiu6;  // ../RTL/cortexm0ds_logic.v(744)
  wire Gyxhu6;  // ../RTL/cortexm0ds_logic.v(276)
  wire Gyxow6;  // ../RTL/cortexm0ds_logic.v(1300)
  wire Gyxpw6;  // ../RTL/cortexm0ds_logic.v(1613)
  wire Gz2ju6;  // ../RTL/cortexm0ds_logic.v(825)
  wire Gz3iu6;  // ../RTL/cortexm0ds_logic.v(357)
  wire Gz3pw6;  // ../RTL/cortexm0ds_logic.v(1381)
  wire Gz6ax6;  // ../RTL/cortexm0ds_logic.v(1625)
  wire Gz9ju6;  // ../RTL/cortexm0ds_logic.v(918)
  wire Gzaiu6;  // ../RTL/cortexm0ds_logic.v(450)
  wire Gzapw6;  // ../RTL/cortexm0ds_logic.v(1475)
  wire Gzbow6;  // ../RTL/cortexm0ds_logic.v(1007)
  wire Gzeax6;  // ../RTL/cortexm0ds_logic.v(1641)
  wire Gzhiu6;  // ../RTL/cortexm0ds_logic.v(544)
  wire Gziow6;  // ../RTL/cortexm0ds_logic.v(1100)
  wire Gzoiu6;  // ../RTL/cortexm0ds_logic.v(637)
  wire Gzphu6;  // ../RTL/cortexm0ds_logic.v(169)
  wire Gzpow6;  // ../RTL/cortexm0ds_logic.v(1194)
  wire Gzviu6;  // ../RTL/cortexm0ds_logic.v(731)
  wire Gzwhu6;  // ../RTL/cortexm0ds_logic.v(263)
  wire Gzwow6;  // ../RTL/cortexm0ds_logic.v(1287)
  wire H00iu6;  // ../RTL/cortexm0ds_logic.v(303)
  wire H00pw6;  // ../RTL/cortexm0ds_logic.v(1328)
  wire H06ju6;  // ../RTL/cortexm0ds_logic.v(865)
  wire H07iu6;  // ../RTL/cortexm0ds_logic.v(397)
  wire H07pw6;  // ../RTL/cortexm0ds_logic.v(1421)
  wire H08ow6;  // ../RTL/cortexm0ds_logic.v(953)
  wire H0ebx6;  // ../RTL/cortexm0ds_logic.v(1705)
  wire H0eiu6;  // ../RTL/cortexm0ds_logic.v(491)
  wire H0epw6;  // ../RTL/cortexm0ds_logic.v(1515)
  wire H0fow6;  // ../RTL/cortexm0ds_logic.v(1047)
  wire H0liu6;  // ../RTL/cortexm0ds_logic.v(584)
  wire H0mow6;  // ../RTL/cortexm0ds_logic.v(1141)
  wire H0siu6;  // ../RTL/cortexm0ds_logic.v(678)
  wire H0thu6;  // ../RTL/cortexm0ds_logic.v(210)
  wire H0tow6;  // ../RTL/cortexm0ds_logic.v(1234)
  wire H0ziu6;  // ../RTL/cortexm0ds_logic.v(771)
  wire H15ju6;  // ../RTL/cortexm0ds_logic.v(852)
  wire H16iu6;  // ../RTL/cortexm0ds_logic.v(384)
  wire H16pw6;  // ../RTL/cortexm0ds_logic.v(1408)
  wire H17ow6;  // ../RTL/cortexm0ds_logic.v(940)
  wire H1diu6;  // ../RTL/cortexm0ds_logic.v(478)
  wire H1dpw6;  // ../RTL/cortexm0ds_logic.v(1502)
  wire H1eow6;  // ../RTL/cortexm0ds_logic.v(1034)
  wire H1kiu6;  // ../RTL/cortexm0ds_logic.v(571)
  wire H1low6;  // ../RTL/cortexm0ds_logic.v(1128)
  wire H1riu6;  // ../RTL/cortexm0ds_logic.v(665)
  wire H1shu6;  // ../RTL/cortexm0ds_logic.v(197)
  wire H1sow6;  // ../RTL/cortexm0ds_logic.v(1221)
  wire H1yiu6;  // ../RTL/cortexm0ds_logic.v(758)
  wire H1zhu6;  // ../RTL/cortexm0ds_logic.v(290)
  wire H1zow6;  // ../RTL/cortexm0ds_logic.v(1315)
  wire H24ju6;  // ../RTL/cortexm0ds_logic.v(839)
  wire H25iu6;  // ../RTL/cortexm0ds_logic.v(371)
  wire H25pw6;  // ../RTL/cortexm0ds_logic.v(1395)
  wire H2ciu6;  // ../RTL/cortexm0ds_logic.v(465)
  wire H2cpw6;  // ../RTL/cortexm0ds_logic.v(1489)
  wire H2dow6;  // ../RTL/cortexm0ds_logic.v(1021)
  wire H2hhu6;  // ../RTL/cortexm0ds_logic.v(127)
  wire H2jiu6;  // ../RTL/cortexm0ds_logic.v(558)
  wire H2kow6;  // ../RTL/cortexm0ds_logic.v(1115)
  wire H2qiu6;  // ../RTL/cortexm0ds_logic.v(652)
  wire H2rhu6;  // ../RTL/cortexm0ds_logic.v(184)
  wire H2row6;  // ../RTL/cortexm0ds_logic.v(1208)
  wire H2xiu6;  // ../RTL/cortexm0ds_logic.v(745)
  wire H2yhu6;  // ../RTL/cortexm0ds_logic.v(277)
  wire H2yow6;  // ../RTL/cortexm0ds_logic.v(1302)
  wire H33ju6;  // ../RTL/cortexm0ds_logic.v(826)
  wire H34iu6;  // ../RTL/cortexm0ds_logic.v(358)
  wire H34pw6;  // ../RTL/cortexm0ds_logic.v(1382)
  wire H3aju6;  // ../RTL/cortexm0ds_logic.v(920)
  wire H3biu6;  // ../RTL/cortexm0ds_logic.v(452)
  wire H3bpw6;  // ../RTL/cortexm0ds_logic.v(1476)
  wire H3cow6;  // ../RTL/cortexm0ds_logic.v(1008)
  wire H3iiu6;  // ../RTL/cortexm0ds_logic.v(545)
  wire H3jow6;  // ../RTL/cortexm0ds_logic.v(1102)
  wire H3lpw6;  // ../RTL/cortexm0ds_logic.v(1590)
  wire H3piu6;  // ../RTL/cortexm0ds_logic.v(639)
  wire H3qhu6;  // ../RTL/cortexm0ds_logic.v(171)
  wire H3qow6;  // ../RTL/cortexm0ds_logic.v(1195)
  wire H3wiu6;  // ../RTL/cortexm0ds_logic.v(732)
  wire H3xhu6;  // ../RTL/cortexm0ds_logic.v(264)
  wire H3xow6;  // ../RTL/cortexm0ds_logic.v(1289)
  wire H42ju6;  // ../RTL/cortexm0ds_logic.v(813)
  wire H43iu6;  // ../RTL/cortexm0ds_logic.v(345)
  wire H43pw6;  // ../RTL/cortexm0ds_logic.v(1369)
  wire H49ju6;  // ../RTL/cortexm0ds_logic.v(907)
  wire H4aiu6;  // ../RTL/cortexm0ds_logic.v(439)
  wire H4apw6;  // ../RTL/cortexm0ds_logic.v(1463)
  wire H4bax6;  // ../RTL/cortexm0ds_logic.v(1633)
  wire H4bow6;  // ../RTL/cortexm0ds_logic.v(995)
  wire H4ghu6;  // ../RTL/cortexm0ds_logic.v(125)
  wire H4hiu6;  // ../RTL/cortexm0ds_logic.v(532)
  wire H4iow6;  // ../RTL/cortexm0ds_logic.v(1089)
  wire H4oiu6;  // ../RTL/cortexm0ds_logic.v(626)
  wire H4phu6;  // ../RTL/cortexm0ds_logic.v(158)
  wire H4pow6;  // ../RTL/cortexm0ds_logic.v(1182)
  wire H4viu6;  // ../RTL/cortexm0ds_logic.v(719)
  wire H4whu6;  // ../RTL/cortexm0ds_logic.v(251)
  wire H4wow6;  // ../RTL/cortexm0ds_logic.v(1276)
  wire H4ypw6;  // ../RTL/cortexm0ds_logic.v(1613)
  wire H4zax6;  // ../RTL/cortexm0ds_logic.v(1678)
  wire H51ju6;  // ../RTL/cortexm0ds_logic.v(800)
  wire H52iu6;  // ../RTL/cortexm0ds_logic.v(332)
  wire H52pw6;  // ../RTL/cortexm0ds_logic.v(1356)
  wire H58ju6;  // ../RTL/cortexm0ds_logic.v(894)
  wire H59iu6;  // ../RTL/cortexm0ds_logic.v(426)
  wire H59pw6;  // ../RTL/cortexm0ds_logic.v(1450)
  wire H5aow6;  // ../RTL/cortexm0ds_logic.v(982)
  wire H5giu6;  // ../RTL/cortexm0ds_logic.v(519)
  wire H5how6;  // ../RTL/cortexm0ds_logic.v(1076)
  wire H5niu6;  // ../RTL/cortexm0ds_logic.v(613)
  wire H5oow6;  // ../RTL/cortexm0ds_logic.v(1169)
  wire H5uiu6;  // ../RTL/cortexm0ds_logic.v(706)
  wire H5vhu6;  // ../RTL/cortexm0ds_logic.v(238)
  wire H5vow6;  // ../RTL/cortexm0ds_logic.v(1263)
  wire H60ju6;  // ../RTL/cortexm0ds_logic.v(787)
  wire H61iu6;  // ../RTL/cortexm0ds_logic.v(319)
  wire H61pw6;  // ../RTL/cortexm0ds_logic.v(1343)
  wire H67ju6;  // ../RTL/cortexm0ds_logic.v(881)
  wire H68iu6;  // ../RTL/cortexm0ds_logic.v(413)
  wire H68pw6;  // ../RTL/cortexm0ds_logic.v(1437)
  wire H69ow6;  // ../RTL/cortexm0ds_logic.v(969)
  wire H6fiu6;  // ../RTL/cortexm0ds_logic.v(506)
  wire H6ghu6;  // ../RTL/cortexm0ds_logic.v(126)
  wire H6gow6;  // ../RTL/cortexm0ds_logic.v(1063)
  wire H6miu6;  // ../RTL/cortexm0ds_logic.v(600)
  wire H6now6;  // ../RTL/cortexm0ds_logic.v(1156)
  wire H6tiu6;  // ../RTL/cortexm0ds_logic.v(693)
  wire H6uhu6;  // ../RTL/cortexm0ds_logic.v(225)
  wire H6uow6;  // ../RTL/cortexm0ds_logic.v(1250)
  wire H70iu6;  // ../RTL/cortexm0ds_logic.v(306)
  wire H70pw6;  // ../RTL/cortexm0ds_logic.v(1330)
  wire H76ju6;  // ../RTL/cortexm0ds_logic.v(868)
  wire H77iu6;  // ../RTL/cortexm0ds_logic.v(400)
  wire H77pw6;  // ../RTL/cortexm0ds_logic.v(1424)
  wire H78ow6;  // ../RTL/cortexm0ds_logic.v(956)
  wire H7eiu6;  // ../RTL/cortexm0ds_logic.v(493)
  wire H7fow6;  // ../RTL/cortexm0ds_logic.v(1050)
  wire H7hbx6;  // ../RTL/cortexm0ds_logic.v(1710)
  wire H7liu6;  // ../RTL/cortexm0ds_logic.v(587)
  wire H7mow6;  // ../RTL/cortexm0ds_logic.v(1143)
  wire H7siu6;  // ../RTL/cortexm0ds_logic.v(680)
  wire H7thu6;  // ../RTL/cortexm0ds_logic.v(212)
  wire H7tow6;  // ../RTL/cortexm0ds_logic.v(1237)
  wire H7ziu6;  // ../RTL/cortexm0ds_logic.v(774)
  wire H85ju6;  // ../RTL/cortexm0ds_logic.v(855)
  wire H86iu6;  // ../RTL/cortexm0ds_logic.v(387)
  wire H86pw6;  // ../RTL/cortexm0ds_logic.v(1411)
  wire H87ow6;  // ../RTL/cortexm0ds_logic.v(943)
  wire H8diu6;  // ../RTL/cortexm0ds_logic.v(480)
  wire H8dpw6;  // ../RTL/cortexm0ds_logic.v(1505)
  wire H8eow6;  // ../RTL/cortexm0ds_logic.v(1037)
  wire H8gax6;  // ../RTL/cortexm0ds_logic.v(1643)
  wire H8kiu6;  // ../RTL/cortexm0ds_logic.v(574)
  wire H8low6;  // ../RTL/cortexm0ds_logic.v(1130)
  wire H8riu6;  // ../RTL/cortexm0ds_logic.v(667)
  wire H8shu6;  // ../RTL/cortexm0ds_logic.v(199)
  wire H8sow6;  // ../RTL/cortexm0ds_logic.v(1224)
  wire H8yiu6;  // ../RTL/cortexm0ds_logic.v(761)
  wire H8zhu6;  // ../RTL/cortexm0ds_logic.v(293)
  wire H8zow6;  // ../RTL/cortexm0ds_logic.v(1317)
  wire H94ju6;  // ../RTL/cortexm0ds_logic.v(842)
  wire H95iu6;  // ../RTL/cortexm0ds_logic.v(374)
  wire H95pw6;  // ../RTL/cortexm0ds_logic.v(1398)
  wire H96ow6;  // ../RTL/cortexm0ds_logic.v(930)
  wire H9ciu6;  // ../RTL/cortexm0ds_logic.v(467)
  wire H9cpw6;  // ../RTL/cortexm0ds_logic.v(1492)
  wire H9dow6;  // ../RTL/cortexm0ds_logic.v(1024)
  wire H9jiu6;  // ../RTL/cortexm0ds_logic.v(561)
  wire H9kow6;  // ../RTL/cortexm0ds_logic.v(1117)
  wire H9qiu6;  // ../RTL/cortexm0ds_logic.v(654)
  wire H9rhu6;  // ../RTL/cortexm0ds_logic.v(186)
  wire H9row6;  // ../RTL/cortexm0ds_logic.v(1211)
  wire H9xiu6;  // ../RTL/cortexm0ds_logic.v(748)
  wire H9yhu6;  // ../RTL/cortexm0ds_logic.v(280)
  wire H9yow6;  // ../RTL/cortexm0ds_logic.v(1304)
  wire Ha3ju6;  // ../RTL/cortexm0ds_logic.v(829)
  wire Ha4iu6;  // ../RTL/cortexm0ds_logic.v(361)
  wire Ha4pw6;  // ../RTL/cortexm0ds_logic.v(1385)
  wire Haaju6;  // ../RTL/cortexm0ds_logic.v(922)
  wire Habiu6;  // ../RTL/cortexm0ds_logic.v(454)
  wire Habpw6;  // ../RTL/cortexm0ds_logic.v(1479)
  wire Hacow6;  // ../RTL/cortexm0ds_logic.v(1011)
  wire Haiiu6;  // ../RTL/cortexm0ds_logic.v(548)
  wire Hajow6;  // ../RTL/cortexm0ds_logic.v(1104)
  wire Halax6;  // ../RTL/cortexm0ds_logic.v(1653)
  wire Hapiu6;  // ../RTL/cortexm0ds_logic.v(641)
  wire Haqhu6;  // ../RTL/cortexm0ds_logic.v(173)
  wire Haqow6;  // ../RTL/cortexm0ds_logic.v(1198)
  wire Hawiu6;  // ../RTL/cortexm0ds_logic.v(735)
  wire Haxhu6;  // ../RTL/cortexm0ds_logic.v(267)
  wire Haxow6;  // ../RTL/cortexm0ds_logic.v(1291)
  wire Hb2ju6;  // ../RTL/cortexm0ds_logic.v(816)
  wire Hb3iu6;  // ../RTL/cortexm0ds_logic.v(348)
  wire Hb3pw6;  // ../RTL/cortexm0ds_logic.v(1372)
  wire Hb9ju6;  // ../RTL/cortexm0ds_logic.v(909)
  wire Hbaiu6;  // ../RTL/cortexm0ds_logic.v(441)
  wire Hbapw6;  // ../RTL/cortexm0ds_logic.v(1466)
  wire Hbbow6;  // ../RTL/cortexm0ds_logic.v(998)
  wire Hbgbx6;  // ../RTL/cortexm0ds_logic.v(1709)
  wire Hbhhu6;  // ../RTL/cortexm0ds_logic.v(128)
  wire Hbhiu6;  // ../RTL/cortexm0ds_logic.v(535)
  wire Hbiow6;  // ../RTL/cortexm0ds_logic.v(1091)
  wire Hboiu6;  // ../RTL/cortexm0ds_logic.v(628)
  wire Hbphu6;  // ../RTL/cortexm0ds_logic.v(160)
  wire Hbpow6;  // ../RTL/cortexm0ds_logic.v(1185)
  wire Hbviu6;  // ../RTL/cortexm0ds_logic.v(722)
  wire Hbwhu6;  // ../RTL/cortexm0ds_logic.v(254)
  wire Hbwow6;  // ../RTL/cortexm0ds_logic.v(1278)
  wire Hc1ju6;  // ../RTL/cortexm0ds_logic.v(803)
  wire Hc2iu6;  // ../RTL/cortexm0ds_logic.v(335)
  wire Hc2pw6;  // ../RTL/cortexm0ds_logic.v(1359)
  wire Hc8ju6;  // ../RTL/cortexm0ds_logic.v(896)
  wire Hc9iu6;  // ../RTL/cortexm0ds_logic.v(428)
  wire Hc9pw6;  // ../RTL/cortexm0ds_logic.v(1453)
  wire Hcaow6;  // ../RTL/cortexm0ds_logic.v(985)
  wire Hcgiu6;  // ../RTL/cortexm0ds_logic.v(522)
  wire Hchow6;  // ../RTL/cortexm0ds_logic.v(1078)
  wire Hcniu6;  // ../RTL/cortexm0ds_logic.v(615)
  wire Hcohu6;  // ../RTL/cortexm0ds_logic.v(147)
  wire Hcoow6;  // ../RTL/cortexm0ds_logic.v(1172)
  wire Hcuiu6;  // ../RTL/cortexm0ds_logic.v(709)
  wire Hcvhu6;  // ../RTL/cortexm0ds_logic.v(241)
  wire Hcvow6;  // ../RTL/cortexm0ds_logic.v(1265)
  wire Hd0ju6;  // ../RTL/cortexm0ds_logic.v(790)
  wire Hd1iu6;  // ../RTL/cortexm0ds_logic.v(322)
  wire Hd1pw6;  // ../RTL/cortexm0ds_logic.v(1346)
  wire Hd7ju6;  // ../RTL/cortexm0ds_logic.v(883)
  wire Hd8iu6;  // ../RTL/cortexm0ds_logic.v(415)
  wire Hd8pw6;  // ../RTL/cortexm0ds_logic.v(1440)
  wire Hd9ow6;  // ../RTL/cortexm0ds_logic.v(972)
  wire Hdbax6;  // ../RTL/cortexm0ds_logic.v(1634)
  wire Hdfax6;  // ../RTL/cortexm0ds_logic.v(1642)
  wire Hdfiu6;  // ../RTL/cortexm0ds_logic.v(509)
  wire Hdgow6;  // ../RTL/cortexm0ds_logic.v(1065)
  wire Hdmiu6;  // ../RTL/cortexm0ds_logic.v(602)
  wire Hdnow6;  // ../RTL/cortexm0ds_logic.v(1159)
  wire Hdtiu6;  // ../RTL/cortexm0ds_logic.v(696)
  wire Hduhu6;  // ../RTL/cortexm0ds_logic.v(228)
  wire Hduow6;  // ../RTL/cortexm0ds_logic.v(1252)
  wire He0iu6;  // ../RTL/cortexm0ds_logic.v(309)
  wire He0pw6;  // ../RTL/cortexm0ds_logic.v(1333)
  wire He6ju6;  // ../RTL/cortexm0ds_logic.v(870)
  wire He7iu6;  // ../RTL/cortexm0ds_logic.v(402)
  wire He7pw6;  // ../RTL/cortexm0ds_logic.v(1427)
  wire He8ow6;  // ../RTL/cortexm0ds_logic.v(959)
  wire Heaax6;  // ../RTL/cortexm0ds_logic.v(1632)
  wire Heeiu6;  // ../RTL/cortexm0ds_logic.v(496)
  wire Hefow6;  // ../RTL/cortexm0ds_logic.v(1052)
  wire Heliu6;  // ../RTL/cortexm0ds_logic.v(589)
  wire Hemow6;  // ../RTL/cortexm0ds_logic.v(1146)
  wire Hesiu6;  // ../RTL/cortexm0ds_logic.v(683)
  wire Hethu6;  // ../RTL/cortexm0ds_logic.v(215)
  wire Hetow6;  // ../RTL/cortexm0ds_logic.v(1239)
  wire Heziu6;  // ../RTL/cortexm0ds_logic.v(777)
  wire Hf0bx6;  // ../RTL/cortexm0ds_logic.v(1680)
  wire Hf5ju6;  // ../RTL/cortexm0ds_logic.v(857)
  wire Hf6iu6;  // ../RTL/cortexm0ds_logic.v(389)
  wire Hf6pw6;  // ../RTL/cortexm0ds_logic.v(1414)
  wire Hf7ow6;  // ../RTL/cortexm0ds_logic.v(946)
  wire Hfdiu6;  // ../RTL/cortexm0ds_logic.v(483)
  wire Hfdpw6;  // ../RTL/cortexm0ds_logic.v(1507)
  wire Hfeow6;  // ../RTL/cortexm0ds_logic.v(1039)
  wire Hfkiu6;  // ../RTL/cortexm0ds_logic.v(576)
  wire Hflow6;  // ../RTL/cortexm0ds_logic.v(1133)
  wire Hfriu6;  // ../RTL/cortexm0ds_logic.v(670)
  wire Hfshu6;  // ../RTL/cortexm0ds_logic.v(202)
  wire Hfsow6;  // ../RTL/cortexm0ds_logic.v(1226)
  wire Hfyiu6;  // ../RTL/cortexm0ds_logic.v(764)
  wire Hfzhu6;  // ../RTL/cortexm0ds_logic.v(296)
  wire Hfzow6;  // ../RTL/cortexm0ds_logic.v(1320)
  wire Hg3bx6;  // ../RTL/cortexm0ds_logic.v(1685)
  wire Hg4ju6;  // ../RTL/cortexm0ds_logic.v(844)
  wire Hg5iu6;  // ../RTL/cortexm0ds_logic.v(376)
  wire Hg5pw6;  // ../RTL/cortexm0ds_logic.v(1401)
  wire Hg6ow6;  // ../RTL/cortexm0ds_logic.v(933)
  wire Hg7ax6;  // ../RTL/cortexm0ds_logic.v(1626)
  wire Hgciu6;  // ../RTL/cortexm0ds_logic.v(470)
  wire Hgcpw6;  // ../RTL/cortexm0ds_logic.v(1494)
  wire Hgdow6;  // ../RTL/cortexm0ds_logic.v(1026)
  wire Hgjiu6;  // ../RTL/cortexm0ds_logic.v(563)
  wire Hgkow6;  // ../RTL/cortexm0ds_logic.v(1120)
  wire Hgqiu6;  // ../RTL/cortexm0ds_logic.v(657)
  wire Hgrhu6;  // ../RTL/cortexm0ds_logic.v(189)
  wire Hgrow6;  // ../RTL/cortexm0ds_logic.v(1213)
  wire Hgrpw6;  // ../RTL/cortexm0ds_logic.v(1601)
  wire Hgxiu6;  // ../RTL/cortexm0ds_logic.v(751)
  wire Hgyhu6;  // ../RTL/cortexm0ds_logic.v(283)
  wire Hgyow6;  // ../RTL/cortexm0ds_logic.v(1307)
  wire Hh3ju6;  // ../RTL/cortexm0ds_logic.v(831)
  wire Hh4iu6;  // ../RTL/cortexm0ds_logic.v(363)
  wire Hh4pw6;  // ../RTL/cortexm0ds_logic.v(1388)
  wire Hhaju6;  // ../RTL/cortexm0ds_logic.v(925)
  wire Hhbiu6;  // ../RTL/cortexm0ds_logic.v(457)
  wire Hhbpw6;  // ../RTL/cortexm0ds_logic.v(1481)
  wire Hhcow6;  // ../RTL/cortexm0ds_logic.v(1013)
  wire Hhiiu6;  // ../RTL/cortexm0ds_logic.v(550)
  wire Hhjow6;  // ../RTL/cortexm0ds_logic.v(1107)
  wire Hhpiu6;  // ../RTL/cortexm0ds_logic.v(644)
  wire Hhqhu6;  // ../RTL/cortexm0ds_logic.v(176)
  wire Hhqow6;  // ../RTL/cortexm0ds_logic.v(1200)
  wire Hhvpw6;  // ../RTL/cortexm0ds_logic.v(1609)
  wire Hhwiu6;  // ../RTL/cortexm0ds_logic.v(738)
  wire Hhxhu6;  // ../RTL/cortexm0ds_logic.v(270)
  wire Hhxow6;  // ../RTL/cortexm0ds_logic.v(1294)
  wire Hi2ju6;  // ../RTL/cortexm0ds_logic.v(818)
  wire Hi3iu6;  // ../RTL/cortexm0ds_logic.v(350)
  wire Hi3pw6;  // ../RTL/cortexm0ds_logic.v(1375)
  wire Hi9bx6;  // ../RTL/cortexm0ds_logic.v(1696)
  wire Hi9ju6;  // ../RTL/cortexm0ds_logic.v(912)
  wire Hiaiu6;  // ../RTL/cortexm0ds_logic.v(444)
  wire Hiapw6;  // ../RTL/cortexm0ds_logic.v(1468)
  wire Hibow6;  // ../RTL/cortexm0ds_logic.v(1000)
  wire Hihiu6;  // ../RTL/cortexm0ds_logic.v(537)
  wire Hiiow6;  // ../RTL/cortexm0ds_logic.v(1094)
  wire Hioiu6;  // ../RTL/cortexm0ds_logic.v(631)
  wire Hiphu6;  // ../RTL/cortexm0ds_logic.v(163)
  wire Hipow6;  // ../RTL/cortexm0ds_logic.v(1187)
  wire Hirpw6;  // ../RTL/cortexm0ds_logic.v(1601)
  wire Hiviu6;  // ../RTL/cortexm0ds_logic.v(725)
  wire Hiwhu6;  // ../RTL/cortexm0ds_logic.v(257)
  wire Hiwow6;  // ../RTL/cortexm0ds_logic.v(1281)
  wire Hj1ju6;  // ../RTL/cortexm0ds_logic.v(805)
  wire Hj2iu6;  // ../RTL/cortexm0ds_logic.v(337)
  wire Hj2pw6;  // ../RTL/cortexm0ds_logic.v(1362)
  wire Hj8ju6;  // ../RTL/cortexm0ds_logic.v(899)
  wire Hj9iu6;  // ../RTL/cortexm0ds_logic.v(431)
  wire Hj9pw6;  // ../RTL/cortexm0ds_logic.v(1455)
  wire Hjaow6;  // ../RTL/cortexm0ds_logic.v(987)
  wire Hjgax6;  // ../RTL/cortexm0ds_logic.v(1644)
  wire Hjgiu6;  // ../RTL/cortexm0ds_logic.v(524)
  wire Hjhow6;  // ../RTL/cortexm0ds_logic.v(1081)
  wire Hjniu6;  // ../RTL/cortexm0ds_logic.v(618)
  wire Hjohu6;  // ../RTL/cortexm0ds_logic.v(150)
  wire Hjoow6;  // ../RTL/cortexm0ds_logic.v(1174)
  wire Hjuiu6;  // ../RTL/cortexm0ds_logic.v(712)
  wire Hjvhu6;  // ../RTL/cortexm0ds_logic.v(244)
  wire Hjvow6;  // ../RTL/cortexm0ds_logic.v(1268)
  wire Hk0ju6;  // ../RTL/cortexm0ds_logic.v(792)
  wire Hk1iu6;  // ../RTL/cortexm0ds_logic.v(324)
  wire Hk1pw6;  // ../RTL/cortexm0ds_logic.v(1349)
  wire Hk7ju6;  // ../RTL/cortexm0ds_logic.v(886)
  wire Hk8iu6;  // ../RTL/cortexm0ds_logic.v(418)
  wire Hk8pw6;  // ../RTL/cortexm0ds_logic.v(1442)
  wire Hk9ow6;  // ../RTL/cortexm0ds_logic.v(974)
  wire Hkfiu6;  // ../RTL/cortexm0ds_logic.v(511)
  wire Hkgow6;  // ../RTL/cortexm0ds_logic.v(1068)
  wire Hkmiu6;  // ../RTL/cortexm0ds_logic.v(605)
  wire Hknhu6;  // ../RTL/cortexm0ds_logic.v(145)
  wire Hknow6;  // ../RTL/cortexm0ds_logic.v(1161)
  wire Hktiu6;  // ../RTL/cortexm0ds_logic.v(699)
  wire Hkuhu6;  // ../RTL/cortexm0ds_logic.v(231)
  wire Hkuow6;  // ../RTL/cortexm0ds_logic.v(1255)
  wire Hkxpw6;  // ../RTL/cortexm0ds_logic.v(1612)
  wire Hl0iu6;  // ../RTL/cortexm0ds_logic.v(311)
  wire Hl0pw6;  // ../RTL/cortexm0ds_logic.v(1336)
  wire Hl6ju6;  // ../RTL/cortexm0ds_logic.v(873)
  wire Hl7iu6;  // ../RTL/cortexm0ds_logic.v(405)
  wire Hl7pw6;  // ../RTL/cortexm0ds_logic.v(1429)
  wire Hl8ow6;  // ../RTL/cortexm0ds_logic.v(961)
  wire Hlcax6;  // ../RTL/cortexm0ds_logic.v(1636)
  wire Hleiu6;  // ../RTL/cortexm0ds_logic.v(498)
  wire Hlfow6;  // ../RTL/cortexm0ds_logic.v(1055)
  wire Hlliu6;  // ../RTL/cortexm0ds_logic.v(592)
  wire Hlmow6;  // ../RTL/cortexm0ds_logic.v(1148)
  wire Hlsiu6;  // ../RTL/cortexm0ds_logic.v(686)
  wire Hlthu6;  // ../RTL/cortexm0ds_logic.v(218)
  wire Hltow6;  // ../RTL/cortexm0ds_logic.v(1242)
  wire Hlwpw6;  // ../RTL/cortexm0ds_logic.v(1611)
  wire Hlziu6;  // ../RTL/cortexm0ds_logic.v(779)
  wire Hm5ju6;  // ../RTL/cortexm0ds_logic.v(860)
  wire Hm6iu6;  // ../RTL/cortexm0ds_logic.v(392)
  wire Hm6pw6;  // ../RTL/cortexm0ds_logic.v(1416)
  wire Hm7ow6;  // ../RTL/cortexm0ds_logic.v(948)
  wire Hmbax6;  // ../RTL/cortexm0ds_logic.v(1634)
  wire Hmdiu6;  // ../RTL/cortexm0ds_logic.v(485)
  wire Hmdpw6;  // ../RTL/cortexm0ds_logic.v(1510)
  wire Hmeow6;  // ../RTL/cortexm0ds_logic.v(1042)
  wire Hmkiu6;  // ../RTL/cortexm0ds_logic.v(579)
  wire Hmlow6;  // ../RTL/cortexm0ds_logic.v(1135)
  wire Hmriu6;  // ../RTL/cortexm0ds_logic.v(673)
  wire Hmshu6;  // ../RTL/cortexm0ds_logic.v(205)
  wire Hmsow6;  // ../RTL/cortexm0ds_logic.v(1229)
  wire Hmxpw6;  // ../RTL/cortexm0ds_logic.v(1613)
  wire Hmyiu6;  // ../RTL/cortexm0ds_logic.v(766)
  wire Hmzhu6;  // ../RTL/cortexm0ds_logic.v(298)
  wire Hmzow6;  // ../RTL/cortexm0ds_logic.v(1323)
  wire Hn4ju6;  // ../RTL/cortexm0ds_logic.v(847)
  wire Hn5iu6;  // ../RTL/cortexm0ds_logic.v(379)
  wire Hn5pw6;  // ../RTL/cortexm0ds_logic.v(1403)
  wire Hn6ow6;  // ../RTL/cortexm0ds_logic.v(935)
  wire Hnciu6;  // ../RTL/cortexm0ds_logic.v(472)
  wire Hncpw6;  // ../RTL/cortexm0ds_logic.v(1497)
  wire Hndow6;  // ../RTL/cortexm0ds_logic.v(1029)
  wire Hnjiu6;  // ../RTL/cortexm0ds_logic.v(566)
  wire Hnkow6;  // ../RTL/cortexm0ds_logic.v(1122)
  wire Hnqiu6;  // ../RTL/cortexm0ds_logic.v(660)
  wire Hnrhu6;  // ../RTL/cortexm0ds_logic.v(192)
  wire Hnrow6;  // ../RTL/cortexm0ds_logic.v(1216)
  wire Hnxiu6;  // ../RTL/cortexm0ds_logic.v(753)
  wire Hnyhu6;  // ../RTL/cortexm0ds_logic.v(285)
  wire Hnyow6;  // ../RTL/cortexm0ds_logic.v(1310)
  wire Ho3ju6;  // ../RTL/cortexm0ds_logic.v(834)
  wire Ho4iu6;  // ../RTL/cortexm0ds_logic.v(366)
  wire Ho4pw6;  // ../RTL/cortexm0ds_logic.v(1390)
  wire Hoaju6;  // ../RTL/cortexm0ds_logic.v(927)
  wire Hobiu6;  // ../RTL/cortexm0ds_logic.v(459)
  wire Hobpw6;  // ../RTL/cortexm0ds_logic.v(1484)
  wire Hocow6;  // ../RTL/cortexm0ds_logic.v(1016)
  wire Hoiiu6;  // ../RTL/cortexm0ds_logic.v(553)
  wire Hojow6;  // ../RTL/cortexm0ds_logic.v(1109)
  wire Hopiu6;  // ../RTL/cortexm0ds_logic.v(647)
  wire Hoqhu6;  // ../RTL/cortexm0ds_logic.v(179)
  wire Hoqow6;  // ../RTL/cortexm0ds_logic.v(1203)
  wire Howiu6;  // ../RTL/cortexm0ds_logic.v(740)
  wire Hoxhu6;  // ../RTL/cortexm0ds_logic.v(272)
  wire Hoxow6;  // ../RTL/cortexm0ds_logic.v(1297)
  wire Hoxpw6;  // ../RTL/cortexm0ds_logic.v(1613)
  wire Hp2ju6;  // ../RTL/cortexm0ds_logic.v(821)
  wire Hp3iu6;  // ../RTL/cortexm0ds_logic.v(353)
  wire Hp3pw6;  // ../RTL/cortexm0ds_logic.v(1377)
  wire Hp9ju6;  // ../RTL/cortexm0ds_logic.v(914)
  wire Hpaiu6;  // ../RTL/cortexm0ds_logic.v(446)
  wire Hpapw6;  // ../RTL/cortexm0ds_logic.v(1471)
  wire Hpbbx6;  // ../RTL/cortexm0ds_logic.v(1700)
  wire Hpbow6;  // ../RTL/cortexm0ds_logic.v(1003)
  wire Hpcbx6;  // ../RTL/cortexm0ds_logic.v(1702)
  wire Hphax6;  // ../RTL/cortexm0ds_logic.v(1646)
  wire Hphiu6;  // ../RTL/cortexm0ds_logic.v(540)
  wire Hpiow6;  // ../RTL/cortexm0ds_logic.v(1096)
  wire Hpoiu6;  // ../RTL/cortexm0ds_logic.v(634)
  wire Hpphu6;  // ../RTL/cortexm0ds_logic.v(166)
  wire Hppow6;  // ../RTL/cortexm0ds_logic.v(1190)
  wire Hpviu6;  // ../RTL/cortexm0ds_logic.v(727)
  wire Hpwhu6;  // ../RTL/cortexm0ds_logic.v(259)
  wire Hpwow6;  // ../RTL/cortexm0ds_logic.v(1284)
  wire Hq1ju6;  // ../RTL/cortexm0ds_logic.v(808)
  wire Hq2iu6;  // ../RTL/cortexm0ds_logic.v(340)
  wire Hq2pw6;  // ../RTL/cortexm0ds_logic.v(1364)
  wire Hq8ju6;  // ../RTL/cortexm0ds_logic.v(901)
  wire Hq9iu6;  // ../RTL/cortexm0ds_logic.v(433)
  wire Hq9pw6;  // ../RTL/cortexm0ds_logic.v(1458)
  wire Hqabx6;  // ../RTL/cortexm0ds_logic.v(1698)
  wire Hqaow6;  // ../RTL/cortexm0ds_logic.v(990)
  wire Hqgiu6;  // ../RTL/cortexm0ds_logic.v(527)
  wire Hqhow6;  // ../RTL/cortexm0ds_logic.v(1083)
  wire Hqniu6;  // ../RTL/cortexm0ds_logic.v(621)
  wire Hqohu6;  // ../RTL/cortexm0ds_logic.v(153)
  wire Hqoow6;  // ../RTL/cortexm0ds_logic.v(1177)
  wire Hquiu6;  // ../RTL/cortexm0ds_logic.v(714)
  wire Hqvhu6;  // ../RTL/cortexm0ds_logic.v(246)
  wire Hqvow6;  // ../RTL/cortexm0ds_logic.v(1271)
  wire Hqxpw6;  // ../RTL/cortexm0ds_logic.v(1613)
  wire Hr0ju6;  // ../RTL/cortexm0ds_logic.v(795)
  wire Hr1iu6;  // ../RTL/cortexm0ds_logic.v(327)
  wire Hr1pw6;  // ../RTL/cortexm0ds_logic.v(1351)
  wire Hr7ju6;  // ../RTL/cortexm0ds_logic.v(888)
  wire Hr8iu6;  // ../RTL/cortexm0ds_logic.v(420)
  wire Hr8pw6;  // ../RTL/cortexm0ds_logic.v(1445)
  wire Hr9ow6;  // ../RTL/cortexm0ds_logic.v(977)
  wire Hrfbx6;  // ../RTL/cortexm0ds_logic.v(1708)
  wire Hrfiu6;  // ../RTL/cortexm0ds_logic.v(514)
  wire Hrgow6;  // ../RTL/cortexm0ds_logic.v(1070)
  wire Hrmiu6;  // ../RTL/cortexm0ds_logic.v(608)
  wire Hrnow6;  // ../RTL/cortexm0ds_logic.v(1164)
  wire Hroax6;  // ../RTL/cortexm0ds_logic.v(1659)
  wire Hrtiu6;  // ../RTL/cortexm0ds_logic.v(701)
  wire Hruhu6;  // ../RTL/cortexm0ds_logic.v(233)
  wire Hruow6;  // ../RTL/cortexm0ds_logic.v(1258)
  wire Hs0iu6;  // ../RTL/cortexm0ds_logic.v(314)
  wire Hs0pw6;  // ../RTL/cortexm0ds_logic.v(1338)
  wire Hs6ju6;  // ../RTL/cortexm0ds_logic.v(875)
  wire Hs7iu6;  // ../RTL/cortexm0ds_logic.v(407)
  wire Hs7pw6;  // ../RTL/cortexm0ds_logic.v(1432)
  wire Hs8ow6;  // ../RTL/cortexm0ds_logic.v(964)
  wire Hsdax6;  // ../RTL/cortexm0ds_logic.v(1639)
  wire Hseiu6;  // ../RTL/cortexm0ds_logic.v(501)
  wire Hsfow6;  // ../RTL/cortexm0ds_logic.v(1057)
  wire Hsliu6;  // ../RTL/cortexm0ds_logic.v(595)
  wire Hsmow6;  // ../RTL/cortexm0ds_logic.v(1151)
  wire Hssiu6;  // ../RTL/cortexm0ds_logic.v(688)
  wire Hsthu6;  // ../RTL/cortexm0ds_logic.v(220)
  wire Hstow6;  // ../RTL/cortexm0ds_logic.v(1245)
  wire Hsxpw6;  // ../RTL/cortexm0ds_logic.v(1613)
  wire Hsziu6;  // ../RTL/cortexm0ds_logic.v(782)
  wire Ht1qw6;  // ../RTL/cortexm0ds_logic.v(1620)
  wire Ht5ju6;  // ../RTL/cortexm0ds_logic.v(862)
  wire Ht6iu6;  // ../RTL/cortexm0ds_logic.v(394)
  wire Ht6pw6;  // ../RTL/cortexm0ds_logic.v(1419)
  wire Ht7ow6;  // ../RTL/cortexm0ds_logic.v(951)
  wire Htbax6;  // ../RTL/cortexm0ds_logic.v(1635)
  wire Htdiu6;  // ../RTL/cortexm0ds_logic.v(488)
  wire Htdpw6;  // ../RTL/cortexm0ds_logic.v(1512)
  wire Hteow6;  // ../RTL/cortexm0ds_logic.v(1044)
  wire Htkiu6;  // ../RTL/cortexm0ds_logic.v(582)
  wire Htlow6;  // ../RTL/cortexm0ds_logic.v(1138)
  wire Htmpw6;  // ../RTL/cortexm0ds_logic.v(1593)
  wire Htriu6;  // ../RTL/cortexm0ds_logic.v(675)
  wire Htshu6;  // ../RTL/cortexm0ds_logic.v(207)
  wire Htsow6;  // ../RTL/cortexm0ds_logic.v(1232)
  wire Htyiu6;  // ../RTL/cortexm0ds_logic.v(769)
  wire Htzhu6;  // ../RTL/cortexm0ds_logic.v(301)
  wire Htzow6;  // ../RTL/cortexm0ds_logic.v(1325)
  wire Hu4ju6;  // ../RTL/cortexm0ds_logic.v(849)
  wire Hu5iu6;  // ../RTL/cortexm0ds_logic.v(381)
  wire Hu5pw6;  // ../RTL/cortexm0ds_logic.v(1406)
  wire Hu6ow6;  // ../RTL/cortexm0ds_logic.v(938)
  wire Huciu6;  // ../RTL/cortexm0ds_logic.v(475)
  wire Hucpw6;  // ../RTL/cortexm0ds_logic.v(1499)
  wire Hudow6;  // ../RTL/cortexm0ds_logic.v(1031)
  wire Hujiu6;  // ../RTL/cortexm0ds_logic.v(569)
  wire Hukow6;  // ../RTL/cortexm0ds_logic.v(1125)
  wire Huqiu6;  // ../RTL/cortexm0ds_logic.v(662)
  wire Hurhu6;  // ../RTL/cortexm0ds_logic.v(194)
  wire Hurow6;  // ../RTL/cortexm0ds_logic.v(1219)
  wire Huxiu6;  // ../RTL/cortexm0ds_logic.v(756)
  wire Huxpw6;  // ../RTL/cortexm0ds_logic.v(1613)
  wire Huyhu6;  // ../RTL/cortexm0ds_logic.v(288)
  wire Huyow6;  // ../RTL/cortexm0ds_logic.v(1312)
  wire Hv3ju6;  // ../RTL/cortexm0ds_logic.v(836)
  wire Hv4pw6;  // ../RTL/cortexm0ds_logic.v(1393)
  wire Hvbiu6;  // ../RTL/cortexm0ds_logic.v(462)
  wire Hvbpw6;  // ../RTL/cortexm0ds_logic.v(1486)
  wire Hvcow6;  // ../RTL/cortexm0ds_logic.v(1018)
  wire Hviiu6;  // ../RTL/cortexm0ds_logic.v(556)
  wire Hvjow6;  // ../RTL/cortexm0ds_logic.v(1112)
  wire Hvpiu6;  // ../RTL/cortexm0ds_logic.v(649)
  wire Hvqhu6;  // ../RTL/cortexm0ds_logic.v(181)
  wire Hvqow6;  // ../RTL/cortexm0ds_logic.v(1206)
  wire Hvwiu6;  // ../RTL/cortexm0ds_logic.v(743)
  wire Hvxhu6;  // ../RTL/cortexm0ds_logic.v(275)
  wire Hvxow6;  // ../RTL/cortexm0ds_logic.v(1299)
  wire Hw2ju6;  // ../RTL/cortexm0ds_logic.v(823)
  wire Hw3iu6;  // ../RTL/cortexm0ds_logic.v(355)
  wire Hw3pw6;  // ../RTL/cortexm0ds_logic.v(1380)
  wire Hw8ax6;  // ../RTL/cortexm0ds_logic.v(1629)
  wire Hw9ju6;  // ../RTL/cortexm0ds_logic.v(917)
  wire Hwaiu6;  // ../RTL/cortexm0ds_logic.v(449)
  wire Hwapw6;  // ../RTL/cortexm0ds_logic.v(1473)
  wire Hwbow6;  // ../RTL/cortexm0ds_logic.v(1005)
  wire Hwhiu6;  // ../RTL/cortexm0ds_logic.v(543)
  wire Hwhpw6;  // ../RTL/cortexm0ds_logic.v(1584)
  wire Hwiow6;  // ../RTL/cortexm0ds_logic.v(1099)
  wire Hwmhu6;  // ../RTL/cortexm0ds_logic.v(143)
  wire Hwoiu6;  // ../RTL/cortexm0ds_logic.v(636)
  wire Hwphu6;  // ../RTL/cortexm0ds_logic.v(168)
  wire Hwpow6;  // ../RTL/cortexm0ds_logic.v(1193)
  wire Hwviu6;  // ../RTL/cortexm0ds_logic.v(730)
  wire Hwwhu6;  // ../RTL/cortexm0ds_logic.v(262)
  wire Hwwow6;  // ../RTL/cortexm0ds_logic.v(1286)
  wire Hx1ju6;  // ../RTL/cortexm0ds_logic.v(810)
  wire Hx2iu6;  // ../RTL/cortexm0ds_logic.v(342)
  wire Hx2pw6;  // ../RTL/cortexm0ds_logic.v(1367)
  wire Hx8ju6;  // ../RTL/cortexm0ds_logic.v(904)
  wire Hx9iu6;  // ../RTL/cortexm0ds_logic.v(436)
  wire Hx9pw6;  // ../RTL/cortexm0ds_logic.v(1460)
  wire Hxaow6;  // ../RTL/cortexm0ds_logic.v(992)
  wire Hxgiu6;  // ../RTL/cortexm0ds_logic.v(530)
  wire Hxhow6;  // ../RTL/cortexm0ds_logic.v(1086)
  wire Hxniu6;  // ../RTL/cortexm0ds_logic.v(623)
  wire Hxohu6;  // ../RTL/cortexm0ds_logic.v(155)
  wire Hxoow6;  // ../RTL/cortexm0ds_logic.v(1180)
  wire Hxuiu6;  // ../RTL/cortexm0ds_logic.v(717)
  wire Hxvhu6;  // ../RTL/cortexm0ds_logic.v(249)
  wire Hxvow6;  // ../RTL/cortexm0ds_logic.v(1273)
  wire Hy0ju6;  // ../RTL/cortexm0ds_logic.v(797)
  wire Hy1iu6;  // ../RTL/cortexm0ds_logic.v(329)
  wire Hy1pw6;  // ../RTL/cortexm0ds_logic.v(1354)
  wire Hy7ju6;  // ../RTL/cortexm0ds_logic.v(891)
  wire Hy8iu6;  // ../RTL/cortexm0ds_logic.v(423)
  wire Hy8pw6;  // ../RTL/cortexm0ds_logic.v(1447)
  wire Hy9ow6;  // ../RTL/cortexm0ds_logic.v(979)
  wire Hyfiu6;  // ../RTL/cortexm0ds_logic.v(517)
  wire Hygow6;  // ../RTL/cortexm0ds_logic.v(1073)
  wire Hymiu6;  // ../RTL/cortexm0ds_logic.v(610)
  wire Hynow6;  // ../RTL/cortexm0ds_logic.v(1167)
  wire Hysax6;  // ../RTL/cortexm0ds_logic.v(1667)
  wire Hytiu6;  // ../RTL/cortexm0ds_logic.v(704)
  wire Hyuhu6;  // ../RTL/cortexm0ds_logic.v(236)
  wire Hyuow6;  // ../RTL/cortexm0ds_logic.v(1260)
  wire Hz0iu6;  // ../RTL/cortexm0ds_logic.v(316)
  wire Hz0pw6;  // ../RTL/cortexm0ds_logic.v(1341)
  wire Hz6ju6;  // ../RTL/cortexm0ds_logic.v(878)
  wire Hz7iu6;  // ../RTL/cortexm0ds_logic.v(410)
  wire Hz7pw6;  // ../RTL/cortexm0ds_logic.v(1434)
  wire Hz8ow6;  // ../RTL/cortexm0ds_logic.v(966)
  wire Hz9ax6;  // ../RTL/cortexm0ds_logic.v(1631)
  wire Hzeiu6;  // ../RTL/cortexm0ds_logic.v(504)
  wire Hzfow6;  // ../RTL/cortexm0ds_logic.v(1060)
  wire Hzlhu6;  // ../RTL/cortexm0ds_logic.v(141)
  wire Hzliu6;  // ../RTL/cortexm0ds_logic.v(597)
  wire Hzmow6;  // ../RTL/cortexm0ds_logic.v(1154)
  wire Hzsiu6;  // ../RTL/cortexm0ds_logic.v(691)
  wire Hzthu6;  // ../RTL/cortexm0ds_logic.v(223)
  wire Hztow6;  // ../RTL/cortexm0ds_logic.v(1247)
  wire Hzziu6;  // ../RTL/cortexm0ds_logic.v(784)
  wire I03ju6;  // ../RTL/cortexm0ds_logic.v(825)
  wire I04iu6;  // ../RTL/cortexm0ds_logic.v(357)
  wire I04pw6;  // ../RTL/cortexm0ds_logic.v(1381)
  wire I0aju6;  // ../RTL/cortexm0ds_logic.v(919)
  wire I0biu6;  // ../RTL/cortexm0ds_logic.v(451)
  wire I0bpw6;  // ../RTL/cortexm0ds_logic.v(1475)
  wire I0cow6;  // ../RTL/cortexm0ds_logic.v(1007)
  wire I0dax6;  // ../RTL/cortexm0ds_logic.v(1637)
  wire I0iiu6;  // ../RTL/cortexm0ds_logic.v(544)
  wire I0jow6;  // ../RTL/cortexm0ds_logic.v(1101)
  wire I0opw6;  // ../RTL/cortexm0ds_logic.v(1595)
  wire I0piu6;  // ../RTL/cortexm0ds_logic.v(638)
  wire I0qhu6;  // ../RTL/cortexm0ds_logic.v(170)
  wire I0qow6;  // ../RTL/cortexm0ds_logic.v(1194)
  wire I0wiu6;  // ../RTL/cortexm0ds_logic.v(731)
  wire I0xhu6;  // ../RTL/cortexm0ds_logic.v(263)
  wire I0xow6;  // ../RTL/cortexm0ds_logic.v(1288)
  wire I12ju6;  // ../RTL/cortexm0ds_logic.v(812)
  wire I13iu6;  // ../RTL/cortexm0ds_logic.v(344)
  wire I13pw6;  // ../RTL/cortexm0ds_logic.v(1368)
  wire I19ju6;  // ../RTL/cortexm0ds_logic.v(906)
  wire I1aiu6;  // ../RTL/cortexm0ds_logic.v(438)
  wire I1apw6;  // ../RTL/cortexm0ds_logic.v(1462)
  wire I1bow6;  // ../RTL/cortexm0ds_logic.v(994)
  wire I1hiu6;  // ../RTL/cortexm0ds_logic.v(531)
  wire I1iow6;  // ../RTL/cortexm0ds_logic.v(1088)
  wire I1lpw6;  // ../RTL/cortexm0ds_logic.v(1589)
  wire I1oiu6;  // ../RTL/cortexm0ds_logic.v(625)
  wire I1phu6;  // ../RTL/cortexm0ds_logic.v(157)
  wire I1pow6;  // ../RTL/cortexm0ds_logic.v(1181)
  wire I1qpw6;  // ../RTL/cortexm0ds_logic.v(1599)
  wire I1viu6;  // ../RTL/cortexm0ds_logic.v(718)
  wire I1whu6;  // ../RTL/cortexm0ds_logic.v(250)
  wire I1wow6;  // ../RTL/cortexm0ds_logic.v(1275)
  wire I21ju6;  // ../RTL/cortexm0ds_logic.v(799)
  wire I22iu6;  // ../RTL/cortexm0ds_logic.v(331)
  wire I22pw6;  // ../RTL/cortexm0ds_logic.v(1355)
  wire I28ju6;  // ../RTL/cortexm0ds_logic.v(893)
  wire I29iu6;  // ../RTL/cortexm0ds_logic.v(425)
  wire I29pw6;  // ../RTL/cortexm0ds_logic.v(1449)
  wire I2aow6;  // ../RTL/cortexm0ds_logic.v(981)
  wire I2giu6;  // ../RTL/cortexm0ds_logic.v(518)
  wire I2how6;  // ../RTL/cortexm0ds_logic.v(1075)
  wire I2niu6;  // ../RTL/cortexm0ds_logic.v(612)
  wire I2oow6;  // ../RTL/cortexm0ds_logic.v(1168)
  wire I2uiu6;  // ../RTL/cortexm0ds_logic.v(705)
  wire I2vhu6;  // ../RTL/cortexm0ds_logic.v(237)
  wire I2vow6;  // ../RTL/cortexm0ds_logic.v(1262)
  wire I2zax6;  // ../RTL/cortexm0ds_logic.v(1678)
  wire I30ju6;  // ../RTL/cortexm0ds_logic.v(786)
  wire I31iu6;  // ../RTL/cortexm0ds_logic.v(318)
  wire I31pw6;  // ../RTL/cortexm0ds_logic.v(1342)
  wire I37ju6;  // ../RTL/cortexm0ds_logic.v(880)
  wire I38iu6;  // ../RTL/cortexm0ds_logic.v(412)
  wire I38pw6;  // ../RTL/cortexm0ds_logic.v(1436)
  wire I39ow6;  // ../RTL/cortexm0ds_logic.v(968)
  wire I3fhu6;  // ../RTL/cortexm0ds_logic.v(123)
  wire I3fiu6;  // ../RTL/cortexm0ds_logic.v(505)
  wire I3gow6;  // ../RTL/cortexm0ds_logic.v(1062)
  wire I3lhu6;  // ../RTL/cortexm0ds_logic.v(138)
  wire I3miu6;  // ../RTL/cortexm0ds_logic.v(599)
  wire I3now6;  // ../RTL/cortexm0ds_logic.v(1155)
  wire I3qpw6;  // ../RTL/cortexm0ds_logic.v(1599)
  wire I3tiu6;  // ../RTL/cortexm0ds_logic.v(692)
  wire I3uhu6;  // ../RTL/cortexm0ds_logic.v(224)
  wire I3uow6;  // ../RTL/cortexm0ds_logic.v(1249)
  wire I40iu6;  // ../RTL/cortexm0ds_logic.v(305)
  wire I40pw6;  // ../RTL/cortexm0ds_logic.v(1329)
  wire I45bx6;  // ../RTL/cortexm0ds_logic.v(1688)
  wire I46ju6;  // ../RTL/cortexm0ds_logic.v(867)
  wire I47iu6;  // ../RTL/cortexm0ds_logic.v(399)
  wire I47pw6;  // ../RTL/cortexm0ds_logic.v(1423)
  wire I48ow6;  // ../RTL/cortexm0ds_logic.v(955)
  wire I4eiu6;  // ../RTL/cortexm0ds_logic.v(492)
  wire I4epw6;  // ../RTL/cortexm0ds_logic.v(1517)
  wire I4fow6;  // ../RTL/cortexm0ds_logic.v(1049)
  wire I4liu6;  // ../RTL/cortexm0ds_logic.v(586)
  wire I4mow6;  // ../RTL/cortexm0ds_logic.v(1142)
  wire I4rpw6;  // ../RTL/cortexm0ds_logic.v(1601)
  wire I4siu6;  // ../RTL/cortexm0ds_logic.v(679)
  wire I4thu6;  // ../RTL/cortexm0ds_logic.v(211)
  wire I4tow6;  // ../RTL/cortexm0ds_logic.v(1236)
  wire I4ziu6;  // ../RTL/cortexm0ds_logic.v(773)
  wire I55ju6;  // ../RTL/cortexm0ds_logic.v(854)
  wire I56iu6;  // ../RTL/cortexm0ds_logic.v(386)
  wire I56pw6;  // ../RTL/cortexm0ds_logic.v(1410)
  wire I57ow6;  // ../RTL/cortexm0ds_logic.v(942)
  wire I5diu6;  // ../RTL/cortexm0ds_logic.v(479)
  wire I5dpw6;  // ../RTL/cortexm0ds_logic.v(1504)
  wire I5eow6;  // ../RTL/cortexm0ds_logic.v(1036)
  wire I5khu6;  // ../RTL/cortexm0ds_logic.v(136)
  wire I5kiu6;  // ../RTL/cortexm0ds_logic.v(573)
  wire I5low6;  // ../RTL/cortexm0ds_logic.v(1129)
  wire I5nhu6;  // ../RTL/cortexm0ds_logic.v(144)
  wire I5qpw6;  // ../RTL/cortexm0ds_logic.v(1599)
  wire I5riu6;  // ../RTL/cortexm0ds_logic.v(666)
  wire I5shu6;  // ../RTL/cortexm0ds_logic.v(198)
  wire I5sow6;  // ../RTL/cortexm0ds_logic.v(1223)
  wire I5xax6;  // ../RTL/cortexm0ds_logic.v(1674)
  wire I5yiu6;  // ../RTL/cortexm0ds_logic.v(760)
  wire I5zhu6;  // ../RTL/cortexm0ds_logic.v(292)
  wire I5zow6;  // ../RTL/cortexm0ds_logic.v(1316)
  wire I64ju6;  // ../RTL/cortexm0ds_logic.v(841)
  wire I65iu6;  // ../RTL/cortexm0ds_logic.v(373)
  wire I65pw6;  // ../RTL/cortexm0ds_logic.v(1397)
  wire I6ciu6;  // ../RTL/cortexm0ds_logic.v(466)
  wire I6cpw6;  // ../RTL/cortexm0ds_logic.v(1491)
  wire I6dow6;  // ../RTL/cortexm0ds_logic.v(1023)
  wire I6jiu6;  // ../RTL/cortexm0ds_logic.v(560)
  wire I6kow6;  // ../RTL/cortexm0ds_logic.v(1116)
  wire I6qiu6;  // ../RTL/cortexm0ds_logic.v(653)
  wire I6rhu6;  // ../RTL/cortexm0ds_logic.v(185)
  wire I6row6;  // ../RTL/cortexm0ds_logic.v(1210)
  wire I6xiu6;  // ../RTL/cortexm0ds_logic.v(747)
  wire I6yhu6;  // ../RTL/cortexm0ds_logic.v(279)
  wire I6yow6;  // ../RTL/cortexm0ds_logic.v(1303)
  wire I73ju6;  // ../RTL/cortexm0ds_logic.v(828)
  wire I74bx6;  // ../RTL/cortexm0ds_logic.v(1687)
  wire I74iu6;  // ../RTL/cortexm0ds_logic.v(360)
  wire I74pw6;  // ../RTL/cortexm0ds_logic.v(1384)
  wire I7aju6;  // ../RTL/cortexm0ds_logic.v(921)
  wire I7biu6;  // ../RTL/cortexm0ds_logic.v(453)
  wire I7bpw6;  // ../RTL/cortexm0ds_logic.v(1478)
  wire I7cow6;  // ../RTL/cortexm0ds_logic.v(1010)
  wire I7iiu6;  // ../RTL/cortexm0ds_logic.v(547)
  wire I7jhu6;  // ../RTL/cortexm0ds_logic.v(133)
  wire I7jow6;  // ../RTL/cortexm0ds_logic.v(1103)
  wire I7piu6;  // ../RTL/cortexm0ds_logic.v(640)
  wire I7qhu6;  // ../RTL/cortexm0ds_logic.v(172)
  wire I7qow6;  // ../RTL/cortexm0ds_logic.v(1197)
  wire I7qpw6;  // ../RTL/cortexm0ds_logic.v(1599)
  wire I7wiu6;  // ../RTL/cortexm0ds_logic.v(734)
  wire I7xhu6;  // ../RTL/cortexm0ds_logic.v(266)
  wire I7xow6;  // ../RTL/cortexm0ds_logic.v(1290)
  wire I82ju6;  // ../RTL/cortexm0ds_logic.v(815)
  wire I83iu6;  // ../RTL/cortexm0ds_logic.v(347)
  wire I83pw6;  // ../RTL/cortexm0ds_logic.v(1371)
  wire I89ju6;  // ../RTL/cortexm0ds_logic.v(908)
  wire I8aiu6;  // ../RTL/cortexm0ds_logic.v(440)
  wire I8apw6;  // ../RTL/cortexm0ds_logic.v(1465)
  wire I8bow6;  // ../RTL/cortexm0ds_logic.v(997)
  wire I8hax6;  // ../RTL/cortexm0ds_logic.v(1645)
  wire I8hiu6;  // ../RTL/cortexm0ds_logic.v(534)
  wire I8iow6;  // ../RTL/cortexm0ds_logic.v(1090)
  wire I8lax6;  // ../RTL/cortexm0ds_logic.v(1653)
  wire I8oiu6;  // ../RTL/cortexm0ds_logic.v(627)
  wire I8phu6;  // ../RTL/cortexm0ds_logic.v(159)
  wire I8pow6;  // ../RTL/cortexm0ds_logic.v(1184)
  wire I8viu6;  // ../RTL/cortexm0ds_logic.v(721)
  wire I8whu6;  // ../RTL/cortexm0ds_logic.v(253)
  wire I8wow6;  // ../RTL/cortexm0ds_logic.v(1277)
  wire I91ju6;  // ../RTL/cortexm0ds_logic.v(802)
  wire I92iu6;  // ../RTL/cortexm0ds_logic.v(334)
  wire I92pw6;  // ../RTL/cortexm0ds_logic.v(1358)
  wire I98ju6;  // ../RTL/cortexm0ds_logic.v(895)
  wire I99iu6;  // ../RTL/cortexm0ds_logic.v(427)
  wire I99pw6;  // ../RTL/cortexm0ds_logic.v(1452)
  wire I9aow6;  // ../RTL/cortexm0ds_logic.v(984)
  wire I9giu6;  // ../RTL/cortexm0ds_logic.v(521)
  wire I9how6;  // ../RTL/cortexm0ds_logic.v(1077)
  wire I9ihu6;  // ../RTL/cortexm0ds_logic.v(130)
  wire I9niu6;  // ../RTL/cortexm0ds_logic.v(614)
  wire I9oow6;  // ../RTL/cortexm0ds_logic.v(1171)
  wire I9qpw6;  // ../RTL/cortexm0ds_logic.v(1599)
  wire I9uiu6;  // ../RTL/cortexm0ds_logic.v(708)
  wire I9vhu6;  // ../RTL/cortexm0ds_logic.v(240)
  wire I9vow6;  // ../RTL/cortexm0ds_logic.v(1264)
  wire Ia0ju6;  // ../RTL/cortexm0ds_logic.v(789)
  wire Ia1iu6;  // ../RTL/cortexm0ds_logic.v(321)
  wire Ia1pw6;  // ../RTL/cortexm0ds_logic.v(1345)
  wire Ia7ju6;  // ../RTL/cortexm0ds_logic.v(882)
  wire Ia8iu6;  // ../RTL/cortexm0ds_logic.v(414)
  wire Ia8pw6;  // ../RTL/cortexm0ds_logic.v(1439)
  wire Ia9ow6;  // ../RTL/cortexm0ds_logic.v(971)
  wire Iafiu6;  // ../RTL/cortexm0ds_logic.v(508)
  wire Iagow6;  // ../RTL/cortexm0ds_logic.v(1064)
  wire Iamiu6;  // ../RTL/cortexm0ds_logic.v(601)
  wire Ianow6;  // ../RTL/cortexm0ds_logic.v(1158)
  wire Iatiu6;  // ../RTL/cortexm0ds_logic.v(695)
  wire Iauhu6;  // ../RTL/cortexm0ds_logic.v(227)
  wire Iauow6;  // ../RTL/cortexm0ds_logic.v(1251)
  wire Ib0iu6;  // ../RTL/cortexm0ds_logic.v(308)
  wire Ib0pw6;  // ../RTL/cortexm0ds_logic.v(1332)
  wire Ib6ju6;  // ../RTL/cortexm0ds_logic.v(869)
  wire Ib7iu6;  // ../RTL/cortexm0ds_logic.v(401)
  wire Ib7pw6;  // ../RTL/cortexm0ds_logic.v(1426)
  wire Ib8ow6;  // ../RTL/cortexm0ds_logic.v(958)
  wire Ibeiu6;  // ../RTL/cortexm0ds_logic.v(495)
  wire Ibfow6;  // ../RTL/cortexm0ds_logic.v(1051)
  wire Ibliu6;  // ../RTL/cortexm0ds_logic.v(588)
  wire Ibmow6;  // ../RTL/cortexm0ds_logic.v(1145)
  wire Ibqpw6;  // ../RTL/cortexm0ds_logic.v(1599)
  wire Ibsiu6;  // ../RTL/cortexm0ds_logic.v(682)
  wire Ibthu6;  // ../RTL/cortexm0ds_logic.v(214)
  wire Ibtow6;  // ../RTL/cortexm0ds_logic.v(1238)
  wire Ibziu6;  // ../RTL/cortexm0ds_logic.v(776)
  wire Ic5ju6;  // ../RTL/cortexm0ds_logic.v(856)
  wire Ic6iu6;  // ../RTL/cortexm0ds_logic.v(388)
  wire Ic6pw6;  // ../RTL/cortexm0ds_logic.v(1413)
  wire Ic7ow6;  // ../RTL/cortexm0ds_logic.v(945)
  wire Icdiu6;  // ../RTL/cortexm0ds_logic.v(482)
  wire Icdpw6;  // ../RTL/cortexm0ds_logic.v(1506)
  wire Iceow6;  // ../RTL/cortexm0ds_logic.v(1038)
  wire Ickiu6;  // ../RTL/cortexm0ds_logic.v(575)
  wire Iclow6;  // ../RTL/cortexm0ds_logic.v(1132)
  wire Icriu6;  // ../RTL/cortexm0ds_logic.v(669)
  wire Icshu6;  // ../RTL/cortexm0ds_logic.v(201)
  wire Icsow6;  // ../RTL/cortexm0ds_logic.v(1225)
  wire Icyiu6;  // ../RTL/cortexm0ds_logic.v(763)
  wire Iczhu6;  // ../RTL/cortexm0ds_logic.v(295)
  wire Iczow6;  // ../RTL/cortexm0ds_logic.v(1319)
  wire Id4ju6;  // ../RTL/cortexm0ds_logic.v(843)
  wire Id5iu6;  // ../RTL/cortexm0ds_logic.v(375)
  wire Id5pw6;  // ../RTL/cortexm0ds_logic.v(1400)
  wire Id6ow6;  // ../RTL/cortexm0ds_logic.v(932)
  wire Idciu6;  // ../RTL/cortexm0ds_logic.v(469)
  wire Idcpw6;  // ../RTL/cortexm0ds_logic.v(1493)
  wire Iddax6;  // ../RTL/cortexm0ds_logic.v(1638)
  wire Iddow6;  // ../RTL/cortexm0ds_logic.v(1025)
  wire Idjiu6;  // ../RTL/cortexm0ds_logic.v(562)
  wire Idkow6;  // ../RTL/cortexm0ds_logic.v(1119)
  wire Idqiu6;  // ../RTL/cortexm0ds_logic.v(656)
  wire Idqpw6;  // ../RTL/cortexm0ds_logic.v(1599)
  wire Idrhu6;  // ../RTL/cortexm0ds_logic.v(188)
  wire Idrow6;  // ../RTL/cortexm0ds_logic.v(1212)
  wire Idxiu6;  // ../RTL/cortexm0ds_logic.v(750)
  wire Idyhu6;  // ../RTL/cortexm0ds_logic.v(282)
  wire Idyow6;  // ../RTL/cortexm0ds_logic.v(1306)
  wire Ie1bx6;  // ../RTL/cortexm0ds_logic.v(1682)
  wire Ie3ju6;  // ../RTL/cortexm0ds_logic.v(830)
  wire Ie4iu6;  // ../RTL/cortexm0ds_logic.v(362)
  wire Ie4pw6;  // ../RTL/cortexm0ds_logic.v(1387)
  wire Ieaju6;  // ../RTL/cortexm0ds_logic.v(924)
  wire Iebiu6;  // ../RTL/cortexm0ds_logic.v(456)
  wire Iebpw6;  // ../RTL/cortexm0ds_logic.v(1480)
  wire Iecow6;  // ../RTL/cortexm0ds_logic.v(1012)
  wire Ieiiu6;  // ../RTL/cortexm0ds_logic.v(549)
  wire Iejow6;  // ../RTL/cortexm0ds_logic.v(1106)
  wire Iekax6;  // ../RTL/cortexm0ds_logic.v(1651)
  wire Iepiu6;  // ../RTL/cortexm0ds_logic.v(643)
  wire Ieqhu6;  // ../RTL/cortexm0ds_logic.v(175)
  wire Ieqow6;  // ../RTL/cortexm0ds_logic.v(1199)
  wire Iewiu6;  // ../RTL/cortexm0ds_logic.v(737)
  wire Iexhu6;  // ../RTL/cortexm0ds_logic.v(269)
  wire Iexow6;  // ../RTL/cortexm0ds_logic.v(1293)
  wire If2ju6;  // ../RTL/cortexm0ds_logic.v(817)
  wire If3iu6;  // ../RTL/cortexm0ds_logic.v(349)
  wire If3pw6;  // ../RTL/cortexm0ds_logic.v(1374)
  wire If9ju6;  // ../RTL/cortexm0ds_logic.v(911)
  wire Ifaiu6;  // ../RTL/cortexm0ds_logic.v(443)
  wire Ifapw6;  // ../RTL/cortexm0ds_logic.v(1467)
  wire Ifbow6;  // ../RTL/cortexm0ds_logic.v(999)
  wire Ifhiu6;  // ../RTL/cortexm0ds_logic.v(536)
  wire Ifiow6;  // ../RTL/cortexm0ds_logic.v(1093)
  wire Ifoiu6;  // ../RTL/cortexm0ds_logic.v(630)
  wire Ifphu6;  // ../RTL/cortexm0ds_logic.v(162)
  wire Ifpow6;  // ../RTL/cortexm0ds_logic.v(1186)
  wire Ifviu6;  // ../RTL/cortexm0ds_logic.v(724)
  wire Ifwhu6;  // ../RTL/cortexm0ds_logic.v(256)
  wire Ifwow6;  // ../RTL/cortexm0ds_logic.v(1280)
  wire Ig1ju6;  // ../RTL/cortexm0ds_logic.v(804)
  wire Ig2bx6;  // ../RTL/cortexm0ds_logic.v(1684)
  wire Ig2iu6;  // ../RTL/cortexm0ds_logic.v(336)
  wire Ig2pw6;  // ../RTL/cortexm0ds_logic.v(1361)
  wire Ig8ju6;  // ../RTL/cortexm0ds_logic.v(898)
  wire Ig9iu6;  // ../RTL/cortexm0ds_logic.v(430)
  wire Ig9pw6;  // ../RTL/cortexm0ds_logic.v(1454)
  wire Igaow6;  // ../RTL/cortexm0ds_logic.v(986)
  wire Iggiu6;  // ../RTL/cortexm0ds_logic.v(523)
  wire Ighow6;  // ../RTL/cortexm0ds_logic.v(1080)
  wire Igniu6;  // ../RTL/cortexm0ds_logic.v(617)
  wire Igohu6;  // ../RTL/cortexm0ds_logic.v(149)
  wire Igoow6;  // ../RTL/cortexm0ds_logic.v(1173)
  wire Iguiu6;  // ../RTL/cortexm0ds_logic.v(711)
  wire Igvhu6;  // ../RTL/cortexm0ds_logic.v(243)
  wire Igvow6;  // ../RTL/cortexm0ds_logic.v(1267)
  wire Ih0bx6;  // ../RTL/cortexm0ds_logic.v(1680)
  wire Ih0ju6;  // ../RTL/cortexm0ds_logic.v(791)
  wire Ih1iu6;  // ../RTL/cortexm0ds_logic.v(323)
  wire Ih1pw6;  // ../RTL/cortexm0ds_logic.v(1348)
  wire Ih7ju6;  // ../RTL/cortexm0ds_logic.v(885)
  wire Ih8iu6;  // ../RTL/cortexm0ds_logic.v(417)
  wire Ih8pw6;  // ../RTL/cortexm0ds_logic.v(1441)
  wire Ih9ow6;  // ../RTL/cortexm0ds_logic.v(973)
  wire Ihfiu6;  // ../RTL/cortexm0ds_logic.v(510)
  wire Ihmiu6;  // ../RTL/cortexm0ds_logic.v(604)
  wire Ihnow6;  // ../RTL/cortexm0ds_logic.v(1160)
  wire Ihtiu6;  // ../RTL/cortexm0ds_logic.v(698)
  wire Ihuhu6;  // ../RTL/cortexm0ds_logic.v(230)
  wire Ihuow6;  // ../RTL/cortexm0ds_logic.v(1254)
  wire Ii0iu6;  // ../RTL/cortexm0ds_logic.v(310)
  wire Ii0pw6;  // ../RTL/cortexm0ds_logic.v(1335)
  wire Ii6ju6;  // ../RTL/cortexm0ds_logic.v(872)
  wire Ii7iu6;  // ../RTL/cortexm0ds_logic.v(404)
  wire Ii7pw6;  // ../RTL/cortexm0ds_logic.v(1428)
  wire Ii8ow6;  // ../RTL/cortexm0ds_logic.v(960)
  wire Iieiu6;  // ../RTL/cortexm0ds_logic.v(497)
  wire Iifow6;  // ../RTL/cortexm0ds_logic.v(1054)
  wire Iiliu6;  // ../RTL/cortexm0ds_logic.v(591)
  wire Iimhu6;  // ../RTL/cortexm0ds_logic.v(142)
  wire Iimow6;  // ../RTL/cortexm0ds_logic.v(1147)
  wire Iisiu6;  // ../RTL/cortexm0ds_logic.v(685)
  wire Iithu6;  // ../RTL/cortexm0ds_logic.v(217)
  wire Iitow6;  // ../RTL/cortexm0ds_logic.v(1241)
  wire Iixpw6;  // ../RTL/cortexm0ds_logic.v(1612)
  wire Iiziu6;  // ../RTL/cortexm0ds_logic.v(778)
  wire Ij5ju6;  // ../RTL/cortexm0ds_logic.v(859)
  wire Ij6iu6;  // ../RTL/cortexm0ds_logic.v(391)
  wire Ij6pw6;  // ../RTL/cortexm0ds_logic.v(1415)
  wire Ij7ow6;  // ../RTL/cortexm0ds_logic.v(947)
  wire Ijdiu6;  // ../RTL/cortexm0ds_logic.v(484)
  wire Ijdpw6;  // ../RTL/cortexm0ds_logic.v(1509)
  wire Ijehu6;  // ../RTL/cortexm0ds_logic.v(122)
  wire Ijeow6;  // ../RTL/cortexm0ds_logic.v(1041)
  wire Ijhhu6;  // ../RTL/cortexm0ds_logic.v(128)
  wire Ijiax6;  // ../RTL/cortexm0ds_logic.v(1648)
  wire Ijkiu6;  // ../RTL/cortexm0ds_logic.v(578)
  wire Ijlow6;  // ../RTL/cortexm0ds_logic.v(1134)
  wire Ijriu6;  // ../RTL/cortexm0ds_logic.v(672)
  wire Ijshu6;  // ../RTL/cortexm0ds_logic.v(204)
  wire Ijsow6;  // ../RTL/cortexm0ds_logic.v(1228)
  wire Ijyiu6;  // ../RTL/cortexm0ds_logic.v(765)
  wire Ijzhu6;  // ../RTL/cortexm0ds_logic.v(297)
  wire Ijzow6;  // ../RTL/cortexm0ds_logic.v(1322)
  wire Ik4ju6;  // ../RTL/cortexm0ds_logic.v(846)
  wire Ik5iu6;  // ../RTL/cortexm0ds_logic.v(378)
  wire Ik5pw6;  // ../RTL/cortexm0ds_logic.v(1402)
  wire Ik6ow6;  // ../RTL/cortexm0ds_logic.v(934)
  wire Ikciu6;  // ../RTL/cortexm0ds_logic.v(471)
  wire Ikcpw6;  // ../RTL/cortexm0ds_logic.v(1496)
  wire Ikdow6;  // ../RTL/cortexm0ds_logic.v(1028)
  wire Ikghu6;  // ../RTL/cortexm0ds_logic.v(126)
  wire Ikhbx6;  // ../RTL/cortexm0ds_logic.v(1711)
  wire Ikjiu6;  // ../RTL/cortexm0ds_logic.v(565)
  wire Ikkow6;  // ../RTL/cortexm0ds_logic.v(1121)
  wire Ikqiu6;  // ../RTL/cortexm0ds_logic.v(659)
  wire Ikrhu6;  // ../RTL/cortexm0ds_logic.v(191)
  wire Ikrow6;  // ../RTL/cortexm0ds_logic.v(1215)
  wire Ikxiu6;  // ../RTL/cortexm0ds_logic.v(752)
  wire Ikyhu6;  // ../RTL/cortexm0ds_logic.v(284)
  wire Ikyow6;  // ../RTL/cortexm0ds_logic.v(1309)
  wire Il3ju6;  // ../RTL/cortexm0ds_logic.v(833)
  wire Il4iu6;  // ../RTL/cortexm0ds_logic.v(365)
  wire Il4pw6;  // ../RTL/cortexm0ds_logic.v(1389)
  wire Ilaju6;  // ../RTL/cortexm0ds_logic.v(926)
  wire Ilbiu6;  // ../RTL/cortexm0ds_logic.v(458)
  wire Ilbpw6;  // ../RTL/cortexm0ds_logic.v(1483)
  wire Ilcow6;  // ../RTL/cortexm0ds_logic.v(1015)
  wire Iliiu6;  // ../RTL/cortexm0ds_logic.v(552)
  wire Iljow6;  // ../RTL/cortexm0ds_logic.v(1108)
  wire Illhu6;  // ../RTL/cortexm0ds_logic.v(140)
  wire Ilpiu6;  // ../RTL/cortexm0ds_logic.v(646)
  wire Ilqhu6;  // ../RTL/cortexm0ds_logic.v(178)
  wire Ilqow6;  // ../RTL/cortexm0ds_logic.v(1202)
  wire Ilwiu6;  // ../RTL/cortexm0ds_logic.v(739)
  wire Ilxhu6;  // ../RTL/cortexm0ds_logic.v(271)
  wire Ilxow6;  // ../RTL/cortexm0ds_logic.v(1296)
  wire Im2ju6;  // ../RTL/cortexm0ds_logic.v(820)
  wire Im3iu6;  // ../RTL/cortexm0ds_logic.v(352)
  wire Im3pw6;  // ../RTL/cortexm0ds_logic.v(1376)
  wire Im9ax6;  // ../RTL/cortexm0ds_logic.v(1630)
  wire Im9ju6;  // ../RTL/cortexm0ds_logic.v(913)
  wire Imaiu6;  // ../RTL/cortexm0ds_logic.v(445)
  wire Imapw6;  // ../RTL/cortexm0ds_logic.v(1470)
  wire Imbow6;  // ../RTL/cortexm0ds_logic.v(1002)
  wire Imhbx6;  // ../RTL/cortexm0ds_logic.v(1711)
  wire Imhiu6;  // ../RTL/cortexm0ds_logic.v(539)
  wire Imiow6;  // ../RTL/cortexm0ds_logic.v(1095)
  wire Imkhu6;  // ../RTL/cortexm0ds_logic.v(137)
  wire Imoiu6;  // ../RTL/cortexm0ds_logic.v(633)
  wire Imphu6;  // ../RTL/cortexm0ds_logic.v(165)
  wire Impow6;  // ../RTL/cortexm0ds_logic.v(1189)
  wire Imviu6;  // ../RTL/cortexm0ds_logic.v(726)
  wire Imwhu6;  // ../RTL/cortexm0ds_logic.v(258)
  wire Imwow6;  // ../RTL/cortexm0ds_logic.v(1283)
  wire In1ju6;  // ../RTL/cortexm0ds_logic.v(807)
  wire In2iu6;  // ../RTL/cortexm0ds_logic.v(339)
  wire In2pw6;  // ../RTL/cortexm0ds_logic.v(1363)
  wire In8ju6;  // ../RTL/cortexm0ds_logic.v(900)
  wire In9iu6;  // ../RTL/cortexm0ds_logic.v(432)
  wire In9pw6;  // ../RTL/cortexm0ds_logic.v(1457)
  wire Inaow6;  // ../RTL/cortexm0ds_logic.v(989)
  wire Ingiu6;  // ../RTL/cortexm0ds_logic.v(526)
  wire Inhow6;  // ../RTL/cortexm0ds_logic.v(1082)
  wire Inniu6;  // ../RTL/cortexm0ds_logic.v(620)
  wire Inohu6;  // ../RTL/cortexm0ds_logic.v(152)
  wire Inoow6;  // ../RTL/cortexm0ds_logic.v(1176)
  wire Inuiu6;  // ../RTL/cortexm0ds_logic.v(713)
  wire Invhu6;  // ../RTL/cortexm0ds_logic.v(245)
  wire Invow6;  // ../RTL/cortexm0ds_logic.v(1270)
  wire Io0ju6;  // ../RTL/cortexm0ds_logic.v(794)
  wire Io1iu6;  // ../RTL/cortexm0ds_logic.v(326)
  wire Io1pw6;  // ../RTL/cortexm0ds_logic.v(1350)
  wire Io7ju6;  // ../RTL/cortexm0ds_logic.v(887)
  wire Io8iu6;  // ../RTL/cortexm0ds_logic.v(419)
  wire Io8pw6;  // ../RTL/cortexm0ds_logic.v(1444)
  wire Io9ow6;  // ../RTL/cortexm0ds_logic.v(976)
  wire Iofiu6;  // ../RTL/cortexm0ds_logic.v(513)
  wire Iogow6;  // ../RTL/cortexm0ds_logic.v(1069)
  wire Iojhu6;  // ../RTL/cortexm0ds_logic.v(134)
  wire Iomiu6;  // ../RTL/cortexm0ds_logic.v(607)
  wire Ionow6;  // ../RTL/cortexm0ds_logic.v(1163)
  wire Iotiu6;  // ../RTL/cortexm0ds_logic.v(700)
  wire Iouhu6;  // ../RTL/cortexm0ds_logic.v(232)
  wire Iouow6;  // ../RTL/cortexm0ds_logic.v(1257)
  wire Ip0iu6;  // ../RTL/cortexm0ds_logic.v(313)
  wire Ip0pw6;  // ../RTL/cortexm0ds_logic.v(1337)
  wire Ip6ju6;  // ../RTL/cortexm0ds_logic.v(874)
  wire Ip7iu6;  // ../RTL/cortexm0ds_logic.v(406)
  wire Ip7pw6;  // ../RTL/cortexm0ds_logic.v(1431)
  wire Ip8ow6;  // ../RTL/cortexm0ds_logic.v(963)
  wire Ipeiu6;  // ../RTL/cortexm0ds_logic.v(500)
  wire Ipfow6;  // ../RTL/cortexm0ds_logic.v(1056)
  wire Ipliu6;  // ../RTL/cortexm0ds_logic.v(594)
  wire Ipmow6;  // ../RTL/cortexm0ds_logic.v(1150)
  wire Ipoax6;  // ../RTL/cortexm0ds_logic.v(1659)
  wire Ipsiu6;  // ../RTL/cortexm0ds_logic.v(687)
  wire Ipthu6;  // ../RTL/cortexm0ds_logic.v(219)
  wire Iptow6;  // ../RTL/cortexm0ds_logic.v(1244)
  wire Ipziu6;  // ../RTL/cortexm0ds_logic.v(781)
  wire Iq5ju6;  // ../RTL/cortexm0ds_logic.v(861)
  wire Iq6iu6;  // ../RTL/cortexm0ds_logic.v(393)
  wire Iq6pw6;  // ../RTL/cortexm0ds_logic.v(1418)
  wire Iq7ow6;  // ../RTL/cortexm0ds_logic.v(950)
  wire Iqdiu6;  // ../RTL/cortexm0ds_logic.v(487)
  wire Iqdpw6;  // ../RTL/cortexm0ds_logic.v(1511)
  wire Iqeow6;  // ../RTL/cortexm0ds_logic.v(1043)
  wire Iqihu6;  // ../RTL/cortexm0ds_logic.v(132)
  wire Iqkiu6;  // ../RTL/cortexm0ds_logic.v(581)
  wire Iqlow6;  // ../RTL/cortexm0ds_logic.v(1137)
  wire Iqnhu6;  // ../RTL/cortexm0ds_logic.v(145)
  wire Iqriu6;  // ../RTL/cortexm0ds_logic.v(674)
  wire Iqshu6;  // ../RTL/cortexm0ds_logic.v(206)
  wire Iqsow6;  // ../RTL/cortexm0ds_logic.v(1231)
  wire Iqyiu6;  // ../RTL/cortexm0ds_logic.v(768)
  wire Iqzhu6;  // ../RTL/cortexm0ds_logic.v(300)
  wire Iqzow6;  // ../RTL/cortexm0ds_logic.v(1324)
  wire Ir1qw6;  // ../RTL/cortexm0ds_logic.v(1620)
  wire Ir4ju6;  // ../RTL/cortexm0ds_logic.v(848)
  wire Ir5iu6;  // ../RTL/cortexm0ds_logic.v(380)
  wire Ir5pw6;  // ../RTL/cortexm0ds_logic.v(1405)
  wire Ir6ow6;  // ../RTL/cortexm0ds_logic.v(937)
  wire Irciu6;  // ../RTL/cortexm0ds_logic.v(474)
  wire Ircpw6;  // ../RTL/cortexm0ds_logic.v(1498)
  wire Irdow6;  // ../RTL/cortexm0ds_logic.v(1030)
  wire Irjiu6;  // ../RTL/cortexm0ds_logic.v(568)
  wire Irkow6;  // ../RTL/cortexm0ds_logic.v(1124)
  wire Irmpw6;  // ../RTL/cortexm0ds_logic.v(1593)
  wire Irqiu6;  // ../RTL/cortexm0ds_logic.v(661)
  wire Irrhu6;  // ../RTL/cortexm0ds_logic.v(193)
  wire Irrow6;  // ../RTL/cortexm0ds_logic.v(1218)
  wire Irxiu6;  // ../RTL/cortexm0ds_logic.v(755)
  wire Iryhu6;  // ../RTL/cortexm0ds_logic.v(287)
  wire Iryow6;  // ../RTL/cortexm0ds_logic.v(1311)
  wire Is3ju6;  // ../RTL/cortexm0ds_logic.v(835)
  wire Is4iu6;  // ../RTL/cortexm0ds_logic.v(367)
  wire Is4pw6;  // ../RTL/cortexm0ds_logic.v(1392)
  wire Isaju6;  // ../RTL/cortexm0ds_logic.v(929)
  wire Isbiu6;  // ../RTL/cortexm0ds_logic.v(461)
  wire Isbpw6;  // ../RTL/cortexm0ds_logic.v(1485)
  wire Iscow6;  // ../RTL/cortexm0ds_logic.v(1017)
  wire Isiiu6;  // ../RTL/cortexm0ds_logic.v(555)
  wire Isjow6;  // ../RTL/cortexm0ds_logic.v(1111)
  wire Isjpw6;  // ../RTL/cortexm0ds_logic.v(1587)
  wire Ispiu6;  // ../RTL/cortexm0ds_logic.v(648)
  wire Isqhu6;  // ../RTL/cortexm0ds_logic.v(180)
  wire Isqow6;  // ../RTL/cortexm0ds_logic.v(1205)
  wire Iswiu6;  // ../RTL/cortexm0ds_logic.v(742)
  wire Isxhu6;  // ../RTL/cortexm0ds_logic.v(274)
  wire Isxow6;  // ../RTL/cortexm0ds_logic.v(1298)
  wire It2ju6;  // ../RTL/cortexm0ds_logic.v(822)
  wire It3iu6;  // ../RTL/cortexm0ds_logic.v(354)
  wire It3pw6;  // ../RTL/cortexm0ds_logic.v(1379)
  wire It9ju6;  // ../RTL/cortexm0ds_logic.v(916)
  wire Itaiu6;  // ../RTL/cortexm0ds_logic.v(448)
  wire Itapw6;  // ../RTL/cortexm0ds_logic.v(1472)
  wire Itbow6;  // ../RTL/cortexm0ds_logic.v(1004)
  wire Itcbx6;  // ../RTL/cortexm0ds_logic.v(1702)
  wire Ithiu6;  // ../RTL/cortexm0ds_logic.v(542)
  wire Itiow6;  // ../RTL/cortexm0ds_logic.v(1098)
  wire Itoiu6;  // ../RTL/cortexm0ds_logic.v(635)
  wire Itphu6;  // ../RTL/cortexm0ds_logic.v(167)
  wire Itpow6;  // ../RTL/cortexm0ds_logic.v(1192)
  wire Itviu6;  // ../RTL/cortexm0ds_logic.v(729)
  wire Itwhu6;  // ../RTL/cortexm0ds_logic.v(261)
  wire Itwow6;  // ../RTL/cortexm0ds_logic.v(1285)
  wire Iu1ju6;  // ../RTL/cortexm0ds_logic.v(809)
  wire Iu2iu6;  // ../RTL/cortexm0ds_logic.v(341)
  wire Iu2pw6;  // ../RTL/cortexm0ds_logic.v(1366)
  wire Iu8ju6;  // ../RTL/cortexm0ds_logic.v(903)
  wire Iu9iu6;  // ../RTL/cortexm0ds_logic.v(435)
  wire Iu9pw6;  // ../RTL/cortexm0ds_logic.v(1459)
  wire Iuaow6;  // ../RTL/cortexm0ds_logic.v(991)
  wire Iugiu6;  // ../RTL/cortexm0ds_logic.v(529)
  wire Iuhow6;  // ../RTL/cortexm0ds_logic.v(1085)
  wire Iuniu6;  // ../RTL/cortexm0ds_logic.v(622)
  wire Iuohu6;  // ../RTL/cortexm0ds_logic.v(154)
  wire Iuoow6;  // ../RTL/cortexm0ds_logic.v(1179)
  wire Iuuiu6;  // ../RTL/cortexm0ds_logic.v(716)
  wire Iuvhu6;  // ../RTL/cortexm0ds_logic.v(248)
  wire Iuvow6;  // ../RTL/cortexm0ds_logic.v(1272)
  wire Iv0ju6;  // ../RTL/cortexm0ds_logic.v(796)
  wire Iv1iu6;  // ../RTL/cortexm0ds_logic.v(328)
  wire Iv1pw6;  // ../RTL/cortexm0ds_logic.v(1353)
  wire Iv7ju6;  // ../RTL/cortexm0ds_logic.v(890)
  wire Iv8iu6;  // ../RTL/cortexm0ds_logic.v(422)
  wire Iv8pw6;  // ../RTL/cortexm0ds_logic.v(1446)
  wire Iv9ow6;  // ../RTL/cortexm0ds_logic.v(978)
  wire Ivfhu6;  // ../RTL/cortexm0ds_logic.v(125)
  wire Ivfiu6;  // ../RTL/cortexm0ds_logic.v(516)
  wire Ivgow6;  // ../RTL/cortexm0ds_logic.v(1072)
  wire Ivmiu6;  // ../RTL/cortexm0ds_logic.v(609)
  wire Ivnow6;  // ../RTL/cortexm0ds_logic.v(1166)
  wire Ivtiu6;  // ../RTL/cortexm0ds_logic.v(703)
  wire Ivuhu6;  // ../RTL/cortexm0ds_logic.v(235)
  wire Ivuow6;  // ../RTL/cortexm0ds_logic.v(1259)
  wire Iw0iu6;  // ../RTL/cortexm0ds_logic.v(315)
  wire Iw0pw6;  // ../RTL/cortexm0ds_logic.v(1340)
  wire Iw6ju6;  // ../RTL/cortexm0ds_logic.v(877)
  wire Iw7iu6;  // ../RTL/cortexm0ds_logic.v(409)
  wire Iw7pw6;  // ../RTL/cortexm0ds_logic.v(1433)
  wire Iw8ow6;  // ../RTL/cortexm0ds_logic.v(965)
  wire Iweiu6;  // ../RTL/cortexm0ds_logic.v(503)
  wire Iwfow6;  // ../RTL/cortexm0ds_logic.v(1059)
  wire Iwliu6;  // ../RTL/cortexm0ds_logic.v(596)
  wire Iwmow6;  // ../RTL/cortexm0ds_logic.v(1153)
  wire Iwsax6;  // ../RTL/cortexm0ds_logic.v(1667)
  wire Iwsiu6;  // ../RTL/cortexm0ds_logic.v(690)
  wire Iwthu6;  // ../RTL/cortexm0ds_logic.v(222)
  wire Iwtow6;  // ../RTL/cortexm0ds_logic.v(1246)
  wire Iwziu6;  // ../RTL/cortexm0ds_logic.v(783)
  wire Ix5ju6;  // ../RTL/cortexm0ds_logic.v(864)
  wire Ix6iu6;  // ../RTL/cortexm0ds_logic.v(396)
  wire Ix6pw6;  // ../RTL/cortexm0ds_logic.v(1420)
  wire Ix7ow6;  // ../RTL/cortexm0ds_logic.v(952)
  wire Ixdiu6;  // ../RTL/cortexm0ds_logic.v(490)
  wire Ixdpw6;  // ../RTL/cortexm0ds_logic.v(1514)
  wire Ixeow6;  // ../RTL/cortexm0ds_logic.v(1046)
  wire Ixkiu6;  // ../RTL/cortexm0ds_logic.v(583)
  wire Ixlow6;  // ../RTL/cortexm0ds_logic.v(1140)
  wire Ixppw6;  // ../RTL/cortexm0ds_logic.v(1599)
  wire Ixriu6;  // ../RTL/cortexm0ds_logic.v(677)
  wire Ixshu6;  // ../RTL/cortexm0ds_logic.v(209)
  wire Ixsow6;  // ../RTL/cortexm0ds_logic.v(1233)
  wire Ixyiu6;  // ../RTL/cortexm0ds_logic.v(770)
  wire Ixzhu6;  // ../RTL/cortexm0ds_logic.v(302)
  wire Ixzow6;  // ../RTL/cortexm0ds_logic.v(1327)
  wire Iy4ju6;  // ../RTL/cortexm0ds_logic.v(851)
  wire Iy5iu6;  // ../RTL/cortexm0ds_logic.v(383)
  wire Iy5pw6;  // ../RTL/cortexm0ds_logic.v(1407)
  wire Iy6ow6;  // ../RTL/cortexm0ds_logic.v(939)
  wire Iyciu6;  // ../RTL/cortexm0ds_logic.v(477)
  wire Iycpw6;  // ../RTL/cortexm0ds_logic.v(1501)
  wire Iydow6;  // ../RTL/cortexm0ds_logic.v(1033)
  wire Iyjiu6;  // ../RTL/cortexm0ds_logic.v(570)
  wire Iykow6;  // ../RTL/cortexm0ds_logic.v(1127)
  wire Iyqiu6;  // ../RTL/cortexm0ds_logic.v(664)
  wire Iyrhu6;  // ../RTL/cortexm0ds_logic.v(196)
  wire Iyrow6;  // ../RTL/cortexm0ds_logic.v(1220)
  wire Iyxiu6;  // ../RTL/cortexm0ds_logic.v(757)
  wire Iyyhu6;  // ../RTL/cortexm0ds_logic.v(289)
  wire Iyyow6;  // ../RTL/cortexm0ds_logic.v(1314)
  wire Iz3ju6;  // ../RTL/cortexm0ds_logic.v(838)
  wire Iz4iu6;  // ../RTL/cortexm0ds_logic.v(370)
  wire Iz4pw6;  // ../RTL/cortexm0ds_logic.v(1394)
  wire Izbiu6;  // ../RTL/cortexm0ds_logic.v(464)
  wire Izbpw6;  // ../RTL/cortexm0ds_logic.v(1488)
  wire Izcow6;  // ../RTL/cortexm0ds_logic.v(1020)
  wire Iziiu6;  // ../RTL/cortexm0ds_logic.v(557)
  wire Izjow6;  // ../RTL/cortexm0ds_logic.v(1114)
  wire Izpiu6;  // ../RTL/cortexm0ds_logic.v(651)
  wire Izppw6;  // ../RTL/cortexm0ds_logic.v(1599)
  wire Izqhu6;  // ../RTL/cortexm0ds_logic.v(183)
  wire Izqow6;  // ../RTL/cortexm0ds_logic.v(1207)
  wire Izwiu6;  // ../RTL/cortexm0ds_logic.v(744)
  wire Izxhu6;  // ../RTL/cortexm0ds_logic.v(276)
  wire Izxow6;  // ../RTL/cortexm0ds_logic.v(1301)
  wire J00ju6;  // ../RTL/cortexm0ds_logic.v(785)
  wire J01iu6;  // ../RTL/cortexm0ds_logic.v(317)
  wire J01pw6;  // ../RTL/cortexm0ds_logic.v(1341)
  wire J06bx6;  // ../RTL/cortexm0ds_logic.v(1690)
  wire J07ju6;  // ../RTL/cortexm0ds_logic.v(878)
  wire J08iu6;  // ../RTL/cortexm0ds_logic.v(410)
  wire J08pw6;  // ../RTL/cortexm0ds_logic.v(1435)
  wire J09ow6;  // ../RTL/cortexm0ds_logic.v(967)
  wire J0fiu6;  // ../RTL/cortexm0ds_logic.v(504)
  wire J0gax6;  // ../RTL/cortexm0ds_logic.v(1643)
  wire J0gow6;  // ../RTL/cortexm0ds_logic.v(1060)
  wire J0iax6;  // ../RTL/cortexm0ds_logic.v(1647)
  wire J0miu6;  // ../RTL/cortexm0ds_logic.v(598)
  wire J0now6;  // ../RTL/cortexm0ds_logic.v(1154)
  wire J0tiu6;  // ../RTL/cortexm0ds_logic.v(691)
  wire J0uhu6;  // ../RTL/cortexm0ds_logic.v(223)
  wire J0uow6;  // ../RTL/cortexm0ds_logic.v(1248)
  wire J10iu6;  // ../RTL/cortexm0ds_logic.v(304)
  wire J10pw6;  // ../RTL/cortexm0ds_logic.v(1328)
  wire J16ju6;  // ../RTL/cortexm0ds_logic.v(865)
  wire J17iu6;  // ../RTL/cortexm0ds_logic.v(397)
  wire J17pw6;  // ../RTL/cortexm0ds_logic.v(1422)
  wire J18ow6;  // ../RTL/cortexm0ds_logic.v(954)
  wire J1eiu6;  // ../RTL/cortexm0ds_logic.v(491)
  wire J1epw6;  // ../RTL/cortexm0ds_logic.v(1515)
  wire J1fow6;  // ../RTL/cortexm0ds_logic.v(1047)
  wire J1liu6;  // ../RTL/cortexm0ds_logic.v(585)
  wire J1mow6;  // ../RTL/cortexm0ds_logic.v(1141)
  wire J1siu6;  // ../RTL/cortexm0ds_logic.v(678)
  wire J1thu6;  // ../RTL/cortexm0ds_logic.v(210)
  wire J1tow6;  // ../RTL/cortexm0ds_logic.v(1235)
  wire J1ziu6;  // ../RTL/cortexm0ds_logic.v(772)
  wire J25ju6;  // ../RTL/cortexm0ds_logic.v(852)
  wire J26iu6;  // ../RTL/cortexm0ds_logic.v(384)
  wire J26pw6;  // ../RTL/cortexm0ds_logic.v(1409)
  wire J27ow6;  // ../RTL/cortexm0ds_logic.v(941)
  wire J2diu6;  // ../RTL/cortexm0ds_logic.v(478)
  wire J2dpw6;  // ../RTL/cortexm0ds_logic.v(1502)
  wire J2eow6;  // ../RTL/cortexm0ds_logic.v(1034)
  wire J2kiu6;  // ../RTL/cortexm0ds_logic.v(572)
  wire J2low6;  // ../RTL/cortexm0ds_logic.v(1128)
  wire J2riu6;  // ../RTL/cortexm0ds_logic.v(665)
  wire J2shu6;  // ../RTL/cortexm0ds_logic.v(197)
  wire J2sow6;  // ../RTL/cortexm0ds_logic.v(1222)
  wire J2yiu6;  // ../RTL/cortexm0ds_logic.v(759)
  wire J2zhu6;  // ../RTL/cortexm0ds_logic.v(291)
  wire J2zow6;  // ../RTL/cortexm0ds_logic.v(1315)
  wire J34ju6;  // ../RTL/cortexm0ds_logic.v(839)
  wire J35iu6;  // ../RTL/cortexm0ds_logic.v(371)
  wire J35pw6;  // ../RTL/cortexm0ds_logic.v(1396)
  wire J39bx6;  // ../RTL/cortexm0ds_logic.v(1695)
  wire J3ciu6;  // ../RTL/cortexm0ds_logic.v(465)
  wire J3cpw6;  // ../RTL/cortexm0ds_logic.v(1489)
  wire J3dow6;  // ../RTL/cortexm0ds_logic.v(1021)
  wire J3jiu6;  // ../RTL/cortexm0ds_logic.v(559)
  wire J3kow6;  // ../RTL/cortexm0ds_logic.v(1115)
  wire J3qiu6;  // ../RTL/cortexm0ds_logic.v(652)
  wire J3rhu6;  // ../RTL/cortexm0ds_logic.v(184)
  wire J3row6;  // ../RTL/cortexm0ds_logic.v(1209)
  wire J3xax6;  // ../RTL/cortexm0ds_logic.v(1674)
  wire J3xiu6;  // ../RTL/cortexm0ds_logic.v(746)
  wire J3yhu6;  // ../RTL/cortexm0ds_logic.v(278)
  wire J3yow6;  // ../RTL/cortexm0ds_logic.v(1302)
  wire J43ju6;  // ../RTL/cortexm0ds_logic.v(826)
  wire J44iu6;  // ../RTL/cortexm0ds_logic.v(358)
  wire J44pw6;  // ../RTL/cortexm0ds_logic.v(1383)
  wire J4aju6;  // ../RTL/cortexm0ds_logic.v(920)
  wire J4biu6;  // ../RTL/cortexm0ds_logic.v(452)
  wire J4bpw6;  // ../RTL/cortexm0ds_logic.v(1476)
  wire J4cbx6;  // ../RTL/cortexm0ds_logic.v(1701)
  wire J4cow6;  // ../RTL/cortexm0ds_logic.v(1008)
  wire J4iiu6;  // ../RTL/cortexm0ds_logic.v(546)
  wire J4jow6;  // ../RTL/cortexm0ds_logic.v(1102)
  wire J4mhu6;  // ../RTL/cortexm0ds_logic.v(141)
  wire J4piu6;  // ../RTL/cortexm0ds_logic.v(639)
  wire J4qhu6;  // ../RTL/cortexm0ds_logic.v(171)
  wire J4qow6;  // ../RTL/cortexm0ds_logic.v(1196)
  wire J4wiu6;  // ../RTL/cortexm0ds_logic.v(733)
  wire J4xhu6;  // ../RTL/cortexm0ds_logic.v(265)
  wire J4xow6;  // ../RTL/cortexm0ds_logic.v(1289)
  wire J52ju6;  // ../RTL/cortexm0ds_logic.v(813)
  wire J53pw6;  // ../RTL/cortexm0ds_logic.v(1370)
  wire J59ax6;  // ../RTL/cortexm0ds_logic.v(1630)
  wire J59ju6;  // ../RTL/cortexm0ds_logic.v(907)
  wire J5aiu6;  // ../RTL/cortexm0ds_logic.v(439)
  wire J5apw6;  // ../RTL/cortexm0ds_logic.v(1463)
  wire J5bow6;  // ../RTL/cortexm0ds_logic.v(995)
  wire J5eax6;  // ../RTL/cortexm0ds_logic.v(1639)
  wire J5hiu6;  // ../RTL/cortexm0ds_logic.v(533)
  wire J5iow6;  // ../RTL/cortexm0ds_logic.v(1089)
  wire J5jbx6;  // ../RTL/cortexm0ds_logic.v(1714)
  wire J5oiu6;  // ../RTL/cortexm0ds_logic.v(626)
  wire J5phu6;  // ../RTL/cortexm0ds_logic.v(158)
  wire J5pow6;  // ../RTL/cortexm0ds_logic.v(1183)
  wire J5viu6;  // ../RTL/cortexm0ds_logic.v(720)
  wire J5whu6;  // ../RTL/cortexm0ds_logic.v(252)
  wire J5wow6;  // ../RTL/cortexm0ds_logic.v(1276)
  wire J61ju6;  // ../RTL/cortexm0ds_logic.v(800)
  wire J62iu6;  // ../RTL/cortexm0ds_logic.v(332)
  wire J62pw6;  // ../RTL/cortexm0ds_logic.v(1357)
  wire J68ju6;  // ../RTL/cortexm0ds_logic.v(894)
  wire J69iu6;  // ../RTL/cortexm0ds_logic.v(426)
  wire J69pw6;  // ../RTL/cortexm0ds_logic.v(1450)
  wire J6aow6;  // ../RTL/cortexm0ds_logic.v(982)
  wire J6ebx6;  // ../RTL/cortexm0ds_logic.v(1705)
  wire J6giu6;  // ../RTL/cortexm0ds_logic.v(520)
  wire J6how6;  // ../RTL/cortexm0ds_logic.v(1076)
  wire J6niu6;  // ../RTL/cortexm0ds_logic.v(613)
  wire J6oow6;  // ../RTL/cortexm0ds_logic.v(1170)
  wire J6uiu6;  // ../RTL/cortexm0ds_logic.v(707)
  wire J6vhu6;  // ../RTL/cortexm0ds_logic.v(239)
  wire J6vow6;  // ../RTL/cortexm0ds_logic.v(1263)
  wire J6zax6;  // ../RTL/cortexm0ds_logic.v(1678)
  wire J70ju6;  // ../RTL/cortexm0ds_logic.v(787)
  wire J71iu6;  // ../RTL/cortexm0ds_logic.v(319)
  wire J71pw6;  // ../RTL/cortexm0ds_logic.v(1344)
  wire J77ju6;  // ../RTL/cortexm0ds_logic.v(881)
  wire J78iu6;  // ../RTL/cortexm0ds_logic.v(413)
  wire J78pw6;  // ../RTL/cortexm0ds_logic.v(1437)
  wire J79ow6;  // ../RTL/cortexm0ds_logic.v(969)
  wire J7fiu6;  // ../RTL/cortexm0ds_logic.v(507)
  wire J7gow6;  // ../RTL/cortexm0ds_logic.v(1063)
  wire J7miu6;  // ../RTL/cortexm0ds_logic.v(600)
  wire J7now6;  // ../RTL/cortexm0ds_logic.v(1157)
  wire J7tiu6;  // ../RTL/cortexm0ds_logic.v(694)
  wire J7uhu6;  // ../RTL/cortexm0ds_logic.v(226)
  wire J7uow6;  // ../RTL/cortexm0ds_logic.v(1250)
  wire J7xax6;  // ../RTL/cortexm0ds_logic.v(1674)
  wire J80iu6;  // ../RTL/cortexm0ds_logic.v(306)
  wire J80pw6;  // ../RTL/cortexm0ds_logic.v(1331)
  wire J86ju6;  // ../RTL/cortexm0ds_logic.v(868)
  wire J87iu6;  // ../RTL/cortexm0ds_logic.v(400)
  wire J87pw6;  // ../RTL/cortexm0ds_logic.v(1424)
  wire J88ow6;  // ../RTL/cortexm0ds_logic.v(956)
  wire J8cax6;  // ../RTL/cortexm0ds_logic.v(1636)
  wire J8eiu6;  // ../RTL/cortexm0ds_logic.v(494)
  wire J8fow6;  // ../RTL/cortexm0ds_logic.v(1050)
  wire J8liu6;  // ../RTL/cortexm0ds_logic.v(587)
  wire J8mow6;  // ../RTL/cortexm0ds_logic.v(1144)
  wire J8siu6;  // ../RTL/cortexm0ds_logic.v(681)
  wire J8thu6;  // ../RTL/cortexm0ds_logic.v(213)
  wire J8tow6;  // ../RTL/cortexm0ds_logic.v(1237)
  wire J8ziu6;  // ../RTL/cortexm0ds_logic.v(774)
  wire J95ju6;  // ../RTL/cortexm0ds_logic.v(855)
  wire J96iu6;  // ../RTL/cortexm0ds_logic.v(387)
  wire J96pw6;  // ../RTL/cortexm0ds_logic.v(1411)
  wire J97ow6;  // ../RTL/cortexm0ds_logic.v(943)
  wire J9diu6;  // ../RTL/cortexm0ds_logic.v(481)
  wire J9dpw6;  // ../RTL/cortexm0ds_logic.v(1505)
  wire J9eow6;  // ../RTL/cortexm0ds_logic.v(1037)
  wire J9kiu6;  // ../RTL/cortexm0ds_logic.v(574)
  wire J9low6;  // ../RTL/cortexm0ds_logic.v(1131)
  wire J9riu6;  // ../RTL/cortexm0ds_logic.v(668)
  wire J9shu6;  // ../RTL/cortexm0ds_logic.v(200)
  wire J9sow6;  // ../RTL/cortexm0ds_logic.v(1224)
  wire J9yiu6;  // ../RTL/cortexm0ds_logic.v(761)
  wire J9zhu6;  // ../RTL/cortexm0ds_logic.v(293)
  wire J9zow6;  // ../RTL/cortexm0ds_logic.v(1318)
  wire Ja4ju6;  // ../RTL/cortexm0ds_logic.v(842)
  wire Ja5iu6;  // ../RTL/cortexm0ds_logic.v(374)
  wire Ja5pw6;  // ../RTL/cortexm0ds_logic.v(1398)
  wire Ja6ow6;  // ../RTL/cortexm0ds_logic.v(930)
  wire Jaciu6;  // ../RTL/cortexm0ds_logic.v(468)
  wire Jacpw6;  // ../RTL/cortexm0ds_logic.v(1492)
  wire Jadow6;  // ../RTL/cortexm0ds_logic.v(1024)
  wire Jajiu6;  // ../RTL/cortexm0ds_logic.v(561)
  wire Jakow6;  // ../RTL/cortexm0ds_logic.v(1118)
  wire Jaqiu6;  // ../RTL/cortexm0ds_logic.v(655)
  wire Jarhu6;  // ../RTL/cortexm0ds_logic.v(187)
  wire Jarow6;  // ../RTL/cortexm0ds_logic.v(1211)
  wire Jaxiu6;  // ../RTL/cortexm0ds_logic.v(748)
  wire Jayhu6;  // ../RTL/cortexm0ds_logic.v(280)
  wire Jayow6;  // ../RTL/cortexm0ds_logic.v(1305)
  wire Jb3ju6;  // ../RTL/cortexm0ds_logic.v(829)
  wire Jb4iu6;  // ../RTL/cortexm0ds_logic.v(361)
  wire Jb4pw6;  // ../RTL/cortexm0ds_logic.v(1385)
  wire Jbaju6;  // ../RTL/cortexm0ds_logic.v(923)
  wire Jbbiu6;  // ../RTL/cortexm0ds_logic.v(455)
  wire Jbbpw6;  // ../RTL/cortexm0ds_logic.v(1479)
  wire Jbcow6;  // ../RTL/cortexm0ds_logic.v(1011)
  wire Jbiiu6;  // ../RTL/cortexm0ds_logic.v(548)
  wire Jbjow6;  // ../RTL/cortexm0ds_logic.v(1105)
  wire Jbpiu6;  // ../RTL/cortexm0ds_logic.v(642)
  wire Jbqhu6;  // ../RTL/cortexm0ds_logic.v(174)
  wire Jbqow6;  // ../RTL/cortexm0ds_logic.v(1198)
  wire Jbwiu6;  // ../RTL/cortexm0ds_logic.v(735)
  wire Jbxhu6;  // ../RTL/cortexm0ds_logic.v(267)
  wire Jbxow6;  // ../RTL/cortexm0ds_logic.v(1292)
  wire Jc2ju6;  // ../RTL/cortexm0ds_logic.v(816)
  wire Jc3iu6;  // ../RTL/cortexm0ds_logic.v(348)
  wire Jc3pw6;  // ../RTL/cortexm0ds_logic.v(1372)
  wire Jc9ju6;  // ../RTL/cortexm0ds_logic.v(910)
  wire Jcaiu6;  // ../RTL/cortexm0ds_logic.v(442)
  wire Jcapw6;  // ../RTL/cortexm0ds_logic.v(1466)
  wire Jcbow6;  // ../RTL/cortexm0ds_logic.v(998)
  wire Jchiu6;  // ../RTL/cortexm0ds_logic.v(535)
  wire Jciow6;  // ../RTL/cortexm0ds_logic.v(1092)
  wire Jckax6;  // ../RTL/cortexm0ds_logic.v(1651)
  wire Jcoiu6;  // ../RTL/cortexm0ds_logic.v(629)
  wire Jcphu6;  // ../RTL/cortexm0ds_logic.v(161)
  wire Jcpow6;  // ../RTL/cortexm0ds_logic.v(1185)
  wire Jcviu6;  // ../RTL/cortexm0ds_logic.v(722)
  wire Jcwhu6;  // ../RTL/cortexm0ds_logic.v(254)
  wire Jcwow6;  // ../RTL/cortexm0ds_logic.v(1279)
  wire Jd1ju6;  // ../RTL/cortexm0ds_logic.v(803)
  wire Jd2iu6;  // ../RTL/cortexm0ds_logic.v(335)
  wire Jd2pw6;  // ../RTL/cortexm0ds_logic.v(1359)
  wire Jd8ju6;  // ../RTL/cortexm0ds_logic.v(897)
  wire Jd9iu6;  // ../RTL/cortexm0ds_logic.v(429)
  wire Jd9pw6;  // ../RTL/cortexm0ds_logic.v(1453)
  wire Jdaow6;  // ../RTL/cortexm0ds_logic.v(985)
  wire Jdgbx6;  // ../RTL/cortexm0ds_logic.v(1709)
  wire Jdgiu6;  // ../RTL/cortexm0ds_logic.v(522)
  wire Jdhow6;  // ../RTL/cortexm0ds_logic.v(1079)
  wire Jdnhu6;  // ../RTL/cortexm0ds_logic.v(144)
  wire Jdniu6;  // ../RTL/cortexm0ds_logic.v(616)
  wire Jdohu6;  // ../RTL/cortexm0ds_logic.v(148)
  wire Jdoow6;  // ../RTL/cortexm0ds_logic.v(1172)
  wire Jduiu6;  // ../RTL/cortexm0ds_logic.v(709)
  wire Jdvhu6;  // ../RTL/cortexm0ds_logic.v(241)
  wire Jdvow6;  // ../RTL/cortexm0ds_logic.v(1266)
  wire Je0ju6;  // ../RTL/cortexm0ds_logic.v(790)
  wire Je1iu6;  // ../RTL/cortexm0ds_logic.v(322)
  wire Je1pw6;  // ../RTL/cortexm0ds_logic.v(1346)
  wire Je7ju6;  // ../RTL/cortexm0ds_logic.v(884)
  wire Je8iu6;  // ../RTL/cortexm0ds_logic.v(416)
  wire Je8pw6;  // ../RTL/cortexm0ds_logic.v(1440)
  wire Je9ow6;  // ../RTL/cortexm0ds_logic.v(972)
  wire Jefiu6;  // ../RTL/cortexm0ds_logic.v(509)
  wire Jegow6;  // ../RTL/cortexm0ds_logic.v(1066)
  wire Jehhu6;  // ../RTL/cortexm0ds_logic.v(128)
  wire Jemiu6;  // ../RTL/cortexm0ds_logic.v(603)
  wire Jenow6;  // ../RTL/cortexm0ds_logic.v(1159)
  wire Jetiu6;  // ../RTL/cortexm0ds_logic.v(696)
  wire Jeuhu6;  // ../RTL/cortexm0ds_logic.v(228)
  wire Jeuow6;  // ../RTL/cortexm0ds_logic.v(1253)
  wire Jf0iu6;  // ../RTL/cortexm0ds_logic.v(309)
  wire Jf0pw6;  // ../RTL/cortexm0ds_logic.v(1333)
  wire Jf6ju6;  // ../RTL/cortexm0ds_logic.v(871)
  wire Jf7iu6;  // ../RTL/cortexm0ds_logic.v(403)
  wire Jf7pw6;  // ../RTL/cortexm0ds_logic.v(1427)
  wire Jf8ow6;  // ../RTL/cortexm0ds_logic.v(959)
  wire Jfdbx6;  // ../RTL/cortexm0ds_logic.v(1703)
  wire Jfeiu6;  // ../RTL/cortexm0ds_logic.v(496)
  wire Jffow6;  // ../RTL/cortexm0ds_logic.v(1053)
  wire Jfliu6;  // ../RTL/cortexm0ds_logic.v(590)
  wire Jflpw6;  // ../RTL/cortexm0ds_logic.v(1590)
  wire Jfmow6;  // ../RTL/cortexm0ds_logic.v(1146)
  wire Jfsiu6;  // ../RTL/cortexm0ds_logic.v(683)
  wire Jfthu6;  // ../RTL/cortexm0ds_logic.v(215)
  wire Jftow6;  // ../RTL/cortexm0ds_logic.v(1240)
  wire Jfziu6;  // ../RTL/cortexm0ds_logic.v(777)
  wire Jg5ju6;  // ../RTL/cortexm0ds_logic.v(858)
  wire Jg6iu6;  // ../RTL/cortexm0ds_logic.v(390)
  wire Jg6pw6;  // ../RTL/cortexm0ds_logic.v(1414)
  wire Jg7ow6;  // ../RTL/cortexm0ds_logic.v(946)
  wire Jgdiu6;  // ../RTL/cortexm0ds_logic.v(483)
  wire Jgdpw6;  // ../RTL/cortexm0ds_logic.v(1508)
  wire Jgeow6;  // ../RTL/cortexm0ds_logic.v(1040)
  wire Jgkiu6;  // ../RTL/cortexm0ds_logic.v(577)
  wire Jglow6;  // ../RTL/cortexm0ds_logic.v(1133)
  wire Jgriu6;  // ../RTL/cortexm0ds_logic.v(670)
  wire Jgshu6;  // ../RTL/cortexm0ds_logic.v(202)
  wire Jgsow6;  // ../RTL/cortexm0ds_logic.v(1227)
  wire Jgxpw6;  // ../RTL/cortexm0ds_logic.v(1612)
  wire Jgyiu6;  // ../RTL/cortexm0ds_logic.v(764)
  wire Jgzhu6;  // ../RTL/cortexm0ds_logic.v(296)
  wire Jgzow6;  // ../RTL/cortexm0ds_logic.v(1320)
  wire Jh4ju6;  // ../RTL/cortexm0ds_logic.v(845)
  wire Jh5iu6;  // ../RTL/cortexm0ds_logic.v(377)
  wire Jh5pw6;  // ../RTL/cortexm0ds_logic.v(1401)
  wire Jh6ow6;  // ../RTL/cortexm0ds_logic.v(933)
  wire Jhciu6;  // ../RTL/cortexm0ds_logic.v(470)
  wire Jhcpw6;  // ../RTL/cortexm0ds_logic.v(1495)
  wire Jhdow6;  // ../RTL/cortexm0ds_logic.v(1027)
  wire Jhebx6;  // ../RTL/cortexm0ds_logic.v(1705)
  wire Jhjiu6;  // ../RTL/cortexm0ds_logic.v(564)
  wire Jhkow6;  // ../RTL/cortexm0ds_logic.v(1120)
  wire Jhqiu6;  // ../RTL/cortexm0ds_logic.v(657)
  wire Jhrhu6;  // ../RTL/cortexm0ds_logic.v(189)
  wire Jhrow6;  // ../RTL/cortexm0ds_logic.v(1214)
  wire Jhxiu6;  // ../RTL/cortexm0ds_logic.v(751)
  wire Jhyhu6;  // ../RTL/cortexm0ds_logic.v(283)
  wire Jhyow6;  // ../RTL/cortexm0ds_logic.v(1307)
  wire Ji3ju6;  // ../RTL/cortexm0ds_logic.v(832)
  wire Ji4iu6;  // ../RTL/cortexm0ds_logic.v(364)
  wire Ji4pw6;  // ../RTL/cortexm0ds_logic.v(1388)
  wire Jiaju6;  // ../RTL/cortexm0ds_logic.v(925)
  wire Jibiu6;  // ../RTL/cortexm0ds_logic.v(457)
  wire Jibpw6;  // ../RTL/cortexm0ds_logic.v(1482)
  wire Jicow6;  // ../RTL/cortexm0ds_logic.v(1014)
  wire Jieax6;  // ../RTL/cortexm0ds_logic.v(1640)
  wire Jiiiu6;  // ../RTL/cortexm0ds_logic.v(551)
  wire Jijow6;  // ../RTL/cortexm0ds_logic.v(1107)
  wire Jipiu6;  // ../RTL/cortexm0ds_logic.v(644)
  wire Jiqhu6;  // ../RTL/cortexm0ds_logic.v(176)
  wire Jiqow6;  // ../RTL/cortexm0ds_logic.v(1201)
  wire Jiwiu6;  // ../RTL/cortexm0ds_logic.v(738)
  wire Jixhu6;  // ../RTL/cortexm0ds_logic.v(270)
  wire Jixow6;  // ../RTL/cortexm0ds_logic.v(1294)
  wire Jj0bx6;  // ../RTL/cortexm0ds_logic.v(1680)
  wire Jj2ju6;  // ../RTL/cortexm0ds_logic.v(819)
  wire Jj3iu6;  // ../RTL/cortexm0ds_logic.v(351)
  wire Jj3pw6;  // ../RTL/cortexm0ds_logic.v(1375)
  wire Jj9ju6;  // ../RTL/cortexm0ds_logic.v(912)
  wire Jjaiu6;  // ../RTL/cortexm0ds_logic.v(444)
  wire Jjapw6;  // ../RTL/cortexm0ds_logic.v(1469)
  wire Jjbow6;  // ../RTL/cortexm0ds_logic.v(1001)
  wire Jjhiu6;  // ../RTL/cortexm0ds_logic.v(538)
  wire Jjiow6;  // ../RTL/cortexm0ds_logic.v(1094)
  wire Jjoiu6;  // ../RTL/cortexm0ds_logic.v(631)
  wire Jjphu6;  // ../RTL/cortexm0ds_logic.v(163)
  wire Jjpow6;  // ../RTL/cortexm0ds_logic.v(1188)
  wire Jjviu6;  // ../RTL/cortexm0ds_logic.v(725)
  wire Jjvpw6;  // ../RTL/cortexm0ds_logic.v(1609)
  wire Jjwhu6;  // ../RTL/cortexm0ds_logic.v(257)
  wire Jjwow6;  // ../RTL/cortexm0ds_logic.v(1281)
  wire Jk1ju6;  // ../RTL/cortexm0ds_logic.v(806)
  wire Jk2iu6;  // ../RTL/cortexm0ds_logic.v(338)
  wire Jk2pw6;  // ../RTL/cortexm0ds_logic.v(1362)
  wire Jk8ju6;  // ../RTL/cortexm0ds_logic.v(899)
  wire Jk9iu6;  // ../RTL/cortexm0ds_logic.v(431)
  wire Jk9pw6;  // ../RTL/cortexm0ds_logic.v(1456)
  wire Jkaow6;  // ../RTL/cortexm0ds_logic.v(988)
  wire Jkgiu6;  // ../RTL/cortexm0ds_logic.v(525)
  wire Jkhow6;  // ../RTL/cortexm0ds_logic.v(1081)
  wire Jkniu6;  // ../RTL/cortexm0ds_logic.v(618)
  wire Jkohu6;  // ../RTL/cortexm0ds_logic.v(150)
  wire Jkoow6;  // ../RTL/cortexm0ds_logic.v(1175)
  wire Jkuiu6;  // ../RTL/cortexm0ds_logic.v(712)
  wire Jkvhu6;  // ../RTL/cortexm0ds_logic.v(244)
  wire Jkvow6;  // ../RTL/cortexm0ds_logic.v(1268)
  wire Jl0ju6;  // ../RTL/cortexm0ds_logic.v(793)
  wire Jl1iu6;  // ../RTL/cortexm0ds_logic.v(325)
  wire Jl1pw6;  // ../RTL/cortexm0ds_logic.v(1349)
  wire Jl3qw6;  // ../RTL/cortexm0ds_logic.v(1624)
  wire Jl7ju6;  // ../RTL/cortexm0ds_logic.v(886)
  wire Jl8iu6;  // ../RTL/cortexm0ds_logic.v(418)
  wire Jl8pw6;  // ../RTL/cortexm0ds_logic.v(1443)
  wire Jl9ow6;  // ../RTL/cortexm0ds_logic.v(975)
  wire Jlfiu6;  // ../RTL/cortexm0ds_logic.v(512)
  wire Jlgow6;  // ../RTL/cortexm0ds_logic.v(1068)
  wire Jlmiu6;  // ../RTL/cortexm0ds_logic.v(605)
  wire Jlnow6;  // ../RTL/cortexm0ds_logic.v(1162)
  wire Jltiu6;  // ../RTL/cortexm0ds_logic.v(699)
  wire Jluhu6;  // ../RTL/cortexm0ds_logic.v(231)
  wire Jluow6;  // ../RTL/cortexm0ds_logic.v(1255)
  wire Jlvpw6;  // ../RTL/cortexm0ds_logic.v(1609)
  wire Jm0iu6;  // ../RTL/cortexm0ds_logic.v(312)
  wire Jm0pw6;  // ../RTL/cortexm0ds_logic.v(1336)
  wire Jm6ju6;  // ../RTL/cortexm0ds_logic.v(873)
  wire Jm7iu6;  // ../RTL/cortexm0ds_logic.v(405)
  wire Jm7pw6;  // ../RTL/cortexm0ds_logic.v(1430)
  wire Jm8ow6;  // ../RTL/cortexm0ds_logic.v(962)
  wire Jmeiu6;  // ../RTL/cortexm0ds_logic.v(499)
  wire Jmfow6;  // ../RTL/cortexm0ds_logic.v(1055)
  wire Jmliu6;  // ../RTL/cortexm0ds_logic.v(592)
  wire Jmmow6;  // ../RTL/cortexm0ds_logic.v(1149)
  wire Jmsiu6;  // ../RTL/cortexm0ds_logic.v(686)
  wire Jmthu6;  // ../RTL/cortexm0ds_logic.v(218)
  wire Jmtow6;  // ../RTL/cortexm0ds_logic.v(1242)
  wire Jmziu6;  // ../RTL/cortexm0ds_logic.v(780)
  wire Jn5ju6;  // ../RTL/cortexm0ds_logic.v(860)
  wire Jn6iu6;  // ../RTL/cortexm0ds_logic.v(392)
  wire Jn6pw6;  // ../RTL/cortexm0ds_logic.v(1417)
  wire Jn7ow6;  // ../RTL/cortexm0ds_logic.v(949)
  wire Jndiu6;  // ../RTL/cortexm0ds_logic.v(486)
  wire Jndpw6;  // ../RTL/cortexm0ds_logic.v(1510)
  wire Jneow6;  // ../RTL/cortexm0ds_logic.v(1042)
  wire Jnkiu6;  // ../RTL/cortexm0ds_logic.v(579)
  wire Jnlow6;  // ../RTL/cortexm0ds_logic.v(1136)
  wire Jnoax6;  // ../RTL/cortexm0ds_logic.v(1659)
  wire Jnriu6;  // ../RTL/cortexm0ds_logic.v(673)
  wire Jnshu6;  // ../RTL/cortexm0ds_logic.v(205)
  wire Jnsow6;  // ../RTL/cortexm0ds_logic.v(1229)
  wire Jnvpw6;  // ../RTL/cortexm0ds_logic.v(1609)
  wire Jnyiu6;  // ../RTL/cortexm0ds_logic.v(767)
  wire Jnzhu6;  // ../RTL/cortexm0ds_logic.v(299)
  wire Jnzow6;  // ../RTL/cortexm0ds_logic.v(1323)
  wire Jo4ju6;  // ../RTL/cortexm0ds_logic.v(847)
  wire Jo5iu6;  // ../RTL/cortexm0ds_logic.v(379)
  wire Jo5pw6;  // ../RTL/cortexm0ds_logic.v(1404)
  wire Jo6ow6;  // ../RTL/cortexm0ds_logic.v(936)
  wire Jociu6;  // ../RTL/cortexm0ds_logic.v(473)
  wire Jocpw6;  // ../RTL/cortexm0ds_logic.v(1497)
  wire Jodow6;  // ../RTL/cortexm0ds_logic.v(1029)
  wire Johbx6;  // ../RTL/cortexm0ds_logic.v(1711)
  wire Jojiu6;  // ../RTL/cortexm0ds_logic.v(566)
  wire Jokow6;  // ../RTL/cortexm0ds_logic.v(1123)
  wire Joqiu6;  // ../RTL/cortexm0ds_logic.v(660)
  wire Jorhu6;  // ../RTL/cortexm0ds_logic.v(192)
  wire Jorow6;  // ../RTL/cortexm0ds_logic.v(1216)
  wire Joxiu6;  // ../RTL/cortexm0ds_logic.v(754)
  wire Joyhu6;  // ../RTL/cortexm0ds_logic.v(286)
  wire Joyow6;  // ../RTL/cortexm0ds_logic.v(1310)
  wire Jp1qw6;  // ../RTL/cortexm0ds_logic.v(1620)
  wire Jp3ju6;  // ../RTL/cortexm0ds_logic.v(834)
  wire Jp4iu6;  // ../RTL/cortexm0ds_logic.v(366)
  wire Jp4pw6;  // ../RTL/cortexm0ds_logic.v(1391)
  wire Jp9bx6;  // ../RTL/cortexm0ds_logic.v(1697)
  wire Jpaju6;  // ../RTL/cortexm0ds_logic.v(928)
  wire Jpbiu6;  // ../RTL/cortexm0ds_logic.v(460)
  wire Jpbpw6;  // ../RTL/cortexm0ds_logic.v(1484)
  wire Jpcow6;  // ../RTL/cortexm0ds_logic.v(1016)
  wire Jpiiu6;  // ../RTL/cortexm0ds_logic.v(553)
  wire Jpjow6;  // ../RTL/cortexm0ds_logic.v(1110)
  wire Jpmpw6;  // ../RTL/cortexm0ds_logic.v(1593)
  wire Jppiu6;  // ../RTL/cortexm0ds_logic.v(647)
  wire Jpqhu6;  // ../RTL/cortexm0ds_logic.v(179)
  wire Jpqow6;  // ../RTL/cortexm0ds_logic.v(1203)
  wire Jpvpw6;  // ../RTL/cortexm0ds_logic.v(1609)
  wire Jpwiu6;  // ../RTL/cortexm0ds_logic.v(741)
  wire Jpxhu6;  // ../RTL/cortexm0ds_logic.v(273)
  wire Jpxow6;  // ../RTL/cortexm0ds_logic.v(1297)
  wire Jq2ju6;  // ../RTL/cortexm0ds_logic.v(821)
  wire Jq3iu6;  // ../RTL/cortexm0ds_logic.v(353)
  wire Jq3pw6;  // ../RTL/cortexm0ds_logic.v(1378)
  wire Jq9ju6;  // ../RTL/cortexm0ds_logic.v(915)
  wire Jqaiu6;  // ../RTL/cortexm0ds_logic.v(447)
  wire Jqapw6;  // ../RTL/cortexm0ds_logic.v(1471)
  wire Jqbow6;  // ../RTL/cortexm0ds_logic.v(1003)
  wire Jqhiu6;  // ../RTL/cortexm0ds_logic.v(540)
  wire Jqiow6;  // ../RTL/cortexm0ds_logic.v(1097)
  wire Jqoiu6;  // ../RTL/cortexm0ds_logic.v(634)
  wire Jqphu6;  // ../RTL/cortexm0ds_logic.v(166)
  wire Jqpow6;  // ../RTL/cortexm0ds_logic.v(1190)
  wire Jqviu6;  // ../RTL/cortexm0ds_logic.v(728)
  wire Jqwhu6;  // ../RTL/cortexm0ds_logic.v(260)
  wire Jqwow6;  // ../RTL/cortexm0ds_logic.v(1284)
  wire Jr1ju6;  // ../RTL/cortexm0ds_logic.v(808)
  wire Jr2iu6;  // ../RTL/cortexm0ds_logic.v(340)
  wire Jr2pw6;  // ../RTL/cortexm0ds_logic.v(1365)
  wire Jr8ju6;  // ../RTL/cortexm0ds_logic.v(902)
  wire Jr9iu6;  // ../RTL/cortexm0ds_logic.v(434)
  wire Jr9pw6;  // ../RTL/cortexm0ds_logic.v(1458)
  wire Jraax6;  // ../RTL/cortexm0ds_logic.v(1633)
  wire Jraow6;  // ../RTL/cortexm0ds_logic.v(990)
  wire Jrgiu6;  // ../RTL/cortexm0ds_logic.v(527)
  wire Jrhow6;  // ../RTL/cortexm0ds_logic.v(1084)
  wire Jrniu6;  // ../RTL/cortexm0ds_logic.v(621)
  wire Jrohu6;  // ../RTL/cortexm0ds_logic.v(153)
  wire Jroow6;  // ../RTL/cortexm0ds_logic.v(1177)
  wire Jruiu6;  // ../RTL/cortexm0ds_logic.v(715)
  wire Jrvhu6;  // ../RTL/cortexm0ds_logic.v(247)
  wire Jrvow6;  // ../RTL/cortexm0ds_logic.v(1271)
  wire Jrvpw6;  // ../RTL/cortexm0ds_logic.v(1609)
  wire Jrypw6;  // ../RTL/cortexm0ds_logic.v(1615)
  wire Js0ju6;  // ../RTL/cortexm0ds_logic.v(795)
  wire Js1iu6;  // ../RTL/cortexm0ds_logic.v(327)
  wire Js1pw6;  // ../RTL/cortexm0ds_logic.v(1352)
  wire Js7ju6;  // ../RTL/cortexm0ds_logic.v(889)
  wire Js8iu6;  // ../RTL/cortexm0ds_logic.v(421)
  wire Js8pw6;  // ../RTL/cortexm0ds_logic.v(1445)
  wire Js9ow6;  // ../RTL/cortexm0ds_logic.v(977)
  wire Jsfiu6;  // ../RTL/cortexm0ds_logic.v(514)
  wire Jsgow6;  // ../RTL/cortexm0ds_logic.v(1071)
  wire Jsmiu6;  // ../RTL/cortexm0ds_logic.v(608)
  wire Jsnow6;  // ../RTL/cortexm0ds_logic.v(1164)
  wire Jstiu6;  // ../RTL/cortexm0ds_logic.v(702)
  wire Jsuhu6;  // ../RTL/cortexm0ds_logic.v(234)
  wire Jsuow6;  // ../RTL/cortexm0ds_logic.v(1258)
  wire Jt0iu6;  // ../RTL/cortexm0ds_logic.v(314)
  wire Jt0pw6;  // ../RTL/cortexm0ds_logic.v(1339)
  wire Jt6ju6;  // ../RTL/cortexm0ds_logic.v(876)
  wire Jt7iu6;  // ../RTL/cortexm0ds_logic.v(408)
  wire Jt7pw6;  // ../RTL/cortexm0ds_logic.v(1432)
  wire Jt8ow6;  // ../RTL/cortexm0ds_logic.v(964)
  wire Jteiu6;  // ../RTL/cortexm0ds_logic.v(501)
  wire Jtfow6;  // ../RTL/cortexm0ds_logic.v(1058)
  wire Jtliu6;  // ../RTL/cortexm0ds_logic.v(595)
  wire Jtmow6;  // ../RTL/cortexm0ds_logic.v(1151)
  wire Jtsiu6;  // ../RTL/cortexm0ds_logic.v(689)
  wire Jtthu6;  // ../RTL/cortexm0ds_logic.v(221)
  wire Jttow6;  // ../RTL/cortexm0ds_logic.v(1245)
  wire Jtvpw6;  // ../RTL/cortexm0ds_logic.v(1609)
  wire Jtziu6;  // ../RTL/cortexm0ds_logic.v(782)
  wire Ju5ju6;  // ../RTL/cortexm0ds_logic.v(863)
  wire Ju6iu6;  // ../RTL/cortexm0ds_logic.v(395)
  wire Ju6pw6;  // ../RTL/cortexm0ds_logic.v(1419)
  wire Ju7ow6;  // ../RTL/cortexm0ds_logic.v(951)
  wire Judiu6;  // ../RTL/cortexm0ds_logic.v(488)
  wire Judpw6;  // ../RTL/cortexm0ds_logic.v(1513)
  wire Jueow6;  // ../RTL/cortexm0ds_logic.v(1045)
  wire Jukiu6;  // ../RTL/cortexm0ds_logic.v(582)
  wire Julow6;  // ../RTL/cortexm0ds_logic.v(1138)
  wire Juriu6;  // ../RTL/cortexm0ds_logic.v(676)
  wire Jusax6;  // ../RTL/cortexm0ds_logic.v(1666)
  wire Jushu6;  // ../RTL/cortexm0ds_logic.v(208)
  wire Jusow6;  // ../RTL/cortexm0ds_logic.v(1232)
  wire Juyiu6;  // ../RTL/cortexm0ds_logic.v(769)
  wire Juzhu6;  // ../RTL/cortexm0ds_logic.v(301)
  wire Juzow6;  // ../RTL/cortexm0ds_logic.v(1326)
  wire Jv4ju6;  // ../RTL/cortexm0ds_logic.v(850)
  wire Jv5iu6;  // ../RTL/cortexm0ds_logic.v(382)
  wire Jv5pw6;  // ../RTL/cortexm0ds_logic.v(1406)
  wire Jv6ow6;  // ../RTL/cortexm0ds_logic.v(938)
  wire Jvciu6;  // ../RTL/cortexm0ds_logic.v(475)
  wire Jvcpw6;  // ../RTL/cortexm0ds_logic.v(1500)
  wire Jvdow6;  // ../RTL/cortexm0ds_logic.v(1032)
  wire Jvjiu6;  // ../RTL/cortexm0ds_logic.v(569)
  wire Jvkow6;  // ../RTL/cortexm0ds_logic.v(1125)
  wire Jvkpw6;  // ../RTL/cortexm0ds_logic.v(1589)
  wire Jvppw6;  // ../RTL/cortexm0ds_logic.v(1599)
  wire Jvqiu6;  // ../RTL/cortexm0ds_logic.v(663)
  wire Jvrhu6;  // ../RTL/cortexm0ds_logic.v(195)
  wire Jvrow6;  // ../RTL/cortexm0ds_logic.v(1219)
  wire Jvvpw6;  // ../RTL/cortexm0ds_logic.v(1609)
  wire Jvxiu6;  // ../RTL/cortexm0ds_logic.v(756)
  wire Jvyhu6;  // ../RTL/cortexm0ds_logic.v(288)
  wire Jvyow6;  // ../RTL/cortexm0ds_logic.v(1313)
  wire Jw3ju6;  // ../RTL/cortexm0ds_logic.v(837)
  wire Jw4iu6;  // ../RTL/cortexm0ds_logic.v(369)
  wire Jw4pw6;  // ../RTL/cortexm0ds_logic.v(1393)
  wire Jwbiu6;  // ../RTL/cortexm0ds_logic.v(462)
  wire Jwbpw6;  // ../RTL/cortexm0ds_logic.v(1487)
  wire Jwcow6;  // ../RTL/cortexm0ds_logic.v(1019)
  wire Jwiiu6;  // ../RTL/cortexm0ds_logic.v(556)
  wire Jwjow6;  // ../RTL/cortexm0ds_logic.v(1112)
  wire Jwpiu6;  // ../RTL/cortexm0ds_logic.v(650)
  wire Jwqhu6;  // ../RTL/cortexm0ds_logic.v(182)
  wire Jwqow6;  // ../RTL/cortexm0ds_logic.v(1206)
  wire Jwwiu6;  // ../RTL/cortexm0ds_logic.v(743)
  wire Jwxhu6;  // ../RTL/cortexm0ds_logic.v(275)
  wire Jwxow6;  // ../RTL/cortexm0ds_logic.v(1300)
  wire Jx1bx6;  // ../RTL/cortexm0ds_logic.v(1683)
  wire Jx2ju6;  // ../RTL/cortexm0ds_logic.v(824)
  wire Jx3iu6;  // ../RTL/cortexm0ds_logic.v(356)
  wire Jx3pw6;  // ../RTL/cortexm0ds_logic.v(1380)
  wire Jx9ju6;  // ../RTL/cortexm0ds_logic.v(917)
  wire Jxaiu6;  // ../RTL/cortexm0ds_logic.v(449)
  wire Jxapw6;  // ../RTL/cortexm0ds_logic.v(1474)
  wire Jxbow6;  // ../RTL/cortexm0ds_logic.v(1006)
  wire Jxgax6;  // ../RTL/cortexm0ds_logic.v(1645)
  wire Jxhiu6;  // ../RTL/cortexm0ds_logic.v(543)
  wire Jxiow6;  // ../RTL/cortexm0ds_logic.v(1099)
  wire Jxoiu6;  // ../RTL/cortexm0ds_logic.v(637)
  wire Jxphu6;  // ../RTL/cortexm0ds_logic.v(169)
  wire Jxpow6;  // ../RTL/cortexm0ds_logic.v(1193)
  wire Jxviu6;  // ../RTL/cortexm0ds_logic.v(730)
  wire Jxwhu6;  // ../RTL/cortexm0ds_logic.v(262)
  wire Jxwow6;  // ../RTL/cortexm0ds_logic.v(1287)
  wire Jy1ju6;  // ../RTL/cortexm0ds_logic.v(811)
  wire Jy2iu6;  // ../RTL/cortexm0ds_logic.v(343)
  wire Jy2pw6;  // ../RTL/cortexm0ds_logic.v(1367)
  wire Jy5bx6;  // ../RTL/cortexm0ds_logic.v(1690)
  wire Jy8ju6;  // ../RTL/cortexm0ds_logic.v(904)
  wire Jy9iu6;  // ../RTL/cortexm0ds_logic.v(436)
  wire Jy9pw6;  // ../RTL/cortexm0ds_logic.v(1461)
  wire Jyaow6;  // ../RTL/cortexm0ds_logic.v(993)
  wire Jydhu6;  // ../RTL/cortexm0ds_logic.v(121)
  wire Jygiu6;  // ../RTL/cortexm0ds_logic.v(530)
  wire Jyhow6;  // ../RTL/cortexm0ds_logic.v(1086)
  wire Jyniu6;  // ../RTL/cortexm0ds_logic.v(624)
  wire Jyohu6;  // ../RTL/cortexm0ds_logic.v(156)
  wire Jyoow6;  // ../RTL/cortexm0ds_logic.v(1180)
  wire Jyuiu6;  // ../RTL/cortexm0ds_logic.v(717)
  wire Jyvhu6;  // ../RTL/cortexm0ds_logic.v(249)
  wire Jyvow6;  // ../RTL/cortexm0ds_logic.v(1274)
  wire Jz0ju6;  // ../RTL/cortexm0ds_logic.v(798)
  wire Jz1iu6;  // ../RTL/cortexm0ds_logic.v(330)
  wire Jz1pw6;  // ../RTL/cortexm0ds_logic.v(1354)
  wire Jz2bx6;  // ../RTL/cortexm0ds_logic.v(1684)
  wire Jz7ju6;  // ../RTL/cortexm0ds_logic.v(891)
  wire Jz8iu6;  // ../RTL/cortexm0ds_logic.v(423)
  wire Jz8pw6;  // ../RTL/cortexm0ds_logic.v(1448)
  wire Jz9ow6;  // ../RTL/cortexm0ds_logic.v(980)
  wire Jzfiu6;  // ../RTL/cortexm0ds_logic.v(517)
  wire Jzgow6;  // ../RTL/cortexm0ds_logic.v(1073)
  wire Jzmhu6;  // ../RTL/cortexm0ds_logic.v(143)
  wire Jzmiu6;  // ../RTL/cortexm0ds_logic.v(611)
  wire Jznow6;  // ../RTL/cortexm0ds_logic.v(1167)
  wire Jztiu6;  // ../RTL/cortexm0ds_logic.v(704)
  wire Jzuhu6;  // ../RTL/cortexm0ds_logic.v(236)
  wire Jzuow6;  // ../RTL/cortexm0ds_logic.v(1261)
  wire K04ju6;  // ../RTL/cortexm0ds_logic.v(838)
  wire K05iu6;  // ../RTL/cortexm0ds_logic.v(370)
  wire K05pw6;  // ../RTL/cortexm0ds_logic.v(1395)
  wire K0ciu6;  // ../RTL/cortexm0ds_logic.v(464)
  wire K0cpw6;  // ../RTL/cortexm0ds_logic.v(1488)
  wire K0dow6;  // ../RTL/cortexm0ds_logic.v(1020)
  wire K0jiu6;  // ../RTL/cortexm0ds_logic.v(558)
  wire K0kow6;  // ../RTL/cortexm0ds_logic.v(1114)
  wire K0qiu6;  // ../RTL/cortexm0ds_logic.v(651)
  wire K0rhu6;  // ../RTL/cortexm0ds_logic.v(183)
  wire K0row6;  // ../RTL/cortexm0ds_logic.v(1208)
  wire K0xiu6;  // ../RTL/cortexm0ds_logic.v(745)
  wire K0yhu6;  // ../RTL/cortexm0ds_logic.v(277)
  wire K0yow6;  // ../RTL/cortexm0ds_logic.v(1301)
  wire K13ju6;  // ../RTL/cortexm0ds_logic.v(825)
  wire K14iu6;  // ../RTL/cortexm0ds_logic.v(357)
  wire K14pw6;  // ../RTL/cortexm0ds_logic.v(1382)
  wire K1aju6;  // ../RTL/cortexm0ds_logic.v(919)
  wire K1biu6;  // ../RTL/cortexm0ds_logic.v(451)
  wire K1bpw6;  // ../RTL/cortexm0ds_logic.v(1475)
  wire K1cow6;  // ../RTL/cortexm0ds_logic.v(1007)
  wire K1iiu6;  // ../RTL/cortexm0ds_logic.v(545)
  wire K1jow6;  // ../RTL/cortexm0ds_logic.v(1101)
  wire K1khu6;  // ../RTL/cortexm0ds_logic.v(135)
  wire K1piu6;  // ../RTL/cortexm0ds_logic.v(638)
  wire K1qhu6;  // ../RTL/cortexm0ds_logic.v(170)
  wire K1qow6;  // ../RTL/cortexm0ds_logic.v(1195)
  wire K1wiu6;  // ../RTL/cortexm0ds_logic.v(732)
  wire K1xax6;  // ../RTL/cortexm0ds_logic.v(1674)
  wire K1xhu6;  // ../RTL/cortexm0ds_logic.v(264)
  wire K1xow6;  // ../RTL/cortexm0ds_logic.v(1288)
  wire K22ju6;  // ../RTL/cortexm0ds_logic.v(812)
  wire K23iu6;  // ../RTL/cortexm0ds_logic.v(344)
  wire K23pw6;  // ../RTL/cortexm0ds_logic.v(1369)
  wire K29ju6;  // ../RTL/cortexm0ds_logic.v(906)
  wire K2aiu6;  // ../RTL/cortexm0ds_logic.v(438)
  wire K2apw6;  // ../RTL/cortexm0ds_logic.v(1462)
  wire K2bow6;  // ../RTL/cortexm0ds_logic.v(994)
  wire K2hiu6;  // ../RTL/cortexm0ds_logic.v(532)
  wire K2iow6;  // ../RTL/cortexm0ds_logic.v(1088)
  wire K2oiu6;  // ../RTL/cortexm0ds_logic.v(625)
  wire K2phu6;  // ../RTL/cortexm0ds_logic.v(157)
  wire K2pow6;  // ../RTL/cortexm0ds_logic.v(1182)
  wire K2viu6;  // ../RTL/cortexm0ds_logic.v(719)
  wire K2whu6;  // ../RTL/cortexm0ds_logic.v(251)
  wire K2wow6;  // ../RTL/cortexm0ds_logic.v(1275)
  wire K31ju6;  // ../RTL/cortexm0ds_logic.v(799)
  wire K32iu6;  // ../RTL/cortexm0ds_logic.v(331)
  wire K32pw6;  // ../RTL/cortexm0ds_logic.v(1356)
  wire K38ju6;  // ../RTL/cortexm0ds_logic.v(893)
  wire K39iu6;  // ../RTL/cortexm0ds_logic.v(425)
  wire K39pw6;  // ../RTL/cortexm0ds_logic.v(1449)
  wire K3aow6;  // ../RTL/cortexm0ds_logic.v(981)
  wire K3giu6;  // ../RTL/cortexm0ds_logic.v(519)
  wire K3how6;  // ../RTL/cortexm0ds_logic.v(1075)
  wire K3jhu6;  // ../RTL/cortexm0ds_logic.v(133)
  wire K3niu6;  // ../RTL/cortexm0ds_logic.v(612)
  wire K3oow6;  // ../RTL/cortexm0ds_logic.v(1169)
  wire K3uiu6;  // ../RTL/cortexm0ds_logic.v(706)
  wire K3vhu6;  // ../RTL/cortexm0ds_logic.v(238)
  wire K3vow6;  // ../RTL/cortexm0ds_logic.v(1262)
  wire K40ju6;  // ../RTL/cortexm0ds_logic.v(786)
  wire K41iu6;  // ../RTL/cortexm0ds_logic.v(318)
  wire K41pw6;  // ../RTL/cortexm0ds_logic.v(1343)
  wire K47ju6;  // ../RTL/cortexm0ds_logic.v(880)
  wire K48iu6;  // ../RTL/cortexm0ds_logic.v(412)
  wire K48pw6;  // ../RTL/cortexm0ds_logic.v(1436)
  wire K49ow6;  // ../RTL/cortexm0ds_logic.v(968)
  wire K4fiu6;  // ../RTL/cortexm0ds_logic.v(506)
  wire K4gow6;  // ../RTL/cortexm0ds_logic.v(1062)
  wire K4miu6;  // ../RTL/cortexm0ds_logic.v(599)
  wire K4now6;  // ../RTL/cortexm0ds_logic.v(1156)
  wire K4tiu6;  // ../RTL/cortexm0ds_logic.v(693)
  wire K4uhu6;  // ../RTL/cortexm0ds_logic.v(225)
  wire K4uow6;  // ../RTL/cortexm0ds_logic.v(1249)
  wire K50iu6;  // ../RTL/cortexm0ds_logic.v(305)
  wire K50pw6;  // ../RTL/cortexm0ds_logic.v(1330)
  wire K56ju6;  // ../RTL/cortexm0ds_logic.v(867)
  wire K57iu6;  // ../RTL/cortexm0ds_logic.v(399)
  wire K57pw6;  // ../RTL/cortexm0ds_logic.v(1423)
  wire K58ow6;  // ../RTL/cortexm0ds_logic.v(955)
  wire K5eiu6;  // ../RTL/cortexm0ds_logic.v(493)
  wire K5fow6;  // ../RTL/cortexm0ds_logic.v(1049)
  wire K5hbx6;  // ../RTL/cortexm0ds_logic.v(1710)
  wire K5ihu6;  // ../RTL/cortexm0ds_logic.v(130)
  wire K5liu6;  // ../RTL/cortexm0ds_logic.v(586)
  wire K5mow6;  // ../RTL/cortexm0ds_logic.v(1143)
  wire K5siu6;  // ../RTL/cortexm0ds_logic.v(680)
  wire K5thu6;  // ../RTL/cortexm0ds_logic.v(212)
  wire K5tow6;  // ../RTL/cortexm0ds_logic.v(1236)
  wire K5ziu6;  // ../RTL/cortexm0ds_logic.v(773)
  wire K65bx6;  // ../RTL/cortexm0ds_logic.v(1688)
  wire K65ju6;  // ../RTL/cortexm0ds_logic.v(854)
  wire K66iu6;  // ../RTL/cortexm0ds_logic.v(386)
  wire K66pw6;  // ../RTL/cortexm0ds_logic.v(1410)
  wire K67ow6;  // ../RTL/cortexm0ds_logic.v(942)
  wire K6diu6;  // ../RTL/cortexm0ds_logic.v(480)
  wire K6dpw6;  // ../RTL/cortexm0ds_logic.v(1504)
  wire K6eow6;  // ../RTL/cortexm0ds_logic.v(1036)
  wire K6fhu6;  // ../RTL/cortexm0ds_logic.v(123)
  wire K6gax6;  // ../RTL/cortexm0ds_logic.v(1643)
  wire K6kiu6;  // ../RTL/cortexm0ds_logic.v(573)
  wire K6low6;  // ../RTL/cortexm0ds_logic.v(1130)
  wire K6riu6;  // ../RTL/cortexm0ds_logic.v(667)
  wire K6shu6;  // ../RTL/cortexm0ds_logic.v(199)
  wire K6sow6;  // ../RTL/cortexm0ds_logic.v(1223)
  wire K6yiu6;  // ../RTL/cortexm0ds_logic.v(760)
  wire K6zhu6;  // ../RTL/cortexm0ds_logic.v(292)
  wire K6zow6;  // ../RTL/cortexm0ds_logic.v(1317)
  wire K74ju6;  // ../RTL/cortexm0ds_logic.v(841)
  wire K75iu6;  // ../RTL/cortexm0ds_logic.v(373)
  wire K75pw6;  // ../RTL/cortexm0ds_logic.v(1397)
  wire K76ow6;  // ../RTL/cortexm0ds_logic.v(929)
  wire K7ciu6;  // ../RTL/cortexm0ds_logic.v(467)
  wire K7cpw6;  // ../RTL/cortexm0ds_logic.v(1491)
  wire K7dow6;  // ../RTL/cortexm0ds_logic.v(1023)
  wire K7jiu6;  // ../RTL/cortexm0ds_logic.v(560)
  wire K7kow6;  // ../RTL/cortexm0ds_logic.v(1117)
  wire K7qiu6;  // ../RTL/cortexm0ds_logic.v(654)
  wire K7rhu6;  // ../RTL/cortexm0ds_logic.v(186)
  wire K7row6;  // ../RTL/cortexm0ds_logic.v(1210)
  wire K7vpw6;  // ../RTL/cortexm0ds_logic.v(1608)
  wire K7xiu6;  // ../RTL/cortexm0ds_logic.v(747)
  wire K7yhu6;  // ../RTL/cortexm0ds_logic.v(279)
  wire K7yow6;  // ../RTL/cortexm0ds_logic.v(1304)
  wire K83ju6;  // ../RTL/cortexm0ds_logic.v(828)
  wire K84iu6;  // ../RTL/cortexm0ds_logic.v(360)
  wire K84pw6;  // ../RTL/cortexm0ds_logic.v(1384)
  wire K8aju6;  // ../RTL/cortexm0ds_logic.v(922)
  wire K8biu6;  // ../RTL/cortexm0ds_logic.v(454)
  wire K8bpw6;  // ../RTL/cortexm0ds_logic.v(1478)
  wire K8cow6;  // ../RTL/cortexm0ds_logic.v(1010)
  wire K8iiu6;  // ../RTL/cortexm0ds_logic.v(547)
  wire K8jow6;  // ../RTL/cortexm0ds_logic.v(1104)
  wire K8piu6;  // ../RTL/cortexm0ds_logic.v(641)
  wire K8qhu6;  // ../RTL/cortexm0ds_logic.v(173)
  wire K8qow6;  // ../RTL/cortexm0ds_logic.v(1197)
  wire K8wiu6;  // ../RTL/cortexm0ds_logic.v(734)
  wire K8xhu6;  // ../RTL/cortexm0ds_logic.v(266)
  wire K8xow6;  // ../RTL/cortexm0ds_logic.v(1291)
  wire K92ju6;  // ../RTL/cortexm0ds_logic.v(815)
  wire K93iu6;  // ../RTL/cortexm0ds_logic.v(347)
  wire K93pw6;  // ../RTL/cortexm0ds_logic.v(1371)
  wire K94bx6;  // ../RTL/cortexm0ds_logic.v(1687)
  wire K99ju6;  // ../RTL/cortexm0ds_logic.v(909)
  wire K9aiu6;  // ../RTL/cortexm0ds_logic.v(441)
  wire K9apw6;  // ../RTL/cortexm0ds_logic.v(1465)
  wire K9bow6;  // ../RTL/cortexm0ds_logic.v(997)
  wire K9hiu6;  // ../RTL/cortexm0ds_logic.v(534)
  wire K9iow6;  // ../RTL/cortexm0ds_logic.v(1091)
  wire K9oiu6;  // ../RTL/cortexm0ds_logic.v(628)
  wire K9phu6;  // ../RTL/cortexm0ds_logic.v(160)
  wire K9pow6;  // ../RTL/cortexm0ds_logic.v(1184)
  wire K9viu6;  // ../RTL/cortexm0ds_logic.v(721)
  wire K9whu6;  // ../RTL/cortexm0ds_logic.v(253)
  wire K9wow6;  // ../RTL/cortexm0ds_logic.v(1278)
  wire Ka1ju6;  // ../RTL/cortexm0ds_logic.v(802)
  wire Ka2iu6;  // ../RTL/cortexm0ds_logic.v(334)
  wire Ka2pw6;  // ../RTL/cortexm0ds_logic.v(1358)
  wire Ka8ju6;  // ../RTL/cortexm0ds_logic.v(896)
  wire Ka9iu6;  // ../RTL/cortexm0ds_logic.v(428)
  wire Ka9pw6;  // ../RTL/cortexm0ds_logic.v(1452)
  wire Kaaow6;  // ../RTL/cortexm0ds_logic.v(984)
  wire Kadbx6;  // ../RTL/cortexm0ds_logic.v(1703)
  wire Kagiu6;  // ../RTL/cortexm0ds_logic.v(521)
  wire Kahow6;  // ../RTL/cortexm0ds_logic.v(1078)
  wire Kakax6;  // ../RTL/cortexm0ds_logic.v(1651)
  wire Kalpw6;  // ../RTL/cortexm0ds_logic.v(1590)
  wire Kaniu6;  // ../RTL/cortexm0ds_logic.v(615)
  wire Kaohu6;  // ../RTL/cortexm0ds_logic.v(147)
  wire Kaoow6;  // ../RTL/cortexm0ds_logic.v(1171)
  wire Kauiu6;  // ../RTL/cortexm0ds_logic.v(708)
  wire Kavhu6;  // ../RTL/cortexm0ds_logic.v(240)
  wire Kavow6;  // ../RTL/cortexm0ds_logic.v(1265)
  wire Kb0ju6;  // ../RTL/cortexm0ds_logic.v(789)
  wire Kb1iu6;  // ../RTL/cortexm0ds_logic.v(321)
  wire Kb1pw6;  // ../RTL/cortexm0ds_logic.v(1345)
  wire Kb7ju6;  // ../RTL/cortexm0ds_logic.v(883)
  wire Kb8iu6;  // ../RTL/cortexm0ds_logic.v(415)
  wire Kb8pw6;  // ../RTL/cortexm0ds_logic.v(1439)
  wire Kb9ow6;  // ../RTL/cortexm0ds_logic.v(971)
  wire Kbfiu6;  // ../RTL/cortexm0ds_logic.v(508)
  wire Kbgow6;  // ../RTL/cortexm0ds_logic.v(1065)
  wire Kbmiu6;  // ../RTL/cortexm0ds_logic.v(602)
  wire Kbnow6;  // ../RTL/cortexm0ds_logic.v(1158)
  wire Kbtiu6;  // ../RTL/cortexm0ds_logic.v(695)
  wire Kbuhu6;  // ../RTL/cortexm0ds_logic.v(227)
  wire Kbuow6;  // ../RTL/cortexm0ds_logic.v(1252)
  wire Kc0iu6;  // ../RTL/cortexm0ds_logic.v(308)
  wire Kc0pw6;  // ../RTL/cortexm0ds_logic.v(1332)
  wire Kc6ju6;  // ../RTL/cortexm0ds_logic.v(870)
  wire Kc7iu6;  // ../RTL/cortexm0ds_logic.v(402)
  wire Kc7pw6;  // ../RTL/cortexm0ds_logic.v(1426)
  wire Kc8ow6;  // ../RTL/cortexm0ds_logic.v(958)
  wire Kcaax6;  // ../RTL/cortexm0ds_logic.v(1632)
  wire Kceiu6;  // ../RTL/cortexm0ds_logic.v(495)
  wire Kcfow6;  // ../RTL/cortexm0ds_logic.v(1052)
  wire Kcliu6;  // ../RTL/cortexm0ds_logic.v(589)
  wire Kcmow6;  // ../RTL/cortexm0ds_logic.v(1145)
  wire Kcsiu6;  // ../RTL/cortexm0ds_logic.v(682)
  wire Kcthu6;  // ../RTL/cortexm0ds_logic.v(214)
  wire Kctow6;  // ../RTL/cortexm0ds_logic.v(1239)
  wire Kcziu6;  // ../RTL/cortexm0ds_logic.v(776)
  wire Kd5ju6;  // ../RTL/cortexm0ds_logic.v(857)
  wire Kd6iu6;  // ../RTL/cortexm0ds_logic.v(389)
  wire Kd6pw6;  // ../RTL/cortexm0ds_logic.v(1413)
  wire Kd7ow6;  // ../RTL/cortexm0ds_logic.v(945)
  wire Kddiu6;  // ../RTL/cortexm0ds_logic.v(482)
  wire Kddpw6;  // ../RTL/cortexm0ds_logic.v(1507)
  wire Kdeow6;  // ../RTL/cortexm0ds_logic.v(1039)
  wire Kdkiu6;  // ../RTL/cortexm0ds_logic.v(576)
  wire Kdlow6;  // ../RTL/cortexm0ds_logic.v(1132)
  wire Kdriu6;  // ../RTL/cortexm0ds_logic.v(669)
  wire Kdshu6;  // ../RTL/cortexm0ds_logic.v(201)
  wire Kdsow6;  // ../RTL/cortexm0ds_logic.v(1226)
  wire Kdyiu6;  // ../RTL/cortexm0ds_logic.v(763)
  wire Kdzhu6;  // ../RTL/cortexm0ds_logic.v(295)
  wire Kdzow6;  // ../RTL/cortexm0ds_logic.v(1319)
  wire Ke1qw6;  // ../RTL/cortexm0ds_logic.v(1619)
  wire Ke4ju6;  // ../RTL/cortexm0ds_logic.v(844)
  wire Ke5iu6;  // ../RTL/cortexm0ds_logic.v(376)
  wire Ke5pw6;  // ../RTL/cortexm0ds_logic.v(1400)
  wire Ke6ow6;  // ../RTL/cortexm0ds_logic.v(932)
  wire Keciu6;  // ../RTL/cortexm0ds_logic.v(469)
  wire Kecpw6;  // ../RTL/cortexm0ds_logic.v(1494)
  wire Kedow6;  // ../RTL/cortexm0ds_logic.v(1026)
  wire Kejiu6;  // ../RTL/cortexm0ds_logic.v(563)
  wire Kekow6;  // ../RTL/cortexm0ds_logic.v(1119)
  wire Keqiu6;  // ../RTL/cortexm0ds_logic.v(656)
  wire Kerhu6;  // ../RTL/cortexm0ds_logic.v(188)
  wire Kerow6;  // ../RTL/cortexm0ds_logic.v(1213)
  wire Kexiu6;  // ../RTL/cortexm0ds_logic.v(750)
  wire Keyhu6;  // ../RTL/cortexm0ds_logic.v(282)
  wire Keyow6;  // ../RTL/cortexm0ds_logic.v(1306)
  wire Kf3ju6;  // ../RTL/cortexm0ds_logic.v(831)
  wire Kf4iu6;  // ../RTL/cortexm0ds_logic.v(363)
  wire Kf4pw6;  // ../RTL/cortexm0ds_logic.v(1387)
  wire Kfaju6;  // ../RTL/cortexm0ds_logic.v(924)
  wire Kfbiu6;  // ../RTL/cortexm0ds_logic.v(456)
  wire Kfbpw6;  // ../RTL/cortexm0ds_logic.v(1481)
  wire Kfcow6;  // ../RTL/cortexm0ds_logic.v(1013)
  wire Kfiiu6;  // ../RTL/cortexm0ds_logic.v(550)
  wire Kfjow6;  // ../RTL/cortexm0ds_logic.v(1106)
  wire Kfoax6;  // ../RTL/cortexm0ds_logic.v(1658)
  wire Kfpiu6;  // ../RTL/cortexm0ds_logic.v(643)
  wire Kfqhu6;  // ../RTL/cortexm0ds_logic.v(175)
  wire Kfqow6;  // ../RTL/cortexm0ds_logic.v(1200)
  wire Kfwiu6;  // ../RTL/cortexm0ds_logic.v(737)
  wire Kfxhu6;  // ../RTL/cortexm0ds_logic.v(269)
  wire Kfxow6;  // ../RTL/cortexm0ds_logic.v(1293)
  wire Kg2ju6;  // ../RTL/cortexm0ds_logic.v(818)
  wire Kg3iu6;  // ../RTL/cortexm0ds_logic.v(350)
  wire Kg3pw6;  // ../RTL/cortexm0ds_logic.v(1374)
  wire Kg9ju6;  // ../RTL/cortexm0ds_logic.v(911)
  wire Kgaiu6;  // ../RTL/cortexm0ds_logic.v(443)
  wire Kgapw6;  // ../RTL/cortexm0ds_logic.v(1468)
  wire Kgbow6;  // ../RTL/cortexm0ds_logic.v(1000)
  wire Kghiu6;  // ../RTL/cortexm0ds_logic.v(537)
  wire Kgiow6;  // ../RTL/cortexm0ds_logic.v(1093)
  wire Kgoiu6;  // ../RTL/cortexm0ds_logic.v(630)
  wire Kgphu6;  // ../RTL/cortexm0ds_logic.v(162)
  wire Kgpow6;  // ../RTL/cortexm0ds_logic.v(1187)
  wire Kgviu6;  // ../RTL/cortexm0ds_logic.v(724)
  wire Kgwhu6;  // ../RTL/cortexm0ds_logic.v(256)
  wire Kgwow6;  // ../RTL/cortexm0ds_logic.v(1280)
  wire Kh1ju6;  // ../RTL/cortexm0ds_logic.v(805)
  wire Kh2iu6;  // ../RTL/cortexm0ds_logic.v(337)
  wire Kh2pw6;  // ../RTL/cortexm0ds_logic.v(1361)
  wire Kh8ju6;  // ../RTL/cortexm0ds_logic.v(898)
  wire Kh9iu6;  // ../RTL/cortexm0ds_logic.v(430)
  wire Kh9pw6;  // ../RTL/cortexm0ds_logic.v(1455)
  wire Khaow6;  // ../RTL/cortexm0ds_logic.v(987)
  wire Khgax6;  // ../RTL/cortexm0ds_logic.v(1644)
  wire Khgiu6;  // ../RTL/cortexm0ds_logic.v(524)
  wire Khhow6;  // ../RTL/cortexm0ds_logic.v(1080)
  wire Khniu6;  // ../RTL/cortexm0ds_logic.v(617)
  wire Khoax6;  // ../RTL/cortexm0ds_logic.v(1659)
  wire Khohu6;  // ../RTL/cortexm0ds_logic.v(149)
  wire Khoow6;  // ../RTL/cortexm0ds_logic.v(1174)
  wire Khuiu6;  // ../RTL/cortexm0ds_logic.v(711)
  wire Khvhu6;  // ../RTL/cortexm0ds_logic.v(243)
  wire Khvow6;  // ../RTL/cortexm0ds_logic.v(1267)
  wire Ki0ju6;  // ../RTL/cortexm0ds_logic.v(792)
  wire Ki1iu6;  // ../RTL/cortexm0ds_logic.v(324)
  wire Ki1pw6;  // ../RTL/cortexm0ds_logic.v(1348)
  wire Ki3bx6;  // ../RTL/cortexm0ds_logic.v(1685)
  wire Ki7ju6;  // ../RTL/cortexm0ds_logic.v(885)
  wire Ki8iu6;  // ../RTL/cortexm0ds_logic.v(417)
  wire Ki8pw6;  // ../RTL/cortexm0ds_logic.v(1442)
  wire Ki9ow6;  // ../RTL/cortexm0ds_logic.v(974)
  wire Kifiu6;  // ../RTL/cortexm0ds_logic.v(511)
  wire Kigow6;  // ../RTL/cortexm0ds_logic.v(1067)
  wire Kikhu6;  // ../RTL/cortexm0ds_logic.v(137)
  wire Kimiu6;  // ../RTL/cortexm0ds_logic.v(604)
  wire Kinow6;  // ../RTL/cortexm0ds_logic.v(1161)
  wire Kitiu6;  // ../RTL/cortexm0ds_logic.v(698)
  wire Kiuhu6;  // ../RTL/cortexm0ds_logic.v(230)
  wire Kiuow6;  // ../RTL/cortexm0ds_logic.v(1254)
  wire Kj0iu6;  // ../RTL/cortexm0ds_logic.v(311)
  wire Kj0pw6;  // ../RTL/cortexm0ds_logic.v(1335)
  wire Kj6ju6;  // ../RTL/cortexm0ds_logic.v(872)
  wire Kj7iu6;  // ../RTL/cortexm0ds_logic.v(404)
  wire Kj7pw6;  // ../RTL/cortexm0ds_logic.v(1429)
  wire Kj8ow6;  // ../RTL/cortexm0ds_logic.v(961)
  wire Kjeiu6;  // ../RTL/cortexm0ds_logic.v(498)
  wire Kjfow6;  // ../RTL/cortexm0ds_logic.v(1054)
  wire Kjliu6;  // ../RTL/cortexm0ds_logic.v(591)
  wire Kjmow6;  // ../RTL/cortexm0ds_logic.v(1148)
  wire Kjoax6;  // ../RTL/cortexm0ds_logic.v(1659)
  wire Kjsiu6;  // ../RTL/cortexm0ds_logic.v(685)
  wire Kjthu6;  // ../RTL/cortexm0ds_logic.v(217)
  wire Kjtow6;  // ../RTL/cortexm0ds_logic.v(1241)
  wire Kjziu6;  // ../RTL/cortexm0ds_logic.v(779)
  wire Kk5ju6;  // ../RTL/cortexm0ds_logic.v(859)
  wire Kk6iu6;  // ../RTL/cortexm0ds_logic.v(391)
  wire Kk6pw6;  // ../RTL/cortexm0ds_logic.v(1416)
  wire Kk7ow6;  // ../RTL/cortexm0ds_logic.v(948)
  wire Kkdiu6;  // ../RTL/cortexm0ds_logic.v(485)
  wire Kkdpw6;  // ../RTL/cortexm0ds_logic.v(1509)
  wire Kkeow6;  // ../RTL/cortexm0ds_logic.v(1041)
  wire Kkjhu6;  // ../RTL/cortexm0ds_logic.v(134)
  wire Kkjpw6;  // ../RTL/cortexm0ds_logic.v(1587)
  wire Kkkiu6;  // ../RTL/cortexm0ds_logic.v(578)
  wire Kklow6;  // ../RTL/cortexm0ds_logic.v(1135)
  wire Kkriu6;  // ../RTL/cortexm0ds_logic.v(672)
  wire Kkshu6;  // ../RTL/cortexm0ds_logic.v(204)
  wire Kksow6;  // ../RTL/cortexm0ds_logic.v(1228)
  wire Kkyiu6;  // ../RTL/cortexm0ds_logic.v(766)
  wire Kkzhu6;  // ../RTL/cortexm0ds_logic.v(298)
  wire Kkzow6;  // ../RTL/cortexm0ds_logic.v(1322)
  wire Kl0bx6;  // ../RTL/cortexm0ds_logic.v(1680)
  wire Kl4ju6;  // ../RTL/cortexm0ds_logic.v(846)
  wire Kl5iu6;  // ../RTL/cortexm0ds_logic.v(378)
  wire Kl5pw6;  // ../RTL/cortexm0ds_logic.v(1403)
  wire Kl6ow6;  // ../RTL/cortexm0ds_logic.v(935)
  wire Kl8ax6;  // ../RTL/cortexm0ds_logic.v(1628)
  wire Klciu6;  // ../RTL/cortexm0ds_logic.v(472)
  wire Klcpw6;  // ../RTL/cortexm0ds_logic.v(1496)
  wire Kldow6;  // ../RTL/cortexm0ds_logic.v(1028)
  wire Kljiu6;  // ../RTL/cortexm0ds_logic.v(565)
  wire Klkow6;  // ../RTL/cortexm0ds_logic.v(1122)
  wire Kloax6;  // ../RTL/cortexm0ds_logic.v(1659)
  wire Klqiu6;  // ../RTL/cortexm0ds_logic.v(659)
  wire Klrhu6;  // ../RTL/cortexm0ds_logic.v(191)
  wire Klrow6;  // ../RTL/cortexm0ds_logic.v(1215)
  wire Klxiu6;  // ../RTL/cortexm0ds_logic.v(753)
  wire Klyhu6;  // ../RTL/cortexm0ds_logic.v(285)
  wire Klyow6;  // ../RTL/cortexm0ds_logic.v(1309)
  wire Km3ju6;  // ../RTL/cortexm0ds_logic.v(833)
  wire Km4iu6;  // ../RTL/cortexm0ds_logic.v(365)
  wire Km4pw6;  // ../RTL/cortexm0ds_logic.v(1390)
  wire Kmaju6;  // ../RTL/cortexm0ds_logic.v(927)
  wire Kmbiu6;  // ../RTL/cortexm0ds_logic.v(459)
  wire Kmbpw6;  // ../RTL/cortexm0ds_logic.v(1483)
  wire Kmcow6;  // ../RTL/cortexm0ds_logic.v(1015)
  wire Kmehu6;  // ../RTL/cortexm0ds_logic.v(122)
  wire Kmihu6;  // ../RTL/cortexm0ds_logic.v(131)
  wire Kmiiu6;  // ../RTL/cortexm0ds_logic.v(552)
  wire Kmjow6;  // ../RTL/cortexm0ds_logic.v(1109)
  wire Kmjpw6;  // ../RTL/cortexm0ds_logic.v(1587)
  wire Kmpiu6;  // ../RTL/cortexm0ds_logic.v(646)
  wire Kmqhu6;  // ../RTL/cortexm0ds_logic.v(178)
  wire Kmqow6;  // ../RTL/cortexm0ds_logic.v(1202)
  wire Kmsax6;  // ../RTL/cortexm0ds_logic.v(1666)
  wire Kmwiu6;  // ../RTL/cortexm0ds_logic.v(740)
  wire Kmxhu6;  // ../RTL/cortexm0ds_logic.v(272)
  wire Kmxow6;  // ../RTL/cortexm0ds_logic.v(1296)
  wire Kn1qw6;  // ../RTL/cortexm0ds_logic.v(1620)
  wire Kn2ju6;  // ../RTL/cortexm0ds_logic.v(820)
  wire Kn2qw6;  // ../RTL/cortexm0ds_logic.v(1622)
  wire Kn3iu6;  // ../RTL/cortexm0ds_logic.v(352)
  wire Kn3pw6;  // ../RTL/cortexm0ds_logic.v(1377)
  wire Kn9ju6;  // ../RTL/cortexm0ds_logic.v(914)
  wire Knaiu6;  // ../RTL/cortexm0ds_logic.v(446)
  wire Knapw6;  // ../RTL/cortexm0ds_logic.v(1470)
  wire Knbbx6;  // ../RTL/cortexm0ds_logic.v(1700)
  wire Knbow6;  // ../RTL/cortexm0ds_logic.v(1002)
  wire Knhax6;  // ../RTL/cortexm0ds_logic.v(1646)
  wire Knhiu6;  // ../RTL/cortexm0ds_logic.v(539)
  wire Kniow6;  // ../RTL/cortexm0ds_logic.v(1096)
  wire Knmhu6;  // ../RTL/cortexm0ds_logic.v(143)
  wire Knoiu6;  // ../RTL/cortexm0ds_logic.v(633)
  wire Knphu6;  // ../RTL/cortexm0ds_logic.v(165)
  wire Knpow6;  // ../RTL/cortexm0ds_logic.v(1189)
  wire Knviu6;  // ../RTL/cortexm0ds_logic.v(727)
  wire Knwhu6;  // ../RTL/cortexm0ds_logic.v(259)
  wire Knwow6;  // ../RTL/cortexm0ds_logic.v(1283)
  wire Ko1ju6;  // ../RTL/cortexm0ds_logic.v(807)
  wire Ko2iu6;  // ../RTL/cortexm0ds_logic.v(339)
  wire Ko2pw6;  // ../RTL/cortexm0ds_logic.v(1364)
  wire Ko8ju6;  // ../RTL/cortexm0ds_logic.v(901)
  wire Ko9iu6;  // ../RTL/cortexm0ds_logic.v(433)
  wire Ko9pw6;  // ../RTL/cortexm0ds_logic.v(1457)
  wire Koabx6;  // ../RTL/cortexm0ds_logic.v(1698)
  wire Koaow6;  // ../RTL/cortexm0ds_logic.v(989)
  wire Kogiu6;  // ../RTL/cortexm0ds_logic.v(526)
  wire Kohhu6;  // ../RTL/cortexm0ds_logic.v(129)
  wire Kohow6;  // ../RTL/cortexm0ds_logic.v(1083)
  wire Kojpw6;  // ../RTL/cortexm0ds_logic.v(1587)
  wire Koniu6;  // ../RTL/cortexm0ds_logic.v(620)
  wire Koohu6;  // ../RTL/cortexm0ds_logic.v(152)
  wire Kooow6;  // ../RTL/cortexm0ds_logic.v(1176)
  wire Kosax6;  // ../RTL/cortexm0ds_logic.v(1666)
  wire Kouiu6;  // ../RTL/cortexm0ds_logic.v(714)
  wire Kovhu6;  // ../RTL/cortexm0ds_logic.v(246)
  wire Kovow6;  // ../RTL/cortexm0ds_logic.v(1270)
  wire Kp0ju6;  // ../RTL/cortexm0ds_logic.v(794)
  wire Kp1iu6;  // ../RTL/cortexm0ds_logic.v(326)
  wire Kp1pw6;  // ../RTL/cortexm0ds_logic.v(1351)
  wire Kp7ju6;  // ../RTL/cortexm0ds_logic.v(888)
  wire Kp8iu6;  // ../RTL/cortexm0ds_logic.v(420)
  wire Kp8pw6;  // ../RTL/cortexm0ds_logic.v(1444)
  wire Kp9ow6;  // ../RTL/cortexm0ds_logic.v(976)
  wire Kpfbx6;  // ../RTL/cortexm0ds_logic.v(1708)
  wire Kpfiu6;  // ../RTL/cortexm0ds_logic.v(513)
  wire Kpgow6;  // ../RTL/cortexm0ds_logic.v(1070)
  wire Kpmiu6;  // ../RTL/cortexm0ds_logic.v(607)
  wire Kpnow6;  // ../RTL/cortexm0ds_logic.v(1163)
  wire Kptiu6;  // ../RTL/cortexm0ds_logic.v(701)
  wire Kpuhu6;  // ../RTL/cortexm0ds_logic.v(233)
  wire Kpuow6;  // ../RTL/cortexm0ds_logic.v(1257)
  wire Kq0iu6;  // ../RTL/cortexm0ds_logic.v(313)
  wire Kq0pw6;  // ../RTL/cortexm0ds_logic.v(1338)
  wire Kq6ju6;  // ../RTL/cortexm0ds_logic.v(875)
  wire Kq7iu6;  // ../RTL/cortexm0ds_logic.v(407)
  wire Kq7pw6;  // ../RTL/cortexm0ds_logic.v(1431)
  wire Kq8ow6;  // ../RTL/cortexm0ds_logic.v(963)
  wire Kqdax6;  // ../RTL/cortexm0ds_logic.v(1638)
  wire Kqeiu6;  // ../RTL/cortexm0ds_logic.v(500)
  wire Kqfow6;  // ../RTL/cortexm0ds_logic.v(1057)
  wire Kqhbx6;  // ../RTL/cortexm0ds_logic.v(1711)
  wire Kqlhu6;  // ../RTL/cortexm0ds_logic.v(140)
  wire Kqliu6;  // ../RTL/cortexm0ds_logic.v(594)
  wire Kqmow6;  // ../RTL/cortexm0ds_logic.v(1150)
  wire Kqsax6;  // ../RTL/cortexm0ds_logic.v(1666)
  wire Kqsiu6;  // ../RTL/cortexm0ds_logic.v(688)
  wire Kqthu6;  // ../RTL/cortexm0ds_logic.v(220)
  wire Kqtow6;  // ../RTL/cortexm0ds_logic.v(1244)
  wire Kqziu6;  // ../RTL/cortexm0ds_logic.v(781)
  wire Kr5ju6;  // ../RTL/cortexm0ds_logic.v(862)
  wire Kr6iu6;  // ../RTL/cortexm0ds_logic.v(394)
  wire Kr6pw6;  // ../RTL/cortexm0ds_logic.v(1418)
  wire Kr7ow6;  // ../RTL/cortexm0ds_logic.v(950)
  wire Krbax6;  // ../RTL/cortexm0ds_logic.v(1635)
  wire Krdiu6;  // ../RTL/cortexm0ds_logic.v(487)
  wire Krdpw6;  // ../RTL/cortexm0ds_logic.v(1512)
  wire Kreow6;  // ../RTL/cortexm0ds_logic.v(1044)
  wire Krghu6;  // ../RTL/cortexm0ds_logic.v(127)
  wire Krkiu6;  // ../RTL/cortexm0ds_logic.v(581)
  wire Krlow6;  // ../RTL/cortexm0ds_logic.v(1137)
  wire Krlpw6;  // ../RTL/cortexm0ds_logic.v(1591)
  wire Krriu6;  // ../RTL/cortexm0ds_logic.v(675)
  wire Krshu6;  // ../RTL/cortexm0ds_logic.v(207)
  wire Krsow6;  // ../RTL/cortexm0ds_logic.v(1231)
  wire Kryiu6;  // ../RTL/cortexm0ds_logic.v(768)
  wire Krzhu6;  // ../RTL/cortexm0ds_logic.v(300)
  wire Krzow6;  // ../RTL/cortexm0ds_logic.v(1325)
  wire Ks4ju6;  // ../RTL/cortexm0ds_logic.v(849)
  wire Ks5iu6;  // ../RTL/cortexm0ds_logic.v(381)
  wire Ks5pw6;  // ../RTL/cortexm0ds_logic.v(1405)
  wire Ks6ow6;  // ../RTL/cortexm0ds_logic.v(937)
  wire Ksciu6;  // ../RTL/cortexm0ds_logic.v(474)
  wire Kscpw6;  // ../RTL/cortexm0ds_logic.v(1499)
  wire Ksdow6;  // ../RTL/cortexm0ds_logic.v(1031)
  wire Ksgax6;  // ../RTL/cortexm0ds_logic.v(1644)
  wire Kshbx6;  // ../RTL/cortexm0ds_logic.v(1711)
  wire Kshhu6;  // ../RTL/cortexm0ds_logic.v(129)
  wire Ksjiu6;  // ../RTL/cortexm0ds_logic.v(568)
  wire Kskow6;  // ../RTL/cortexm0ds_logic.v(1124)
  wire Ksqiu6;  // ../RTL/cortexm0ds_logic.v(662)
  wire Ksrhu6;  // ../RTL/cortexm0ds_logic.v(194)
  wire Ksrow6;  // ../RTL/cortexm0ds_logic.v(1218)
  wire Kssax6;  // ../RTL/cortexm0ds_logic.v(1666)
  wire Kswpw6;  // ../RTL/cortexm0ds_logic.v(1611)
  wire Ksxiu6;  // ../RTL/cortexm0ds_logic.v(755)
  wire Ksyhu6;  // ../RTL/cortexm0ds_logic.v(287)
  wire Ksyow6;  // ../RTL/cortexm0ds_logic.v(1312)
  wire Kt3ju6;  // ../RTL/cortexm0ds_logic.v(836)
  wire Kt4iu6;  // ../RTL/cortexm0ds_logic.v(368)
  wire Kt4pw6;  // ../RTL/cortexm0ds_logic.v(1392)
  wire Ktbiu6;  // ../RTL/cortexm0ds_logic.v(461)
  wire Ktbpw6;  // ../RTL/cortexm0ds_logic.v(1486)
  wire Ktcow6;  // ../RTL/cortexm0ds_logic.v(1018)
  wire Ktiiu6;  // ../RTL/cortexm0ds_logic.v(555)
  wire Ktjow6;  // ../RTL/cortexm0ds_logic.v(1111)
  wire Ktpiu6;  // ../RTL/cortexm0ds_logic.v(649)
  wire Ktppw6;  // ../RTL/cortexm0ds_logic.v(1598)
  wire Ktqhu6;  // ../RTL/cortexm0ds_logic.v(181)
  wire Ktqow6;  // ../RTL/cortexm0ds_logic.v(1205)
  wire Ktwiu6;  // ../RTL/cortexm0ds_logic.v(742)
  wire Ktxhu6;  // ../RTL/cortexm0ds_logic.v(274)
  wire Ktxow6;  // ../RTL/cortexm0ds_logic.v(1299)
  wire Ku2ju6;  // ../RTL/cortexm0ds_logic.v(823)
  wire Ku3iu6;  // ../RTL/cortexm0ds_logic.v(355)
  wire Ku3pw6;  // ../RTL/cortexm0ds_logic.v(1379)
  wire Ku9ju6;  // ../RTL/cortexm0ds_logic.v(916)
  wire Kuaiu6;  // ../RTL/cortexm0ds_logic.v(448)
  wire Kuapw6;  // ../RTL/cortexm0ds_logic.v(1473)
  wire Kubow6;  // ../RTL/cortexm0ds_logic.v(1005)
  wire Kuhiu6;  // ../RTL/cortexm0ds_logic.v(542)
  wire Kuiow6;  // ../RTL/cortexm0ds_logic.v(1098)
  wire Kuoiu6;  // ../RTL/cortexm0ds_logic.v(636)
  wire Kuphu6;  // ../RTL/cortexm0ds_logic.v(168)
  wire Kupow6;  // ../RTL/cortexm0ds_logic.v(1192)
  wire Kuviu6;  // ../RTL/cortexm0ds_logic.v(729)
  wire Kuwhu6;  // ../RTL/cortexm0ds_logic.v(261)
  wire Kuwow6;  // ../RTL/cortexm0ds_logic.v(1286)
  wire Kv1ju6;  // ../RTL/cortexm0ds_logic.v(810)
  wire Kv2iu6;  // ../RTL/cortexm0ds_logic.v(342)
  wire Kv2pw6;  // ../RTL/cortexm0ds_logic.v(1366)
  wire Kv8ju6;  // ../RTL/cortexm0ds_logic.v(903)
  wire Kv9iu6;  // ../RTL/cortexm0ds_logic.v(435)
  wire Kv9pw6;  // ../RTL/cortexm0ds_logic.v(1460)
  wire Kvaow6;  // ../RTL/cortexm0ds_logic.v(992)
  wire Kvgiu6;  // ../RTL/cortexm0ds_logic.v(529)
  wire Kvhow6;  // ../RTL/cortexm0ds_logic.v(1085)
  wire Kvniu6;  // ../RTL/cortexm0ds_logic.v(623)
  wire Kvohu6;  // ../RTL/cortexm0ds_logic.v(155)
  wire Kvoow6;  // ../RTL/cortexm0ds_logic.v(1179)
  wire Kvuiu6;  // ../RTL/cortexm0ds_logic.v(716)
  wire Kvvhu6;  // ../RTL/cortexm0ds_logic.v(248)
  wire Kvvow6;  // ../RTL/cortexm0ds_logic.v(1273)
  wire Kw0ju6;  // ../RTL/cortexm0ds_logic.v(797)
  wire Kw1iu6;  // ../RTL/cortexm0ds_logic.v(329)
  wire Kw1pw6;  // ../RTL/cortexm0ds_logic.v(1353)
  wire Kw7ju6;  // ../RTL/cortexm0ds_logic.v(890)
  wire Kw8iu6;  // ../RTL/cortexm0ds_logic.v(422)
  wire Kw8pw6;  // ../RTL/cortexm0ds_logic.v(1447)
  wire Kw9ow6;  // ../RTL/cortexm0ds_logic.v(979)
  wire Kwfiu6;  // ../RTL/cortexm0ds_logic.v(516)
  wire Kwgow6;  // ../RTL/cortexm0ds_logic.v(1072)
  wire Kwlpw6;  // ../RTL/cortexm0ds_logic.v(1591)
  wire Kwmiu6;  // ../RTL/cortexm0ds_logic.v(610)
  wire Kwnow6;  // ../RTL/cortexm0ds_logic.v(1166)
  wire Kwtiu6;  // ../RTL/cortexm0ds_logic.v(703)
  wire Kwuhu6;  // ../RTL/cortexm0ds_logic.v(235)
  wire Kwuow6;  // ../RTL/cortexm0ds_logic.v(1260)
  wire Kx0iu6;  // ../RTL/cortexm0ds_logic.v(316)
  wire Kx0pw6;  // ../RTL/cortexm0ds_logic.v(1340)
  wire Kx6ju6;  // ../RTL/cortexm0ds_logic.v(877)
  wire Kx7iu6;  // ../RTL/cortexm0ds_logic.v(409)
  wire Kx7pw6;  // ../RTL/cortexm0ds_logic.v(1434)
  wire Kx8ow6;  // ../RTL/cortexm0ds_logic.v(966)
  wire Kxeax6;  // ../RTL/cortexm0ds_logic.v(1641)
  wire Kxeiu6;  // ../RTL/cortexm0ds_logic.v(503)
  wire Kxfow6;  // ../RTL/cortexm0ds_logic.v(1059)
  wire Kxhpw6;  // ../RTL/cortexm0ds_logic.v(1584)
  wire Kxliu6;  // ../RTL/cortexm0ds_logic.v(597)
  wire Kxmow6;  // ../RTL/cortexm0ds_logic.v(1153)
  wire Kxsiu6;  // ../RTL/cortexm0ds_logic.v(690)
  wire Kxthu6;  // ../RTL/cortexm0ds_logic.v(222)
  wire Kxziu6;  // ../RTL/cortexm0ds_logic.v(784)
  wire Ky5ju6;  // ../RTL/cortexm0ds_logic.v(864)
  wire Ky6iu6;  // ../RTL/cortexm0ds_logic.v(396)
  wire Ky6pw6;  // ../RTL/cortexm0ds_logic.v(1421)
  wire Ky7ow6;  // ../RTL/cortexm0ds_logic.v(953)
  wire Kydiu6;  // ../RTL/cortexm0ds_logic.v(490)
  wire Kydpw6;  // ../RTL/cortexm0ds_logic.v(1514)
  wire Kyeow6;  // ../RTL/cortexm0ds_logic.v(1046)
  wire Kykiu6;  // ../RTL/cortexm0ds_logic.v(584)
  wire Kylow6;  // ../RTL/cortexm0ds_logic.v(1140)
  wire Kyriu6;  // ../RTL/cortexm0ds_logic.v(677)
  wire Kyshu6;  // ../RTL/cortexm0ds_logic.v(209)
  wire Kysow6;  // ../RTL/cortexm0ds_logic.v(1234)
  wire Kyyiu6;  // ../RTL/cortexm0ds_logic.v(771)
  wire Kyzhu6;  // ../RTL/cortexm0ds_logic.v(303)
  wire Kyzow6;  // ../RTL/cortexm0ds_logic.v(1327)
  wire Kz4ju6;  // ../RTL/cortexm0ds_logic.v(851)
  wire Kz5iu6;  // ../RTL/cortexm0ds_logic.v(383)
  wire Kz5pw6;  // ../RTL/cortexm0ds_logic.v(1408)
  wire Kz6ow6;  // ../RTL/cortexm0ds_logic.v(940)
  wire Kzabx6;  // ../RTL/cortexm0ds_logic.v(1699)
  wire Kzciu6;  // ../RTL/cortexm0ds_logic.v(477)
  wire Kzcpw6;  // ../RTL/cortexm0ds_logic.v(1501)
  wire Kzdow6;  // ../RTL/cortexm0ds_logic.v(1033)
  wire Kzjiu6;  // ../RTL/cortexm0ds_logic.v(571)
  wire Kzkhu6;  // ../RTL/cortexm0ds_logic.v(138)
  wire Kzkow6;  // ../RTL/cortexm0ds_logic.v(1127)
  wire Kzqiu6;  // ../RTL/cortexm0ds_logic.v(664)
  wire Kzrhu6;  // ../RTL/cortexm0ds_logic.v(196)
  wire Kzrow6;  // ../RTL/cortexm0ds_logic.v(1221)
  wire Kzxiu6;  // ../RTL/cortexm0ds_logic.v(758)
  wire Kzyhu6;  // ../RTL/cortexm0ds_logic.v(290)
  wire Kzyow6;  // ../RTL/cortexm0ds_logic.v(1314)
  wire L01ju6;  // ../RTL/cortexm0ds_logic.v(798)
  wire L02iu6;  // ../RTL/cortexm0ds_logic.v(330)
  wire L02pw6;  // ../RTL/cortexm0ds_logic.v(1355)
  wire L03qw6;  // ../RTL/cortexm0ds_logic.v(1623)
  wire L08ju6;  // ../RTL/cortexm0ds_logic.v(892)
  wire L09iu6;  // ../RTL/cortexm0ds_logic.v(424)
  wire L09pw6;  // ../RTL/cortexm0ds_logic.v(1448)
  wire L0aow6;  // ../RTL/cortexm0ds_logic.v(980)
  wire L0giu6;  // ../RTL/cortexm0ds_logic.v(517)
  wire L0how6;  // ../RTL/cortexm0ds_logic.v(1074)
  wire L0niu6;  // ../RTL/cortexm0ds_logic.v(611)
  wire L0oow6;  // ../RTL/cortexm0ds_logic.v(1167)
  wire L0uiu6;  // ../RTL/cortexm0ds_logic.v(705)
  wire L0vhu6;  // ../RTL/cortexm0ds_logic.v(237)
  wire L0vow6;  // ../RTL/cortexm0ds_logic.v(1261)
  wire L0ypw6;  // ../RTL/cortexm0ds_logic.v(1613)
  wire L10ju6;  // ../RTL/cortexm0ds_logic.v(785)
  wire L11iu6;  // ../RTL/cortexm0ds_logic.v(317)
  wire L11pw6;  // ../RTL/cortexm0ds_logic.v(1342)
  wire L17ju6;  // ../RTL/cortexm0ds_logic.v(879)
  wire L18iu6;  // ../RTL/cortexm0ds_logic.v(411)
  wire L18pw6;  // ../RTL/cortexm0ds_logic.v(1435)
  wire L19ow6;  // ../RTL/cortexm0ds_logic.v(967)
  wire L1bbx6;  // ../RTL/cortexm0ds_logic.v(1699)
  wire L1fiu6;  // ../RTL/cortexm0ds_logic.v(504)
  wire L1gow6;  // ../RTL/cortexm0ds_logic.v(1061)
  wire L1miu6;  // ../RTL/cortexm0ds_logic.v(598)
  wire L1now6;  // ../RTL/cortexm0ds_logic.v(1154)
  wire L1tiu6;  // ../RTL/cortexm0ds_logic.v(692)
  wire L1uhu6;  // ../RTL/cortexm0ds_logic.v(224)
  wire L1uow6;  // ../RTL/cortexm0ds_logic.v(1248)
  wire L20iu6;  // ../RTL/cortexm0ds_logic.v(304)
  wire L20pw6;  // ../RTL/cortexm0ds_logic.v(1329)
  wire L26ju6;  // ../RTL/cortexm0ds_logic.v(866)
  wire L27iu6;  // ../RTL/cortexm0ds_logic.v(398)
  wire L27pw6;  // ../RTL/cortexm0ds_logic.v(1422)
  wire L28ow6;  // ../RTL/cortexm0ds_logic.v(954)
  wire L2bax6;  // ../RTL/cortexm0ds_logic.v(1633)
  wire L2eiu6;  // ../RTL/cortexm0ds_logic.v(491)
  wire L2epw6;  // ../RTL/cortexm0ds_logic.v(1516)
  wire L2fow6;  // ../RTL/cortexm0ds_logic.v(1048)
  wire L2liu6;  // ../RTL/cortexm0ds_logic.v(585)
  wire L2mow6;  // ../RTL/cortexm0ds_logic.v(1141)
  wire L2siu6;  // ../RTL/cortexm0ds_logic.v(679)
  wire L2thu6;  // ../RTL/cortexm0ds_logic.v(211)
  wire L2tow6;  // ../RTL/cortexm0ds_logic.v(1235)
  wire L2ziu6;  // ../RTL/cortexm0ds_logic.v(772)
  wire L35ju6;  // ../RTL/cortexm0ds_logic.v(853)
  wire L36iu6;  // ../RTL/cortexm0ds_logic.v(385)
  wire L36pw6;  // ../RTL/cortexm0ds_logic.v(1409)
  wire L37ow6;  // ../RTL/cortexm0ds_logic.v(941)
  wire L3bbx6;  // ../RTL/cortexm0ds_logic.v(1699)
  wire L3diu6;  // ../RTL/cortexm0ds_logic.v(478)
  wire L3dpw6;  // ../RTL/cortexm0ds_logic.v(1503)
  wire L3ehu6;  // ../RTL/cortexm0ds_logic.v(121)
  wire L3eow6;  // ../RTL/cortexm0ds_logic.v(1035)
  wire L3kiu6;  // ../RTL/cortexm0ds_logic.v(572)
  wire L3low6;  // ../RTL/cortexm0ds_logic.v(1128)
  wire L3riu6;  // ../RTL/cortexm0ds_logic.v(666)
  wire L3shu6;  // ../RTL/cortexm0ds_logic.v(198)
  wire L3sow6;  // ../RTL/cortexm0ds_logic.v(1222)
  wire L3yiu6;  // ../RTL/cortexm0ds_logic.v(759)
  wire L3zhu6;  // ../RTL/cortexm0ds_logic.v(291)
  wire L3zow6;  // ../RTL/cortexm0ds_logic.v(1316)
  wire L44ju6;  // ../RTL/cortexm0ds_logic.v(840)
  wire L45iu6;  // ../RTL/cortexm0ds_logic.v(372)
  wire L45pw6;  // ../RTL/cortexm0ds_logic.v(1396)
  wire L4ciu6;  // ../RTL/cortexm0ds_logic.v(465)
  wire L4cpw6;  // ../RTL/cortexm0ds_logic.v(1490)
  wire L4dow6;  // ../RTL/cortexm0ds_logic.v(1022)
  wire L4jiu6;  // ../RTL/cortexm0ds_logic.v(559)
  wire L4kow6;  // ../RTL/cortexm0ds_logic.v(1115)
  wire L4lax6;  // ../RTL/cortexm0ds_logic.v(1652)
  wire L4qiu6;  // ../RTL/cortexm0ds_logic.v(653)
  wire L4rhu6;  // ../RTL/cortexm0ds_logic.v(185)
  wire L4row6;  // ../RTL/cortexm0ds_logic.v(1209)
  wire L4xiu6;  // ../RTL/cortexm0ds_logic.v(746)
  wire L4yhu6;  // ../RTL/cortexm0ds_logic.v(278)
  wire L4yow6;  // ../RTL/cortexm0ds_logic.v(1303)
  wire L53ju6;  // ../RTL/cortexm0ds_logic.v(827)
  wire L54iu6;  // ../RTL/cortexm0ds_logic.v(359)
  wire L54pw6;  // ../RTL/cortexm0ds_logic.v(1383)
  wire L5aju6;  // ../RTL/cortexm0ds_logic.v(920)
  wire L5biu6;  // ../RTL/cortexm0ds_logic.v(452)
  wire L5bpw6;  // ../RTL/cortexm0ds_logic.v(1477)
  wire L5cow6;  // ../RTL/cortexm0ds_logic.v(1009)
  wire L5iiu6;  // ../RTL/cortexm0ds_logic.v(546)
  wire L5jow6;  // ../RTL/cortexm0ds_logic.v(1102)
  wire L5lpw6;  // ../RTL/cortexm0ds_logic.v(1590)
  wire L5piu6;  // ../RTL/cortexm0ds_logic.v(640)
  wire L5qhu6;  // ../RTL/cortexm0ds_logic.v(172)
  wire L5qow6;  // ../RTL/cortexm0ds_logic.v(1196)
  wire L5wiu6;  // ../RTL/cortexm0ds_logic.v(733)
  wire L5xhu6;  // ../RTL/cortexm0ds_logic.v(265)
  wire L5xow6;  // ../RTL/cortexm0ds_logic.v(1290)
  wire L62ju6;  // ../RTL/cortexm0ds_logic.v(814)
  wire L63iu6;  // ../RTL/cortexm0ds_logic.v(346)
  wire L63pw6;  // ../RTL/cortexm0ds_logic.v(1370)
  wire L69ju6;  // ../RTL/cortexm0ds_logic.v(907)
  wire L6aiu6;  // ../RTL/cortexm0ds_logic.v(439)
  wire L6apw6;  // ../RTL/cortexm0ds_logic.v(1464)
  wire L6bow6;  // ../RTL/cortexm0ds_logic.v(996)
  wire L6hax6;  // ../RTL/cortexm0ds_logic.v(1645)
  wire L6hiu6;  // ../RTL/cortexm0ds_logic.v(533)
  wire L6iow6;  // ../RTL/cortexm0ds_logic.v(1089)
  wire L6lax6;  // ../RTL/cortexm0ds_logic.v(1653)
  wire L6oiu6;  // ../RTL/cortexm0ds_logic.v(627)
  wire L6phu6;  // ../RTL/cortexm0ds_logic.v(159)
  wire L6pow6;  // ../RTL/cortexm0ds_logic.v(1183)
  wire L6viu6;  // ../RTL/cortexm0ds_logic.v(720)
  wire L6whu6;  // ../RTL/cortexm0ds_logic.v(252)
  wire L6wow6;  // ../RTL/cortexm0ds_logic.v(1277)
  wire L71ju6;  // ../RTL/cortexm0ds_logic.v(801)
  wire L72iu6;  // ../RTL/cortexm0ds_logic.v(333)
  wire L72pw6;  // ../RTL/cortexm0ds_logic.v(1357)
  wire L78ju6;  // ../RTL/cortexm0ds_logic.v(894)
  wire L79iu6;  // ../RTL/cortexm0ds_logic.v(426)
  wire L79pw6;  // ../RTL/cortexm0ds_logic.v(1451)
  wire L7aow6;  // ../RTL/cortexm0ds_logic.v(983)
  wire L7giu6;  // ../RTL/cortexm0ds_logic.v(520)
  wire L7how6;  // ../RTL/cortexm0ds_logic.v(1076)
  wire L7niu6;  // ../RTL/cortexm0ds_logic.v(614)
  wire L7oow6;  // ../RTL/cortexm0ds_logic.v(1170)
  wire L7uiu6;  // ../RTL/cortexm0ds_logic.v(707)
  wire L7vhu6;  // ../RTL/cortexm0ds_logic.v(239)
  wire L7vow6;  // ../RTL/cortexm0ds_logic.v(1264)
  wire L80ju6;  // ../RTL/cortexm0ds_logic.v(788)
  wire L81iu6;  // ../RTL/cortexm0ds_logic.v(320)
  wire L81pw6;  // ../RTL/cortexm0ds_logic.v(1344)
  wire L87ju6;  // ../RTL/cortexm0ds_logic.v(881)
  wire L88iu6;  // ../RTL/cortexm0ds_logic.v(413)
  wire L88pw6;  // ../RTL/cortexm0ds_logic.v(1438)
  wire L89ow6;  // ../RTL/cortexm0ds_logic.v(970)
  wire L8ehu6;  // ../RTL/cortexm0ds_logic.v(121)
  wire L8fiu6;  // ../RTL/cortexm0ds_logic.v(507)
  wire L8gow6;  // ../RTL/cortexm0ds_logic.v(1063)
  wire L8kax6;  // ../RTL/cortexm0ds_logic.v(1651)
  wire L8miu6;  // ../RTL/cortexm0ds_logic.v(601)
  wire L8now6;  // ../RTL/cortexm0ds_logic.v(1157)
  wire L8tiu6;  // ../RTL/cortexm0ds_logic.v(694)
  wire L8uhu6;  // ../RTL/cortexm0ds_logic.v(226)
  wire L8uow6;  // ../RTL/cortexm0ds_logic.v(1251)
  wire L8zax6;  // ../RTL/cortexm0ds_logic.v(1678)
  wire L90iu6;  // ../RTL/cortexm0ds_logic.v(307)
  wire L90pw6;  // ../RTL/cortexm0ds_logic.v(1331)
  wire L96ju6;  // ../RTL/cortexm0ds_logic.v(868)
  wire L97iu6;  // ../RTL/cortexm0ds_logic.v(400)
  wire L97pw6;  // ../RTL/cortexm0ds_logic.v(1425)
  wire L98ow6;  // ../RTL/cortexm0ds_logic.v(957)
  wire L9bbx6;  // ../RTL/cortexm0ds_logic.v(1699)
  wire L9eiu6;  // ../RTL/cortexm0ds_logic.v(494)
  wire L9fow6;  // ../RTL/cortexm0ds_logic.v(1050)
  wire L9liu6;  // ../RTL/cortexm0ds_logic.v(588)
  wire L9mhu6;  // ../RTL/cortexm0ds_logic.v(141)
  wire L9mow6;  // ../RTL/cortexm0ds_logic.v(1144)
  wire L9siu6;  // ../RTL/cortexm0ds_logic.v(681)
  wire L9thu6;  // ../RTL/cortexm0ds_logic.v(213)
  wire L9tow6;  // ../RTL/cortexm0ds_logic.v(1238)
  wire L9xax6;  // ../RTL/cortexm0ds_logic.v(1674)
  wire L9ziu6;  // ../RTL/cortexm0ds_logic.v(775)
  wire La5ju6;  // ../RTL/cortexm0ds_logic.v(855)
  wire La6iu6;  // ../RTL/cortexm0ds_logic.v(387)
  wire La6pw6;  // ../RTL/cortexm0ds_logic.v(1412)
  wire La7ow6;  // ../RTL/cortexm0ds_logic.v(944)
  wire Ladiu6;  // ../RTL/cortexm0ds_logic.v(481)
  wire Ladpw6;  // ../RTL/cortexm0ds_logic.v(1505)
  wire Laeow6;  // ../RTL/cortexm0ds_logic.v(1037)
  wire Lakiu6;  // ../RTL/cortexm0ds_logic.v(575)
  wire Lalow6;  // ../RTL/cortexm0ds_logic.v(1131)
  wire Lariu6;  // ../RTL/cortexm0ds_logic.v(668)
  wire Lashu6;  // ../RTL/cortexm0ds_logic.v(200)
  wire Lasow6;  // ../RTL/cortexm0ds_logic.v(1225)
  wire Layiu6;  // ../RTL/cortexm0ds_logic.v(762)
  wire Lazhu6;  // ../RTL/cortexm0ds_logic.v(294)
  wire Lazow6;  // ../RTL/cortexm0ds_logic.v(1318)
  wire Lb4ju6;  // ../RTL/cortexm0ds_logic.v(842)
  wire Lb5iu6;  // ../RTL/cortexm0ds_logic.v(374)
  wire Lb5pw6;  // ../RTL/cortexm0ds_logic.v(1399)
  wire Lb6ow6;  // ../RTL/cortexm0ds_logic.v(931)
  wire Lbbax6;  // ../RTL/cortexm0ds_logic.v(1634)
  wire Lbciu6;  // ../RTL/cortexm0ds_logic.v(468)
  wire Lbcpw6;  // ../RTL/cortexm0ds_logic.v(1492)
  wire Lbdow6;  // ../RTL/cortexm0ds_logic.v(1024)
  wire Lbjiu6;  // ../RTL/cortexm0ds_logic.v(562)
  wire Lbkow6;  // ../RTL/cortexm0ds_logic.v(1118)
  wire Lbqiu6;  // ../RTL/cortexm0ds_logic.v(655)
  wire Lbrhu6;  // ../RTL/cortexm0ds_logic.v(187)
  wire Lbrow6;  // ../RTL/cortexm0ds_logic.v(1212)
  wire Lbxiu6;  // ../RTL/cortexm0ds_logic.v(749)
  wire Lbyhu6;  // ../RTL/cortexm0ds_logic.v(281)
  wire Lbyow6;  // ../RTL/cortexm0ds_logic.v(1305)
  wire Lc3ju6;  // ../RTL/cortexm0ds_logic.v(829)
  wire Lc4iu6;  // ../RTL/cortexm0ds_logic.v(361)
  wire Lc4pw6;  // ../RTL/cortexm0ds_logic.v(1386)
  wire Lcaju6;  // ../RTL/cortexm0ds_logic.v(923)
  wire Lcbiu6;  // ../RTL/cortexm0ds_logic.v(455)
  wire Lcbpw6;  // ../RTL/cortexm0ds_logic.v(1479)
  wire Lccow6;  // ../RTL/cortexm0ds_logic.v(1011)
  wire Lciiu6;  // ../RTL/cortexm0ds_logic.v(549)
  wire Lcjow6;  // ../RTL/cortexm0ds_logic.v(1105)
  wire Lclhu6;  // ../RTL/cortexm0ds_logic.v(139)
  wire Lcpiu6;  // ../RTL/cortexm0ds_logic.v(642)
  wire Lcqhu6;  // ../RTL/cortexm0ds_logic.v(174)
  wire Lcqow6;  // ../RTL/cortexm0ds_logic.v(1199)
  wire Lcwiu6;  // ../RTL/cortexm0ds_logic.v(736)
  wire Lcxhu6;  // ../RTL/cortexm0ds_logic.v(268)
  wire Lcxow6;  // ../RTL/cortexm0ds_logic.v(1292)
  wire Ld2ju6;  // ../RTL/cortexm0ds_logic.v(816)
  wire Ld3iu6;  // ../RTL/cortexm0ds_logic.v(348)
  wire Ld3pw6;  // ../RTL/cortexm0ds_logic.v(1373)
  wire Ld9ju6;  // ../RTL/cortexm0ds_logic.v(910)
  wire Ldaiu6;  // ../RTL/cortexm0ds_logic.v(442)
  wire Ldapw6;  // ../RTL/cortexm0ds_logic.v(1466)
  wire Ldbow6;  // ../RTL/cortexm0ds_logic.v(998)
  wire Ldhiu6;  // ../RTL/cortexm0ds_logic.v(536)
  wire Ldiow6;  // ../RTL/cortexm0ds_logic.v(1092)
  wire Ldoax6;  // ../RTL/cortexm0ds_logic.v(1658)
  wire Ldoiu6;  // ../RTL/cortexm0ds_logic.v(629)
  wire Ldphu6;  // ../RTL/cortexm0ds_logic.v(161)
  wire Ldpow6;  // ../RTL/cortexm0ds_logic.v(1186)
  wire Ldviu6;  // ../RTL/cortexm0ds_logic.v(723)
  wire Ldvpw6;  // ../RTL/cortexm0ds_logic.v(1608)
  wire Ldwax6;  // ../RTL/cortexm0ds_logic.v(1673)
  wire Ldwhu6;  // ../RTL/cortexm0ds_logic.v(255)
  wire Ldwow6;  // ../RTL/cortexm0ds_logic.v(1279)
  wire Le1ju6;  // ../RTL/cortexm0ds_logic.v(803)
  wire Le2iu6;  // ../RTL/cortexm0ds_logic.v(335)
  wire Le2pw6;  // ../RTL/cortexm0ds_logic.v(1360)
  wire Le2qw6;  // ../RTL/cortexm0ds_logic.v(1621)
  wire Le8ju6;  // ../RTL/cortexm0ds_logic.v(897)
  wire Le9iu6;  // ../RTL/cortexm0ds_logic.v(429)
  wire Le9pw6;  // ../RTL/cortexm0ds_logic.v(1453)
  wire Leaow6;  // ../RTL/cortexm0ds_logic.v(985)
  wire Legiu6;  // ../RTL/cortexm0ds_logic.v(523)
  wire Lehow6;  // ../RTL/cortexm0ds_logic.v(1079)
  wire Leniu6;  // ../RTL/cortexm0ds_logic.v(616)
  wire Leohu6;  // ../RTL/cortexm0ds_logic.v(148)
  wire Leoow6;  // ../RTL/cortexm0ds_logic.v(1173)
  wire Lerpw6;  // ../RTL/cortexm0ds_logic.v(1601)
  wire Leuiu6;  // ../RTL/cortexm0ds_logic.v(710)
  wire Levhu6;  // ../RTL/cortexm0ds_logic.v(242)
  wire Levow6;  // ../RTL/cortexm0ds_logic.v(1266)
  wire Lf0ju6;  // ../RTL/cortexm0ds_logic.v(790)
  wire Lf1iu6;  // ../RTL/cortexm0ds_logic.v(322)
  wire Lf1pw6;  // ../RTL/cortexm0ds_logic.v(1347)
  wire Lf7ju6;  // ../RTL/cortexm0ds_logic.v(884)
  wire Lf8iu6;  // ../RTL/cortexm0ds_logic.v(416)
  wire Lf8pw6;  // ../RTL/cortexm0ds_logic.v(1440)
  wire Lf9ow6;  // ../RTL/cortexm0ds_logic.v(972)
  wire Lffiu6;  // ../RTL/cortexm0ds_logic.v(510)
  wire Lfgbx6;  // ../RTL/cortexm0ds_logic.v(1709)
  wire Lfgow6;  // ../RTL/cortexm0ds_logic.v(1066)
  wire Lfmiu6;  // ../RTL/cortexm0ds_logic.v(603)
  wire Lfnow6;  // ../RTL/cortexm0ds_logic.v(1160)
  wire Lfppw6;  // ../RTL/cortexm0ds_logic.v(1598)
  wire Lftiu6;  // ../RTL/cortexm0ds_logic.v(697)
  wire Lfuhu6;  // ../RTL/cortexm0ds_logic.v(229)
  wire Lfuow6;  // ../RTL/cortexm0ds_logic.v(1253)
  wire Lfwax6;  // ../RTL/cortexm0ds_logic.v(1673)
  wire Lg0iu6;  // ../RTL/cortexm0ds_logic.v(309)
  wire Lg0pw6;  // ../RTL/cortexm0ds_logic.v(1334)
  wire Lg1bx6;  // ../RTL/cortexm0ds_logic.v(1682)
  wire Lg6ju6;  // ../RTL/cortexm0ds_logic.v(871)
  wire Lg7iu6;  // ../RTL/cortexm0ds_logic.v(403)
  wire Lg7pw6;  // ../RTL/cortexm0ds_logic.v(1427)
  wire Lg8ow6;  // ../RTL/cortexm0ds_logic.v(959)
  wire Lg9bx6;  // ../RTL/cortexm0ds_logic.v(1696)
  wire Lgeiu6;  // ../RTL/cortexm0ds_logic.v(497)
  wire Lgfow6;  // ../RTL/cortexm0ds_logic.v(1053)
  wire Lgkax6;  // ../RTL/cortexm0ds_logic.v(1651)
  wire Lgliu6;  // ../RTL/cortexm0ds_logic.v(590)
  wire Lgmow6;  // ../RTL/cortexm0ds_logic.v(1147)
  wire Lgsiu6;  // ../RTL/cortexm0ds_logic.v(684)
  wire Lgthu6;  // ../RTL/cortexm0ds_logic.v(216)
  wire Lgtow6;  // ../RTL/cortexm0ds_logic.v(1240)
  wire Lgziu6;  // ../RTL/cortexm0ds_logic.v(777)
  wire Lh5ju6;  // ../RTL/cortexm0ds_logic.v(858)
  wire Lh6iu6;  // ../RTL/cortexm0ds_logic.v(390)
  wire Lh6pw6;  // ../RTL/cortexm0ds_logic.v(1414)
  wire Lh7ow6;  // ../RTL/cortexm0ds_logic.v(946)
  wire Lhbbx6;  // ../RTL/cortexm0ds_logic.v(1700)
  wire Lhdiu6;  // ../RTL/cortexm0ds_logic.v(484)
  wire Lhdpw6;  // ../RTL/cortexm0ds_logic.v(1508)
  wire Lheow6;  // ../RTL/cortexm0ds_logic.v(1040)
  wire Lhkiu6;  // ../RTL/cortexm0ds_logic.v(577)
  wire Lhlow6;  // ../RTL/cortexm0ds_logic.v(1134)
  wire Lhppw6;  // ../RTL/cortexm0ds_logic.v(1598)
  wire Lhriu6;  // ../RTL/cortexm0ds_logic.v(671)
  wire Lhshu6;  // ../RTL/cortexm0ds_logic.v(203)
  wire Lhsow6;  // ../RTL/cortexm0ds_logic.v(1227)
  wire Lhwax6;  // ../RTL/cortexm0ds_logic.v(1673)
  wire Lhyiu6;  // ../RTL/cortexm0ds_logic.v(764)
  wire Lhzhu6;  // ../RTL/cortexm0ds_logic.v(296)
  wire Lhzow6;  // ../RTL/cortexm0ds_logic.v(1321)
  wire Li2bx6;  // ../RTL/cortexm0ds_logic.v(1684)
  wire Li4ju6;  // ../RTL/cortexm0ds_logic.v(845)
  wire Li5iu6;  // ../RTL/cortexm0ds_logic.v(377)
  wire Li5pw6;  // ../RTL/cortexm0ds_logic.v(1401)
  wire Li6ow6;  // ../RTL/cortexm0ds_logic.v(933)
  wire Li7ax6;  // ../RTL/cortexm0ds_logic.v(1626)
  wire Liabx6;  // ../RTL/cortexm0ds_logic.v(1698)
  wire Liciu6;  // ../RTL/cortexm0ds_logic.v(471)
  wire Licpw6;  // ../RTL/cortexm0ds_logic.v(1495)
  wire Lidow6;  // ../RTL/cortexm0ds_logic.v(1027)
  wire Lijiu6;  // ../RTL/cortexm0ds_logic.v(564)
  wire Likow6;  // ../RTL/cortexm0ds_logic.v(1121)
  wire Liqiu6;  // ../RTL/cortexm0ds_logic.v(658)
  wire Lirhu6;  // ../RTL/cortexm0ds_logic.v(190)
  wire Lirow6;  // ../RTL/cortexm0ds_logic.v(1214)
  wire Lixiu6;  // ../RTL/cortexm0ds_logic.v(751)
  wire Liyhu6;  // ../RTL/cortexm0ds_logic.v(283)
  wire Liyow6;  // ../RTL/cortexm0ds_logic.v(1308)
  wire Lj3ju6;  // ../RTL/cortexm0ds_logic.v(832)
  wire Lj4iu6;  // ../RTL/cortexm0ds_logic.v(364)
  wire Lj4pw6;  // ../RTL/cortexm0ds_logic.v(1388)
  wire Ljaju6;  // ../RTL/cortexm0ds_logic.v(926)
  wire Ljbiu6;  // ../RTL/cortexm0ds_logic.v(458)
  wire Ljbpw6;  // ../RTL/cortexm0ds_logic.v(1482)
  wire Ljcax6;  // ../RTL/cortexm0ds_logic.v(1636)
  wire Ljcow6;  // ../RTL/cortexm0ds_logic.v(1014)
  wire Ljiiu6;  // ../RTL/cortexm0ds_logic.v(551)
  wire Ljjow6;  // ../RTL/cortexm0ds_logic.v(1108)
  wire Ljpiu6;  // ../RTL/cortexm0ds_logic.v(645)
  wire Ljppw6;  // ../RTL/cortexm0ds_logic.v(1598)
  wire Ljqhu6;  // ../RTL/cortexm0ds_logic.v(177)
  wire Ljqow6;  // ../RTL/cortexm0ds_logic.v(1201)
  wire Ljwax6;  // ../RTL/cortexm0ds_logic.v(1673)
  wire Ljwiu6;  // ../RTL/cortexm0ds_logic.v(738)
  wire Ljxhu6;  // ../RTL/cortexm0ds_logic.v(270)
  wire Ljxow6;  // ../RTL/cortexm0ds_logic.v(1295)
  wire Lk2ju6;  // ../RTL/cortexm0ds_logic.v(819)
  wire Lk3iu6;  // ../RTL/cortexm0ds_logic.v(351)
  wire Lk3pw6;  // ../RTL/cortexm0ds_logic.v(1375)
  wire Lk9ax6;  // ../RTL/cortexm0ds_logic.v(1630)
  wire Lk9ju6;  // ../RTL/cortexm0ds_logic.v(913)
  wire Lkaiu6;  // ../RTL/cortexm0ds_logic.v(445)
  wire Lkapw6;  // ../RTL/cortexm0ds_logic.v(1469)
  wire Lkbow6;  // ../RTL/cortexm0ds_logic.v(1001)
  wire Lkhiu6;  // ../RTL/cortexm0ds_logic.v(538)
  wire Lkiow6;  // ../RTL/cortexm0ds_logic.v(1095)
  wire Lkoiu6;  // ../RTL/cortexm0ds_logic.v(632)
  wire Lkphu6;  // ../RTL/cortexm0ds_logic.v(164)
  wire Lkpow6;  // ../RTL/cortexm0ds_logic.v(1188)
  wire Lksax6;  // ../RTL/cortexm0ds_logic.v(1666)
  wire Lkviu6;  // ../RTL/cortexm0ds_logic.v(725)
  wire Lkwhu6;  // ../RTL/cortexm0ds_logic.v(257)
  wire Lkwow6;  // ../RTL/cortexm0ds_logic.v(1282)
  wire Ll1ju6;  // ../RTL/cortexm0ds_logic.v(806)
  wire Ll2iu6;  // ../RTL/cortexm0ds_logic.v(338)
  wire Ll2pw6;  // ../RTL/cortexm0ds_logic.v(1362)
  wire Ll8ju6;  // ../RTL/cortexm0ds_logic.v(900)
  wire Ll9iu6;  // ../RTL/cortexm0ds_logic.v(432)
  wire Ll9pw6;  // ../RTL/cortexm0ds_logic.v(1456)
  wire Llaow6;  // ../RTL/cortexm0ds_logic.v(988)
  wire Llgiu6;  // ../RTL/cortexm0ds_logic.v(525)
  wire Llhow6;  // ../RTL/cortexm0ds_logic.v(1082)
  wire Llniu6;  // ../RTL/cortexm0ds_logic.v(619)
  wire Llohu6;  // ../RTL/cortexm0ds_logic.v(151)
  wire Lloow6;  // ../RTL/cortexm0ds_logic.v(1175)
  wire Llppw6;  // ../RTL/cortexm0ds_logic.v(1598)
  wire Lluiu6;  // ../RTL/cortexm0ds_logic.v(712)
  wire Llvhu6;  // ../RTL/cortexm0ds_logic.v(244)
  wire Llvow6;  // ../RTL/cortexm0ds_logic.v(1269)
  wire Llwax6;  // ../RTL/cortexm0ds_logic.v(1673)
  wire Lm0ju6;  // ../RTL/cortexm0ds_logic.v(793)
  wire Lm1iu6;  // ../RTL/cortexm0ds_logic.v(325)
  wire Lm1pw6;  // ../RTL/cortexm0ds_logic.v(1349)
  wire Lm7ju6;  // ../RTL/cortexm0ds_logic.v(887)
  wire Lm8iu6;  // ../RTL/cortexm0ds_logic.v(419)
  wire Lm8pw6;  // ../RTL/cortexm0ds_logic.v(1443)
  wire Lm9ow6;  // ../RTL/cortexm0ds_logic.v(975)
  wire Lmfiu6;  // ../RTL/cortexm0ds_logic.v(512)
  wire Lmgow6;  // ../RTL/cortexm0ds_logic.v(1069)
  wire Lmkbx6;  // ../RTL/cortexm0ds_logic.v(1717)
  wire Lmmiu6;  // ../RTL/cortexm0ds_logic.v(606)
  wire Lmnow6;  // ../RTL/cortexm0ds_logic.v(1162)
  wire Lmtiu6;  // ../RTL/cortexm0ds_logic.v(699)
  wire Lmuhu6;  // ../RTL/cortexm0ds_logic.v(231)
  wire Lmuow6;  // ../RTL/cortexm0ds_logic.v(1256)
  wire Ln0bx6;  // ../RTL/cortexm0ds_logic.v(1680)
  wire Ln0iu6;  // ../RTL/cortexm0ds_logic.v(312)
  wire Ln0pw6;  // ../RTL/cortexm0ds_logic.v(1336)
  wire Ln6ju6;  // ../RTL/cortexm0ds_logic.v(874)
  wire Ln7iu6;  // ../RTL/cortexm0ds_logic.v(406)
  wire Ln7pw6;  // ../RTL/cortexm0ds_logic.v(1430)
  wire Ln8ow6;  // ../RTL/cortexm0ds_logic.v(962)
  wire Lneiu6;  // ../RTL/cortexm0ds_logic.v(499)
  wire Lnfow6;  // ../RTL/cortexm0ds_logic.v(1056)
  wire Lnliu6;  // ../RTL/cortexm0ds_logic.v(593)
  wire Lnmow6;  // ../RTL/cortexm0ds_logic.v(1149)
  wire Lnppw6;  // ../RTL/cortexm0ds_logic.v(1598)
  wire Lnsiu6;  // ../RTL/cortexm0ds_logic.v(686)
  wire Lnthu6;  // ../RTL/cortexm0ds_logic.v(218)
  wire Lntow6;  // ../RTL/cortexm0ds_logic.v(1243)
  wire Lnwax6;  // ../RTL/cortexm0ds_logic.v(1673)
  wire Lnziu6;  // ../RTL/cortexm0ds_logic.v(780)
  wire Lo5ju6;  // ../RTL/cortexm0ds_logic.v(861)
  wire Lo6iu6;  // ../RTL/cortexm0ds_logic.v(393)
  wire Lo6pw6;  // ../RTL/cortexm0ds_logic.v(1417)
  wire Lo7ow6;  // ../RTL/cortexm0ds_logic.v(949)
  wire Lodiu6;  // ../RTL/cortexm0ds_logic.v(486)
  wire Lodpw6;  // ../RTL/cortexm0ds_logic.v(1511)
  wire Loeow6;  // ../RTL/cortexm0ds_logic.v(1043)
  wire Lokiu6;  // ../RTL/cortexm0ds_logic.v(580)
  wire Lolow6;  // ../RTL/cortexm0ds_logic.v(1136)
  wire Loriu6;  // ../RTL/cortexm0ds_logic.v(673)
  wire Loshu6;  // ../RTL/cortexm0ds_logic.v(205)
  wire Losow6;  // ../RTL/cortexm0ds_logic.v(1230)
  wire Loyiu6;  // ../RTL/cortexm0ds_logic.v(767)
  wire Lozhu6;  // ../RTL/cortexm0ds_logic.v(299)
  wire Lozow6;  // ../RTL/cortexm0ds_logic.v(1323)
  wire Lp4ju6;  // ../RTL/cortexm0ds_logic.v(848)
  wire Lp5iu6;  // ../RTL/cortexm0ds_logic.v(380)
  wire Lp5pw6;  // ../RTL/cortexm0ds_logic.v(1404)
  wire Lp6ow6;  // ../RTL/cortexm0ds_logic.v(936)
  wire Lp7ax6;  // ../RTL/cortexm0ds_logic.v(1627)
  wire Lpciu6;  // ../RTL/cortexm0ds_logic.v(473)
  wire Lpcpw6;  // ../RTL/cortexm0ds_logic.v(1498)
  wire Lpdow6;  // ../RTL/cortexm0ds_logic.v(1030)
  wire Lpjiu6;  // ../RTL/cortexm0ds_logic.v(567)
  wire Lpkow6;  // ../RTL/cortexm0ds_logic.v(1123)
  wire Lpppw6;  // ../RTL/cortexm0ds_logic.v(1598)
  wire Lpqiu6;  // ../RTL/cortexm0ds_logic.v(660)
  wire Lprhu6;  // ../RTL/cortexm0ds_logic.v(192)
  wire Lprow6;  // ../RTL/cortexm0ds_logic.v(1217)
  wire Lpwax6;  // ../RTL/cortexm0ds_logic.v(1673)
  wire Lpxiu6;  // ../RTL/cortexm0ds_logic.v(754)
  wire Lpyhu6;  // ../RTL/cortexm0ds_logic.v(286)
  wire Lpyow6;  // ../RTL/cortexm0ds_logic.v(1310)
  wire Lq3ju6;  // ../RTL/cortexm0ds_logic.v(835)
  wire Lq4iu6;  // ../RTL/cortexm0ds_logic.v(367)
  wire Lq4pw6;  // ../RTL/cortexm0ds_logic.v(1391)
  wire Lqaju6;  // ../RTL/cortexm0ds_logic.v(928)
  wire Lqbiu6;  // ../RTL/cortexm0ds_logic.v(460)
  wire Lqbpw6;  // ../RTL/cortexm0ds_logic.v(1485)
  wire Lqcow6;  // ../RTL/cortexm0ds_logic.v(1017)
  wire Lqiiu6;  // ../RTL/cortexm0ds_logic.v(554)
  wire Lqjow6;  // ../RTL/cortexm0ds_logic.v(1110)
  wire Lqjpw6;  // ../RTL/cortexm0ds_logic.v(1587)
  wire Lqpiu6;  // ../RTL/cortexm0ds_logic.v(647)
  wire Lqqhu6;  // ../RTL/cortexm0ds_logic.v(179)
  wire Lqqow6;  // ../RTL/cortexm0ds_logic.v(1204)
  wire Lqwiu6;  // ../RTL/cortexm0ds_logic.v(741)
  wire Lqxhu6;  // ../RTL/cortexm0ds_logic.v(273)
  wire Lqxow6;  // ../RTL/cortexm0ds_logic.v(1297)
  wire Lr2ju6;  // ../RTL/cortexm0ds_logic.v(822)
  wire Lr3iu6;  // ../RTL/cortexm0ds_logic.v(354)
  wire Lr3pw6;  // ../RTL/cortexm0ds_logic.v(1378)
  wire Lr9bx6;  // ../RTL/cortexm0ds_logic.v(1697)
  wire Lr9ju6;  // ../RTL/cortexm0ds_logic.v(915)
  wire Lraiu6;  // ../RTL/cortexm0ds_logic.v(447)
  wire Lrapw6;  // ../RTL/cortexm0ds_logic.v(1472)
  wire Lrbow6;  // ../RTL/cortexm0ds_logic.v(1004)
  wire Lrhiu6;  // ../RTL/cortexm0ds_logic.v(541)
  wire Lriow6;  // ../RTL/cortexm0ds_logic.v(1097)
  wire Lroiu6;  // ../RTL/cortexm0ds_logic.v(634)
  wire Lrphu6;  // ../RTL/cortexm0ds_logic.v(166)
  wire Lrpow6;  // ../RTL/cortexm0ds_logic.v(1191)
  wire Lrppw6;  // ../RTL/cortexm0ds_logic.v(1598)
  wire Lrviu6;  // ../RTL/cortexm0ds_logic.v(728)
  wire Lrwax6;  // ../RTL/cortexm0ds_logic.v(1674)
  wire Lrwhu6;  // ../RTL/cortexm0ds_logic.v(260)
  wire Lrwow6;  // ../RTL/cortexm0ds_logic.v(1284)
  wire Ls1ju6;  // ../RTL/cortexm0ds_logic.v(809)
  wire Ls2iu6;  // ../RTL/cortexm0ds_logic.v(341)
  wire Ls2pw6;  // ../RTL/cortexm0ds_logic.v(1365)
  wire Ls8ju6;  // ../RTL/cortexm0ds_logic.v(902)
  wire Ls9iu6;  // ../RTL/cortexm0ds_logic.v(434)
  wire Ls9pw6;  // ../RTL/cortexm0ds_logic.v(1459)
  wire Lsaow6;  // ../RTL/cortexm0ds_logic.v(991)
  wire Lsgiu6;  // ../RTL/cortexm0ds_logic.v(528)
  wire Lshow6;  // ../RTL/cortexm0ds_logic.v(1084)
  wire Lsniu6;  // ../RTL/cortexm0ds_logic.v(621)
  wire Lsohu6;  // ../RTL/cortexm0ds_logic.v(153)
  wire Lsoow6;  // ../RTL/cortexm0ds_logic.v(1178)
  wire Lsuiu6;  // ../RTL/cortexm0ds_logic.v(715)
  wire Lsvhu6;  // ../RTL/cortexm0ds_logic.v(247)
  wire Lsvow6;  // ../RTL/cortexm0ds_logic.v(1271)
  wire Lt0ju6;  // ../RTL/cortexm0ds_logic.v(796)
  wire Lt1iu6;  // ../RTL/cortexm0ds_logic.v(328)
  wire Lt1pw6;  // ../RTL/cortexm0ds_logic.v(1352)
  wire Lt7ju6;  // ../RTL/cortexm0ds_logic.v(889)
  wire Lt8iu6;  // ../RTL/cortexm0ds_logic.v(421)
  wire Lt8pw6;  // ../RTL/cortexm0ds_logic.v(1446)
  wire Lt9ow6;  // ../RTL/cortexm0ds_logic.v(978)
  wire Ltfiu6;  // ../RTL/cortexm0ds_logic.v(515)
  wire Ltgow6;  // ../RTL/cortexm0ds_logic.v(1071)
  wire Ltmiu6;  // ../RTL/cortexm0ds_logic.v(608)
  wire Ltnow6;  // ../RTL/cortexm0ds_logic.v(1165)
  wire Lttiu6;  // ../RTL/cortexm0ds_logic.v(702)
  wire Ltuhu6;  // ../RTL/cortexm0ds_logic.v(234)
  wire Ltuow6;  // ../RTL/cortexm0ds_logic.v(1258)
  wire Ltwax6;  // ../RTL/cortexm0ds_logic.v(1674)
  wire Lu0iu6;  // ../RTL/cortexm0ds_logic.v(315)
  wire Lu0pw6;  // ../RTL/cortexm0ds_logic.v(1339)
  wire Lu6ju6;  // ../RTL/cortexm0ds_logic.v(876)
  wire Lu7iu6;  // ../RTL/cortexm0ds_logic.v(408)
  wire Lu7pw6;  // ../RTL/cortexm0ds_logic.v(1433)
  wire Lu8ow6;  // ../RTL/cortexm0ds_logic.v(965)
  wire Lueiu6;  // ../RTL/cortexm0ds_logic.v(502)
  wire Lufow6;  // ../RTL/cortexm0ds_logic.v(1058)
  wire Luliu6;  // ../RTL/cortexm0ds_logic.v(595)
  wire Lumow6;  // ../RTL/cortexm0ds_logic.v(1152)
  wire Lusiu6;  // ../RTL/cortexm0ds_logic.v(689)
  wire Luthu6;  // ../RTL/cortexm0ds_logic.v(221)
  wire Lutow6;  // ../RTL/cortexm0ds_logic.v(1245)
  wire Luziu6;  // ../RTL/cortexm0ds_logic.v(783)
  wire Lv5ju6;  // ../RTL/cortexm0ds_logic.v(863)
  wire Lv6iu6;  // ../RTL/cortexm0ds_logic.v(395)
  wire Lv6pw6;  // ../RTL/cortexm0ds_logic.v(1420)
  wire Lv7ow6;  // ../RTL/cortexm0ds_logic.v(952)
  wire Lvdiu6;  // ../RTL/cortexm0ds_logic.v(489)
  wire Lvdpw6;  // ../RTL/cortexm0ds_logic.v(1513)
  wire Lveow6;  // ../RTL/cortexm0ds_logic.v(1045)
  wire Lvkiu6;  // ../RTL/cortexm0ds_logic.v(582)
  wire Lvlow6;  // ../RTL/cortexm0ds_logic.v(1139)
  wire Lvriu6;  // ../RTL/cortexm0ds_logic.v(676)
  wire Lvshu6;  // ../RTL/cortexm0ds_logic.v(208)
  wire Lvsow6;  // ../RTL/cortexm0ds_logic.v(1232)
  wire Lvwax6;  // ../RTL/cortexm0ds_logic.v(1674)
  wire Lvyiu6;  // ../RTL/cortexm0ds_logic.v(770)
  wire Lvzhu6;  // ../RTL/cortexm0ds_logic.v(302)
  wire Lvzow6;  // ../RTL/cortexm0ds_logic.v(1326)
  wire Lw4ju6;  // ../RTL/cortexm0ds_logic.v(850)
  wire Lw5iu6;  // ../RTL/cortexm0ds_logic.v(382)
  wire Lw5pw6;  // ../RTL/cortexm0ds_logic.v(1407)
  wire Lw6ow6;  // ../RTL/cortexm0ds_logic.v(939)
  wire Lwciu6;  // ../RTL/cortexm0ds_logic.v(476)
  wire Lwcpw6;  // ../RTL/cortexm0ds_logic.v(1500)
  wire Lwdow6;  // ../RTL/cortexm0ds_logic.v(1032)
  wire Lwjiu6;  // ../RTL/cortexm0ds_logic.v(569)
  wire Lwkow6;  // ../RTL/cortexm0ds_logic.v(1126)
  wire Lwqiu6;  // ../RTL/cortexm0ds_logic.v(663)
  wire Lwrhu6;  // ../RTL/cortexm0ds_logic.v(195)
  wire Lwrow6;  // ../RTL/cortexm0ds_logic.v(1219)
  wire Lwxiu6;  // ../RTL/cortexm0ds_logic.v(757)
  wire Lwyhu6;  // ../RTL/cortexm0ds_logic.v(289)
  wire Lwyow6;  // ../RTL/cortexm0ds_logic.v(1313)
  wire Lx3ju6;  // ../RTL/cortexm0ds_logic.v(837)
  wire Lx4iu6;  // ../RTL/cortexm0ds_logic.v(369)
  wire Lx4pw6;  // ../RTL/cortexm0ds_logic.v(1394)
  wire Lx9ax6;  // ../RTL/cortexm0ds_logic.v(1631)
  wire Lxbiu6;  // ../RTL/cortexm0ds_logic.v(463)
  wire Lxbpw6;  // ../RTL/cortexm0ds_logic.v(1487)
  wire Lxcow6;  // ../RTL/cortexm0ds_logic.v(1019)
  wire Lxiiu6;  // ../RTL/cortexm0ds_logic.v(556)
  wire Lxjow6;  // ../RTL/cortexm0ds_logic.v(1113)
  wire Lxpiu6;  // ../RTL/cortexm0ds_logic.v(650)
  wire Lxqhu6;  // ../RTL/cortexm0ds_logic.v(182)
  wire Lxqow6;  // ../RTL/cortexm0ds_logic.v(1206)
  wire Lxwax6;  // ../RTL/cortexm0ds_logic.v(1674)
  wire Lxwiu6;  // ../RTL/cortexm0ds_logic.v(744)
  wire Lxxhu6;  // ../RTL/cortexm0ds_logic.v(276)
  wire Lxxow6;  // ../RTL/cortexm0ds_logic.v(1300)
  wire Ly2ju6;  // ../RTL/cortexm0ds_logic.v(824)
  wire Ly3iu6;  // ../RTL/cortexm0ds_logic.v(356)
  wire Ly3pw6;  // ../RTL/cortexm0ds_logic.v(1381)
  wire Ly9ju6;  // ../RTL/cortexm0ds_logic.v(918)
  wire Lyaiu6;  // ../RTL/cortexm0ds_logic.v(450)
  wire Lyapw6;  // ../RTL/cortexm0ds_logic.v(1474)
  wire Lybow6;  // ../RTL/cortexm0ds_logic.v(1006)
  wire Lycax6;  // ../RTL/cortexm0ds_logic.v(1637)
  wire Lyhiu6;  // ../RTL/cortexm0ds_logic.v(543)
  wire Lyiow6;  // ../RTL/cortexm0ds_logic.v(1100)
  wire Lyoiu6;  // ../RTL/cortexm0ds_logic.v(637)
  wire Lyphu6;  // ../RTL/cortexm0ds_logic.v(169)
  wire Lypow6;  // ../RTL/cortexm0ds_logic.v(1193)
  wire Lyviu6;  // ../RTL/cortexm0ds_logic.v(731)
  wire Lywhu6;  // ../RTL/cortexm0ds_logic.v(263)
  wire Lywow6;  // ../RTL/cortexm0ds_logic.v(1287)
  wire Lywpw6;  // ../RTL/cortexm0ds_logic.v(1611)
  wire Lz1ju6;  // ../RTL/cortexm0ds_logic.v(811)
  wire Lz2iu6;  // ../RTL/cortexm0ds_logic.v(343)
  wire Lz2pw6;  // ../RTL/cortexm0ds_logic.v(1368)
  wire Lz8ju6;  // ../RTL/cortexm0ds_logic.v(905)
  wire Lz9iu6;  // ../RTL/cortexm0ds_logic.v(437)
  wire Lz9pw6;  // ../RTL/cortexm0ds_logic.v(1461)
  wire Lzaow6;  // ../RTL/cortexm0ds_logic.v(993)
  wire Lzgiu6;  // ../RTL/cortexm0ds_logic.v(530)
  wire Lzhow6;  // ../RTL/cortexm0ds_logic.v(1087)
  wire Lznhu6;  // ../RTL/cortexm0ds_logic.v(146)
  wire Lzniu6;  // ../RTL/cortexm0ds_logic.v(624)
  wire Lzohu6;  // ../RTL/cortexm0ds_logic.v(156)
  wire Lzoow6;  // ../RTL/cortexm0ds_logic.v(1180)
  wire Lzuiu6;  // ../RTL/cortexm0ds_logic.v(718)
  wire Lzvhu6;  // ../RTL/cortexm0ds_logic.v(250)
  wire Lzvow6;  // ../RTL/cortexm0ds_logic.v(1274)
  wire Lzwax6;  // ../RTL/cortexm0ds_logic.v(1674)
  wire M05ju6;  // ../RTL/cortexm0ds_logic.v(852)
  wire M06iu6;  // ../RTL/cortexm0ds_logic.v(384)
  wire M06pw6;  // ../RTL/cortexm0ds_logic.v(1408)
  wire M07ow6;  // ../RTL/cortexm0ds_logic.v(940)
  wire M0diu6;  // ../RTL/cortexm0ds_logic.v(477)
  wire M0dpw6;  // ../RTL/cortexm0ds_logic.v(1502)
  wire M0eow6;  // ../RTL/cortexm0ds_logic.v(1034)
  wire M0kiu6;  // ../RTL/cortexm0ds_logic.v(571)
  wire M0low6;  // ../RTL/cortexm0ds_logic.v(1127)
  wire M0riu6;  // ../RTL/cortexm0ds_logic.v(665)
  wire M0shu6;  // ../RTL/cortexm0ds_logic.v(197)
  wire M0sow6;  // ../RTL/cortexm0ds_logic.v(1221)
  wire M0yiu6;  // ../RTL/cortexm0ds_logic.v(758)
  wire M0zhu6;  // ../RTL/cortexm0ds_logic.v(290)
  wire M0zow6;  // ../RTL/cortexm0ds_logic.v(1315)
  wire M13bx6;  // ../RTL/cortexm0ds_logic.v(1685)
  wire M14ju6;  // ../RTL/cortexm0ds_logic.v(839)
  wire M15iu6;  // ../RTL/cortexm0ds_logic.v(371)
  wire M15pw6;  // ../RTL/cortexm0ds_logic.v(1395)
  wire M1ciu6;  // ../RTL/cortexm0ds_logic.v(464)
  wire M1cpw6;  // ../RTL/cortexm0ds_logic.v(1489)
  wire M1dow6;  // ../RTL/cortexm0ds_logic.v(1021)
  wire M1ihu6;  // ../RTL/cortexm0ds_logic.v(130)
  wire M1jiu6;  // ../RTL/cortexm0ds_logic.v(558)
  wire M1kow6;  // ../RTL/cortexm0ds_logic.v(1114)
  wire M1qiu6;  // ../RTL/cortexm0ds_logic.v(652)
  wire M1rhu6;  // ../RTL/cortexm0ds_logic.v(184)
  wire M1row6;  // ../RTL/cortexm0ds_logic.v(1208)
  wire M1xiu6;  // ../RTL/cortexm0ds_logic.v(745)
  wire M1yhu6;  // ../RTL/cortexm0ds_logic.v(277)
  wire M1yow6;  // ../RTL/cortexm0ds_logic.v(1302)
  wire M23ju6;  // ../RTL/cortexm0ds_logic.v(826)
  wire M24iu6;  // ../RTL/cortexm0ds_logic.v(358)
  wire M24pw6;  // ../RTL/cortexm0ds_logic.v(1382)
  wire M2aju6;  // ../RTL/cortexm0ds_logic.v(919)
  wire M2biu6;  // ../RTL/cortexm0ds_logic.v(451)
  wire M2bpw6;  // ../RTL/cortexm0ds_logic.v(1476)
  wire M2cow6;  // ../RTL/cortexm0ds_logic.v(1008)
  wire M2ebx6;  // ../RTL/cortexm0ds_logic.v(1705)
  wire M2iiu6;  // ../RTL/cortexm0ds_logic.v(545)
  wire M2jow6;  // ../RTL/cortexm0ds_logic.v(1101)
  wire M2lax6;  // ../RTL/cortexm0ds_logic.v(1652)
  wire M2piu6;  // ../RTL/cortexm0ds_logic.v(639)
  wire M2qhu6;  // ../RTL/cortexm0ds_logic.v(171)
  wire M2qow6;  // ../RTL/cortexm0ds_logic.v(1195)
  wire M2wiu6;  // ../RTL/cortexm0ds_logic.v(732)
  wire M2xhu6;  // ../RTL/cortexm0ds_logic.v(264)
  wire M2xow6;  // ../RTL/cortexm0ds_logic.v(1289)
  wire M32ju6;  // ../RTL/cortexm0ds_logic.v(813)
  wire M33iu6;  // ../RTL/cortexm0ds_logic.v(345)
  wire M33pw6;  // ../RTL/cortexm0ds_logic.v(1369)
  wire M39ju6;  // ../RTL/cortexm0ds_logic.v(906)
  wire M3aiu6;  // ../RTL/cortexm0ds_logic.v(438)
  wire M3apw6;  // ../RTL/cortexm0ds_logic.v(1463)
  wire M3bow6;  // ../RTL/cortexm0ds_logic.v(995)
  wire M3hiu6;  // ../RTL/cortexm0ds_logic.v(532)
  wire M3iow6;  // ../RTL/cortexm0ds_logic.v(1088)
  wire M3oiu6;  // ../RTL/cortexm0ds_logic.v(626)
  wire M3phu6;  // ../RTL/cortexm0ds_logic.v(158)
  wire M3pow6;  // ../RTL/cortexm0ds_logic.v(1182)
  wire M3viu6;  // ../RTL/cortexm0ds_logic.v(719)
  wire M3wax6;  // ../RTL/cortexm0ds_logic.v(1672)
  wire M3whu6;  // ../RTL/cortexm0ds_logic.v(251)
  wire M3wow6;  // ../RTL/cortexm0ds_logic.v(1276)
  wire M41ju6;  // ../RTL/cortexm0ds_logic.v(800)
  wire M42iu6;  // ../RTL/cortexm0ds_logic.v(332)
  wire M42pw6;  // ../RTL/cortexm0ds_logic.v(1356)
  wire M48ju6;  // ../RTL/cortexm0ds_logic.v(893)
  wire M49iu6;  // ../RTL/cortexm0ds_logic.v(425)
  wire M49pw6;  // ../RTL/cortexm0ds_logic.v(1450)
  wire M4aow6;  // ../RTL/cortexm0ds_logic.v(982)
  wire M4ebx6;  // ../RTL/cortexm0ds_logic.v(1705)
  wire M4giu6;  // ../RTL/cortexm0ds_logic.v(519)
  wire M4how6;  // ../RTL/cortexm0ds_logic.v(1075)
  wire M4niu6;  // ../RTL/cortexm0ds_logic.v(613)
  wire M4oow6;  // ../RTL/cortexm0ds_logic.v(1169)
  wire M4uiu6;  // ../RTL/cortexm0ds_logic.v(706)
  wire M4vhu6;  // ../RTL/cortexm0ds_logic.v(238)
  wire M4vow6;  // ../RTL/cortexm0ds_logic.v(1263)
  wire M50ju6;  // ../RTL/cortexm0ds_logic.v(787)
  wire M51iu6;  // ../RTL/cortexm0ds_logic.v(319)
  wire M51pw6;  // ../RTL/cortexm0ds_logic.v(1343)
  wire M57ju6;  // ../RTL/cortexm0ds_logic.v(880)
  wire M58iu6;  // ../RTL/cortexm0ds_logic.v(412)
  wire M58pw6;  // ../RTL/cortexm0ds_logic.v(1437)
  wire M59ow6;  // ../RTL/cortexm0ds_logic.v(969)
  wire M5fiu6;  // ../RTL/cortexm0ds_logic.v(506)
  wire M5gow6;  // ../RTL/cortexm0ds_logic.v(1062)
  wire M5miu6;  // ../RTL/cortexm0ds_logic.v(600)
  wire M5now6;  // ../RTL/cortexm0ds_logic.v(1156)
  wire M5tiu6;  // ../RTL/cortexm0ds_logic.v(693)
  wire M5uhu6;  // ../RTL/cortexm0ds_logic.v(225)
  wire M5uow6;  // ../RTL/cortexm0ds_logic.v(1250)
  wire M5wax6;  // ../RTL/cortexm0ds_logic.v(1672)
  wire M60iu6;  // ../RTL/cortexm0ds_logic.v(306)
  wire M60pw6;  // ../RTL/cortexm0ds_logic.v(1330)
  wire M66ju6;  // ../RTL/cortexm0ds_logic.v(867)
  wire M67iu6;  // ../RTL/cortexm0ds_logic.v(399)
  wire M67pw6;  // ../RTL/cortexm0ds_logic.v(1424)
  wire M68ow6;  // ../RTL/cortexm0ds_logic.v(956)
  wire M6cax6;  // ../RTL/cortexm0ds_logic.v(1635)
  wire M6eiu6;  // ../RTL/cortexm0ds_logic.v(493)
  wire M6fow6;  // ../RTL/cortexm0ds_logic.v(1049)
  wire M6kax6;  // ../RTL/cortexm0ds_logic.v(1651)
  wire M6liu6;  // ../RTL/cortexm0ds_logic.v(587)
  wire M6mow6;  // ../RTL/cortexm0ds_logic.v(1143)
  wire M6rpw6;  // ../RTL/cortexm0ds_logic.v(1601)
  wire M6siu6;  // ../RTL/cortexm0ds_logic.v(680)
  wire M6thu6;  // ../RTL/cortexm0ds_logic.v(212)
  wire M6tow6;  // ../RTL/cortexm0ds_logic.v(1237)
  wire M6ziu6;  // ../RTL/cortexm0ds_logic.v(774)
  wire M75ju6;  // ../RTL/cortexm0ds_logic.v(854)
  wire M76iu6;  // ../RTL/cortexm0ds_logic.v(386)
  wire M76pw6;  // ../RTL/cortexm0ds_logic.v(1411)
  wire M77ow6;  // ../RTL/cortexm0ds_logic.v(943)
  wire M7diu6;  // ../RTL/cortexm0ds_logic.v(480)
  wire M7dpw6;  // ../RTL/cortexm0ds_logic.v(1504)
  wire M7eow6;  // ../RTL/cortexm0ds_logic.v(1036)
  wire M7kiu6;  // ../RTL/cortexm0ds_logic.v(574)
  wire M7low6;  // ../RTL/cortexm0ds_logic.v(1130)
  wire M7riu6;  // ../RTL/cortexm0ds_logic.v(667)
  wire M7shu6;  // ../RTL/cortexm0ds_logic.v(199)
  wire M7sow6;  // ../RTL/cortexm0ds_logic.v(1224)
  wire M7wax6;  // ../RTL/cortexm0ds_logic.v(1673)
  wire M7yiu6;  // ../RTL/cortexm0ds_logic.v(761)
  wire M7zhu6;  // ../RTL/cortexm0ds_logic.v(293)
  wire M7zow6;  // ../RTL/cortexm0ds_logic.v(1317)
  wire M81qw6;  // ../RTL/cortexm0ds_logic.v(1619)
  wire M84ju6;  // ../RTL/cortexm0ds_logic.v(841)
  wire M85bx6;  // ../RTL/cortexm0ds_logic.v(1688)
  wire M85iu6;  // ../RTL/cortexm0ds_logic.v(373)
  wire M85pw6;  // ../RTL/cortexm0ds_logic.v(1398)
  wire M86ow6;  // ../RTL/cortexm0ds_logic.v(930)
  wire M8ciu6;  // ../RTL/cortexm0ds_logic.v(467)
  wire M8cpw6;  // ../RTL/cortexm0ds_logic.v(1491)
  wire M8dow6;  // ../RTL/cortexm0ds_logic.v(1023)
  wire M8fax6;  // ../RTL/cortexm0ds_logic.v(1641)
  wire M8ipw6;  // ../RTL/cortexm0ds_logic.v(1584)
  wire M8jiu6;  // ../RTL/cortexm0ds_logic.v(561)
  wire M8kow6;  // ../RTL/cortexm0ds_logic.v(1117)
  wire M8qiu6;  // ../RTL/cortexm0ds_logic.v(654)
  wire M8rhu6;  // ../RTL/cortexm0ds_logic.v(186)
  wire M8row6;  // ../RTL/cortexm0ds_logic.v(1211)
  wire M8xiu6;  // ../RTL/cortexm0ds_logic.v(748)
  wire M8yhu6;  // ../RTL/cortexm0ds_logic.v(280)
  wire M8yow6;  // ../RTL/cortexm0ds_logic.v(1304)
  wire M93ju6;  // ../RTL/cortexm0ds_logic.v(828)
  wire M94iu6;  // ../RTL/cortexm0ds_logic.v(360)
  wire M94pw6;  // ../RTL/cortexm0ds_logic.v(1385)
  wire M9aju6;  // ../RTL/cortexm0ds_logic.v(922)
  wire M9biu6;  // ../RTL/cortexm0ds_logic.v(454)
  wire M9bpw6;  // ../RTL/cortexm0ds_logic.v(1478)
  wire M9cow6;  // ../RTL/cortexm0ds_logic.v(1010)
  wire M9fhu6;  // ../RTL/cortexm0ds_logic.v(124)
  wire M9iiu6;  // ../RTL/cortexm0ds_logic.v(548)
  wire M9jow6;  // ../RTL/cortexm0ds_logic.v(1104)
  wire M9ohu6;  // ../RTL/cortexm0ds_logic.v(146)
  wire M9piu6;  // ../RTL/cortexm0ds_logic.v(641)
  wire M9qhu6;  // ../RTL/cortexm0ds_logic.v(173)
  wire M9qow6;  // ../RTL/cortexm0ds_logic.v(1198)
  wire M9wax6;  // ../RTL/cortexm0ds_logic.v(1673)
  wire M9wiu6;  // ../RTL/cortexm0ds_logic.v(735)
  wire M9xhu6;  // ../RTL/cortexm0ds_logic.v(267)
  wire M9xow6;  // ../RTL/cortexm0ds_logic.v(1291)
  wire Ma2ju6;  // ../RTL/cortexm0ds_logic.v(815)
  wire Ma3iu6;  // ../RTL/cortexm0ds_logic.v(347)
  wire Ma3pw6;  // ../RTL/cortexm0ds_logic.v(1372)
  wire Ma9ju6;  // ../RTL/cortexm0ds_logic.v(909)
  wire Maaiu6;  // ../RTL/cortexm0ds_logic.v(441)
  wire Maapw6;  // ../RTL/cortexm0ds_logic.v(1465)
  wire Mabow6;  // ../RTL/cortexm0ds_logic.v(997)
  wire Mahiu6;  // ../RTL/cortexm0ds_logic.v(535)
  wire Maiow6;  // ../RTL/cortexm0ds_logic.v(1091)
  wire Maoiu6;  // ../RTL/cortexm0ds_logic.v(628)
  wire Maphu6;  // ../RTL/cortexm0ds_logic.v(160)
  wire Mapow6;  // ../RTL/cortexm0ds_logic.v(1185)
  wire Maviu6;  // ../RTL/cortexm0ds_logic.v(722)
  wire Mawhu6;  // ../RTL/cortexm0ds_logic.v(254)
  wire Mawow6;  // ../RTL/cortexm0ds_logic.v(1278)
  wire Mb1ju6;  // ../RTL/cortexm0ds_logic.v(802)
  wire Mb2iu6;  // ../RTL/cortexm0ds_logic.v(334)
  wire Mb2pw6;  // ../RTL/cortexm0ds_logic.v(1359)
  wire Mb4bx6;  // ../RTL/cortexm0ds_logic.v(1687)
  wire Mb8ju6;  // ../RTL/cortexm0ds_logic.v(896)
  wire Mb9iu6;  // ../RTL/cortexm0ds_logic.v(428)
  wire Mb9pw6;  // ../RTL/cortexm0ds_logic.v(1452)
  wire Mbaow6;  // ../RTL/cortexm0ds_logic.v(984)
  wire Mbdax6;  // ../RTL/cortexm0ds_logic.v(1638)
  wire Mbgiu6;  // ../RTL/cortexm0ds_logic.v(522)
  wire Mbhow6;  // ../RTL/cortexm0ds_logic.v(1078)
  wire Mbniu6;  // ../RTL/cortexm0ds_logic.v(615)
  wire Mboax6;  // ../RTL/cortexm0ds_logic.v(1658)
  wire Mbohu6;  // ../RTL/cortexm0ds_logic.v(147)
  wire Mboow6;  // ../RTL/cortexm0ds_logic.v(1172)
  wire Mbuiu6;  // ../RTL/cortexm0ds_logic.v(709)
  wire Mbvhu6;  // ../RTL/cortexm0ds_logic.v(241)
  wire Mbvow6;  // ../RTL/cortexm0ds_logic.v(1265)
  wire Mbwax6;  // ../RTL/cortexm0ds_logic.v(1673)
  wire Mc0ju6;  // ../RTL/cortexm0ds_logic.v(789)
  wire Mc1iu6;  // ../RTL/cortexm0ds_logic.v(321)
  wire Mc1pw6;  // ../RTL/cortexm0ds_logic.v(1346)
  wire Mc7ju6;  // ../RTL/cortexm0ds_logic.v(883)
  wire Mc8iu6;  // ../RTL/cortexm0ds_logic.v(415)
  wire Mc8pw6;  // ../RTL/cortexm0ds_logic.v(1439)
  wire Mc9ow6;  // ../RTL/cortexm0ds_logic.v(971)
  wire Mcfiu6;  // ../RTL/cortexm0ds_logic.v(509)
  wire Mcgow6;  // ../RTL/cortexm0ds_logic.v(1065)
  wire Mcmiu6;  // ../RTL/cortexm0ds_logic.v(602)
  wire Mcnow6;  // ../RTL/cortexm0ds_logic.v(1159)
  wire Mctiu6;  // ../RTL/cortexm0ds_logic.v(696)
  wire Mcuhu6;  // ../RTL/cortexm0ds_logic.v(228)
  wire Mcuow6;  // ../RTL/cortexm0ds_logic.v(1252)
  wire Md0iu6;  // ../RTL/cortexm0ds_logic.v(308)
  wire Md0pw6;  // ../RTL/cortexm0ds_logic.v(1333)
  wire Md6ju6;  // ../RTL/cortexm0ds_logic.v(870)
  wire Md7iu6;  // ../RTL/cortexm0ds_logic.v(402)
  wire Md7pw6;  // ../RTL/cortexm0ds_logic.v(1426)
  wire Md8ow6;  // ../RTL/cortexm0ds_logic.v(958)
  wire Mdeiu6;  // ../RTL/cortexm0ds_logic.v(496)
  wire Mdfow6;  // ../RTL/cortexm0ds_logic.v(1052)
  wire Mdliu6;  // ../RTL/cortexm0ds_logic.v(589)
  wire Mdmow6;  // ../RTL/cortexm0ds_logic.v(1146)
  wire Mdppw6;  // ../RTL/cortexm0ds_logic.v(1598)
  wire Mdsiu6;  // ../RTL/cortexm0ds_logic.v(683)
  wire Mdthu6;  // ../RTL/cortexm0ds_logic.v(215)
  wire Mdtow6;  // ../RTL/cortexm0ds_logic.v(1239)
  wire Mdziu6;  // ../RTL/cortexm0ds_logic.v(776)
  wire Me5ju6;  // ../RTL/cortexm0ds_logic.v(857)
  wire Me6iu6;  // ../RTL/cortexm0ds_logic.v(389)
  wire Me6pw6;  // ../RTL/cortexm0ds_logic.v(1413)
  wire Me7ow6;  // ../RTL/cortexm0ds_logic.v(945)
  wire Mediu6;  // ../RTL/cortexm0ds_logic.v(483)
  wire Medpw6;  // ../RTL/cortexm0ds_logic.v(1507)
  wire Meeow6;  // ../RTL/cortexm0ds_logic.v(1039)
  wire Mekhu6;  // ../RTL/cortexm0ds_logic.v(136)
  wire Mekiu6;  // ../RTL/cortexm0ds_logic.v(576)
  wire Melow6;  // ../RTL/cortexm0ds_logic.v(1133)
  wire Meriu6;  // ../RTL/cortexm0ds_logic.v(670)
  wire Meshu6;  // ../RTL/cortexm0ds_logic.v(202)
  wire Mesow6;  // ../RTL/cortexm0ds_logic.v(1226)
  wire Meyiu6;  // ../RTL/cortexm0ds_logic.v(763)
  wire Mezhu6;  // ../RTL/cortexm0ds_logic.v(295)
  wire Mezow6;  // ../RTL/cortexm0ds_logic.v(1320)
  wire Mf4ju6;  // ../RTL/cortexm0ds_logic.v(844)
  wire Mf5iu6;  // ../RTL/cortexm0ds_logic.v(376)
  wire Mf5pw6;  // ../RTL/cortexm0ds_logic.v(1400)
  wire Mf6ow6;  // ../RTL/cortexm0ds_logic.v(932)
  wire Mfciu6;  // ../RTL/cortexm0ds_logic.v(470)
  wire Mfcpw6;  // ../RTL/cortexm0ds_logic.v(1494)
  wire Mfdow6;  // ../RTL/cortexm0ds_logic.v(1026)
  wire Mfjiu6;  // ../RTL/cortexm0ds_logic.v(563)
  wire Mfkow6;  // ../RTL/cortexm0ds_logic.v(1120)
  wire Mfqiu6;  // ../RTL/cortexm0ds_logic.v(657)
  wire Mfrhu6;  // ../RTL/cortexm0ds_logic.v(189)
  wire Mfrow6;  // ../RTL/cortexm0ds_logic.v(1213)
  wire Mfxiu6;  // ../RTL/cortexm0ds_logic.v(750)
  wire Mfyax6;  // ../RTL/cortexm0ds_logic.v(1677)
  wire Mfyhu6;  // ../RTL/cortexm0ds_logic.v(282)
  wire Mfyow6;  // ../RTL/cortexm0ds_logic.v(1307)
  wire Mg3ju6;  // ../RTL/cortexm0ds_logic.v(831)
  wire Mg4iu6;  // ../RTL/cortexm0ds_logic.v(363)
  wire Mg4pw6;  // ../RTL/cortexm0ds_logic.v(1387)
  wire Mgaju6;  // ../RTL/cortexm0ds_logic.v(925)
  wire Mgbiu6;  // ../RTL/cortexm0ds_logic.v(457)
  wire Mgbpw6;  // ../RTL/cortexm0ds_logic.v(1481)
  wire Mgcow6;  // ../RTL/cortexm0ds_logic.v(1013)
  wire Mgeax6;  // ../RTL/cortexm0ds_logic.v(1640)
  wire Mgiiu6;  // ../RTL/cortexm0ds_logic.v(550)
  wire Mgjhu6;  // ../RTL/cortexm0ds_logic.v(134)
  wire Mgjow6;  // ../RTL/cortexm0ds_logic.v(1107)
  wire Mgpiu6;  // ../RTL/cortexm0ds_logic.v(644)
  wire Mgqhu6;  // ../RTL/cortexm0ds_logic.v(176)
  wire Mgqow6;  // ../RTL/cortexm0ds_logic.v(1200)
  wire Mgwiu6;  // ../RTL/cortexm0ds_logic.v(737)
  wire Mgxhu6;  // ../RTL/cortexm0ds_logic.v(269)
  wire Mgxow6;  // ../RTL/cortexm0ds_logic.v(1294)
  wire Mh1qw6;  // ../RTL/cortexm0ds_logic.v(1620)
  wire Mh2ju6;  // ../RTL/cortexm0ds_logic.v(818)
  wire Mh3iu6;  // ../RTL/cortexm0ds_logic.v(350)
  wire Mh3pw6;  // ../RTL/cortexm0ds_logic.v(1374)
  wire Mh9ju6;  // ../RTL/cortexm0ds_logic.v(912)
  wire Mhaiu6;  // ../RTL/cortexm0ds_logic.v(444)
  wire Mhapw6;  // ../RTL/cortexm0ds_logic.v(1468)
  wire Mhbow6;  // ../RTL/cortexm0ds_logic.v(1000)
  wire Mhhiu6;  // ../RTL/cortexm0ds_logic.v(537)
  wire Mhiow6;  // ../RTL/cortexm0ds_logic.v(1094)
  wire Mhoiu6;  // ../RTL/cortexm0ds_logic.v(631)
  wire Mhphu6;  // ../RTL/cortexm0ds_logic.v(163)
  wire Mhpow6;  // ../RTL/cortexm0ds_logic.v(1187)
  wire Mhviu6;  // ../RTL/cortexm0ds_logic.v(724)
  wire Mhwhu6;  // ../RTL/cortexm0ds_logic.v(256)
  wire Mhwow6;  // ../RTL/cortexm0ds_logic.v(1281)
  wire Mi1ju6;  // ../RTL/cortexm0ds_logic.v(805)
  wire Mi2iu6;  // ../RTL/cortexm0ds_logic.v(337)
  wire Mi2pw6;  // ../RTL/cortexm0ds_logic.v(1361)
  wire Mi8ju6;  // ../RTL/cortexm0ds_logic.v(899)
  wire Mi9iu6;  // ../RTL/cortexm0ds_logic.v(431)
  wire Mi9pw6;  // ../RTL/cortexm0ds_logic.v(1455)
  wire Miaow6;  // ../RTL/cortexm0ds_logic.v(987)
  wire Migiu6;  // ../RTL/cortexm0ds_logic.v(524)
  wire Mihow6;  // ../RTL/cortexm0ds_logic.v(1081)
  wire Miihu6;  // ../RTL/cortexm0ds_logic.v(131)
  wire Miniu6;  // ../RTL/cortexm0ds_logic.v(618)
  wire Miohu6;  // ../RTL/cortexm0ds_logic.v(150)
  wire Mioow6;  // ../RTL/cortexm0ds_logic.v(1174)
  wire Misax6;  // ../RTL/cortexm0ds_logic.v(1666)
  wire Miuiu6;  // ../RTL/cortexm0ds_logic.v(711)
  wire Mivhu6;  // ../RTL/cortexm0ds_logic.v(243)
  wire Mivow6;  // ../RTL/cortexm0ds_logic.v(1268)
  wire Mj0ju6;  // ../RTL/cortexm0ds_logic.v(792)
  wire Mj1iu6;  // ../RTL/cortexm0ds_logic.v(324)
  wire Mj1pw6;  // ../RTL/cortexm0ds_logic.v(1348)
  wire Mj7ju6;  // ../RTL/cortexm0ds_logic.v(886)
  wire Mj8iu6;  // ../RTL/cortexm0ds_logic.v(418)
  wire Mj8pw6;  // ../RTL/cortexm0ds_logic.v(1442)
  wire Mj9ow6;  // ../RTL/cortexm0ds_logic.v(974)
  wire Mjfiu6;  // ../RTL/cortexm0ds_logic.v(511)
  wire Mjgow6;  // ../RTL/cortexm0ds_logic.v(1068)
  wire Mjmiu6;  // ../RTL/cortexm0ds_logic.v(605)
  wire Mjmpw6;  // ../RTL/cortexm0ds_logic.v(1592)
  wire Mjnow6;  // ../RTL/cortexm0ds_logic.v(1161)
  wire Mjtiu6;  // ../RTL/cortexm0ds_logic.v(698)
  wire Mjuhu6;  // ../RTL/cortexm0ds_logic.v(230)
  wire Mjuow6;  // ../RTL/cortexm0ds_logic.v(1255)
  wire Mk0iu6;  // ../RTL/cortexm0ds_logic.v(311)
  wire Mk0pw6;  // ../RTL/cortexm0ds_logic.v(1335)
  wire Mk3bx6;  // ../RTL/cortexm0ds_logic.v(1685)
  wire Mk6ju6;  // ../RTL/cortexm0ds_logic.v(873)
  wire Mk7iu6;  // ../RTL/cortexm0ds_logic.v(405)
  wire Mk7pw6;  // ../RTL/cortexm0ds_logic.v(1429)
  wire Mk8ow6;  // ../RTL/cortexm0ds_logic.v(961)
  wire Mkeiu6;  // ../RTL/cortexm0ds_logic.v(498)
  wire Mkfow6;  // ../RTL/cortexm0ds_logic.v(1055)
  wire Mkliu6;  // ../RTL/cortexm0ds_logic.v(592)
  wire Mkmow6;  // ../RTL/cortexm0ds_logic.v(1148)
  wire Mksiu6;  // ../RTL/cortexm0ds_logic.v(685)
  wire Mkthu6;  // ../RTL/cortexm0ds_logic.v(217)
  wire Mktow6;  // ../RTL/cortexm0ds_logic.v(1242)
  wire Mkziu6;  // ../RTL/cortexm0ds_logic.v(779)
  wire Ml5ju6;  // ../RTL/cortexm0ds_logic.v(860)
  wire Ml6iu6;  // ../RTL/cortexm0ds_logic.v(392)
  wire Ml6pw6;  // ../RTL/cortexm0ds_logic.v(1416)
  wire Ml7ow6;  // ../RTL/cortexm0ds_logic.v(948)
  wire Mldiu6;  // ../RTL/cortexm0ds_logic.v(485)
  wire Mldpw6;  // ../RTL/cortexm0ds_logic.v(1510)
  wire Mleow6;  // ../RTL/cortexm0ds_logic.v(1042)
  wire Mlkiu6;  // ../RTL/cortexm0ds_logic.v(579)
  wire Mllow6;  // ../RTL/cortexm0ds_logic.v(1135)
  wire Mlmpw6;  // ../RTL/cortexm0ds_logic.v(1593)
  wire Mlriu6;  // ../RTL/cortexm0ds_logic.v(672)
  wire Mlshu6;  // ../RTL/cortexm0ds_logic.v(204)
  wire Mlsow6;  // ../RTL/cortexm0ds_logic.v(1229)
  wire Mlyiu6;  // ../RTL/cortexm0ds_logic.v(766)
  wire Mlzhu6;  // ../RTL/cortexm0ds_logic.v(298)
  wire Mlzow6;  // ../RTL/cortexm0ds_logic.v(1322)
  wire Mm4ju6;  // ../RTL/cortexm0ds_logic.v(847)
  wire Mm5iu6;  // ../RTL/cortexm0ds_logic.v(379)
  wire Mm5pw6;  // ../RTL/cortexm0ds_logic.v(1403)
  wire Mm6ow6;  // ../RTL/cortexm0ds_logic.v(935)
  wire Mmciu6;  // ../RTL/cortexm0ds_logic.v(472)
  wire Mmcpw6;  // ../RTL/cortexm0ds_logic.v(1497)
  wire Mmdow6;  // ../RTL/cortexm0ds_logic.v(1029)
  wire Mmjiu6;  // ../RTL/cortexm0ds_logic.v(566)
  wire Mmkow6;  // ../RTL/cortexm0ds_logic.v(1122)
  wire Mmqiu6;  // ../RTL/cortexm0ds_logic.v(659)
  wire Mmrhu6;  // ../RTL/cortexm0ds_logic.v(191)
  wire Mmrow6;  // ../RTL/cortexm0ds_logic.v(1216)
  wire Mmxiu6;  // ../RTL/cortexm0ds_logic.v(753)
  wire Mmyhu6;  // ../RTL/cortexm0ds_logic.v(285)
  wire Mmyow6;  // ../RTL/cortexm0ds_logic.v(1309)
  wire Mn3ju6;  // ../RTL/cortexm0ds_logic.v(834)
  wire Mn4iu6;  // ../RTL/cortexm0ds_logic.v(366)
  wire Mn4pw6;  // ../RTL/cortexm0ds_logic.v(1390)
  wire Mnaju6;  // ../RTL/cortexm0ds_logic.v(927)
  wire Mnbiu6;  // ../RTL/cortexm0ds_logic.v(459)
  wire Mnbpw6;  // ../RTL/cortexm0ds_logic.v(1484)
  wire Mncow6;  // ../RTL/cortexm0ds_logic.v(1016)
  wire Mniiu6;  // ../RTL/cortexm0ds_logic.v(553)
  wire Mnjow6;  // ../RTL/cortexm0ds_logic.v(1109)
  wire Mnmpw6;  // ../RTL/cortexm0ds_logic.v(1593)
  wire Mnpiu6;  // ../RTL/cortexm0ds_logic.v(646)
  wire Mnqhu6;  // ../RTL/cortexm0ds_logic.v(178)
  wire Mnqow6;  // ../RTL/cortexm0ds_logic.v(1203)
  wire Mnwiu6;  // ../RTL/cortexm0ds_logic.v(740)
  wire Mnxhu6;  // ../RTL/cortexm0ds_logic.v(272)
  wire Mnxow6;  // ../RTL/cortexm0ds_logic.v(1296)
  wire Mo2ju6;  // ../RTL/cortexm0ds_logic.v(821)
  wire Mo3iu6;  // ../RTL/cortexm0ds_logic.v(353)
  wire Mo3pw6;  // ../RTL/cortexm0ds_logic.v(1377)
  wire Mo9ju6;  // ../RTL/cortexm0ds_logic.v(914)
  wire Moaiu6;  // ../RTL/cortexm0ds_logic.v(446)
  wire Moapw6;  // ../RTL/cortexm0ds_logic.v(1471)
  wire Mobow6;  // ../RTL/cortexm0ds_logic.v(1003)
  wire Mohiu6;  // ../RTL/cortexm0ds_logic.v(540)
  wire Moiow6;  // ../RTL/cortexm0ds_logic.v(1096)
  wire Mooiu6;  // ../RTL/cortexm0ds_logic.v(633)
  wire Mophu6;  // ../RTL/cortexm0ds_logic.v(165)
  wire Mopow6;  // ../RTL/cortexm0ds_logic.v(1190)
  wire Moviu6;  // ../RTL/cortexm0ds_logic.v(727)
  wire Mowhu6;  // ../RTL/cortexm0ds_logic.v(259)
  wire Mowow6;  // ../RTL/cortexm0ds_logic.v(1283)
  wire Mp0bx6;  // ../RTL/cortexm0ds_logic.v(1681)
  wire Mp1ju6;  // ../RTL/cortexm0ds_logic.v(808)
  wire Mp2iu6;  // ../RTL/cortexm0ds_logic.v(340)
  wire Mp2pw6;  // ../RTL/cortexm0ds_logic.v(1364)
  wire Mp8ju6;  // ../RTL/cortexm0ds_logic.v(901)
  wire Mp9iu6;  // ../RTL/cortexm0ds_logic.v(433)
  wire Mp9pw6;  // ../RTL/cortexm0ds_logic.v(1458)
  wire Mpaow6;  // ../RTL/cortexm0ds_logic.v(990)
  wire Mpehu6;  // ../RTL/cortexm0ds_logic.v(122)
  wire Mpgiu6;  // ../RTL/cortexm0ds_logic.v(527)
  wire Mphow6;  // ../RTL/cortexm0ds_logic.v(1083)
  wire Mpniu6;  // ../RTL/cortexm0ds_logic.v(620)
  wire Mpohu6;  // ../RTL/cortexm0ds_logic.v(152)
  wire Mpoow6;  // ../RTL/cortexm0ds_logic.v(1177)
  wire Mpuiu6;  // ../RTL/cortexm0ds_logic.v(714)
  wire Mpvhu6;  // ../RTL/cortexm0ds_logic.v(246)
  wire Mpvow6;  // ../RTL/cortexm0ds_logic.v(1270)
  wire Mq0ju6;  // ../RTL/cortexm0ds_logic.v(795)
  wire Mq1iu6;  // ../RTL/cortexm0ds_logic.v(327)
  wire Mq1pw6;  // ../RTL/cortexm0ds_logic.v(1351)
  wire Mq7ju6;  // ../RTL/cortexm0ds_logic.v(888)
  wire Mq8iu6;  // ../RTL/cortexm0ds_logic.v(420)
  wire Mq8pw6;  // ../RTL/cortexm0ds_logic.v(1445)
  wire Mq9ow6;  // ../RTL/cortexm0ds_logic.v(977)
  wire Mqfiu6;  // ../RTL/cortexm0ds_logic.v(514)
  wire Mqgow6;  // ../RTL/cortexm0ds_logic.v(1070)
  wire Mqmiu6;  // ../RTL/cortexm0ds_logic.v(607)
  wire Mqnow6;  // ../RTL/cortexm0ds_logic.v(1164)
  wire Mqtiu6;  // ../RTL/cortexm0ds_logic.v(701)
  wire Mquhu6;  // ../RTL/cortexm0ds_logic.v(233)
  wire Mquow6;  // ../RTL/cortexm0ds_logic.v(1257)
  wire Mr0iu6;  // ../RTL/cortexm0ds_logic.v(314)
  wire Mr0pw6;  // ../RTL/cortexm0ds_logic.v(1338)
  wire Mr6ju6;  // ../RTL/cortexm0ds_logic.v(875)
  wire Mr7iu6;  // ../RTL/cortexm0ds_logic.v(407)
  wire Mr7pw6;  // ../RTL/cortexm0ds_logic.v(1432)
  wire Mr8ow6;  // ../RTL/cortexm0ds_logic.v(964)
  wire Mreiu6;  // ../RTL/cortexm0ds_logic.v(501)
  wire Mrfow6;  // ../RTL/cortexm0ds_logic.v(1057)
  wire Mrliu6;  // ../RTL/cortexm0ds_logic.v(594)
  wire Mrmow6;  // ../RTL/cortexm0ds_logic.v(1151)
  wire Mrsiu6;  // ../RTL/cortexm0ds_logic.v(688)
  wire Mrthu6;  // ../RTL/cortexm0ds_logic.v(220)
  wire Mrtow6;  // ../RTL/cortexm0ds_logic.v(1244)
  wire Mrziu6;  // ../RTL/cortexm0ds_logic.v(782)
  wire Ms5bx6;  // ../RTL/cortexm0ds_logic.v(1689)
  wire Ms5ju6;  // ../RTL/cortexm0ds_logic.v(862)
  wire Ms6iu6;  // ../RTL/cortexm0ds_logic.v(394)
  wire Ms6pw6;  // ../RTL/cortexm0ds_logic.v(1419)
  wire Ms7ow6;  // ../RTL/cortexm0ds_logic.v(951)
  wire Msdiu6;  // ../RTL/cortexm0ds_logic.v(488)
  wire Msdpw6;  // ../RTL/cortexm0ds_logic.v(1512)
  wire Mseow6;  // ../RTL/cortexm0ds_logic.v(1044)
  wire Mskiu6;  // ../RTL/cortexm0ds_logic.v(581)
  wire Mslow6;  // ../RTL/cortexm0ds_logic.v(1138)
  wire Msmhu6;  // ../RTL/cortexm0ds_logic.v(143)
  wire Msriu6;  // ../RTL/cortexm0ds_logic.v(675)
  wire Msshu6;  // ../RTL/cortexm0ds_logic.v(207)
  wire Mssow6;  // ../RTL/cortexm0ds_logic.v(1231)
  wire Msyiu6;  // ../RTL/cortexm0ds_logic.v(769)
  wire Mszhu6;  // ../RTL/cortexm0ds_logic.v(301)
  wire Mszow6;  // ../RTL/cortexm0ds_logic.v(1325)
  wire Mt4ju6;  // ../RTL/cortexm0ds_logic.v(849)
  wire Mt5iu6;  // ../RTL/cortexm0ds_logic.v(381)
  wire Mt5pw6;  // ../RTL/cortexm0ds_logic.v(1406)
  wire Mt6ow6;  // ../RTL/cortexm0ds_logic.v(938)
  wire Mtciu6;  // ../RTL/cortexm0ds_logic.v(475)
  wire Mtcpw6;  // ../RTL/cortexm0ds_logic.v(1499)
  wire Mtdow6;  // ../RTL/cortexm0ds_logic.v(1031)
  wire Mtjiu6;  // ../RTL/cortexm0ds_logic.v(568)
  wire Mtkow6;  // ../RTL/cortexm0ds_logic.v(1125)
  wire Mtqiu6;  // ../RTL/cortexm0ds_logic.v(662)
  wire Mtrhu6;  // ../RTL/cortexm0ds_logic.v(194)
  wire Mtrow6;  // ../RTL/cortexm0ds_logic.v(1218)
  wire Mtxiu6;  // ../RTL/cortexm0ds_logic.v(756)
  wire Mtyhu6;  // ../RTL/cortexm0ds_logic.v(288)
  wire Mtyow6;  // ../RTL/cortexm0ds_logic.v(1312)
  wire Mu3ju6;  // ../RTL/cortexm0ds_logic.v(836)
  wire Mu4iu6;  // ../RTL/cortexm0ds_logic.v(368)
  wire Mu4pw6;  // ../RTL/cortexm0ds_logic.v(1393)
  wire Mubiu6;  // ../RTL/cortexm0ds_logic.v(462)
  wire Mubpw6;  // ../RTL/cortexm0ds_logic.v(1486)
  wire Mucow6;  // ../RTL/cortexm0ds_logic.v(1018)
  wire Muhbx6;  // ../RTL/cortexm0ds_logic.v(1712)
  wire Muiiu6;  // ../RTL/cortexm0ds_logic.v(555)
  wire Mujow6;  // ../RTL/cortexm0ds_logic.v(1112)
  wire Mupiu6;  // ../RTL/cortexm0ds_logic.v(649)
  wire Muqhu6;  // ../RTL/cortexm0ds_logic.v(181)
  wire Muqow6;  // ../RTL/cortexm0ds_logic.v(1205)
  wire Muwiu6;  // ../RTL/cortexm0ds_logic.v(743)
  wire Muxhu6;  // ../RTL/cortexm0ds_logic.v(275)
  wire Muxow6;  // ../RTL/cortexm0ds_logic.v(1299)
  wire Mv2ju6;  // ../RTL/cortexm0ds_logic.v(823)
  wire Mv3iu6;  // ../RTL/cortexm0ds_logic.v(355)
  wire Mv3pw6;  // ../RTL/cortexm0ds_logic.v(1380)
  wire Mv9ju6;  // ../RTL/cortexm0ds_logic.v(917)
  wire Mvaiu6;  // ../RTL/cortexm0ds_logic.v(449)
  wire Mvapw6;  // ../RTL/cortexm0ds_logic.v(1473)
  wire Mvbow6;  // ../RTL/cortexm0ds_logic.v(1005)
  wire Mvhiu6;  // ../RTL/cortexm0ds_logic.v(542)
  wire Mviow6;  // ../RTL/cortexm0ds_logic.v(1099)
  wire Mvkhu6;  // ../RTL/cortexm0ds_logic.v(138)
  wire Mvlhu6;  // ../RTL/cortexm0ds_logic.v(140)
  wire Mvoiu6;  // ../RTL/cortexm0ds_logic.v(636)
  wire Mvphu6;  // ../RTL/cortexm0ds_logic.v(168)
  wire Mvpow6;  // ../RTL/cortexm0ds_logic.v(1192)
  wire Mvviu6;  // ../RTL/cortexm0ds_logic.v(730)
  wire Mvwhu6;  // ../RTL/cortexm0ds_logic.v(262)
  wire Mvwow6;  // ../RTL/cortexm0ds_logic.v(1286)
  wire Mw1ju6;  // ../RTL/cortexm0ds_logic.v(810)
  wire Mw2iu6;  // ../RTL/cortexm0ds_logic.v(342)
  wire Mw2pw6;  // ../RTL/cortexm0ds_logic.v(1367)
  wire Mw5bx6;  // ../RTL/cortexm0ds_logic.v(1690)
  wire Mw8ju6;  // ../RTL/cortexm0ds_logic.v(904)
  wire Mw9iu6;  // ../RTL/cortexm0ds_logic.v(436)
  wire Mw9pw6;  // ../RTL/cortexm0ds_logic.v(1460)
  wire Mwaow6;  // ../RTL/cortexm0ds_logic.v(992)
  wire Mwgiu6;  // ../RTL/cortexm0ds_logic.v(529)
  wire Mwhow6;  // ../RTL/cortexm0ds_logic.v(1086)
  wire Mwniu6;  // ../RTL/cortexm0ds_logic.v(623)
  wire Mwohu6;  // ../RTL/cortexm0ds_logic.v(155)
  wire Mwoow6;  // ../RTL/cortexm0ds_logic.v(1179)
  wire Mwuiu6;  // ../RTL/cortexm0ds_logic.v(717)
  wire Mwvhu6;  // ../RTL/cortexm0ds_logic.v(249)
  wire Mwvow6;  // ../RTL/cortexm0ds_logic.v(1273)
  wire Mx0ju6;  // ../RTL/cortexm0ds_logic.v(797)
  wire Mx1iu6;  // ../RTL/cortexm0ds_logic.v(329)
  wire Mx1pw6;  // ../RTL/cortexm0ds_logic.v(1354)
  wire Mx7ju6;  // ../RTL/cortexm0ds_logic.v(891)
  wire Mx8iu6;  // ../RTL/cortexm0ds_logic.v(423)
  wire Mx8pw6;  // ../RTL/cortexm0ds_logic.v(1447)
  wire Mx9ow6;  // ../RTL/cortexm0ds_logic.v(979)
  wire Mxfiu6;  // ../RTL/cortexm0ds_logic.v(516)
  wire Mxgow6;  // ../RTL/cortexm0ds_logic.v(1073)
  wire Mxjhu6;  // ../RTL/cortexm0ds_logic.v(135)
  wire Mxmiu6;  // ../RTL/cortexm0ds_logic.v(610)
  wire Mxnow6;  // ../RTL/cortexm0ds_logic.v(1166)
  wire Mxtiu6;  // ../RTL/cortexm0ds_logic.v(704)
  wire Mxuhu6;  // ../RTL/cortexm0ds_logic.v(236)
  wire Mxuow6;  // ../RTL/cortexm0ds_logic.v(1260)
  wire My0iu6;  // ../RTL/cortexm0ds_logic.v(316)
  wire My0pw6;  // ../RTL/cortexm0ds_logic.v(1341)
  wire My6ju6;  // ../RTL/cortexm0ds_logic.v(878)
  wire My7iu6;  // ../RTL/cortexm0ds_logic.v(410)
  wire My7pw6;  // ../RTL/cortexm0ds_logic.v(1434)
  wire My8ow6;  // ../RTL/cortexm0ds_logic.v(966)
  wire Myeiu6;  // ../RTL/cortexm0ds_logic.v(503)
  wire Myfow6;  // ../RTL/cortexm0ds_logic.v(1060)
  wire Myliu6;  // ../RTL/cortexm0ds_logic.v(597)
  wire Mymow6;  // ../RTL/cortexm0ds_logic.v(1153)
  wire Mysiu6;  // ../RTL/cortexm0ds_logic.v(691)
  wire Mythu6;  // ../RTL/cortexm0ds_logic.v(223)
  wire Mytow6;  // ../RTL/cortexm0ds_logic.v(1247)
  wire Myziu6;  // ../RTL/cortexm0ds_logic.v(784)
  wire Mz1bx6;  // ../RTL/cortexm0ds_logic.v(1683)
  wire Mz5ju6;  // ../RTL/cortexm0ds_logic.v(865)
  wire Mz6iu6;  // ../RTL/cortexm0ds_logic.v(397)
  wire Mz6pw6;  // ../RTL/cortexm0ds_logic.v(1421)
  wire Mz7ow6;  // ../RTL/cortexm0ds_logic.v(953)
  wire Mzdiu6;  // ../RTL/cortexm0ds_logic.v(490)
  wire Mzdpw6;  // ../RTL/cortexm0ds_logic.v(1515)
  wire Mzeow6;  // ../RTL/cortexm0ds_logic.v(1047)
  wire Mzihu6;  // ../RTL/cortexm0ds_logic.v(132)
  wire Mzkiu6;  // ../RTL/cortexm0ds_logic.v(584)
  wire Mzlow6;  // ../RTL/cortexm0ds_logic.v(1140)
  wire Mzriu6;  // ../RTL/cortexm0ds_logic.v(678)
  wire Mzshu6;  // ../RTL/cortexm0ds_logic.v(210)
  wire Mzsow6;  // ../RTL/cortexm0ds_logic.v(1234)
  wire Mzyiu6;  // ../RTL/cortexm0ds_logic.v(771)
  wire Mzzhu6;  // ../RTL/cortexm0ds_logic.v(303)
  wire Mzzow6;  // ../RTL/cortexm0ds_logic.v(1328)
  wire N02ju6;  // ../RTL/cortexm0ds_logic.v(812)
  wire N03iu6;  // ../RTL/cortexm0ds_logic.v(344)
  wire N03pw6;  // ../RTL/cortexm0ds_logic.v(1368)
  wire N09ju6;  // ../RTL/cortexm0ds_logic.v(905)
  wire N0aiu6;  // ../RTL/cortexm0ds_logic.v(437)
  wire N0apw6;  // ../RTL/cortexm0ds_logic.v(1462)
  wire N0bow6;  // ../RTL/cortexm0ds_logic.v(994)
  wire N0cbx6;  // ../RTL/cortexm0ds_logic.v(1701)
  wire N0hiu6;  // ../RTL/cortexm0ds_logic.v(531)
  wire N0iow6;  // ../RTL/cortexm0ds_logic.v(1087)
  wire N0lax6;  // ../RTL/cortexm0ds_logic.v(1652)
  wire N0oiu6;  // ../RTL/cortexm0ds_logic.v(624)
  wire N0phu6;  // ../RTL/cortexm0ds_logic.v(156)
  wire N0pow6;  // ../RTL/cortexm0ds_logic.v(1181)
  wire N0viu6;  // ../RTL/cortexm0ds_logic.v(718)
  wire N0whu6;  // ../RTL/cortexm0ds_logic.v(250)
  wire N0wow6;  // ../RTL/cortexm0ds_logic.v(1274)
  wire N0xpw6;  // ../RTL/cortexm0ds_logic.v(1611)
  wire N11ju6;  // ../RTL/cortexm0ds_logic.v(799)
  wire N12iu6;  // ../RTL/cortexm0ds_logic.v(331)
  wire N12pw6;  // ../RTL/cortexm0ds_logic.v(1355)
  wire N18ju6;  // ../RTL/cortexm0ds_logic.v(892)
  wire N19bx6;  // ../RTL/cortexm0ds_logic.v(1695)
  wire N19iu6;  // ../RTL/cortexm0ds_logic.v(424)
  wire N19pw6;  // ../RTL/cortexm0ds_logic.v(1449)
  wire N1aow6;  // ../RTL/cortexm0ds_logic.v(981)
  wire N1giu6;  // ../RTL/cortexm0ds_logic.v(518)
  wire N1how6;  // ../RTL/cortexm0ds_logic.v(1074)
  wire N1niu6;  // ../RTL/cortexm0ds_logic.v(611)
  wire N1oax6;  // ../RTL/cortexm0ds_logic.v(1658)
  wire N1oow6;  // ../RTL/cortexm0ds_logic.v(1168)
  wire N1uiu6;  // ../RTL/cortexm0ds_logic.v(705)
  wire N1vhu6;  // ../RTL/cortexm0ds_logic.v(237)
  wire N1vow6;  // ../RTL/cortexm0ds_logic.v(1261)
  wire N1wax6;  // ../RTL/cortexm0ds_logic.v(1672)
  wire N20ju6;  // ../RTL/cortexm0ds_logic.v(786)
  wire N21iu6;  // ../RTL/cortexm0ds_logic.v(318)
  wire N21pw6;  // ../RTL/cortexm0ds_logic.v(1342)
  wire N27ju6;  // ../RTL/cortexm0ds_logic.v(879)
  wire N28iu6;  // ../RTL/cortexm0ds_logic.v(411)
  wire N28pw6;  // ../RTL/cortexm0ds_logic.v(1436)
  wire N29ow6;  // ../RTL/cortexm0ds_logic.v(968)
  wire N2fiu6;  // ../RTL/cortexm0ds_logic.v(505)
  wire N2ghu6;  // ../RTL/cortexm0ds_logic.v(125)
  wire N2gow6;  // ../RTL/cortexm0ds_logic.v(1061)
  wire N2miu6;  // ../RTL/cortexm0ds_logic.v(598)
  wire N2now6;  // ../RTL/cortexm0ds_logic.v(1155)
  wire N2tiu6;  // ../RTL/cortexm0ds_logic.v(692)
  wire N2uhu6;  // ../RTL/cortexm0ds_logic.v(224)
  wire N2uow6;  // ../RTL/cortexm0ds_logic.v(1248)
  wire N30iu6;  // ../RTL/cortexm0ds_logic.v(305)
  wire N30pw6;  // ../RTL/cortexm0ds_logic.v(1329)
  wire N36ju6;  // ../RTL/cortexm0ds_logic.v(866)
  wire N37iu6;  // ../RTL/cortexm0ds_logic.v(398)
  wire N37pw6;  // ../RTL/cortexm0ds_logic.v(1423)
  wire N38ow6;  // ../RTL/cortexm0ds_logic.v(955)
  wire N39ax6;  // ../RTL/cortexm0ds_logic.v(1629)
  wire N3eax6;  // ../RTL/cortexm0ds_logic.v(1639)
  wire N3eiu6;  // ../RTL/cortexm0ds_logic.v(492)
  wire N3epw6;  // ../RTL/cortexm0ds_logic.v(1516)
  wire N3fow6;  // ../RTL/cortexm0ds_logic.v(1048)
  wire N3hbx6;  // ../RTL/cortexm0ds_logic.v(1710)
  wire N3jbx6;  // ../RTL/cortexm0ds_logic.v(1714)
  wire N3liu6;  // ../RTL/cortexm0ds_logic.v(585)
  wire N3mow6;  // ../RTL/cortexm0ds_logic.v(1142)
  wire N3nhu6;  // ../RTL/cortexm0ds_logic.v(144)
  wire N3oax6;  // ../RTL/cortexm0ds_logic.v(1658)
  wire N3siu6;  // ../RTL/cortexm0ds_logic.v(679)
  wire N3thu6;  // ../RTL/cortexm0ds_logic.v(211)
  wire N3tow6;  // ../RTL/cortexm0ds_logic.v(1235)
  wire N3ziu6;  // ../RTL/cortexm0ds_logic.v(773)
  wire N45ju6;  // ../RTL/cortexm0ds_logic.v(853)
  wire N46iu6;  // ../RTL/cortexm0ds_logic.v(385)
  wire N46pw6;  // ../RTL/cortexm0ds_logic.v(1410)
  wire N47ow6;  // ../RTL/cortexm0ds_logic.v(942)
  wire N4diu6;  // ../RTL/cortexm0ds_logic.v(479)
  wire N4dpw6;  // ../RTL/cortexm0ds_logic.v(1503)
  wire N4eow6;  // ../RTL/cortexm0ds_logic.v(1035)
  wire N4gax6;  // ../RTL/cortexm0ds_logic.v(1643)
  wire N4kax6;  // ../RTL/cortexm0ds_logic.v(1651)
  wire N4kiu6;  // ../RTL/cortexm0ds_logic.v(572)
  wire N4low6;  // ../RTL/cortexm0ds_logic.v(1129)
  wire N4riu6;  // ../RTL/cortexm0ds_logic.v(666)
  wire N4shu6;  // ../RTL/cortexm0ds_logic.v(198)
  wire N4sow6;  // ../RTL/cortexm0ds_logic.v(1222)
  wire N4yiu6;  // ../RTL/cortexm0ds_logic.v(760)
  wire N4zhu6;  // ../RTL/cortexm0ds_logic.v(292)
  wire N4zow6;  // ../RTL/cortexm0ds_logic.v(1316)
  wire N54ju6;  // ../RTL/cortexm0ds_logic.v(840)
  wire N55iu6;  // ../RTL/cortexm0ds_logic.v(372)
  wire N55pw6;  // ../RTL/cortexm0ds_logic.v(1397)
  wire N5bbx6;  // ../RTL/cortexm0ds_logic.v(1699)
  wire N5ciu6;  // ../RTL/cortexm0ds_logic.v(466)
  wire N5cpw6;  // ../RTL/cortexm0ds_logic.v(1490)
  wire N5dow6;  // ../RTL/cortexm0ds_logic.v(1022)
  wire N5jiu6;  // ../RTL/cortexm0ds_logic.v(559)
  wire N5kow6;  // ../RTL/cortexm0ds_logic.v(1116)
  wire N5oax6;  // ../RTL/cortexm0ds_logic.v(1658)
  wire N5qiu6;  // ../RTL/cortexm0ds_logic.v(653)
  wire N5rhu6;  // ../RTL/cortexm0ds_logic.v(185)
  wire N5row6;  // ../RTL/cortexm0ds_logic.v(1209)
  wire N5xiu6;  // ../RTL/cortexm0ds_logic.v(747)
  wire N5yhu6;  // ../RTL/cortexm0ds_logic.v(279)
  wire N5yow6;  // ../RTL/cortexm0ds_logic.v(1303)
  wire N61qw6;  // ../RTL/cortexm0ds_logic.v(1619)
  wire N63ju6;  // ../RTL/cortexm0ds_logic.v(827)
  wire N64iu6;  // ../RTL/cortexm0ds_logic.v(359)
  wire N64pw6;  // ../RTL/cortexm0ds_logic.v(1384)
  wire N6aju6;  // ../RTL/cortexm0ds_logic.v(921)
  wire N6biu6;  // ../RTL/cortexm0ds_logic.v(453)
  wire N6bpw6;  // ../RTL/cortexm0ds_logic.v(1477)
  wire N6cow6;  // ../RTL/cortexm0ds_logic.v(1009)
  wire N6iiu6;  // ../RTL/cortexm0ds_logic.v(546)
  wire N6jow6;  // ../RTL/cortexm0ds_logic.v(1103)
  wire N6piu6;  // ../RTL/cortexm0ds_logic.v(640)
  wire N6qhu6;  // ../RTL/cortexm0ds_logic.v(172)
  wire N6qow6;  // ../RTL/cortexm0ds_logic.v(1196)
  wire N6wiu6;  // ../RTL/cortexm0ds_logic.v(734)
  wire N6xhu6;  // ../RTL/cortexm0ds_logic.v(266)
  wire N6xow6;  // ../RTL/cortexm0ds_logic.v(1290)
  wire N72ju6;  // ../RTL/cortexm0ds_logic.v(814)
  wire N73iu6;  // ../RTL/cortexm0ds_logic.v(346)
  wire N73pw6;  // ../RTL/cortexm0ds_logic.v(1371)
  wire N79ju6;  // ../RTL/cortexm0ds_logic.v(908)
  wire N7aiu6;  // ../RTL/cortexm0ds_logic.v(440)
  wire N7apw6;  // ../RTL/cortexm0ds_logic.v(1464)
  wire N7bow6;  // ../RTL/cortexm0ds_logic.v(996)
  wire N7hiu6;  // ../RTL/cortexm0ds_logic.v(533)
  wire N7iow6;  // ../RTL/cortexm0ds_logic.v(1090)
  wire N7oax6;  // ../RTL/cortexm0ds_logic.v(1658)
  wire N7oiu6;  // ../RTL/cortexm0ds_logic.v(627)
  wire N7phu6;  // ../RTL/cortexm0ds_logic.v(159)
  wire N7pow6;  // ../RTL/cortexm0ds_logic.v(1183)
  wire N7ppw6;  // ../RTL/cortexm0ds_logic.v(1597)
  wire N7viu6;  // ../RTL/cortexm0ds_logic.v(721)
  wire N7whu6;  // ../RTL/cortexm0ds_logic.v(253)
  wire N7wow6;  // ../RTL/cortexm0ds_logic.v(1277)
  wire N81ju6;  // ../RTL/cortexm0ds_logic.v(801)
  wire N82iu6;  // ../RTL/cortexm0ds_logic.v(333)
  wire N82pw6;  // ../RTL/cortexm0ds_logic.v(1358)
  wire N88ju6;  // ../RTL/cortexm0ds_logic.v(895)
  wire N89iu6;  // ../RTL/cortexm0ds_logic.v(427)
  wire N89pw6;  // ../RTL/cortexm0ds_logic.v(1451)
  wire N8aow6;  // ../RTL/cortexm0ds_logic.v(983)
  wire N8giu6;  // ../RTL/cortexm0ds_logic.v(520)
  wire N8how6;  // ../RTL/cortexm0ds_logic.v(1077)
  wire N8niu6;  // ../RTL/cortexm0ds_logic.v(614)
  wire N8oow6;  // ../RTL/cortexm0ds_logic.v(1170)
  wire N8rpw6;  // ../RTL/cortexm0ds_logic.v(1601)
  wire N8uiu6;  // ../RTL/cortexm0ds_logic.v(708)
  wire N8vhu6;  // ../RTL/cortexm0ds_logic.v(240)
  wire N8vow6;  // ../RTL/cortexm0ds_logic.v(1264)
  wire N90ju6;  // ../RTL/cortexm0ds_logic.v(788)
  wire N91iu6;  // ../RTL/cortexm0ds_logic.v(320)
  wire N91pw6;  // ../RTL/cortexm0ds_logic.v(1345)
  wire N97ju6;  // ../RTL/cortexm0ds_logic.v(882)
  wire N98iu6;  // ../RTL/cortexm0ds_logic.v(414)
  wire N98pw6;  // ../RTL/cortexm0ds_logic.v(1438)
  wire N99ow6;  // ../RTL/cortexm0ds_logic.v(970)
  wire N9fiu6;  // ../RTL/cortexm0ds_logic.v(507)
  wire N9gow6;  // ../RTL/cortexm0ds_logic.v(1064)
  wire N9miu6;  // ../RTL/cortexm0ds_logic.v(601)
  wire N9now6;  // ../RTL/cortexm0ds_logic.v(1157)
  wire N9oax6;  // ../RTL/cortexm0ds_logic.v(1658)
  wire N9ppw6;  // ../RTL/cortexm0ds_logic.v(1597)
  wire N9tiu6;  // ../RTL/cortexm0ds_logic.v(695)
  wire N9uhu6;  // ../RTL/cortexm0ds_logic.v(227)
  wire N9uow6;  // ../RTL/cortexm0ds_logic.v(1251)
  wire Na0iu6;  // ../RTL/cortexm0ds_logic.v(307)
  wire Na0pw6;  // ../RTL/cortexm0ds_logic.v(1332)
  wire Na6ju6;  // ../RTL/cortexm0ds_logic.v(869)
  wire Na7iu6;  // ../RTL/cortexm0ds_logic.v(401)
  wire Na7pw6;  // ../RTL/cortexm0ds_logic.v(1425)
  wire Na8ow6;  // ../RTL/cortexm0ds_logic.v(957)
  wire Naaax6;  // ../RTL/cortexm0ds_logic.v(1632)
  wire Naeiu6;  // ../RTL/cortexm0ds_logic.v(494)
  wire Nafow6;  // ../RTL/cortexm0ds_logic.v(1051)
  wire Naliu6;  // ../RTL/cortexm0ds_logic.v(588)
  wire Namow6;  // ../RTL/cortexm0ds_logic.v(1144)
  wire Nasiu6;  // ../RTL/cortexm0ds_logic.v(682)
  wire Nathu6;  // ../RTL/cortexm0ds_logic.v(214)
  wire Natow6;  // ../RTL/cortexm0ds_logic.v(1238)
  wire Nazax6;  // ../RTL/cortexm0ds_logic.v(1678)
  wire Naziu6;  // ../RTL/cortexm0ds_logic.v(775)
  wire Nb5ju6;  // ../RTL/cortexm0ds_logic.v(856)
  wire Nb6iu6;  // ../RTL/cortexm0ds_logic.v(388)
  wire Nb6pw6;  // ../RTL/cortexm0ds_logic.v(1412)
  wire Nb7ow6;  // ../RTL/cortexm0ds_logic.v(944)
  wire Nbdiu6;  // ../RTL/cortexm0ds_logic.v(481)
  wire Nbdpw6;  // ../RTL/cortexm0ds_logic.v(1506)
  wire Nbeow6;  // ../RTL/cortexm0ds_logic.v(1038)
  wire Nbkiu6;  // ../RTL/cortexm0ds_logic.v(575)
  wire Nblow6;  // ../RTL/cortexm0ds_logic.v(1131)
  wire Nbppw6;  // ../RTL/cortexm0ds_logic.v(1598)
  wire Nbriu6;  // ../RTL/cortexm0ds_logic.v(669)
  wire Nbshu6;  // ../RTL/cortexm0ds_logic.v(201)
  wire Nbsow6;  // ../RTL/cortexm0ds_logic.v(1225)
  wire Nbxax6;  // ../RTL/cortexm0ds_logic.v(1675)
  wire Nbyiu6;  // ../RTL/cortexm0ds_logic.v(762)
  wire Nbzhu6;  // ../RTL/cortexm0ds_logic.v(294)
  wire Nbzow6;  // ../RTL/cortexm0ds_logic.v(1319)
  wire Nc4ju6;  // ../RTL/cortexm0ds_logic.v(843)
  wire Nc5iu6;  // ../RTL/cortexm0ds_logic.v(375)
  wire Nc5pw6;  // ../RTL/cortexm0ds_logic.v(1399)
  wire Nc6ow6;  // ../RTL/cortexm0ds_logic.v(931)
  wire Ncciu6;  // ../RTL/cortexm0ds_logic.v(468)
  wire Nccpw6;  // ../RTL/cortexm0ds_logic.v(1493)
  wire Ncdow6;  // ../RTL/cortexm0ds_logic.v(1025)
  wire Ncjiu6;  // ../RTL/cortexm0ds_logic.v(562)
  wire Nckbx6;  // ../RTL/cortexm0ds_logic.v(1716)
  wire Nckow6;  // ../RTL/cortexm0ds_logic.v(1118)
  wire Ncqiu6;  // ../RTL/cortexm0ds_logic.v(656)
  wire Ncrhu6;  // ../RTL/cortexm0ds_logic.v(188)
  wire Ncrow6;  // ../RTL/cortexm0ds_logic.v(1212)
  wire Ncxiu6;  // ../RTL/cortexm0ds_logic.v(749)
  wire Ncyhu6;  // ../RTL/cortexm0ds_logic.v(281)
  wire Ncyow6;  // ../RTL/cortexm0ds_logic.v(1306)
  wire Nd3ju6;  // ../RTL/cortexm0ds_logic.v(830)
  wire Nd3qw6;  // ../RTL/cortexm0ds_logic.v(1623)
  wire Nd4iu6;  // ../RTL/cortexm0ds_logic.v(362)
  wire Nd4pw6;  // ../RTL/cortexm0ds_logic.v(1386)
  wire Ndaju6;  // ../RTL/cortexm0ds_logic.v(923)
  wire Ndbiu6;  // ../RTL/cortexm0ds_logic.v(455)
  wire Ndbpw6;  // ../RTL/cortexm0ds_logic.v(1480)
  wire Ndcow6;  // ../RTL/cortexm0ds_logic.v(1012)
  wire Ndghu6;  // ../RTL/cortexm0ds_logic.v(126)
  wire Ndiiu6;  // ../RTL/cortexm0ds_logic.v(549)
  wire Ndjow6;  // ../RTL/cortexm0ds_logic.v(1105)
  wire Ndpiu6;  // ../RTL/cortexm0ds_logic.v(643)
  wire Ndqhu6;  // ../RTL/cortexm0ds_logic.v(175)
  wire Ndqow6;  // ../RTL/cortexm0ds_logic.v(1199)
  wire Ndwiu6;  // ../RTL/cortexm0ds_logic.v(736)
  wire Ndxhu6;  // ../RTL/cortexm0ds_logic.v(268)
  wire Ndxow6;  // ../RTL/cortexm0ds_logic.v(1293)
  wire Ne2ju6;  // ../RTL/cortexm0ds_logic.v(817)
  wire Ne3iu6;  // ../RTL/cortexm0ds_logic.v(349)
  wire Ne3pw6;  // ../RTL/cortexm0ds_logic.v(1373)
  wire Ne9ju6;  // ../RTL/cortexm0ds_logic.v(910)
  wire Neaiu6;  // ../RTL/cortexm0ds_logic.v(442)
  wire Neapw6;  // ../RTL/cortexm0ds_logic.v(1467)
  wire Nebow6;  // ../RTL/cortexm0ds_logic.v(999)
  wire Nehiu6;  // ../RTL/cortexm0ds_logic.v(536)
  wire Neiow6;  // ../RTL/cortexm0ds_logic.v(1092)
  wire Nemhu6;  // ../RTL/cortexm0ds_logic.v(142)
  wire Neoiu6;  // ../RTL/cortexm0ds_logic.v(630)
  wire Nephu6;  // ../RTL/cortexm0ds_logic.v(162)
  wire Nepow6;  // ../RTL/cortexm0ds_logic.v(1186)
  wire Neviu6;  // ../RTL/cortexm0ds_logic.v(723)
  wire Newhu6;  // ../RTL/cortexm0ds_logic.v(255)
  wire Newow6;  // ../RTL/cortexm0ds_logic.v(1280)
  wire Nf1ju6;  // ../RTL/cortexm0ds_logic.v(804)
  wire Nf2iu6;  // ../RTL/cortexm0ds_logic.v(336)
  wire Nf2pw6;  // ../RTL/cortexm0ds_logic.v(1360)
  wire Nf8ju6;  // ../RTL/cortexm0ds_logic.v(897)
  wire Nf9iu6;  // ../RTL/cortexm0ds_logic.v(429)
  wire Nf9pw6;  // ../RTL/cortexm0ds_logic.v(1454)
  wire Nfaow6;  // ../RTL/cortexm0ds_logic.v(986)
  wire Nfgax6;  // ../RTL/cortexm0ds_logic.v(1644)
  wire Nfgiu6;  // ../RTL/cortexm0ds_logic.v(523)
  wire Nfhow6;  // ../RTL/cortexm0ds_logic.v(1079)
  wire Nfnax6;  // ../RTL/cortexm0ds_logic.v(1657)
  wire Nfniu6;  // ../RTL/cortexm0ds_logic.v(617)
  wire Nfohu6;  // ../RTL/cortexm0ds_logic.v(149)
  wire Nfoow6;  // ../RTL/cortexm0ds_logic.v(1173)
  wire Nfqpw6;  // ../RTL/cortexm0ds_logic.v(1600)
  wire Nfuiu6;  // ../RTL/cortexm0ds_logic.v(710)
  wire Nfvhu6;  // ../RTL/cortexm0ds_logic.v(242)
  wire Nfvow6;  // ../RTL/cortexm0ds_logic.v(1267)
  wire Ng0ju6;  // ../RTL/cortexm0ds_logic.v(791)
  wire Ng1iu6;  // ../RTL/cortexm0ds_logic.v(323)
  wire Ng1pw6;  // ../RTL/cortexm0ds_logic.v(1347)
  wire Ng7ju6;  // ../RTL/cortexm0ds_logic.v(884)
  wire Ng8iu6;  // ../RTL/cortexm0ds_logic.v(416)
  wire Ng8pw6;  // ../RTL/cortexm0ds_logic.v(1441)
  wire Ng9ow6;  // ../RTL/cortexm0ds_logic.v(973)
  wire Ngfiu6;  // ../RTL/cortexm0ds_logic.v(510)
  wire Nggow6;  // ../RTL/cortexm0ds_logic.v(1066)
  wire Ngmiu6;  // ../RTL/cortexm0ds_logic.v(604)
  wire Ngnow6;  // ../RTL/cortexm0ds_logic.v(1160)
  wire Ngsax6;  // ../RTL/cortexm0ds_logic.v(1666)
  wire Ngtiu6;  // ../RTL/cortexm0ds_logic.v(697)
  wire Nguhu6;  // ../RTL/cortexm0ds_logic.v(229)
  wire Nguow6;  // ../RTL/cortexm0ds_logic.v(1254)
  wire Nh0iu6;  // ../RTL/cortexm0ds_logic.v(310)
  wire Nh0pw6;  // ../RTL/cortexm0ds_logic.v(1334)
  wire Nh6ju6;  // ../RTL/cortexm0ds_logic.v(871)
  wire Nh7iu6;  // ../RTL/cortexm0ds_logic.v(403)
  wire Nh7pw6;  // ../RTL/cortexm0ds_logic.v(1428)
  wire Nh8ow6;  // ../RTL/cortexm0ds_logic.v(960)
  wire Nheiu6;  // ../RTL/cortexm0ds_logic.v(497)
  wire Nhfow6;  // ../RTL/cortexm0ds_logic.v(1053)
  wire Nhgbx6;  // ../RTL/cortexm0ds_logic.v(1709)
  wire Nhlhu6;  // ../RTL/cortexm0ds_logic.v(139)
  wire Nhliu6;  // ../RTL/cortexm0ds_logic.v(591)
  wire Nhmow6;  // ../RTL/cortexm0ds_logic.v(1147)
  wire Nhnax6;  // ../RTL/cortexm0ds_logic.v(1657)
  wire Nhsiu6;  // ../RTL/cortexm0ds_logic.v(684)
  wire Nhthu6;  // ../RTL/cortexm0ds_logic.v(216)
  wire Nhtow6;  // ../RTL/cortexm0ds_logic.v(1241)
  wire Nhziu6;  // ../RTL/cortexm0ds_logic.v(778)
  wire Ni5bx6;  // ../RTL/cortexm0ds_logic.v(1689)
  wire Ni5ju6;  // ../RTL/cortexm0ds_logic.v(858)
  wire Ni6iu6;  // ../RTL/cortexm0ds_logic.v(390)
  wire Ni6pw6;  // ../RTL/cortexm0ds_logic.v(1415)
  wire Ni7ow6;  // ../RTL/cortexm0ds_logic.v(947)
  wire Nidiu6;  // ../RTL/cortexm0ds_logic.v(484)
  wire Nidpw6;  // ../RTL/cortexm0ds_logic.v(1508)
  wire Nieow6;  // ../RTL/cortexm0ds_logic.v(1040)
  wire Nikiu6;  // ../RTL/cortexm0ds_logic.v(578)
  wire Nilow6;  // ../RTL/cortexm0ds_logic.v(1134)
  wire Niriu6;  // ../RTL/cortexm0ds_logic.v(671)
  wire Nishu6;  // ../RTL/cortexm0ds_logic.v(203)
  wire Nisow6;  // ../RTL/cortexm0ds_logic.v(1228)
  wire Niyiu6;  // ../RTL/cortexm0ds_logic.v(765)
  wire Nizhu6;  // ../RTL/cortexm0ds_logic.v(297)
  wire Nizow6;  // ../RTL/cortexm0ds_logic.v(1321)
  wire Nj2qw6;  // ../RTL/cortexm0ds_logic.v(1622)
  wire Nj4ju6;  // ../RTL/cortexm0ds_logic.v(845)
  wire Nj5iu6;  // ../RTL/cortexm0ds_logic.v(377)
  wire Nj5pw6;  // ../RTL/cortexm0ds_logic.v(1402)
  wire Nj6ow6;  // ../RTL/cortexm0ds_logic.v(934)
  wire Njciu6;  // ../RTL/cortexm0ds_logic.v(471)
  wire Njcpw6;  // ../RTL/cortexm0ds_logic.v(1495)
  wire Njdow6;  // ../RTL/cortexm0ds_logic.v(1027)
  wire Njjiu6;  // ../RTL/cortexm0ds_logic.v(565)
  wire Njkow6;  // ../RTL/cortexm0ds_logic.v(1121)
  wire Njnax6;  // ../RTL/cortexm0ds_logic.v(1657)
  wire Njqiu6;  // ../RTL/cortexm0ds_logic.v(658)
  wire Njrhu6;  // ../RTL/cortexm0ds_logic.v(190)
  wire Njrow6;  // ../RTL/cortexm0ds_logic.v(1215)
  wire Njxiu6;  // ../RTL/cortexm0ds_logic.v(752)
  wire Njyhu6;  // ../RTL/cortexm0ds_logic.v(284)
  wire Njyow6;  // ../RTL/cortexm0ds_logic.v(1308)
  wire Nk3ju6;  // ../RTL/cortexm0ds_logic.v(832)
  wire Nk4iu6;  // ../RTL/cortexm0ds_logic.v(364)
  wire Nk4pw6;  // ../RTL/cortexm0ds_logic.v(1389)
  wire Nk5bx6;  // ../RTL/cortexm0ds_logic.v(1689)
  wire Nkaju6;  // ../RTL/cortexm0ds_logic.v(926)
  wire Nkbiu6;  // ../RTL/cortexm0ds_logic.v(458)
  wire Nkbpw6;  // ../RTL/cortexm0ds_logic.v(1482)
  wire Nkcow6;  // ../RTL/cortexm0ds_logic.v(1014)
  wire Nkiiu6;  // ../RTL/cortexm0ds_logic.v(552)
  wire Nkjow6;  // ../RTL/cortexm0ds_logic.v(1108)
  wire Nkpiu6;  // ../RTL/cortexm0ds_logic.v(645)
  wire Nkqhu6;  // ../RTL/cortexm0ds_logic.v(177)
  wire Nkqow6;  // ../RTL/cortexm0ds_logic.v(1202)
  wire Nkwiu6;  // ../RTL/cortexm0ds_logic.v(739)
  wire Nkxhu6;  // ../RTL/cortexm0ds_logic.v(271)
  wire Nkxow6;  // ../RTL/cortexm0ds_logic.v(1295)
  wire Nl2ju6;  // ../RTL/cortexm0ds_logic.v(819)
  wire Nl3iu6;  // ../RTL/cortexm0ds_logic.v(351)
  wire Nl3pw6;  // ../RTL/cortexm0ds_logic.v(1376)
  wire Nl9ju6;  // ../RTL/cortexm0ds_logic.v(913)
  wire Nlaiu6;  // ../RTL/cortexm0ds_logic.v(445)
  wire Nlapw6;  // ../RTL/cortexm0ds_logic.v(1469)
  wire Nlbbx6;  // ../RTL/cortexm0ds_logic.v(1700)
  wire Nlbow6;  // ../RTL/cortexm0ds_logic.v(1001)
  wire Nlcbx6;  // ../RTL/cortexm0ds_logic.v(1702)
  wire Nlhax6;  // ../RTL/cortexm0ds_logic.v(1646)
  wire Nlhiu6;  // ../RTL/cortexm0ds_logic.v(539)
  wire Nliow6;  // ../RTL/cortexm0ds_logic.v(1095)
  wire Nlnax6;  // ../RTL/cortexm0ds_logic.v(1657)
  wire Nloiu6;  // ../RTL/cortexm0ds_logic.v(632)
  wire Nlphu6;  // ../RTL/cortexm0ds_logic.v(164)
  wire Nlpow6;  // ../RTL/cortexm0ds_logic.v(1189)
  wire Nlviu6;  // ../RTL/cortexm0ds_logic.v(726)
  wire Nlwhu6;  // ../RTL/cortexm0ds_logic.v(258)
  wire Nlwow6;  // ../RTL/cortexm0ds_logic.v(1282)
  wire Nm1ju6;  // ../RTL/cortexm0ds_logic.v(806)
  wire Nm2iu6;  // ../RTL/cortexm0ds_logic.v(338)
  wire Nm2pw6;  // ../RTL/cortexm0ds_logic.v(1363)
  wire Nm5bx6;  // ../RTL/cortexm0ds_logic.v(1689)
  wire Nm8ju6;  // ../RTL/cortexm0ds_logic.v(900)
  wire Nm9iu6;  // ../RTL/cortexm0ds_logic.v(432)
  wire Nm9pw6;  // ../RTL/cortexm0ds_logic.v(1456)
  wire Nmabx6;  // ../RTL/cortexm0ds_logic.v(1698)
  wire Nmaow6;  // ../RTL/cortexm0ds_logic.v(988)
  wire Nmfax6;  // ../RTL/cortexm0ds_logic.v(1642)
  wire Nmgiu6;  // ../RTL/cortexm0ds_logic.v(526)
  wire Nmhow6;  // ../RTL/cortexm0ds_logic.v(1082)
  wire Nmniu6;  // ../RTL/cortexm0ds_logic.v(619)
  wire Nmohu6;  // ../RTL/cortexm0ds_logic.v(151)
  wire Nmoow6;  // ../RTL/cortexm0ds_logic.v(1176)
  wire Nmuiu6;  // ../RTL/cortexm0ds_logic.v(713)
  wire Nmvhu6;  // ../RTL/cortexm0ds_logic.v(245)
  wire Nmvow6;  // ../RTL/cortexm0ds_logic.v(1269)
  wire Nn0ju6;  // ../RTL/cortexm0ds_logic.v(793)
  wire Nn1iu6;  // ../RTL/cortexm0ds_logic.v(325)
  wire Nn1pw6;  // ../RTL/cortexm0ds_logic.v(1350)
  wire Nn7ju6;  // ../RTL/cortexm0ds_logic.v(887)
  wire Nn8iu6;  // ../RTL/cortexm0ds_logic.v(419)
  wire Nn8pw6;  // ../RTL/cortexm0ds_logic.v(1443)
  wire Nn9ow6;  // ../RTL/cortexm0ds_logic.v(975)
  wire Nnfbx6;  // ../RTL/cortexm0ds_logic.v(1708)
  wire Nnfiu6;  // ../RTL/cortexm0ds_logic.v(513)
  wire Nngow6;  // ../RTL/cortexm0ds_logic.v(1069)
  wire Nnmiu6;  // ../RTL/cortexm0ds_logic.v(606)
  wire Nnnax6;  // ../RTL/cortexm0ds_logic.v(1657)
  wire Nnnow6;  // ../RTL/cortexm0ds_logic.v(1163)
  wire Nntiu6;  // ../RTL/cortexm0ds_logic.v(700)
  wire Nnuhu6;  // ../RTL/cortexm0ds_logic.v(232)
  wire Nnuow6;  // ../RTL/cortexm0ds_logic.v(1256)
  wire No0iu6;  // ../RTL/cortexm0ds_logic.v(312)
  wire No0pw6;  // ../RTL/cortexm0ds_logic.v(1337)
  wire No3qw6;  // ../RTL/cortexm0ds_logic.v(1624)
  wire No5bx6;  // ../RTL/cortexm0ds_logic.v(1689)
  wire No6ju6;  // ../RTL/cortexm0ds_logic.v(874)
  wire No7iu6;  // ../RTL/cortexm0ds_logic.v(406)
  wire No7pw6;  // ../RTL/cortexm0ds_logic.v(1430)
  wire No8ow6;  // ../RTL/cortexm0ds_logic.v(962)
  wire Nodax6;  // ../RTL/cortexm0ds_logic.v(1638)
  wire Noeiu6;  // ../RTL/cortexm0ds_logic.v(500)
  wire Nofow6;  // ../RTL/cortexm0ds_logic.v(1056)
  wire Noliu6;  // ../RTL/cortexm0ds_logic.v(593)
  wire Nomow6;  // ../RTL/cortexm0ds_logic.v(1150)
  wire Nosiu6;  // ../RTL/cortexm0ds_logic.v(687)
  wire Nothu6;  // ../RTL/cortexm0ds_logic.v(219)
  wire Notow6;  // ../RTL/cortexm0ds_logic.v(1243)
  wire Noziu6;  // ../RTL/cortexm0ds_logic.v(780)
  wire Np5ju6;  // ../RTL/cortexm0ds_logic.v(861)
  wire Np6iu6;  // ../RTL/cortexm0ds_logic.v(393)
  wire Np6pw6;  // ../RTL/cortexm0ds_logic.v(1417)
  wire Np7ow6;  // ../RTL/cortexm0ds_logic.v(949)
  wire Npaax6;  // ../RTL/cortexm0ds_logic.v(1633)
  wire Npdhu6;  // ../RTL/cortexm0ds_logic.v(120)
  wire Npdiu6;  // ../RTL/cortexm0ds_logic.v(487)
  wire Npdpw6;  // ../RTL/cortexm0ds_logic.v(1511)
  wire Npeow6;  // ../RTL/cortexm0ds_logic.v(1043)
  wire Npghu6;  // ../RTL/cortexm0ds_logic.v(127)
  wire Npkiu6;  // ../RTL/cortexm0ds_logic.v(580)
  wire Nplow6;  // ../RTL/cortexm0ds_logic.v(1137)
  wire Npnax6;  // ../RTL/cortexm0ds_logic.v(1657)
  wire Npriu6;  // ../RTL/cortexm0ds_logic.v(674)
  wire Npshu6;  // ../RTL/cortexm0ds_logic.v(206)
  wire Npsow6;  // ../RTL/cortexm0ds_logic.v(1230)
  wire Npyiu6;  // ../RTL/cortexm0ds_logic.v(767)
  wire Npypw6;  // ../RTL/cortexm0ds_logic.v(1615)
  wire Npzhu6;  // ../RTL/cortexm0ds_logic.v(299)
  wire Npzow6;  // ../RTL/cortexm0ds_logic.v(1324)
  wire Nq4ju6;  // ../RTL/cortexm0ds_logic.v(848)
  wire Nq5bx6;  // ../RTL/cortexm0ds_logic.v(1689)
  wire Nq5iu6;  // ../RTL/cortexm0ds_logic.v(380)
  wire Nq5pw6;  // ../RTL/cortexm0ds_logic.v(1404)
  wire Nq6ow6;  // ../RTL/cortexm0ds_logic.v(936)
  wire Nqciu6;  // ../RTL/cortexm0ds_logic.v(474)
  wire Nqcpw6;  // ../RTL/cortexm0ds_logic.v(1498)
  wire Nqdow6;  // ../RTL/cortexm0ds_logic.v(1030)
  wire Nqjiu6;  // ../RTL/cortexm0ds_logic.v(567)
  wire Nqkow6;  // ../RTL/cortexm0ds_logic.v(1124)
  wire Nqqiu6;  // ../RTL/cortexm0ds_logic.v(661)
  wire Nqrhu6;  // ../RTL/cortexm0ds_logic.v(193)
  wire Nqrow6;  // ../RTL/cortexm0ds_logic.v(1217)
  wire Nqxiu6;  // ../RTL/cortexm0ds_logic.v(754)
  wire Nqyhu6;  // ../RTL/cortexm0ds_logic.v(286)
  wire Nqyow6;  // ../RTL/cortexm0ds_logic.v(1311)
  wire Nr0bx6;  // ../RTL/cortexm0ds_logic.v(1681)
  wire Nr3ju6;  // ../RTL/cortexm0ds_logic.v(835)
  wire Nr4iu6;  // ../RTL/cortexm0ds_logic.v(367)
  wire Nr4pw6;  // ../RTL/cortexm0ds_logic.v(1391)
  wire Nr7ax6;  // ../RTL/cortexm0ds_logic.v(1627)
  wire Nraju6;  // ../RTL/cortexm0ds_logic.v(929)
  wire Nrbiu6;  // ../RTL/cortexm0ds_logic.v(461)
  wire Nrbpw6;  // ../RTL/cortexm0ds_logic.v(1485)
  wire Nrcow6;  // ../RTL/cortexm0ds_logic.v(1017)
  wire Nriiu6;  // ../RTL/cortexm0ds_logic.v(554)
  wire Nrjow6;  // ../RTL/cortexm0ds_logic.v(1111)
  wire Nrkpw6;  // ../RTL/cortexm0ds_logic.v(1589)
  wire Nrnax6;  // ../RTL/cortexm0ds_logic.v(1657)
  wire Nrpiu6;  // ../RTL/cortexm0ds_logic.v(648)
  wire Nrqhu6;  // ../RTL/cortexm0ds_logic.v(180)
  wire Nrqow6;  // ../RTL/cortexm0ds_logic.v(1204)
  wire Nrqpw6;  // ../RTL/cortexm0ds_logic.v(1600)
  wire Nrwiu6;  // ../RTL/cortexm0ds_logic.v(741)
  wire Nrxhu6;  // ../RTL/cortexm0ds_logic.v(273)
  wire Nrxow6;  // ../RTL/cortexm0ds_logic.v(1298)
  wire Ns2ju6;  // ../RTL/cortexm0ds_logic.v(822)
  wire Ns3iu6;  // ../RTL/cortexm0ds_logic.v(354)
  wire Ns3pw6;  // ../RTL/cortexm0ds_logic.v(1378)
  wire Ns8ax6;  // ../RTL/cortexm0ds_logic.v(1629)
  wire Ns9ju6;  // ../RTL/cortexm0ds_logic.v(916)
  wire Nsaiu6;  // ../RTL/cortexm0ds_logic.v(448)
  wire Nsapw6;  // ../RTL/cortexm0ds_logic.v(1472)
  wire Nsbow6;  // ../RTL/cortexm0ds_logic.v(1004)
  wire Nshiu6;  // ../RTL/cortexm0ds_logic.v(541)
  wire Nsiow6;  // ../RTL/cortexm0ds_logic.v(1098)
  wire Nsoiu6;  // ../RTL/cortexm0ds_logic.v(635)
  wire Nsphu6;  // ../RTL/cortexm0ds_logic.v(167)
  wire Nspow6;  // ../RTL/cortexm0ds_logic.v(1191)
  wire Nsviu6;  // ../RTL/cortexm0ds_logic.v(728)
  wire Nswhu6;  // ../RTL/cortexm0ds_logic.v(260)
  wire Nswow6;  // ../RTL/cortexm0ds_logic.v(1285)
  wire Nt1ju6;  // ../RTL/cortexm0ds_logic.v(809)
  wire Nt2iu6;  // ../RTL/cortexm0ds_logic.v(341)
  wire Nt2pw6;  // ../RTL/cortexm0ds_logic.v(1365)
  wire Nt8ju6;  // ../RTL/cortexm0ds_logic.v(903)
  wire Nt9bx6;  // ../RTL/cortexm0ds_logic.v(1697)
  wire Nt9iu6;  // ../RTL/cortexm0ds_logic.v(435)
  wire Nt9pw6;  // ../RTL/cortexm0ds_logic.v(1459)
  wire Ntaow6;  // ../RTL/cortexm0ds_logic.v(991)
  wire Ntfhu6;  // ../RTL/cortexm0ds_logic.v(125)
  wire Ntgiu6;  // ../RTL/cortexm0ds_logic.v(528)
  wire Nthow6;  // ../RTL/cortexm0ds_logic.v(1085)
  wire Ntnax6;  // ../RTL/cortexm0ds_logic.v(1657)
  wire Ntniu6;  // ../RTL/cortexm0ds_logic.v(622)
  wire Ntohu6;  // ../RTL/cortexm0ds_logic.v(154)
  wire Ntoow6;  // ../RTL/cortexm0ds_logic.v(1178)
  wire Ntuiu6;  // ../RTL/cortexm0ds_logic.v(715)
  wire Ntvhu6;  // ../RTL/cortexm0ds_logic.v(247)
  wire Ntvow6;  // ../RTL/cortexm0ds_logic.v(1272)
  wire Nu0ju6;  // ../RTL/cortexm0ds_logic.v(796)
  wire Nu1iu6;  // ../RTL/cortexm0ds_logic.v(328)
  wire Nu1pw6;  // ../RTL/cortexm0ds_logic.v(1352)
  wire Nu5bx6;  // ../RTL/cortexm0ds_logic.v(1689)
  wire Nu7ju6;  // ../RTL/cortexm0ds_logic.v(890)
  wire Nu8iu6;  // ../RTL/cortexm0ds_logic.v(422)
  wire Nu8pw6;  // ../RTL/cortexm0ds_logic.v(1446)
  wire Nu9ow6;  // ../RTL/cortexm0ds_logic.v(978)
  wire Nufiu6;  // ../RTL/cortexm0ds_logic.v(515)
  wire Nugow6;  // ../RTL/cortexm0ds_logic.v(1072)
  wire Numiu6;  // ../RTL/cortexm0ds_logic.v(609)
  wire Nunow6;  // ../RTL/cortexm0ds_logic.v(1165)
  wire Nutiu6;  // ../RTL/cortexm0ds_logic.v(702)
  wire Nuuhu6;  // ../RTL/cortexm0ds_logic.v(234)
  wire Nuuow6;  // ../RTL/cortexm0ds_logic.v(1259)
  wire Nv0iu6;  // ../RTL/cortexm0ds_logic.v(315)
  wire Nv0pw6;  // ../RTL/cortexm0ds_logic.v(1339)
  wire Nv3qw6;  // ../RTL/cortexm0ds_logic.v(1624)
  wire Nv6ju6;  // ../RTL/cortexm0ds_logic.v(877)
  wire Nv7iu6;  // ../RTL/cortexm0ds_logic.v(409)
  wire Nv7pw6;  // ../RTL/cortexm0ds_logic.v(1433)
  wire Nv8ow6;  // ../RTL/cortexm0ds_logic.v(965)
  wire Nv9bx6;  // ../RTL/cortexm0ds_logic.v(1697)
  wire Nveiu6;  // ../RTL/cortexm0ds_logic.v(502)
  wire Nvfow6;  // ../RTL/cortexm0ds_logic.v(1059)
  wire Nvliu6;  // ../RTL/cortexm0ds_logic.v(596)
  wire Nvmow6;  // ../RTL/cortexm0ds_logic.v(1152)
  wire Nvnax6;  // ../RTL/cortexm0ds_logic.v(1657)
  wire Nvsiu6;  // ../RTL/cortexm0ds_logic.v(689)
  wire Nvthu6;  // ../RTL/cortexm0ds_logic.v(221)
  wire Nvtow6;  // ../RTL/cortexm0ds_logic.v(1246)
  wire Nvziu6;  // ../RTL/cortexm0ds_logic.v(783)
  wire Nw5ju6;  // ../RTL/cortexm0ds_logic.v(864)
  wire Nw6iu6;  // ../RTL/cortexm0ds_logic.v(396)
  wire Nw6pw6;  // ../RTL/cortexm0ds_logic.v(1420)
  wire Nw7ow6;  // ../RTL/cortexm0ds_logic.v(952)
  wire Nwbbx6;  // ../RTL/cortexm0ds_logic.v(1701)
  wire Nwdbx6;  // ../RTL/cortexm0ds_logic.v(1704)
  wire Nwdiu6;  // ../RTL/cortexm0ds_logic.v(489)
  wire Nwdpw6;  // ../RTL/cortexm0ds_logic.v(1514)
  wire Nweow6;  // ../RTL/cortexm0ds_logic.v(1046)
  wire Nwkiu6;  // ../RTL/cortexm0ds_logic.v(583)
  wire Nwlow6;  // ../RTL/cortexm0ds_logic.v(1139)
  wire Nwriu6;  // ../RTL/cortexm0ds_logic.v(676)
  wire Nwshu6;  // ../RTL/cortexm0ds_logic.v(208)
  wire Nwsow6;  // ../RTL/cortexm0ds_logic.v(1233)
  wire Nwyiu6;  // ../RTL/cortexm0ds_logic.v(770)
  wire Nwzhu6;  // ../RTL/cortexm0ds_logic.v(302)
  wire Nwzow6;  // ../RTL/cortexm0ds_logic.v(1326)
  wire Nx4ju6;  // ../RTL/cortexm0ds_logic.v(851)
  wire Nx5iu6;  // ../RTL/cortexm0ds_logic.v(383)
  wire Nx5pw6;  // ../RTL/cortexm0ds_logic.v(1407)
  wire Nx6ow6;  // ../RTL/cortexm0ds_logic.v(939)
  wire Nxabx6;  // ../RTL/cortexm0ds_logic.v(1699)
  wire Nxciu6;  // ../RTL/cortexm0ds_logic.v(476)
  wire Nxcpw6;  // ../RTL/cortexm0ds_logic.v(1501)
  wire Nxdow6;  // ../RTL/cortexm0ds_logic.v(1033)
  wire Nxjiu6;  // ../RTL/cortexm0ds_logic.v(570)
  wire Nxkow6;  // ../RTL/cortexm0ds_logic.v(1126)
  wire Nxnax6;  // ../RTL/cortexm0ds_logic.v(1658)
  wire Nxqiu6;  // ../RTL/cortexm0ds_logic.v(663)
  wire Nxrhu6;  // ../RTL/cortexm0ds_logic.v(195)
  wire Nxrow6;  // ../RTL/cortexm0ds_logic.v(1220)
  wire Nxxiu6;  // ../RTL/cortexm0ds_logic.v(757)
  wire Nxyhu6;  // ../RTL/cortexm0ds_logic.v(289)
  wire Nxyow6;  // ../RTL/cortexm0ds_logic.v(1313)
  wire Ny3ju6;  // ../RTL/cortexm0ds_logic.v(838)
  wire Ny4iu6;  // ../RTL/cortexm0ds_logic.v(370)
  wire Ny4pw6;  // ../RTL/cortexm0ds_logic.v(1394)
  wire Nybbx6;  // ../RTL/cortexm0ds_logic.v(1701)
  wire Nybiu6;  // ../RTL/cortexm0ds_logic.v(463)
  wire Nybpw6;  // ../RTL/cortexm0ds_logic.v(1488)
  wire Nycow6;  // ../RTL/cortexm0ds_logic.v(1020)
  wire Nyhax6;  // ../RTL/cortexm0ds_logic.v(1647)
  wire Nyhpw6;  // ../RTL/cortexm0ds_logic.v(1584)
  wire Nyiiu6;  // ../RTL/cortexm0ds_logic.v(557)
  wire Nyjow6;  // ../RTL/cortexm0ds_logic.v(1113)
  wire Nypiu6;  // ../RTL/cortexm0ds_logic.v(650)
  wire Nyqhu6;  // ../RTL/cortexm0ds_logic.v(182)
  wire Nyqow6;  // ../RTL/cortexm0ds_logic.v(1207)
  wire Nywiu6;  // ../RTL/cortexm0ds_logic.v(744)
  wire Nyxhu6;  // ../RTL/cortexm0ds_logic.v(276)
  wire Nyxow6;  // ../RTL/cortexm0ds_logic.v(1300)
  wire Nz2ju6;  // ../RTL/cortexm0ds_logic.v(825)
  wire Nz3iu6;  // ../RTL/cortexm0ds_logic.v(357)
  wire Nz3pw6;  // ../RTL/cortexm0ds_logic.v(1381)
  wire Nz9ju6;  // ../RTL/cortexm0ds_logic.v(918)
  wire Nzaiu6;  // ../RTL/cortexm0ds_logic.v(450)
  wire Nzapw6;  // ../RTL/cortexm0ds_logic.v(1475)
  wire Nzbow6;  // ../RTL/cortexm0ds_logic.v(1007)
  wire Nzhiu6;  // ../RTL/cortexm0ds_logic.v(544)
  wire Nziow6;  // ../RTL/cortexm0ds_logic.v(1100)
  wire Nznax6;  // ../RTL/cortexm0ds_logic.v(1658)
  wire Nzoiu6;  // ../RTL/cortexm0ds_logic.v(637)
  wire Nzphu6;  // ../RTL/cortexm0ds_logic.v(169)
  wire Nzpow6;  // ../RTL/cortexm0ds_logic.v(1194)
  wire Nzviu6;  // ../RTL/cortexm0ds_logic.v(731)
  wire Nzwhu6;  // ../RTL/cortexm0ds_logic.v(263)
  wire Nzwow6;  // ../RTL/cortexm0ds_logic.v(1287)
  wire O00iu6;  // ../RTL/cortexm0ds_logic.v(304)
  wire O00pw6;  // ../RTL/cortexm0ds_logic.v(1328)
  wire O06ju6;  // ../RTL/cortexm0ds_logic.v(865)
  wire O07iu6;  // ../RTL/cortexm0ds_logic.v(397)
  wire O07pw6;  // ../RTL/cortexm0ds_logic.v(1422)
  wire O08ow6;  // ../RTL/cortexm0ds_logic.v(954)
  wire O0eiu6;  // ../RTL/cortexm0ds_logic.v(491)
  wire O0epw6;  // ../RTL/cortexm0ds_logic.v(1515)
  wire O0fow6;  // ../RTL/cortexm0ds_logic.v(1047)
  wire O0liu6;  // ../RTL/cortexm0ds_logic.v(584)
  wire O0mhu6;  // ../RTL/cortexm0ds_logic.v(141)
  wire O0mow6;  // ../RTL/cortexm0ds_logic.v(1141)
  wire O0sax6;  // ../RTL/cortexm0ds_logic.v(1665)
  wire O0siu6;  // ../RTL/cortexm0ds_logic.v(678)
  wire O0thu6;  // ../RTL/cortexm0ds_logic.v(210)
  wire O0tow6;  // ../RTL/cortexm0ds_logic.v(1234)
  wire O0ziu6;  // ../RTL/cortexm0ds_logic.v(772)
  wire O15ju6;  // ../RTL/cortexm0ds_logic.v(852)
  wire O16iu6;  // ../RTL/cortexm0ds_logic.v(384)
  wire O16pw6;  // ../RTL/cortexm0ds_logic.v(1409)
  wire O17ow6;  // ../RTL/cortexm0ds_logic.v(941)
  wire O1diu6;  // ../RTL/cortexm0ds_logic.v(478)
  wire O1dpw6;  // ../RTL/cortexm0ds_logic.v(1502)
  wire O1eow6;  // ../RTL/cortexm0ds_logic.v(1034)
  wire O1jbx6;  // ../RTL/cortexm0ds_logic.v(1714)
  wire O1kiu6;  // ../RTL/cortexm0ds_logic.v(571)
  wire O1low6;  // ../RTL/cortexm0ds_logic.v(1128)
  wire O1mpw6;  // ../RTL/cortexm0ds_logic.v(1592)
  wire O1ppw6;  // ../RTL/cortexm0ds_logic.v(1597)
  wire O1riu6;  // ../RTL/cortexm0ds_logic.v(665)
  wire O1shu6;  // ../RTL/cortexm0ds_logic.v(197)
  wire O1sow6;  // ../RTL/cortexm0ds_logic.v(1221)
  wire O1yiu6;  // ../RTL/cortexm0ds_logic.v(759)
  wire O1zhu6;  // ../RTL/cortexm0ds_logic.v(291)
  wire O1zow6;  // ../RTL/cortexm0ds_logic.v(1315)
  wire O24ju6;  // ../RTL/cortexm0ds_logic.v(839)
  wire O25iu6;  // ../RTL/cortexm0ds_logic.v(371)
  wire O25pw6;  // ../RTL/cortexm0ds_logic.v(1396)
  wire O2ciu6;  // ../RTL/cortexm0ds_logic.v(465)
  wire O2cpw6;  // ../RTL/cortexm0ds_logic.v(1489)
  wire O2dow6;  // ../RTL/cortexm0ds_logic.v(1021)
  wire O2jiu6;  // ../RTL/cortexm0ds_logic.v(558)
  wire O2kax6;  // ../RTL/cortexm0ds_logic.v(1651)
  wire O2kow6;  // ../RTL/cortexm0ds_logic.v(1115)
  wire O2qiu6;  // ../RTL/cortexm0ds_logic.v(652)
  wire O2rhu6;  // ../RTL/cortexm0ds_logic.v(184)
  wire O2row6;  // ../RTL/cortexm0ds_logic.v(1208)
  wire O2sax6;  // ../RTL/cortexm0ds_logic.v(1665)
  wire O2xiu6;  // ../RTL/cortexm0ds_logic.v(746)
  wire O2yhu6;  // ../RTL/cortexm0ds_logic.v(278)
  wire O2yow6;  // ../RTL/cortexm0ds_logic.v(1302)
  wire O33ju6;  // ../RTL/cortexm0ds_logic.v(826)
  wire O34iu6;  // ../RTL/cortexm0ds_logic.v(358)
  wire O34pw6;  // ../RTL/cortexm0ds_logic.v(1383)
  wire O3aju6;  // ../RTL/cortexm0ds_logic.v(920)
  wire O3biu6;  // ../RTL/cortexm0ds_logic.v(452)
  wire O3bpw6;  // ../RTL/cortexm0ds_logic.v(1476)
  wire O3cow6;  // ../RTL/cortexm0ds_logic.v(1008)
  wire O3iiu6;  // ../RTL/cortexm0ds_logic.v(545)
  wire O3jow6;  // ../RTL/cortexm0ds_logic.v(1102)
  wire O3piu6;  // ../RTL/cortexm0ds_logic.v(639)
  wire O3ppw6;  // ../RTL/cortexm0ds_logic.v(1597)
  wire O3qhu6;  // ../RTL/cortexm0ds_logic.v(171)
  wire O3qow6;  // ../RTL/cortexm0ds_logic.v(1195)
  wire O3wiu6;  // ../RTL/cortexm0ds_logic.v(733)
  wire O3xhu6;  // ../RTL/cortexm0ds_logic.v(265)
  wire O3xow6;  // ../RTL/cortexm0ds_logic.v(1289)
  wire O41qw6;  // ../RTL/cortexm0ds_logic.v(1619)
  wire O42ju6;  // ../RTL/cortexm0ds_logic.v(813)
  wire O43iu6;  // ../RTL/cortexm0ds_logic.v(345)
  wire O43pw6;  // ../RTL/cortexm0ds_logic.v(1370)
  wire O49ju6;  // ../RTL/cortexm0ds_logic.v(907)
  wire O4aiu6;  // ../RTL/cortexm0ds_logic.v(439)
  wire O4apw6;  // ../RTL/cortexm0ds_logic.v(1463)
  wire O4bow6;  // ../RTL/cortexm0ds_logic.v(995)
  wire O4hax6;  // ../RTL/cortexm0ds_logic.v(1645)
  wire O4hiu6;  // ../RTL/cortexm0ds_logic.v(532)
  wire O4iow6;  // ../RTL/cortexm0ds_logic.v(1089)
  wire O4oiu6;  // ../RTL/cortexm0ds_logic.v(626)
  wire O4phu6;  // ../RTL/cortexm0ds_logic.v(158)
  wire O4pow6;  // ../RTL/cortexm0ds_logic.v(1182)
  wire O4sax6;  // ../RTL/cortexm0ds_logic.v(1665)
  wire O4viu6;  // ../RTL/cortexm0ds_logic.v(720)
  wire O4whu6;  // ../RTL/cortexm0ds_logic.v(252)
  wire O4wow6;  // ../RTL/cortexm0ds_logic.v(1276)
  wire O51ju6;  // ../RTL/cortexm0ds_logic.v(800)
  wire O52iu6;  // ../RTL/cortexm0ds_logic.v(332)
  wire O52pw6;  // ../RTL/cortexm0ds_logic.v(1357)
  wire O58ju6;  // ../RTL/cortexm0ds_logic.v(894)
  wire O59iu6;  // ../RTL/cortexm0ds_logic.v(426)
  wire O59pw6;  // ../RTL/cortexm0ds_logic.v(1450)
  wire O5aow6;  // ../RTL/cortexm0ds_logic.v(982)
  wire O5giu6;  // ../RTL/cortexm0ds_logic.v(519)
  wire O5how6;  // ../RTL/cortexm0ds_logic.v(1076)
  wire O5niu6;  // ../RTL/cortexm0ds_logic.v(613)
  wire O5ohu6;  // ../RTL/cortexm0ds_logic.v(146)
  wire O5oow6;  // ../RTL/cortexm0ds_logic.v(1169)
  wire O5ppw6;  // ../RTL/cortexm0ds_logic.v(1597)
  wire O5uiu6;  // ../RTL/cortexm0ds_logic.v(707)
  wire O5vhu6;  // ../RTL/cortexm0ds_logic.v(239)
  wire O5vow6;  // ../RTL/cortexm0ds_logic.v(1263)
  wire O60ju6;  // ../RTL/cortexm0ds_logic.v(787)
  wire O61iu6;  // ../RTL/cortexm0ds_logic.v(319)
  wire O61pw6;  // ../RTL/cortexm0ds_logic.v(1344)
  wire O67ju6;  // ../RTL/cortexm0ds_logic.v(881)
  wire O68iu6;  // ../RTL/cortexm0ds_logic.v(413)
  wire O68pw6;  // ../RTL/cortexm0ds_logic.v(1437)
  wire O69ow6;  // ../RTL/cortexm0ds_logic.v(969)
  wire O6fiu6;  // ../RTL/cortexm0ds_logic.v(506)
  wire O6gow6;  // ../RTL/cortexm0ds_logic.v(1063)
  wire O6miu6;  // ../RTL/cortexm0ds_logic.v(600)
  wire O6now6;  // ../RTL/cortexm0ds_logic.v(1156)
  wire O6sax6;  // ../RTL/cortexm0ds_logic.v(1665)
  wire O6tiu6;  // ../RTL/cortexm0ds_logic.v(694)
  wire O6uhu6;  // ../RTL/cortexm0ds_logic.v(226)
  wire O6uow6;  // ../RTL/cortexm0ds_logic.v(1250)
  wire O70iu6;  // ../RTL/cortexm0ds_logic.v(306)
  wire O70pw6;  // ../RTL/cortexm0ds_logic.v(1331)
  wire O76ju6;  // ../RTL/cortexm0ds_logic.v(868)
  wire O77iu6;  // ../RTL/cortexm0ds_logic.v(400)
  wire O77pw6;  // ../RTL/cortexm0ds_logic.v(1424)
  wire O78ow6;  // ../RTL/cortexm0ds_logic.v(956)
  wire O7eiu6;  // ../RTL/cortexm0ds_logic.v(493)
  wire O7fow6;  // ../RTL/cortexm0ds_logic.v(1050)
  wire O7liu6;  // ../RTL/cortexm0ds_logic.v(587)
  wire O7mow6;  // ../RTL/cortexm0ds_logic.v(1143)
  wire O7siu6;  // ../RTL/cortexm0ds_logic.v(681)
  wire O7thu6;  // ../RTL/cortexm0ds_logic.v(213)
  wire O7tow6;  // ../RTL/cortexm0ds_logic.v(1237)
  wire O7ziu6;  // ../RTL/cortexm0ds_logic.v(774)
  wire O85ju6;  // ../RTL/cortexm0ds_logic.v(855)
  wire O86iu6;  // ../RTL/cortexm0ds_logic.v(387)
  wire O86pw6;  // ../RTL/cortexm0ds_logic.v(1411)
  wire O87ow6;  // ../RTL/cortexm0ds_logic.v(943)
  wire O8diu6;  // ../RTL/cortexm0ds_logic.v(480)
  wire O8dpw6;  // ../RTL/cortexm0ds_logic.v(1505)
  wire O8eow6;  // ../RTL/cortexm0ds_logic.v(1037)
  wire O8kiu6;  // ../RTL/cortexm0ds_logic.v(574)
  wire O8lhu6;  // ../RTL/cortexm0ds_logic.v(139)
  wire O8low6;  // ../RTL/cortexm0ds_logic.v(1130)
  wire O8riu6;  // ../RTL/cortexm0ds_logic.v(668)
  wire O8sax6;  // ../RTL/cortexm0ds_logic.v(1665)
  wire O8shu6;  // ../RTL/cortexm0ds_logic.v(200)
  wire O8sow6;  // ../RTL/cortexm0ds_logic.v(1224)
  wire O8yiu6;  // ../RTL/cortexm0ds_logic.v(761)
  wire O8zhu6;  // ../RTL/cortexm0ds_logic.v(293)
  wire O8zow6;  // ../RTL/cortexm0ds_logic.v(1318)
  wire O94ju6;  // ../RTL/cortexm0ds_logic.v(842)
  wire O95iu6;  // ../RTL/cortexm0ds_logic.v(374)
  wire O95pw6;  // ../RTL/cortexm0ds_logic.v(1398)
  wire O96ow6;  // ../RTL/cortexm0ds_logic.v(930)
  wire O9ciu6;  // ../RTL/cortexm0ds_logic.v(467)
  wire O9cpw6;  // ../RTL/cortexm0ds_logic.v(1492)
  wire O9dow6;  // ../RTL/cortexm0ds_logic.v(1024)
  wire O9jiu6;  // ../RTL/cortexm0ds_logic.v(561)
  wire O9kow6;  // ../RTL/cortexm0ds_logic.v(1117)
  wire O9qiu6;  // ../RTL/cortexm0ds_logic.v(655)
  wire O9rhu6;  // ../RTL/cortexm0ds_logic.v(187)
  wire O9row6;  // ../RTL/cortexm0ds_logic.v(1211)
  wire O9xiu6;  // ../RTL/cortexm0ds_logic.v(748)
  wire O9yhu6;  // ../RTL/cortexm0ds_logic.v(280)
  wire O9yow6;  // ../RTL/cortexm0ds_logic.v(1305)
  wire Oa3ju6;  // ../RTL/cortexm0ds_logic.v(829)
  wire Oa4iu6;  // ../RTL/cortexm0ds_logic.v(361)
  wire Oa4pw6;  // ../RTL/cortexm0ds_logic.v(1385)
  wire Oa5bx6;  // ../RTL/cortexm0ds_logic.v(1688)
  wire Oaaju6;  // ../RTL/cortexm0ds_logic.v(922)
  wire Oabiu6;  // ../RTL/cortexm0ds_logic.v(454)
  wire Oabpw6;  // ../RTL/cortexm0ds_logic.v(1479)
  wire Oacow6;  // ../RTL/cortexm0ds_logic.v(1011)
  wire Oaiiu6;  // ../RTL/cortexm0ds_logic.v(548)
  wire Oajow6;  // ../RTL/cortexm0ds_logic.v(1104)
  wire Oakhu6;  // ../RTL/cortexm0ds_logic.v(136)
  wire Oapiu6;  // ../RTL/cortexm0ds_logic.v(642)
  wire Oaqhu6;  // ../RTL/cortexm0ds_logic.v(174)
  wire Oaqow6;  // ../RTL/cortexm0ds_logic.v(1198)
  wire Oarpw6;  // ../RTL/cortexm0ds_logic.v(1601)
  wire Oasax6;  // ../RTL/cortexm0ds_logic.v(1665)
  wire Oawiu6;  // ../RTL/cortexm0ds_logic.v(735)
  wire Oaxhu6;  // ../RTL/cortexm0ds_logic.v(267)
  wire Oaxow6;  // ../RTL/cortexm0ds_logic.v(1292)
  wire Ob2ju6;  // ../RTL/cortexm0ds_logic.v(816)
  wire Ob3iu6;  // ../RTL/cortexm0ds_logic.v(348)
  wire Ob3pw6;  // ../RTL/cortexm0ds_logic.v(1372)
  wire Ob9ju6;  // ../RTL/cortexm0ds_logic.v(909)
  wire Obaiu6;  // ../RTL/cortexm0ds_logic.v(441)
  wire Obapw6;  // ../RTL/cortexm0ds_logic.v(1466)
  wire Obbow6;  // ../RTL/cortexm0ds_logic.v(998)
  wire Obhiu6;  // ../RTL/cortexm0ds_logic.v(535)
  wire Obiow6;  // ../RTL/cortexm0ds_logic.v(1091)
  wire Oboiu6;  // ../RTL/cortexm0ds_logic.v(629)
  wire Obphu6;  // ../RTL/cortexm0ds_logic.v(161)
  wire Obpow6;  // ../RTL/cortexm0ds_logic.v(1185)
  wire Obviu6;  // ../RTL/cortexm0ds_logic.v(722)
  wire Obwhu6;  // ../RTL/cortexm0ds_logic.v(254)
  wire Obwow6;  // ../RTL/cortexm0ds_logic.v(1279)
  wire Oc1ju6;  // ../RTL/cortexm0ds_logic.v(803)
  wire Oc2iu6;  // ../RTL/cortexm0ds_logic.v(335)
  wire Oc2pw6;  // ../RTL/cortexm0ds_logic.v(1359)
  wire Oc8ju6;  // ../RTL/cortexm0ds_logic.v(896)
  wire Oc9iu6;  // ../RTL/cortexm0ds_logic.v(428)
  wire Oc9pw6;  // ../RTL/cortexm0ds_logic.v(1453)
  wire Ocaow6;  // ../RTL/cortexm0ds_logic.v(985)
  wire Ocfhu6;  // ../RTL/cortexm0ds_logic.v(124)
  wire Ocgiu6;  // ../RTL/cortexm0ds_logic.v(522)
  wire Ochow6;  // ../RTL/cortexm0ds_logic.v(1078)
  wire Ocjhu6;  // ../RTL/cortexm0ds_logic.v(133)
  wire Ocniu6;  // ../RTL/cortexm0ds_logic.v(616)
  wire Ocohu6;  // ../RTL/cortexm0ds_logic.v(148)
  wire Ocoow6;  // ../RTL/cortexm0ds_logic.v(1172)
  wire Ocsax6;  // ../RTL/cortexm0ds_logic.v(1666)
  wire Ocuiu6;  // ../RTL/cortexm0ds_logic.v(709)
  wire Ocvhu6;  // ../RTL/cortexm0ds_logic.v(241)
  wire Ocvow6;  // ../RTL/cortexm0ds_logic.v(1266)
  wire Od0ju6;  // ../RTL/cortexm0ds_logic.v(790)
  wire Od1iu6;  // ../RTL/cortexm0ds_logic.v(322)
  wire Od1pw6;  // ../RTL/cortexm0ds_logic.v(1346)
  wire Od4bx6;  // ../RTL/cortexm0ds_logic.v(1687)
  wire Od7ju6;  // ../RTL/cortexm0ds_logic.v(883)
  wire Od8iu6;  // ../RTL/cortexm0ds_logic.v(415)
  wire Od8pw6;  // ../RTL/cortexm0ds_logic.v(1440)
  wire Od9ow6;  // ../RTL/cortexm0ds_logic.v(972)
  wire Odfiu6;  // ../RTL/cortexm0ds_logic.v(509)
  wire Odgow6;  // ../RTL/cortexm0ds_logic.v(1065)
  wire Odmiu6;  // ../RTL/cortexm0ds_logic.v(603)
  wire Odnax6;  // ../RTL/cortexm0ds_logic.v(1657)
  wire Odnow6;  // ../RTL/cortexm0ds_logic.v(1159)
  wire Odtiu6;  // ../RTL/cortexm0ds_logic.v(696)
  wire Oduhu6;  // ../RTL/cortexm0ds_logic.v(228)
  wire Oduow6;  // ../RTL/cortexm0ds_logic.v(1253)
  wire Oe0iu6;  // ../RTL/cortexm0ds_logic.v(309)
  wire Oe0pw6;  // ../RTL/cortexm0ds_logic.v(1333)
  wire Oe6ju6;  // ../RTL/cortexm0ds_logic.v(870)
  wire Oe7iu6;  // ../RTL/cortexm0ds_logic.v(402)
  wire Oe7pw6;  // ../RTL/cortexm0ds_logic.v(1427)
  wire Oe8ow6;  // ../RTL/cortexm0ds_logic.v(959)
  wire Oeeiu6;  // ../RTL/cortexm0ds_logic.v(496)
  wire Oefow6;  // ../RTL/cortexm0ds_logic.v(1052)
  wire Oeihu6;  // ../RTL/cortexm0ds_logic.v(131)
  wire Oeliu6;  // ../RTL/cortexm0ds_logic.v(590)
  wire Oemow6;  // ../RTL/cortexm0ds_logic.v(1146)
  wire Oesax6;  // ../RTL/cortexm0ds_logic.v(1666)
  wire Oesiu6;  // ../RTL/cortexm0ds_logic.v(683)
  wire Oethu6;  // ../RTL/cortexm0ds_logic.v(215)
  wire Oetow6;  // ../RTL/cortexm0ds_logic.v(1240)
  wire Oeziu6;  // ../RTL/cortexm0ds_logic.v(777)
  wire Of5ju6;  // ../RTL/cortexm0ds_logic.v(857)
  wire Of6iu6;  // ../RTL/cortexm0ds_logic.v(389)
  wire Of6pw6;  // ../RTL/cortexm0ds_logic.v(1414)
  wire Of7ow6;  // ../RTL/cortexm0ds_logic.v(946)
  wire Ofdiu6;  // ../RTL/cortexm0ds_logic.v(483)
  wire Ofdpw6;  // ../RTL/cortexm0ds_logic.v(1507)
  wire Ofeow6;  // ../RTL/cortexm0ds_logic.v(1039)
  wire Ofkiu6;  // ../RTL/cortexm0ds_logic.v(577)
  wire Oflow6;  // ../RTL/cortexm0ds_logic.v(1133)
  wire Ofmpw6;  // ../RTL/cortexm0ds_logic.v(1592)
  wire Ofriu6;  // ../RTL/cortexm0ds_logic.v(670)
  wire Ofshu6;  // ../RTL/cortexm0ds_logic.v(202)
  wire Ofsow6;  // ../RTL/cortexm0ds_logic.v(1227)
  wire Ofyiu6;  // ../RTL/cortexm0ds_logic.v(764)
  wire Ofzhu6;  // ../RTL/cortexm0ds_logic.v(296)
  wire Ofzow6;  // ../RTL/cortexm0ds_logic.v(1320)
  wire Og4ju6;  // ../RTL/cortexm0ds_logic.v(844)
  wire Og5bx6;  // ../RTL/cortexm0ds_logic.v(1689)
  wire Og5iu6;  // ../RTL/cortexm0ds_logic.v(376)
  wire Og5pw6;  // ../RTL/cortexm0ds_logic.v(1401)
  wire Og6ow6;  // ../RTL/cortexm0ds_logic.v(933)
  wire Ogciu6;  // ../RTL/cortexm0ds_logic.v(470)
  wire Ogcpw6;  // ../RTL/cortexm0ds_logic.v(1494)
  wire Ogdow6;  // ../RTL/cortexm0ds_logic.v(1026)
  wire Ogjiu6;  // ../RTL/cortexm0ds_logic.v(564)
  wire Ogkow6;  // ../RTL/cortexm0ds_logic.v(1120)
  wire Ogqiu6;  // ../RTL/cortexm0ds_logic.v(657)
  wire Ogrhu6;  // ../RTL/cortexm0ds_logic.v(189)
  wire Ogrow6;  // ../RTL/cortexm0ds_logic.v(1214)
  wire Ogxiu6;  // ../RTL/cortexm0ds_logic.v(751)
  wire Ogyhu6;  // ../RTL/cortexm0ds_logic.v(283)
  wire Ogyow6;  // ../RTL/cortexm0ds_logic.v(1307)
  wire Oh3ju6;  // ../RTL/cortexm0ds_logic.v(831)
  wire Oh4iu6;  // ../RTL/cortexm0ds_logic.v(363)
  wire Oh4pw6;  // ../RTL/cortexm0ds_logic.v(1388)
  wire Oh8ax6;  // ../RTL/cortexm0ds_logic.v(1628)
  wire Ohaju6;  // ../RTL/cortexm0ds_logic.v(925)
  wire Ohbiu6;  // ../RTL/cortexm0ds_logic.v(457)
  wire Ohbpw6;  // ../RTL/cortexm0ds_logic.v(1481)
  wire Ohcow6;  // ../RTL/cortexm0ds_logic.v(1013)
  wire Ohiiu6;  // ../RTL/cortexm0ds_logic.v(551)
  wire Ohjow6;  // ../RTL/cortexm0ds_logic.v(1107)
  wire Ohpiu6;  // ../RTL/cortexm0ds_logic.v(644)
  wire Ohqhu6;  // ../RTL/cortexm0ds_logic.v(176)
  wire Ohqow6;  // ../RTL/cortexm0ds_logic.v(1201)
  wire Ohwiu6;  // ../RTL/cortexm0ds_logic.v(738)
  wire Ohxhu6;  // ../RTL/cortexm0ds_logic.v(270)
  wire Ohxow6;  // ../RTL/cortexm0ds_logic.v(1294)
  wire Ohyax6;  // ../RTL/cortexm0ds_logic.v(1677)
  wire Oi1bx6;  // ../RTL/cortexm0ds_logic.v(1682)
  wire Oi2ju6;  // ../RTL/cortexm0ds_logic.v(818)
  wire Oi3iu6;  // ../RTL/cortexm0ds_logic.v(350)
  wire Oi3pw6;  // ../RTL/cortexm0ds_logic.v(1375)
  wire Oi9ax6;  // ../RTL/cortexm0ds_logic.v(1630)
  wire Oi9ju6;  // ../RTL/cortexm0ds_logic.v(912)
  wire Oiaiu6;  // ../RTL/cortexm0ds_logic.v(444)
  wire Oiapw6;  // ../RTL/cortexm0ds_logic.v(1468)
  wire Oibow6;  // ../RTL/cortexm0ds_logic.v(1000)
  wire Oihiu6;  // ../RTL/cortexm0ds_logic.v(538)
  wire Oiiow6;  // ../RTL/cortexm0ds_logic.v(1094)
  wire Oikax6;  // ../RTL/cortexm0ds_logic.v(1651)
  wire Oioiu6;  // ../RTL/cortexm0ds_logic.v(631)
  wire Oiphu6;  // ../RTL/cortexm0ds_logic.v(163)
  wire Oipow6;  // ../RTL/cortexm0ds_logic.v(1188)
  wire Oiviu6;  // ../RTL/cortexm0ds_logic.v(725)
  wire Oiwhu6;  // ../RTL/cortexm0ds_logic.v(257)
  wire Oiwow6;  // ../RTL/cortexm0ds_logic.v(1281)
  wire Oj1ju6;  // ../RTL/cortexm0ds_logic.v(805)
  wire Oj2iu6;  // ../RTL/cortexm0ds_logic.v(337)
  wire Oj2pw6;  // ../RTL/cortexm0ds_logic.v(1362)
  wire Oj8ju6;  // ../RTL/cortexm0ds_logic.v(899)
  wire Oj9iu6;  // ../RTL/cortexm0ds_logic.v(431)
  wire Oj9pw6;  // ../RTL/cortexm0ds_logic.v(1455)
  wire Ojaow6;  // ../RTL/cortexm0ds_logic.v(987)
  wire Ojebx6;  // ../RTL/cortexm0ds_logic.v(1706)
  wire Ojgiu6;  // ../RTL/cortexm0ds_logic.v(525)
  wire Ojhow6;  // ../RTL/cortexm0ds_logic.v(1081)
  wire Ojniu6;  // ../RTL/cortexm0ds_logic.v(618)
  wire Ojohu6;  // ../RTL/cortexm0ds_logic.v(150)
  wire Ojoow6;  // ../RTL/cortexm0ds_logic.v(1175)
  wire Ojuiu6;  // ../RTL/cortexm0ds_logic.v(712)
  wire Ojvhu6;  // ../RTL/cortexm0ds_logic.v(244)
  wire Ojvow6;  // ../RTL/cortexm0ds_logic.v(1268)
  wire Ok0ju6;  // ../RTL/cortexm0ds_logic.v(792)
  wire Ok1iu6;  // ../RTL/cortexm0ds_logic.v(324)
  wire Ok1pw6;  // ../RTL/cortexm0ds_logic.v(1349)
  wire Ok2bx6;  // ../RTL/cortexm0ds_logic.v(1684)
  wire Ok7ju6;  // ../RTL/cortexm0ds_logic.v(886)
  wire Ok8iu6;  // ../RTL/cortexm0ds_logic.v(418)
  wire Ok8pw6;  // ../RTL/cortexm0ds_logic.v(1442)
  wire Ok9ow6;  // ../RTL/cortexm0ds_logic.v(974)
  wire Okfax6;  // ../RTL/cortexm0ds_logic.v(1642)
  wire Okfiu6;  // ../RTL/cortexm0ds_logic.v(512)
  wire Okgow6;  // ../RTL/cortexm0ds_logic.v(1068)
  wire Okmiu6;  // ../RTL/cortexm0ds_logic.v(605)
  wire Oknow6;  // ../RTL/cortexm0ds_logic.v(1162)
  wire Oktiu6;  // ../RTL/cortexm0ds_logic.v(699)
  wire Okuhu6;  // ../RTL/cortexm0ds_logic.v(231)
  wire Okuow6;  // ../RTL/cortexm0ds_logic.v(1255)
  wire Ol0iu6;  // ../RTL/cortexm0ds_logic.v(311)
  wire Ol0pw6;  // ../RTL/cortexm0ds_logic.v(1336)
  wire Ol6ju6;  // ../RTL/cortexm0ds_logic.v(873)
  wire Ol7iu6;  // ../RTL/cortexm0ds_logic.v(405)
  wire Ol7pw6;  // ../RTL/cortexm0ds_logic.v(1429)
  wire Ol8ow6;  // ../RTL/cortexm0ds_logic.v(961)
  wire Oleiu6;  // ../RTL/cortexm0ds_logic.v(499)
  wire Olfow6;  // ../RTL/cortexm0ds_logic.v(1055)
  wire Olliu6;  // ../RTL/cortexm0ds_logic.v(592)
  wire Olmow6;  // ../RTL/cortexm0ds_logic.v(1149)
  wire Olsiu6;  // ../RTL/cortexm0ds_logic.v(686)
  wire Olthu6;  // ../RTL/cortexm0ds_logic.v(218)
  wire Oltow6;  // ../RTL/cortexm0ds_logic.v(1242)
  wire Olziu6;  // ../RTL/cortexm0ds_logic.v(779)
  wire Om3bx6;  // ../RTL/cortexm0ds_logic.v(1686)
  wire Om5ju6;  // ../RTL/cortexm0ds_logic.v(860)
  wire Om6iu6;  // ../RTL/cortexm0ds_logic.v(392)
  wire Om6pw6;  // ../RTL/cortexm0ds_logic.v(1416)
  wire Om7ow6;  // ../RTL/cortexm0ds_logic.v(948)
  wire Omdiu6;  // ../RTL/cortexm0ds_logic.v(486)
  wire Omdpw6;  // ../RTL/cortexm0ds_logic.v(1510)
  wire Omeow6;  // ../RTL/cortexm0ds_logic.v(1042)
  wire Omkiu6;  // ../RTL/cortexm0ds_logic.v(579)
  wire Omlow6;  // ../RTL/cortexm0ds_logic.v(1136)
  wire Omriu6;  // ../RTL/cortexm0ds_logic.v(673)
  wire Omshu6;  // ../RTL/cortexm0ds_logic.v(205)
  wire Omsow6;  // ../RTL/cortexm0ds_logic.v(1229)
  wire Omyiu6;  // ../RTL/cortexm0ds_logic.v(766)
  wire Omzhu6;  // ../RTL/cortexm0ds_logic.v(298)
  wire Omzow6;  // ../RTL/cortexm0ds_logic.v(1323)
  wire On4ju6;  // ../RTL/cortexm0ds_logic.v(847)
  wire On5iu6;  // ../RTL/cortexm0ds_logic.v(379)
  wire On5pw6;  // ../RTL/cortexm0ds_logic.v(1403)
  wire On6ow6;  // ../RTL/cortexm0ds_logic.v(935)
  wire Onciu6;  // ../RTL/cortexm0ds_logic.v(473)
  wire Oncpw6;  // ../RTL/cortexm0ds_logic.v(1497)
  wire Ondow6;  // ../RTL/cortexm0ds_logic.v(1029)
  wire Onjiu6;  // ../RTL/cortexm0ds_logic.v(566)
  wire Onkow6;  // ../RTL/cortexm0ds_logic.v(1123)
  wire Onqiu6;  // ../RTL/cortexm0ds_logic.v(660)
  wire Onrhu6;  // ../RTL/cortexm0ds_logic.v(192)
  wire Onrow6;  // ../RTL/cortexm0ds_logic.v(1216)
  wire Onxiu6;  // ../RTL/cortexm0ds_logic.v(753)
  wire Onyhu6;  // ../RTL/cortexm0ds_logic.v(285)
  wire Onyow6;  // ../RTL/cortexm0ds_logic.v(1310)
  wire Onypw6;  // ../RTL/cortexm0ds_logic.v(1614)
  wire Oo3ju6;  // ../RTL/cortexm0ds_logic.v(834)
  wire Oo4iu6;  // ../RTL/cortexm0ds_logic.v(366)
  wire Oo4pw6;  // ../RTL/cortexm0ds_logic.v(1390)
  wire Ooaju6;  // ../RTL/cortexm0ds_logic.v(928)
  wire Oobiu6;  // ../RTL/cortexm0ds_logic.v(460)
  wire Oobpw6;  // ../RTL/cortexm0ds_logic.v(1484)
  wire Oocow6;  // ../RTL/cortexm0ds_logic.v(1016)
  wire Oodhu6;  // ../RTL/cortexm0ds_logic.v(120)
  wire Ooiiu6;  // ../RTL/cortexm0ds_logic.v(553)
  wire Oojow6;  // ../RTL/cortexm0ds_logic.v(1110)
  wire Oopiu6;  // ../RTL/cortexm0ds_logic.v(647)
  wire Ooqhu6;  // ../RTL/cortexm0ds_logic.v(179)
  wire Ooqow6;  // ../RTL/cortexm0ds_logic.v(1203)
  wire Oowiu6;  // ../RTL/cortexm0ds_logic.v(740)
  wire Ooxhu6;  // ../RTL/cortexm0ds_logic.v(272)
  wire Ooxow6;  // ../RTL/cortexm0ds_logic.v(1297)
  wire Op2ju6;  // ../RTL/cortexm0ds_logic.v(821)
  wire Op3iu6;  // ../RTL/cortexm0ds_logic.v(353)
  wire Op3pw6;  // ../RTL/cortexm0ds_logic.v(1377)
  wire Op9ju6;  // ../RTL/cortexm0ds_logic.v(915)
  wire Opaiu6;  // ../RTL/cortexm0ds_logic.v(447)
  wire Opapw6;  // ../RTL/cortexm0ds_logic.v(1471)
  wire Opbax6;  // ../RTL/cortexm0ds_logic.v(1635)
  wire Opbow6;  // ../RTL/cortexm0ds_logic.v(1003)
  wire Ophiu6;  // ../RTL/cortexm0ds_logic.v(540)
  wire Opiow6;  // ../RTL/cortexm0ds_logic.v(1097)
  wire Opoiu6;  // ../RTL/cortexm0ds_logic.v(634)
  wire Opphu6;  // ../RTL/cortexm0ds_logic.v(166)
  wire Oppow6;  // ../RTL/cortexm0ds_logic.v(1190)
  wire Opviu6;  // ../RTL/cortexm0ds_logic.v(727)
  wire Opwhu6;  // ../RTL/cortexm0ds_logic.v(259)
  wire Opwow6;  // ../RTL/cortexm0ds_logic.v(1284)
  wire Oq1ju6;  // ../RTL/cortexm0ds_logic.v(808)
  wire Oq2iu6;  // ../RTL/cortexm0ds_logic.v(340)
  wire Oq2pw6;  // ../RTL/cortexm0ds_logic.v(1364)
  wire Oq8ju6;  // ../RTL/cortexm0ds_logic.v(902)
  wire Oq9iu6;  // ../RTL/cortexm0ds_logic.v(434)
  wire Oq9pw6;  // ../RTL/cortexm0ds_logic.v(1458)
  wire Oqaow6;  // ../RTL/cortexm0ds_logic.v(990)
  wire Oqgiu6;  // ../RTL/cortexm0ds_logic.v(527)
  wire Oqhow6;  // ../RTL/cortexm0ds_logic.v(1084)
  wire Oqniu6;  // ../RTL/cortexm0ds_logic.v(621)
  wire Oqohu6;  // ../RTL/cortexm0ds_logic.v(153)
  wire Oqoow6;  // ../RTL/cortexm0ds_logic.v(1177)
  wire Oquiu6;  // ../RTL/cortexm0ds_logic.v(714)
  wire Oqvhu6;  // ../RTL/cortexm0ds_logic.v(246)
  wire Oqvow6;  // ../RTL/cortexm0ds_logic.v(1271)
  wire Or0ju6;  // ../RTL/cortexm0ds_logic.v(795)
  wire Or1iu6;  // ../RTL/cortexm0ds_logic.v(327)
  wire Or1pw6;  // ../RTL/cortexm0ds_logic.v(1351)
  wire Or7ju6;  // ../RTL/cortexm0ds_logic.v(889)
  wire Or8iu6;  // ../RTL/cortexm0ds_logic.v(421)
  wire Or8pw6;  // ../RTL/cortexm0ds_logic.v(1445)
  wire Or9ow6;  // ../RTL/cortexm0ds_logic.v(977)
  wire Orfiu6;  // ../RTL/cortexm0ds_logic.v(514)
  wire Orgow6;  // ../RTL/cortexm0ds_logic.v(1071)
  wire Orkhu6;  // ../RTL/cortexm0ds_logic.v(137)
  wire Ormiu6;  // ../RTL/cortexm0ds_logic.v(608)
  wire Ornow6;  // ../RTL/cortexm0ds_logic.v(1164)
  wire Ortiu6;  // ../RTL/cortexm0ds_logic.v(701)
  wire Oruhu6;  // ../RTL/cortexm0ds_logic.v(233)
  wire Oruow6;  // ../RTL/cortexm0ds_logic.v(1258)
  wire Os0iu6;  // ../RTL/cortexm0ds_logic.v(314)
  wire Os0pw6;  // ../RTL/cortexm0ds_logic.v(1338)
  wire Os6ju6;  // ../RTL/cortexm0ds_logic.v(876)
  wire Os7iu6;  // ../RTL/cortexm0ds_logic.v(408)
  wire Os7pw6;  // ../RTL/cortexm0ds_logic.v(1432)
  wire Os8ow6;  // ../RTL/cortexm0ds_logic.v(964)
  wire Osehu6;  // ../RTL/cortexm0ds_logic.v(122)
  wire Oseiu6;  // ../RTL/cortexm0ds_logic.v(501)
  wire Osfow6;  // ../RTL/cortexm0ds_logic.v(1058)
  wire Osliu6;  // ../RTL/cortexm0ds_logic.v(595)
  wire Osmow6;  // ../RTL/cortexm0ds_logic.v(1151)
  wire Osrax6;  // ../RTL/cortexm0ds_logic.v(1665)
  wire Ossiu6;  // ../RTL/cortexm0ds_logic.v(688)
  wire Osthu6;  // ../RTL/cortexm0ds_logic.v(220)
  wire Ostow6;  // ../RTL/cortexm0ds_logic.v(1245)
  wire Osziu6;  // ../RTL/cortexm0ds_logic.v(782)
  wire Ot0bx6;  // ../RTL/cortexm0ds_logic.v(1681)
  wire Ot5ju6;  // ../RTL/cortexm0ds_logic.v(863)
  wire Ot6iu6;  // ../RTL/cortexm0ds_logic.v(395)
  wire Ot6pw6;  // ../RTL/cortexm0ds_logic.v(1419)
  wire Ot7ow6;  // ../RTL/cortexm0ds_logic.v(951)
  wire Otdiu6;  // ../RTL/cortexm0ds_logic.v(488)
  wire Otdpw6;  // ../RTL/cortexm0ds_logic.v(1513)
  wire Oteow6;  // ../RTL/cortexm0ds_logic.v(1045)
  wire Otjhu6;  // ../RTL/cortexm0ds_logic.v(135)
  wire Otkiu6;  // ../RTL/cortexm0ds_logic.v(582)
  wire Otlow6;  // ../RTL/cortexm0ds_logic.v(1138)
  wire Otopw6;  // ../RTL/cortexm0ds_logic.v(1597)
  wire Otriu6;  // ../RTL/cortexm0ds_logic.v(675)
  wire Otshu6;  // ../RTL/cortexm0ds_logic.v(207)
  wire Otsow6;  // ../RTL/cortexm0ds_logic.v(1232)
  wire Otyiu6;  // ../RTL/cortexm0ds_logic.v(769)
  wire Otzhu6;  // ../RTL/cortexm0ds_logic.v(301)
  wire Otzow6;  // ../RTL/cortexm0ds_logic.v(1325)
  wire Ou4ju6;  // ../RTL/cortexm0ds_logic.v(850)
  wire Ou5iu6;  // ../RTL/cortexm0ds_logic.v(382)
  wire Ou5pw6;  // ../RTL/cortexm0ds_logic.v(1406)
  wire Ou6ow6;  // ../RTL/cortexm0ds_logic.v(938)
  wire Ouciu6;  // ../RTL/cortexm0ds_logic.v(475)
  wire Oucpw6;  // ../RTL/cortexm0ds_logic.v(1500)
  wire Oudow6;  // ../RTL/cortexm0ds_logic.v(1032)
  wire Oujiu6;  // ../RTL/cortexm0ds_logic.v(569)
  wire Oukow6;  // ../RTL/cortexm0ds_logic.v(1125)
  wire Oulpw6;  // ../RTL/cortexm0ds_logic.v(1591)
  wire Ouqiu6;  // ../RTL/cortexm0ds_logic.v(662)
  wire Ourax6;  // ../RTL/cortexm0ds_logic.v(1665)
  wire Ourhu6;  // ../RTL/cortexm0ds_logic.v(194)
  wire Ourow6;  // ../RTL/cortexm0ds_logic.v(1219)
  wire Ouxiu6;  // ../RTL/cortexm0ds_logic.v(756)
  wire Ouyhu6;  // ../RTL/cortexm0ds_logic.v(288)
  wire Ouyow6;  // ../RTL/cortexm0ds_logic.v(1312)
  wire Ov3ju6;  // ../RTL/cortexm0ds_logic.v(837)
  wire Ov4iu6;  // ../RTL/cortexm0ds_logic.v(369)
  wire Ov4pw6;  // ../RTL/cortexm0ds_logic.v(1393)
  wire Ovbiu6;  // ../RTL/cortexm0ds_logic.v(462)
  wire Ovbpw6;  // ../RTL/cortexm0ds_logic.v(1487)
  wire Ovcow6;  // ../RTL/cortexm0ds_logic.v(1019)
  wire Oveax6;  // ../RTL/cortexm0ds_logic.v(1641)
  wire Ovihu6;  // ../RTL/cortexm0ds_logic.v(132)
  wire Oviiu6;  // ../RTL/cortexm0ds_logic.v(556)
  wire Ovjow6;  // ../RTL/cortexm0ds_logic.v(1112)
  wire Ovopw6;  // ../RTL/cortexm0ds_logic.v(1597)
  wire Ovpiu6;  // ../RTL/cortexm0ds_logic.v(649)
  wire Ovqhu6;  // ../RTL/cortexm0ds_logic.v(181)
  wire Ovqow6;  // ../RTL/cortexm0ds_logic.v(1206)
  wire Ovwiu6;  // ../RTL/cortexm0ds_logic.v(743)
  wire Ovxhu6;  // ../RTL/cortexm0ds_logic.v(275)
  wire Ovxow6;  // ../RTL/cortexm0ds_logic.v(1299)
  wire Ow2ju6;  // ../RTL/cortexm0ds_logic.v(824)
  wire Ow3iu6;  // ../RTL/cortexm0ds_logic.v(356)
  wire Ow3pw6;  // ../RTL/cortexm0ds_logic.v(1380)
  wire Ow9ju6;  // ../RTL/cortexm0ds_logic.v(917)
  wire Owaiu6;  // ../RTL/cortexm0ds_logic.v(449)
  wire Owapw6;  // ../RTL/cortexm0ds_logic.v(1474)
  wire Owbow6;  // ../RTL/cortexm0ds_logic.v(1006)
  wire Owcax6;  // ../RTL/cortexm0ds_logic.v(1637)
  wire Owhbx6;  // ../RTL/cortexm0ds_logic.v(1712)
  wire Owhiu6;  // ../RTL/cortexm0ds_logic.v(543)
  wire Owiow6;  // ../RTL/cortexm0ds_logic.v(1099)
  wire Owoiu6;  // ../RTL/cortexm0ds_logic.v(636)
  wire Owphu6;  // ../RTL/cortexm0ds_logic.v(168)
  wire Owpow6;  // ../RTL/cortexm0ds_logic.v(1193)
  wire Owrax6;  // ../RTL/cortexm0ds_logic.v(1665)
  wire Owviu6;  // ../RTL/cortexm0ds_logic.v(730)
  wire Owwhu6;  // ../RTL/cortexm0ds_logic.v(262)
  wire Owwow6;  // ../RTL/cortexm0ds_logic.v(1286)
  wire Ox1ju6;  // ../RTL/cortexm0ds_logic.v(811)
  wire Ox2iu6;  // ../RTL/cortexm0ds_logic.v(343)
  wire Ox2pw6;  // ../RTL/cortexm0ds_logic.v(1367)
  wire Ox8ju6;  // ../RTL/cortexm0ds_logic.v(904)
  wire Ox9bx6;  // ../RTL/cortexm0ds_logic.v(1697)
  wire Ox9iu6;  // ../RTL/cortexm0ds_logic.v(436)
  wire Ox9pw6;  // ../RTL/cortexm0ds_logic.v(1461)
  wire Oxaow6;  // ../RTL/cortexm0ds_logic.v(993)
  wire Oxgiu6;  // ../RTL/cortexm0ds_logic.v(530)
  wire Oxhhu6;  // ../RTL/cortexm0ds_logic.v(129)
  wire Oxhow6;  // ../RTL/cortexm0ds_logic.v(1086)
  wire Oxkpw6;  // ../RTL/cortexm0ds_logic.v(1589)
  wire Oxniu6;  // ../RTL/cortexm0ds_logic.v(623)
  wire Oxohu6;  // ../RTL/cortexm0ds_logic.v(155)
  wire Oxoow6;  // ../RTL/cortexm0ds_logic.v(1180)
  wire Oxopw6;  // ../RTL/cortexm0ds_logic.v(1597)
  wire Oxuiu6;  // ../RTL/cortexm0ds_logic.v(717)
  wire Oxvhu6;  // ../RTL/cortexm0ds_logic.v(249)
  wire Oxvow6;  // ../RTL/cortexm0ds_logic.v(1273)
  wire Oy0ju6;  // ../RTL/cortexm0ds_logic.v(798)
  wire Oy1iu6;  // ../RTL/cortexm0ds_logic.v(330)
  wire Oy1pw6;  // ../RTL/cortexm0ds_logic.v(1354)
  wire Oy7ju6;  // ../RTL/cortexm0ds_logic.v(891)
  wire Oy8iu6;  // ../RTL/cortexm0ds_logic.v(423)
  wire Oy8pw6;  // ../RTL/cortexm0ds_logic.v(1448)
  wire Oy9ow6;  // ../RTL/cortexm0ds_logic.v(980)
  wire Oyfiu6;  // ../RTL/cortexm0ds_logic.v(517)
  wire Oygow6;  // ../RTL/cortexm0ds_logic.v(1073)
  wire Oyhbx6;  // ../RTL/cortexm0ds_logic.v(1712)
  wire Oykax6;  // ../RTL/cortexm0ds_logic.v(1652)
  wire Oymiu6;  // ../RTL/cortexm0ds_logic.v(610)
  wire Oynow6;  // ../RTL/cortexm0ds_logic.v(1167)
  wire Oyrax6;  // ../RTL/cortexm0ds_logic.v(1665)
  wire Oytiu6;  // ../RTL/cortexm0ds_logic.v(704)
  wire Oyuhu6;  // ../RTL/cortexm0ds_logic.v(236)
  wire Oyuow6;  // ../RTL/cortexm0ds_logic.v(1260)
  wire Oz0iu6;  // ../RTL/cortexm0ds_logic.v(317)
  wire Oz0pw6;  // ../RTL/cortexm0ds_logic.v(1341)
  wire Oz6ju6;  // ../RTL/cortexm0ds_logic.v(878)
  wire Oz7iu6;  // ../RTL/cortexm0ds_logic.v(410)
  wire Oz7pw6;  // ../RTL/cortexm0ds_logic.v(1435)
  wire Oz8ow6;  // ../RTL/cortexm0ds_logic.v(967)
  wire Ozeiu6;  // ../RTL/cortexm0ds_logic.v(504)
  wire Ozfow6;  // ../RTL/cortexm0ds_logic.v(1060)
  wire Ozliu6;  // ../RTL/cortexm0ds_logic.v(597)
  wire Ozmow6;  // ../RTL/cortexm0ds_logic.v(1154)
  wire Ozopw6;  // ../RTL/cortexm0ds_logic.v(1597)
  wire Ozsiu6;  // ../RTL/cortexm0ds_logic.v(691)
  wire Ozthu6;  // ../RTL/cortexm0ds_logic.v(223)
  wire Oztow6;  // ../RTL/cortexm0ds_logic.v(1247)
  wire Ozvax6;  // ../RTL/cortexm0ds_logic.v(1672)
  wire Ozziu6;  // ../RTL/cortexm0ds_logic.v(785)
  wire P03ju6;  // ../RTL/cortexm0ds_logic.v(825)
  wire P04iu6;  // ../RTL/cortexm0ds_logic.v(357)
  wire P04pw6;  // ../RTL/cortexm0ds_logic.v(1381)
  wire P0aju6;  // ../RTL/cortexm0ds_logic.v(919)
  wire P0bax6;  // ../RTL/cortexm0ds_logic.v(1633)
  wire P0biu6;  // ../RTL/cortexm0ds_logic.v(451)
  wire P0bpw6;  // ../RTL/cortexm0ds_logic.v(1475)
  wire P0cow6;  // ../RTL/cortexm0ds_logic.v(1007)
  wire P0ibx6;  // ../RTL/cortexm0ds_logic.v(1712)
  wire P0iiu6;  // ../RTL/cortexm0ds_logic.v(544)
  wire P0jow6;  // ../RTL/cortexm0ds_logic.v(1101)
  wire P0kax6;  // ../RTL/cortexm0ds_logic.v(1650)
  wire P0piu6;  // ../RTL/cortexm0ds_logic.v(638)
  wire P0qhu6;  // ../RTL/cortexm0ds_logic.v(170)
  wire P0qow6;  // ../RTL/cortexm0ds_logic.v(1194)
  wire P0wiu6;  // ../RTL/cortexm0ds_logic.v(731)
  wire P0xhu6;  // ../RTL/cortexm0ds_logic.v(263)
  wire P0xow6;  // ../RTL/cortexm0ds_logic.v(1288)
  wire P12bx6;  // ../RTL/cortexm0ds_logic.v(1683)
  wire P12ju6;  // ../RTL/cortexm0ds_logic.v(812)
  wire P13iu6;  // ../RTL/cortexm0ds_logic.v(344)
  wire P13pw6;  // ../RTL/cortexm0ds_logic.v(1368)
  wire P14qw6;  // ../RTL/cortexm0ds_logic.v(1625)
  wire P19ju6;  // ../RTL/cortexm0ds_logic.v(906)
  wire P1aiu6;  // ../RTL/cortexm0ds_logic.v(438)
  wire P1apw6;  // ../RTL/cortexm0ds_logic.v(1462)
  wire P1bow6;  // ../RTL/cortexm0ds_logic.v(994)
  wire P1hiu6;  // ../RTL/cortexm0ds_logic.v(531)
  wire P1iow6;  // ../RTL/cortexm0ds_logic.v(1088)
  wire P1oiu6;  // ../RTL/cortexm0ds_logic.v(625)
  wire P1phu6;  // ../RTL/cortexm0ds_logic.v(157)
  wire P1pow6;  // ../RTL/cortexm0ds_logic.v(1181)
  wire P1viu6;  // ../RTL/cortexm0ds_logic.v(718)
  wire P1whu6;  // ../RTL/cortexm0ds_logic.v(250)
  wire P1wow6;  // ../RTL/cortexm0ds_logic.v(1275)
  wire P21ju6;  // ../RTL/cortexm0ds_logic.v(799)
  wire P21qw6;  // ../RTL/cortexm0ds_logic.v(1619)
  wire P22iu6;  // ../RTL/cortexm0ds_logic.v(331)
  wire P22pw6;  // ../RTL/cortexm0ds_logic.v(1355)
  wire P23qw6;  // ../RTL/cortexm0ds_logic.v(1623)
  wire P28ju6;  // ../RTL/cortexm0ds_logic.v(893)
  wire P29iu6;  // ../RTL/cortexm0ds_logic.v(425)
  wire P29pw6;  // ../RTL/cortexm0ds_logic.v(1449)
  wire P2aow6;  // ../RTL/cortexm0ds_logic.v(981)
  wire P2giu6;  // ../RTL/cortexm0ds_logic.v(518)
  wire P2how6;  // ../RTL/cortexm0ds_logic.v(1075)
  wire P2niu6;  // ../RTL/cortexm0ds_logic.v(612)
  wire P2oow6;  // ../RTL/cortexm0ds_logic.v(1168)
  wire P2uiu6;  // ../RTL/cortexm0ds_logic.v(705)
  wire P2vhu6;  // ../RTL/cortexm0ds_logic.v(237)
  wire P2vow6;  // ../RTL/cortexm0ds_logic.v(1262)
  wire P2xpw6;  // ../RTL/cortexm0ds_logic.v(1612)
  wire P30ju6;  // ../RTL/cortexm0ds_logic.v(786)
  wire P31iu6;  // ../RTL/cortexm0ds_logic.v(318)
  wire P31pw6;  // ../RTL/cortexm0ds_logic.v(1342)
  wire P33bx6;  // ../RTL/cortexm0ds_logic.v(1685)
  wire P34qw6;  // ../RTL/cortexm0ds_logic.v(1625)
  wire P37ju6;  // ../RTL/cortexm0ds_logic.v(880)
  wire P38iu6;  // ../RTL/cortexm0ds_logic.v(412)
  wire P38pw6;  // ../RTL/cortexm0ds_logic.v(1436)
  wire P39ow6;  // ../RTL/cortexm0ds_logic.v(968)
  wire P3fiu6;  // ../RTL/cortexm0ds_logic.v(505)
  wire P3gow6;  // ../RTL/cortexm0ds_logic.v(1062)
  wire P3miu6;  // ../RTL/cortexm0ds_logic.v(599)
  wire P3now6;  // ../RTL/cortexm0ds_logic.v(1155)
  wire P3tiu6;  // ../RTL/cortexm0ds_logic.v(692)
  wire P3uhu6;  // ../RTL/cortexm0ds_logic.v(224)
  wire P3uow6;  // ../RTL/cortexm0ds_logic.v(1249)
  wire P40iu6;  // ../RTL/cortexm0ds_logic.v(305)
  wire P40pw6;  // ../RTL/cortexm0ds_logic.v(1329)
  wire P46ju6;  // ../RTL/cortexm0ds_logic.v(867)
  wire P47iu6;  // ../RTL/cortexm0ds_logic.v(399)
  wire P47pw6;  // ../RTL/cortexm0ds_logic.v(1423)
  wire P48ow6;  // ../RTL/cortexm0ds_logic.v(955)
  wire P4cax6;  // ../RTL/cortexm0ds_logic.v(1635)
  wire P4eiu6;  // ../RTL/cortexm0ds_logic.v(492)
  wire P4epw6;  // ../RTL/cortexm0ds_logic.v(1517)
  wire P4fow6;  // ../RTL/cortexm0ds_logic.v(1049)
  wire P4liu6;  // ../RTL/cortexm0ds_logic.v(586)
  wire P4mow6;  // ../RTL/cortexm0ds_logic.v(1142)
  wire P4siu6;  // ../RTL/cortexm0ds_logic.v(679)
  wire P4thu6;  // ../RTL/cortexm0ds_logic.v(211)
  wire P4tow6;  // ../RTL/cortexm0ds_logic.v(1236)
  wire P4xpw6;  // ../RTL/cortexm0ds_logic.v(1612)
  wire P4ziu6;  // ../RTL/cortexm0ds_logic.v(773)
  wire P54qw6;  // ../RTL/cortexm0ds_logic.v(1625)
  wire P55ju6;  // ../RTL/cortexm0ds_logic.v(854)
  wire P56iu6;  // ../RTL/cortexm0ds_logic.v(386)
  wire P56pw6;  // ../RTL/cortexm0ds_logic.v(1410)
  wire P57ow6;  // ../RTL/cortexm0ds_logic.v(942)
  wire P5diu6;  // ../RTL/cortexm0ds_logic.v(479)
  wire P5dpw6;  // ../RTL/cortexm0ds_logic.v(1504)
  wire P5eow6;  // ../RTL/cortexm0ds_logic.v(1036)
  wire P5kiu6;  // ../RTL/cortexm0ds_logic.v(573)
  wire P5low6;  // ../RTL/cortexm0ds_logic.v(1129)
  wire P5riu6;  // ../RTL/cortexm0ds_logic.v(666)
  wire P5shu6;  // ../RTL/cortexm0ds_logic.v(198)
  wire P5sow6;  // ../RTL/cortexm0ds_logic.v(1223)
  wire P5vpw6;  // ../RTL/cortexm0ds_logic.v(1608)
  wire P5yiu6;  // ../RTL/cortexm0ds_logic.v(760)
  wire P5zhu6;  // ../RTL/cortexm0ds_logic.v(292)
  wire P5zow6;  // ../RTL/cortexm0ds_logic.v(1316)
  wire P64ju6;  // ../RTL/cortexm0ds_logic.v(841)
  wire P65iu6;  // ../RTL/cortexm0ds_logic.v(373)
  wire P65pw6;  // ../RTL/cortexm0ds_logic.v(1397)
  wire P6ciu6;  // ../RTL/cortexm0ds_logic.v(466)
  wire P6cpw6;  // ../RTL/cortexm0ds_logic.v(1491)
  wire P6dow6;  // ../RTL/cortexm0ds_logic.v(1023)
  wire P6jiu6;  // ../RTL/cortexm0ds_logic.v(560)
  wire P6kow6;  // ../RTL/cortexm0ds_logic.v(1116)
  wire P6qiu6;  // ../RTL/cortexm0ds_logic.v(653)
  wire P6rhu6;  // ../RTL/cortexm0ds_logic.v(185)
  wire P6row6;  // ../RTL/cortexm0ds_logic.v(1210)
  wire P6xiu6;  // ../RTL/cortexm0ds_logic.v(747)
  wire P6xpw6;  // ../RTL/cortexm0ds_logic.v(1612)
  wire P6yhu6;  // ../RTL/cortexm0ds_logic.v(279)
  wire P6yow6;  // ../RTL/cortexm0ds_logic.v(1303)
  wire P73ju6;  // ../RTL/cortexm0ds_logic.v(828)
  wire P74iu6;  // ../RTL/cortexm0ds_logic.v(360)
  wire P74pw6;  // ../RTL/cortexm0ds_logic.v(1384)
  wire P7aju6;  // ../RTL/cortexm0ds_logic.v(921)
  wire P7bbx6;  // ../RTL/cortexm0ds_logic.v(1699)
  wire P7biu6;  // ../RTL/cortexm0ds_logic.v(453)
  wire P7bpw6;  // ../RTL/cortexm0ds_logic.v(1478)
  wire P7iiu6;  // ../RTL/cortexm0ds_logic.v(547)
  wire P7jow6;  // ../RTL/cortexm0ds_logic.v(1103)
  wire P7piu6;  // ../RTL/cortexm0ds_logic.v(640)
  wire P7qhu6;  // ../RTL/cortexm0ds_logic.v(172)
  wire P7qow6;  // ../RTL/cortexm0ds_logic.v(1197)
  wire P7wiu6;  // ../RTL/cortexm0ds_logic.v(734)
  wire P7xhu6;  // ../RTL/cortexm0ds_logic.v(266)
  wire P7xow6;  // ../RTL/cortexm0ds_logic.v(1290)
  wire P82ju6;  // ../RTL/cortexm0ds_logic.v(815)
  wire P83iu6;  // ../RTL/cortexm0ds_logic.v(347)
  wire P83pw6;  // ../RTL/cortexm0ds_logic.v(1371)
  wire P89ju6;  // ../RTL/cortexm0ds_logic.v(908)
  wire P8aiu6;  // ../RTL/cortexm0ds_logic.v(440)
  wire P8apw6;  // ../RTL/cortexm0ds_logic.v(1465)
  wire P8bow6;  // ../RTL/cortexm0ds_logic.v(997)
  wire P8hiu6;  // ../RTL/cortexm0ds_logic.v(534)
  wire P8iow6;  // ../RTL/cortexm0ds_logic.v(1090)
  wire P8oiu6;  // ../RTL/cortexm0ds_logic.v(627)
  wire P8phu6;  // ../RTL/cortexm0ds_logic.v(159)
  wire P8pow6;  // ../RTL/cortexm0ds_logic.v(1184)
  wire P8viu6;  // ../RTL/cortexm0ds_logic.v(721)
  wire P8whu6;  // ../RTL/cortexm0ds_logic.v(253)
  wire P8wow6;  // ../RTL/cortexm0ds_logic.v(1277)
  wire P8xpw6;  // ../RTL/cortexm0ds_logic.v(1612)
  wire P91ju6;  // ../RTL/cortexm0ds_logic.v(802)
  wire P92iu6;  // ../RTL/cortexm0ds_logic.v(334)
  wire P92pw6;  // ../RTL/cortexm0ds_logic.v(1358)
  wire P93qw6;  // ../RTL/cortexm0ds_logic.v(1623)
  wire P98ju6;  // ../RTL/cortexm0ds_logic.v(895)
  wire P99iu6;  // ../RTL/cortexm0ds_logic.v(427)
  wire P99pw6;  // ../RTL/cortexm0ds_logic.v(1452)
  wire P9aow6;  // ../RTL/cortexm0ds_logic.v(984)
  wire P9bax6;  // ../RTL/cortexm0ds_logic.v(1634)
  wire P9giu6;  // ../RTL/cortexm0ds_logic.v(521)
  wire P9hhu6;  // ../RTL/cortexm0ds_logic.v(128)
  wire P9how6;  // ../RTL/cortexm0ds_logic.v(1077)
  wire P9niu6;  // ../RTL/cortexm0ds_logic.v(614)
  wire P9oow6;  // ../RTL/cortexm0ds_logic.v(1171)
  wire P9uiu6;  // ../RTL/cortexm0ds_logic.v(708)
  wire P9vhu6;  // ../RTL/cortexm0ds_logic.v(240)
  wire P9vow6;  // ../RTL/cortexm0ds_logic.v(1264)
  wire Pa0ju6;  // ../RTL/cortexm0ds_logic.v(789)
  wire Pa1iu6;  // ../RTL/cortexm0ds_logic.v(321)
  wire Pa1pw6;  // ../RTL/cortexm0ds_logic.v(1345)
  wire Pa7ju6;  // ../RTL/cortexm0ds_logic.v(882)
  wire Pa8iu6;  // ../RTL/cortexm0ds_logic.v(414)
  wire Pa8pw6;  // ../RTL/cortexm0ds_logic.v(1439)
  wire Pa9ow6;  // ../RTL/cortexm0ds_logic.v(971)
  wire Pafiu6;  // ../RTL/cortexm0ds_logic.v(508)
  wire Pagow6;  // ../RTL/cortexm0ds_logic.v(1064)
  wire Pamiu6;  // ../RTL/cortexm0ds_logic.v(601)
  wire Panow6;  // ../RTL/cortexm0ds_logic.v(1158)
  wire Patiu6;  // ../RTL/cortexm0ds_logic.v(695)
  wire Pauhu6;  // ../RTL/cortexm0ds_logic.v(227)
  wire Pauow6;  // ../RTL/cortexm0ds_logic.v(1251)
  wire Paxpw6;  // ../RTL/cortexm0ds_logic.v(1612)
  wire Pb0iu6;  // ../RTL/cortexm0ds_logic.v(308)
  wire Pb0pw6;  // ../RTL/cortexm0ds_logic.v(1332)
  wire Pb6ju6;  // ../RTL/cortexm0ds_logic.v(869)
  wire Pb7iu6;  // ../RTL/cortexm0ds_logic.v(401)
  wire Pb7pw6;  // ../RTL/cortexm0ds_logic.v(1426)
  wire Pb8ow6;  // ../RTL/cortexm0ds_logic.v(958)
  wire Pbbbx6;  // ../RTL/cortexm0ds_logic.v(1699)
  wire Pbeiu6;  // ../RTL/cortexm0ds_logic.v(495)
  wire Pbfow6;  // ../RTL/cortexm0ds_logic.v(1051)
  wire Pbliu6;  // ../RTL/cortexm0ds_logic.v(588)
  wire Pbmow6;  // ../RTL/cortexm0ds_logic.v(1145)
  wire Pbnax6;  // ../RTL/cortexm0ds_logic.v(1656)
  wire Pbsiu6;  // ../RTL/cortexm0ds_logic.v(682)
  wire Pbthu6;  // ../RTL/cortexm0ds_logic.v(214)
  wire Pbtow6;  // ../RTL/cortexm0ds_logic.v(1238)
  wire Pbziu6;  // ../RTL/cortexm0ds_logic.v(776)
  wire Pc5ju6;  // ../RTL/cortexm0ds_logic.v(856)
  wire Pc6iu6;  // ../RTL/cortexm0ds_logic.v(388)
  wire Pc6pw6;  // ../RTL/cortexm0ds_logic.v(1413)
  wire Pc7ow6;  // ../RTL/cortexm0ds_logic.v(945)
  wire Pcdiu6;  // ../RTL/cortexm0ds_logic.v(482)
  wire Pcdpw6;  // ../RTL/cortexm0ds_logic.v(1506)
  wire Pceow6;  // ../RTL/cortexm0ds_logic.v(1038)
  wire Pckiu6;  // ../RTL/cortexm0ds_logic.v(575)
  wire Pclow6;  // ../RTL/cortexm0ds_logic.v(1132)
  wire Pcriu6;  // ../RTL/cortexm0ds_logic.v(669)
  wire Pcrpw6;  // ../RTL/cortexm0ds_logic.v(1601)
  wire Pcshu6;  // ../RTL/cortexm0ds_logic.v(201)
  wire Pcsow6;  // ../RTL/cortexm0ds_logic.v(1225)
  wire Pcxpw6;  // ../RTL/cortexm0ds_logic.v(1612)
  wire Pcyiu6;  // ../RTL/cortexm0ds_logic.v(763)
  wire Pczax6;  // ../RTL/cortexm0ds_logic.v(1678)
  wire Pczhu6;  // ../RTL/cortexm0ds_logic.v(295)
  wire Pczow6;  // ../RTL/cortexm0ds_logic.v(1319)
  wire Pd4ju6;  // ../RTL/cortexm0ds_logic.v(843)
  wire Pd5iu6;  // ../RTL/cortexm0ds_logic.v(375)
  wire Pd5pw6;  // ../RTL/cortexm0ds_logic.v(1400)
  wire Pd6ow6;  // ../RTL/cortexm0ds_logic.v(932)
  wire Pdbbx6;  // ../RTL/cortexm0ds_logic.v(1700)
  wire Pdciu6;  // ../RTL/cortexm0ds_logic.v(469)
  wire Pdcpw6;  // ../RTL/cortexm0ds_logic.v(1493)
  wire Pddow6;  // ../RTL/cortexm0ds_logic.v(1025)
  wire Pdjiu6;  // ../RTL/cortexm0ds_logic.v(562)
  wire Pdkow6;  // ../RTL/cortexm0ds_logic.v(1119)
  wire Pdmpw6;  // ../RTL/cortexm0ds_logic.v(1592)
  wire Pdqiu6;  // ../RTL/cortexm0ds_logic.v(656)
  wire Pdrhu6;  // ../RTL/cortexm0ds_logic.v(188)
  wire Pdrow6;  // ../RTL/cortexm0ds_logic.v(1212)
  wire Pdxax6;  // ../RTL/cortexm0ds_logic.v(1675)
  wire Pdxiu6;  // ../RTL/cortexm0ds_logic.v(750)
  wire Pdyax6;  // ../RTL/cortexm0ds_logic.v(1676)
  wire Pdyhu6;  // ../RTL/cortexm0ds_logic.v(282)
  wire Pdyow6;  // ../RTL/cortexm0ds_logic.v(1306)
  wire Pe3ju6;  // ../RTL/cortexm0ds_logic.v(830)
  wire Pe4iu6;  // ../RTL/cortexm0ds_logic.v(362)
  wire Pe4pw6;  // ../RTL/cortexm0ds_logic.v(1387)
  wire Pe5bx6;  // ../RTL/cortexm0ds_logic.v(1689)
  wire Pe7ax6;  // ../RTL/cortexm0ds_logic.v(1626)
  wire Pe9bx6;  // ../RTL/cortexm0ds_logic.v(1696)
  wire Peaju6;  // ../RTL/cortexm0ds_logic.v(924)
  wire Pebiu6;  // ../RTL/cortexm0ds_logic.v(456)
  wire Pebpw6;  // ../RTL/cortexm0ds_logic.v(1480)
  wire Pecow6;  // ../RTL/cortexm0ds_logic.v(1012)
  wire Peeax6;  // ../RTL/cortexm0ds_logic.v(1640)
  wire Peiiu6;  // ../RTL/cortexm0ds_logic.v(549)
  wire Pejbx6;  // ../RTL/cortexm0ds_logic.v(1714)
  wire Pejow6;  // ../RTL/cortexm0ds_logic.v(1106)
  wire Pepiu6;  // ../RTL/cortexm0ds_logic.v(643)
  wire Peqhu6;  // ../RTL/cortexm0ds_logic.v(175)
  wire Peqow6;  // ../RTL/cortexm0ds_logic.v(1199)
  wire Pewiu6;  // ../RTL/cortexm0ds_logic.v(737)
  wire Pexhu6;  // ../RTL/cortexm0ds_logic.v(269)
  wire Pexow6;  // ../RTL/cortexm0ds_logic.v(1293)
  wire Pexpw6;  // ../RTL/cortexm0ds_logic.v(1612)
  wire Pf2ju6;  // ../RTL/cortexm0ds_logic.v(817)
  wire Pf3iu6;  // ../RTL/cortexm0ds_logic.v(349)
  wire Pf3pw6;  // ../RTL/cortexm0ds_logic.v(1374)
  wire Pf9ju6;  // ../RTL/cortexm0ds_logic.v(911)
  wire Pfaiu6;  // ../RTL/cortexm0ds_logic.v(443)
  wire Pfapw6;  // ../RTL/cortexm0ds_logic.v(1467)
  wire Pfbow6;  // ../RTL/cortexm0ds_logic.v(999)
  wire Pfhiu6;  // ../RTL/cortexm0ds_logic.v(536)
  wire Pfiow6;  // ../RTL/cortexm0ds_logic.v(1093)
  wire Pfoiu6;  // ../RTL/cortexm0ds_logic.v(630)
  wire Pfphu6;  // ../RTL/cortexm0ds_logic.v(162)
  wire Pfpow6;  // ../RTL/cortexm0ds_logic.v(1186)
  wire Pfviu6;  // ../RTL/cortexm0ds_logic.v(724)
  wire Pfwhu6;  // ../RTL/cortexm0ds_logic.v(256)
  wire Pfwow6;  // ../RTL/cortexm0ds_logic.v(1280)
  wire Pg1ju6;  // ../RTL/cortexm0ds_logic.v(804)
  wire Pg2iu6;  // ../RTL/cortexm0ds_logic.v(336)
  wire Pg2pw6;  // ../RTL/cortexm0ds_logic.v(1361)
  wire Pg3qw6;  // ../RTL/cortexm0ds_logic.v(1623)
  wire Pg8ju6;  // ../RTL/cortexm0ds_logic.v(898)
  wire Pg9iu6;  // ../RTL/cortexm0ds_logic.v(430)
  wire Pg9pw6;  // ../RTL/cortexm0ds_logic.v(1454)
  wire Pgaow6;  // ../RTL/cortexm0ds_logic.v(986)
  wire Pggiu6;  // ../RTL/cortexm0ds_logic.v(523)
  wire Pghow6;  // ../RTL/cortexm0ds_logic.v(1080)
  wire Pgjbx6;  // ../RTL/cortexm0ds_logic.v(1715)
  wire Pgniu6;  // ../RTL/cortexm0ds_logic.v(617)
  wire Pgohu6;  // ../RTL/cortexm0ds_logic.v(149)
  wire Pgoow6;  // ../RTL/cortexm0ds_logic.v(1173)
  wire Pguiu6;  // ../RTL/cortexm0ds_logic.v(711)
  wire Pgvhu6;  // ../RTL/cortexm0ds_logic.v(243)
  wire Pgvow6;  // ../RTL/cortexm0ds_logic.v(1267)
  wire Ph0ju6;  // ../RTL/cortexm0ds_logic.v(791)
  wire Ph1iu6;  // ../RTL/cortexm0ds_logic.v(323)
  wire Ph1pw6;  // ../RTL/cortexm0ds_logic.v(1348)
  wire Ph7ju6;  // ../RTL/cortexm0ds_logic.v(885)
  wire Ph8iu6;  // ../RTL/cortexm0ds_logic.v(417)
  wire Ph8pw6;  // ../RTL/cortexm0ds_logic.v(1441)
  wire Ph9ow6;  // ../RTL/cortexm0ds_logic.v(973)
  wire Phcax6;  // ../RTL/cortexm0ds_logic.v(1636)
  wire Phfiu6;  // ../RTL/cortexm0ds_logic.v(510)
  wire Phgow6;  // ../RTL/cortexm0ds_logic.v(1067)
  wire Phmiu6;  // ../RTL/cortexm0ds_logic.v(604)
  wire Phnow6;  // ../RTL/cortexm0ds_logic.v(1160)
  wire Phtiu6;  // ../RTL/cortexm0ds_logic.v(698)
  wire Phuhu6;  // ../RTL/cortexm0ds_logic.v(230)
  wire Phuow6;  // ../RTL/cortexm0ds_logic.v(1254)
  wire Pi0iu6;  // ../RTL/cortexm0ds_logic.v(310)
  wire Pi0pw6;  // ../RTL/cortexm0ds_logic.v(1335)
  wire Pi6ju6;  // ../RTL/cortexm0ds_logic.v(872)
  wire Pi7iu6;  // ../RTL/cortexm0ds_logic.v(404)
  wire Pi7pw6;  // ../RTL/cortexm0ds_logic.v(1428)
  wire Pi8ow6;  // ../RTL/cortexm0ds_logic.v(960)
  wire Pieiu6;  // ../RTL/cortexm0ds_logic.v(497)
  wire Pifax6;  // ../RTL/cortexm0ds_logic.v(1642)
  wire Pifow6;  // ../RTL/cortexm0ds_logic.v(1054)
  wire Piliu6;  // ../RTL/cortexm0ds_logic.v(591)
  wire Pimow6;  // ../RTL/cortexm0ds_logic.v(1147)
  wire Pinhu6;  // ../RTL/cortexm0ds_logic.v(145)
  wire Pisiu6;  // ../RTL/cortexm0ds_logic.v(685)
  wire Pithu6;  // ../RTL/cortexm0ds_logic.v(217)
  wire Pitow6;  // ../RTL/cortexm0ds_logic.v(1241)
  wire Piziu6;  // ../RTL/cortexm0ds_logic.v(778)
  wire Pj5ju6;  // ../RTL/cortexm0ds_logic.v(859)
  wire Pj6iu6;  // ../RTL/cortexm0ds_logic.v(391)
  wire Pj6pw6;  // ../RTL/cortexm0ds_logic.v(1415)
  wire Pj7ow6;  // ../RTL/cortexm0ds_logic.v(947)
  wire Pjdiu6;  // ../RTL/cortexm0ds_logic.v(484)
  wire Pjdpw6;  // ../RTL/cortexm0ds_logic.v(1509)
  wire Pjeow6;  // ../RTL/cortexm0ds_logic.v(1041)
  wire Pjgbx6;  // ../RTL/cortexm0ds_logic.v(1709)
  wire Pjkiu6;  // ../RTL/cortexm0ds_logic.v(578)
  wire Pjlow6;  // ../RTL/cortexm0ds_logic.v(1134)
  wire Pjmhu6;  // ../RTL/cortexm0ds_logic.v(142)
  wire Pjriu6;  // ../RTL/cortexm0ds_logic.v(672)
  wire Pjshu6;  // ../RTL/cortexm0ds_logic.v(204)
  wire Pjsow6;  // ../RTL/cortexm0ds_logic.v(1228)
  wire Pjyiu6;  // ../RTL/cortexm0ds_logic.v(765)
  wire Pjzhu6;  // ../RTL/cortexm0ds_logic.v(297)
  wire Pjzow6;  // ../RTL/cortexm0ds_logic.v(1322)
  wire Pk4ju6;  // ../RTL/cortexm0ds_logic.v(846)
  wire Pk5iu6;  // ../RTL/cortexm0ds_logic.v(378)
  wire Pk5pw6;  // ../RTL/cortexm0ds_logic.v(1402)
  wire Pk6ow6;  // ../RTL/cortexm0ds_logic.v(934)
  wire Pkciu6;  // ../RTL/cortexm0ds_logic.v(471)
  wire Pkcpw6;  // ../RTL/cortexm0ds_logic.v(1496)
  wire Pkdow6;  // ../RTL/cortexm0ds_logic.v(1028)
  wire Pkjiu6;  // ../RTL/cortexm0ds_logic.v(565)
  wire Pkkbx6;  // ../RTL/cortexm0ds_logic.v(1717)
  wire Pkkow6;  // ../RTL/cortexm0ds_logic.v(1121)
  wire Pkqiu6;  // ../RTL/cortexm0ds_logic.v(659)
  wire Pkrhu6;  // ../RTL/cortexm0ds_logic.v(191)
  wire Pkrow6;  // ../RTL/cortexm0ds_logic.v(1215)
  wire Pkxiu6;  // ../RTL/cortexm0ds_logic.v(752)
  wire Pkyhu6;  // ../RTL/cortexm0ds_logic.v(284)
  wire Pkyow6;  // ../RTL/cortexm0ds_logic.v(1309)
  wire Pl3ju6;  // ../RTL/cortexm0ds_logic.v(833)
  wire Pl4iu6;  // ../RTL/cortexm0ds_logic.v(365)
  wire Pl4pw6;  // ../RTL/cortexm0ds_logic.v(1389)
  wire Plaju6;  // ../RTL/cortexm0ds_logic.v(926)
  wire Plbiu6;  // ../RTL/cortexm0ds_logic.v(458)
  wire Plbpw6;  // ../RTL/cortexm0ds_logic.v(1483)
  wire Plcow6;  // ../RTL/cortexm0ds_logic.v(1015)
  wire Pliiu6;  // ../RTL/cortexm0ds_logic.v(552)
  wire Pljow6;  // ../RTL/cortexm0ds_logic.v(1108)
  wire Plpiu6;  // ../RTL/cortexm0ds_logic.v(646)
  wire Plqhu6;  // ../RTL/cortexm0ds_logic.v(178)
  wire Plqow6;  // ../RTL/cortexm0ds_logic.v(1202)
  wire Plwiu6;  // ../RTL/cortexm0ds_logic.v(739)
  wire Plxhu6;  // ../RTL/cortexm0ds_logic.v(271)
  wire Plxow6;  // ../RTL/cortexm0ds_logic.v(1296)
  wire Plypw6;  // ../RTL/cortexm0ds_logic.v(1614)
  wire Pm2ju6;  // ../RTL/cortexm0ds_logic.v(820)
  wire Pm3iu6;  // ../RTL/cortexm0ds_logic.v(352)
  wire Pm3pw6;  // ../RTL/cortexm0ds_logic.v(1376)
  wire Pm9ju6;  // ../RTL/cortexm0ds_logic.v(913)
  wire Pmaiu6;  // ../RTL/cortexm0ds_logic.v(445)
  wire Pmapw6;  // ../RTL/cortexm0ds_logic.v(1470)
  wire Pmbow6;  // ../RTL/cortexm0ds_logic.v(1002)
  wire Pmhiu6;  // ../RTL/cortexm0ds_logic.v(539)
  wire Pmiow6;  // ../RTL/cortexm0ds_logic.v(1095)
  wire Pmlhu6;  // ../RTL/cortexm0ds_logic.v(140)
  wire Pmlpw6;  // ../RTL/cortexm0ds_logic.v(1591)
  wire Pmoiu6;  // ../RTL/cortexm0ds_logic.v(633)
  wire Pmphu6;  // ../RTL/cortexm0ds_logic.v(165)
  wire Pmpow6;  // ../RTL/cortexm0ds_logic.v(1189)
  wire Pmviu6;  // ../RTL/cortexm0ds_logic.v(726)
  wire Pmwhu6;  // ../RTL/cortexm0ds_logic.v(258)
  wire Pmwow6;  // ../RTL/cortexm0ds_logic.v(1283)
  wire Pn1ju6;  // ../RTL/cortexm0ds_logic.v(807)
  wire Pn2iu6;  // ../RTL/cortexm0ds_logic.v(339)
  wire Pn2pw6;  // ../RTL/cortexm0ds_logic.v(1363)
  wire Pn8ju6;  // ../RTL/cortexm0ds_logic.v(900)
  wire Pn9iu6;  // ../RTL/cortexm0ds_logic.v(432)
  wire Pn9pw6;  // ../RTL/cortexm0ds_logic.v(1457)
  wire Pnaow6;  // ../RTL/cortexm0ds_logic.v(989)
  wire Pndhu6;  // ../RTL/cortexm0ds_logic.v(120)
  wire Pngiu6;  // ../RTL/cortexm0ds_logic.v(526)
  wire Pnhow6;  // ../RTL/cortexm0ds_logic.v(1082)
  wire Pnniu6;  // ../RTL/cortexm0ds_logic.v(620)
  wire Pnohu6;  // ../RTL/cortexm0ds_logic.v(152)
  wire Pnoow6;  // ../RTL/cortexm0ds_logic.v(1176)
  wire Pnuiu6;  // ../RTL/cortexm0ds_logic.v(713)
  wire Pnvhu6;  // ../RTL/cortexm0ds_logic.v(245)
  wire Pnvow6;  // ../RTL/cortexm0ds_logic.v(1270)
  wire Po0ju6;  // ../RTL/cortexm0ds_logic.v(794)
  wire Po1iu6;  // ../RTL/cortexm0ds_logic.v(326)
  wire Po1pw6;  // ../RTL/cortexm0ds_logic.v(1350)
  wire Po7ju6;  // ../RTL/cortexm0ds_logic.v(887)
  wire Po8iu6;  // ../RTL/cortexm0ds_logic.v(419)
  wire Po8pw6;  // ../RTL/cortexm0ds_logic.v(1444)
  wire Po9ow6;  // ../RTL/cortexm0ds_logic.v(976)
  wire Pofiu6;  // ../RTL/cortexm0ds_logic.v(513)
  wire Pogow6;  // ../RTL/cortexm0ds_logic.v(1069)
  wire Pomiu6;  // ../RTL/cortexm0ds_logic.v(607)
  wire Ponow6;  // ../RTL/cortexm0ds_logic.v(1163)
  wire Potiu6;  // ../RTL/cortexm0ds_logic.v(700)
  wire Pouhu6;  // ../RTL/cortexm0ds_logic.v(232)
  wire Pouow6;  // ../RTL/cortexm0ds_logic.v(1257)
  wire Pp0iu6;  // ../RTL/cortexm0ds_logic.v(313)
  wire Pp0pw6;  // ../RTL/cortexm0ds_logic.v(1337)
  wire Pp6ju6;  // ../RTL/cortexm0ds_logic.v(874)
  wire Pp7iu6;  // ../RTL/cortexm0ds_logic.v(406)
  wire Pp7pw6;  // ../RTL/cortexm0ds_logic.v(1431)
  wire Pp8ow6;  // ../RTL/cortexm0ds_logic.v(963)
  wire Ppeiu6;  // ../RTL/cortexm0ds_logic.v(500)
  wire Ppfow6;  // ../RTL/cortexm0ds_logic.v(1056)
  wire Ppliu6;  // ../RTL/cortexm0ds_logic.v(594)
  wire Ppmow6;  // ../RTL/cortexm0ds_logic.v(1150)
  wire Ppsiu6;  // ../RTL/cortexm0ds_logic.v(687)
  wire Ppthu6;  // ../RTL/cortexm0ds_logic.v(219)
  wire Pptow6;  // ../RTL/cortexm0ds_logic.v(1244)
  wire Ppziu6;  // ../RTL/cortexm0ds_logic.v(781)
  wire Pq5ju6;  // ../RTL/cortexm0ds_logic.v(861)
  wire Pq6iu6;  // ../RTL/cortexm0ds_logic.v(393)
  wire Pq6pw6;  // ../RTL/cortexm0ds_logic.v(1418)
  wire Pq7ow6;  // ../RTL/cortexm0ds_logic.v(950)
  wire Pqdiu6;  // ../RTL/cortexm0ds_logic.v(487)
  wire Pqdpw6;  // ../RTL/cortexm0ds_logic.v(1511)
  wire Pqeow6;  // ../RTL/cortexm0ds_logic.v(1043)
  wire Pqkiu6;  // ../RTL/cortexm0ds_logic.v(581)
  wire Pqlow6;  // ../RTL/cortexm0ds_logic.v(1137)
  wire Pqrax6;  // ../RTL/cortexm0ds_logic.v(1664)
  wire Pqriu6;  // ../RTL/cortexm0ds_logic.v(674)
  wire Pqshu6;  // ../RTL/cortexm0ds_logic.v(206)
  wire Pqsow6;  // ../RTL/cortexm0ds_logic.v(1231)
  wire Pqyiu6;  // ../RTL/cortexm0ds_logic.v(768)
  wire Pqzhu6;  // ../RTL/cortexm0ds_logic.v(300)
  wire Pqzow6;  // ../RTL/cortexm0ds_logic.v(1324)
  wire Pr4ju6;  // ../RTL/cortexm0ds_logic.v(848)
  wire Pr5iu6;  // ../RTL/cortexm0ds_logic.v(380)
  wire Pr5pw6;  // ../RTL/cortexm0ds_logic.v(1405)
  wire Pr6ow6;  // ../RTL/cortexm0ds_logic.v(937)
  wire Prciu6;  // ../RTL/cortexm0ds_logic.v(474)
  wire Prcpw6;  // ../RTL/cortexm0ds_logic.v(1498)
  wire Prdow6;  // ../RTL/cortexm0ds_logic.v(1030)
  wire Prjiu6;  // ../RTL/cortexm0ds_logic.v(568)
  wire Prkow6;  // ../RTL/cortexm0ds_logic.v(1124)
  wire Propw6;  // ../RTL/cortexm0ds_logic.v(1597)
  wire Prqiu6;  // ../RTL/cortexm0ds_logic.v(661)
  wire Prrhu6;  // ../RTL/cortexm0ds_logic.v(193)
  wire Prrow6;  // ../RTL/cortexm0ds_logic.v(1218)
  wire Prxiu6;  // ../RTL/cortexm0ds_logic.v(755)
  wire Pryhu6;  // ../RTL/cortexm0ds_logic.v(287)
  wire Pryow6;  // ../RTL/cortexm0ds_logic.v(1311)
  wire Ps3ju6;  // ../RTL/cortexm0ds_logic.v(835)
  wire Ps4iu6;  // ../RTL/cortexm0ds_logic.v(367)
  wire Ps4pw6;  // ../RTL/cortexm0ds_logic.v(1392)
  wire Psaju6;  // ../RTL/cortexm0ds_logic.v(929)
  wire Psbiu6;  // ../RTL/cortexm0ds_logic.v(461)
  wire Psbpw6;  // ../RTL/cortexm0ds_logic.v(1485)
  wire Pscow6;  // ../RTL/cortexm0ds_logic.v(1017)
  wire Psiiu6;  // ../RTL/cortexm0ds_logic.v(555)
  wire Psjow6;  // ../RTL/cortexm0ds_logic.v(1111)
  wire Pspiu6;  // ../RTL/cortexm0ds_logic.v(648)
  wire Psqhu6;  // ../RTL/cortexm0ds_logic.v(180)
  wire Psqow6;  // ../RTL/cortexm0ds_logic.v(1205)
  wire Pswiu6;  // ../RTL/cortexm0ds_logic.v(742)
  wire Psxhu6;  // ../RTL/cortexm0ds_logic.v(274)
  wire Psxow6;  // ../RTL/cortexm0ds_logic.v(1298)
  wire Pt2ju6;  // ../RTL/cortexm0ds_logic.v(822)
  wire Pt3iu6;  // ../RTL/cortexm0ds_logic.v(354)
  wire Pt3pw6;  // ../RTL/cortexm0ds_logic.v(1379)
  wire Pt7ax6;  // ../RTL/cortexm0ds_logic.v(1627)
  wire Pt9ju6;  // ../RTL/cortexm0ds_logic.v(916)
  wire Ptaiu6;  // ../RTL/cortexm0ds_logic.v(448)
  wire Ptapw6;  // ../RTL/cortexm0ds_logic.v(1472)
  wire Ptbow6;  // ../RTL/cortexm0ds_logic.v(1004)
  wire Pthiu6;  // ../RTL/cortexm0ds_logic.v(542)
  wire Ptiow6;  // ../RTL/cortexm0ds_logic.v(1098)
  wire Ptoiu6;  // ../RTL/cortexm0ds_logic.v(635)
  wire Ptphu6;  // ../RTL/cortexm0ds_logic.v(167)
  wire Ptpow6;  // ../RTL/cortexm0ds_logic.v(1192)
  wire Ptviu6;  // ../RTL/cortexm0ds_logic.v(729)
  wire Ptwhu6;  // ../RTL/cortexm0ds_logic.v(261)
  wire Ptwow6;  // ../RTL/cortexm0ds_logic.v(1285)
  wire Pu1ju6;  // ../RTL/cortexm0ds_logic.v(809)
  wire Pu2iu6;  // ../RTL/cortexm0ds_logic.v(341)
  wire Pu2pw6;  // ../RTL/cortexm0ds_logic.v(1366)
  wire Pu8ju6;  // ../RTL/cortexm0ds_logic.v(903)
  wire Pu9iu6;  // ../RTL/cortexm0ds_logic.v(435)
  wire Pu9pw6;  // ../RTL/cortexm0ds_logic.v(1459)
  wire Puaow6;  // ../RTL/cortexm0ds_logic.v(991)
  wire Pugiu6;  // ../RTL/cortexm0ds_logic.v(529)
  wire Puhow6;  // ../RTL/cortexm0ds_logic.v(1085)
  wire Punhu6;  // ../RTL/cortexm0ds_logic.v(145)
  wire Puniu6;  // ../RTL/cortexm0ds_logic.v(622)
  wire Puohu6;  // ../RTL/cortexm0ds_logic.v(154)
  wire Puoow6;  // ../RTL/cortexm0ds_logic.v(1179)
  wire Puuiu6;  // ../RTL/cortexm0ds_logic.v(716)
  wire Puvhu6;  // ../RTL/cortexm0ds_logic.v(248)
  wire Puvow6;  // ../RTL/cortexm0ds_logic.v(1272)
  wire Puwpw6;  // ../RTL/cortexm0ds_logic.v(1611)
  wire Pv0bx6;  // ../RTL/cortexm0ds_logic.v(1681)
  wire Pv0ju6;  // ../RTL/cortexm0ds_logic.v(796)
  wire Pv1iu6;  // ../RTL/cortexm0ds_logic.v(328)
  wire Pv1pw6;  // ../RTL/cortexm0ds_logic.v(1353)
  wire Pv7ju6;  // ../RTL/cortexm0ds_logic.v(890)
  wire Pv8iu6;  // ../RTL/cortexm0ds_logic.v(422)
  wire Pv8pw6;  // ../RTL/cortexm0ds_logic.v(1446)
  wire Pv9ax6;  // ../RTL/cortexm0ds_logic.v(1631)
  wire Pv9ow6;  // ../RTL/cortexm0ds_logic.v(978)
  wire Pvfiu6;  // ../RTL/cortexm0ds_logic.v(516)
  wire Pvgow6;  // ../RTL/cortexm0ds_logic.v(1072)
  wire Pvmiu6;  // ../RTL/cortexm0ds_logic.v(609)
  wire Pvnow6;  // ../RTL/cortexm0ds_logic.v(1166)
  wire Pvtiu6;  // ../RTL/cortexm0ds_logic.v(703)
  wire Pvuhu6;  // ../RTL/cortexm0ds_logic.v(235)
  wire Pvuow6;  // ../RTL/cortexm0ds_logic.v(1259)
  wire Pw0iu6;  // ../RTL/cortexm0ds_logic.v(315)
  wire Pw0pw6;  // ../RTL/cortexm0ds_logic.v(1340)
  wire Pw6ju6;  // ../RTL/cortexm0ds_logic.v(877)
  wire Pw7iu6;  // ../RTL/cortexm0ds_logic.v(409)
  wire Pw7pw6;  // ../RTL/cortexm0ds_logic.v(1433)
  wire Pw8ow6;  // ../RTL/cortexm0ds_logic.v(965)
  wire Pweiu6;  // ../RTL/cortexm0ds_logic.v(503)
  wire Pwfow6;  // ../RTL/cortexm0ds_logic.v(1059)
  wire Pwkax6;  // ../RTL/cortexm0ds_logic.v(1652)
  wire Pwliu6;  // ../RTL/cortexm0ds_logic.v(596)
  wire Pwmow6;  // ../RTL/cortexm0ds_logic.v(1153)
  wire Pwsiu6;  // ../RTL/cortexm0ds_logic.v(690)
  wire Pwthu6;  // ../RTL/cortexm0ds_logic.v(222)
  wire Pwtow6;  // ../RTL/cortexm0ds_logic.v(1246)
  wire Pwziu6;  // ../RTL/cortexm0ds_logic.v(783)
  wire Px5ju6;  // ../RTL/cortexm0ds_logic.v(864)
  wire Px6iu6;  // ../RTL/cortexm0ds_logic.v(396)
  wire Px6pw6;  // ../RTL/cortexm0ds_logic.v(1420)
  wire Px7ow6;  // ../RTL/cortexm0ds_logic.v(952)
  wire Pxdiu6;  // ../RTL/cortexm0ds_logic.v(490)
  wire Pxdpw6;  // ../RTL/cortexm0ds_logic.v(1514)
  wire Pxeow6;  // ../RTL/cortexm0ds_logic.v(1046)
  wire Pxkiu6;  // ../RTL/cortexm0ds_logic.v(583)
  wire Pxlow6;  // ../RTL/cortexm0ds_logic.v(1140)
  wire Pxriu6;  // ../RTL/cortexm0ds_logic.v(677)
  wire Pxshu6;  // ../RTL/cortexm0ds_logic.v(209)
  wire Pxsow6;  // ../RTL/cortexm0ds_logic.v(1233)
  wire Pxvax6;  // ../RTL/cortexm0ds_logic.v(1672)
  wire Pxyiu6;  // ../RTL/cortexm0ds_logic.v(770)
  wire Pxzhu6;  // ../RTL/cortexm0ds_logic.v(302)
  wire Pxzow6;  // ../RTL/cortexm0ds_logic.v(1327)
  wire Py4ju6;  // ../RTL/cortexm0ds_logic.v(851)
  wire Py5iu6;  // ../RTL/cortexm0ds_logic.v(383)
  wire Py5pw6;  // ../RTL/cortexm0ds_logic.v(1407)
  wire Py6ow6;  // ../RTL/cortexm0ds_logic.v(939)
  wire Pyciu6;  // ../RTL/cortexm0ds_logic.v(477)
  wire Pycpw6;  // ../RTL/cortexm0ds_logic.v(1501)
  wire Pydow6;  // ../RTL/cortexm0ds_logic.v(1033)
  wire Pyjiu6;  // ../RTL/cortexm0ds_logic.v(570)
  wire Pykow6;  // ../RTL/cortexm0ds_logic.v(1127)
  wire Pyqiu6;  // ../RTL/cortexm0ds_logic.v(664)
  wire Pyrhu6;  // ../RTL/cortexm0ds_logic.v(196)
  wire Pyrow6;  // ../RTL/cortexm0ds_logic.v(1220)
  wire Pyxiu6;  // ../RTL/cortexm0ds_logic.v(757)
  wire Pyyhu6;  // ../RTL/cortexm0ds_logic.v(289)
  wire Pyyow6;  // ../RTL/cortexm0ds_logic.v(1314)
  wire Pz3ju6;  // ../RTL/cortexm0ds_logic.v(838)
  wire Pz4iu6;  // ../RTL/cortexm0ds_logic.v(370)
  wire Pz4pw6;  // ../RTL/cortexm0ds_logic.v(1394)
  wire Pz9bx6;  // ../RTL/cortexm0ds_logic.v(1697)
  wire Pzbiu6;  // ../RTL/cortexm0ds_logic.v(464)
  wire Pzbpw6;  // ../RTL/cortexm0ds_logic.v(1488)
  wire Pzcow6;  // ../RTL/cortexm0ds_logic.v(1020)
  wire Pzibx6;  // ../RTL/cortexm0ds_logic.v(1714)
  wire Pziiu6;  // ../RTL/cortexm0ds_logic.v(557)
  wire Pzjow6;  // ../RTL/cortexm0ds_logic.v(1114)
  wire Pzkpw6;  // ../RTL/cortexm0ds_logic.v(1589)
  wire Pzpiu6;  // ../RTL/cortexm0ds_logic.v(651)
  wire Pzqhu6;  // ../RTL/cortexm0ds_logic.v(183)
  wire Pzqow6;  // ../RTL/cortexm0ds_logic.v(1207)
  wire Pzwiu6;  // ../RTL/cortexm0ds_logic.v(744)
  wire Pzxhu6;  // ../RTL/cortexm0ds_logic.v(276)
  wire Pzxow6;  // ../RTL/cortexm0ds_logic.v(1301)
  wire Q00ju6;  // ../RTL/cortexm0ds_logic.v(785)
  wire Q01iu6;  // ../RTL/cortexm0ds_logic.v(317)
  wire Q01pw6;  // ../RTL/cortexm0ds_logic.v(1341)
  wire Q01qw6;  // ../RTL/cortexm0ds_logic.v(1619)
  wire Q07ju6;  // ../RTL/cortexm0ds_logic.v(879)
  wire Q08iu6;  // ../RTL/cortexm0ds_logic.v(411)
  wire Q08pw6;  // ../RTL/cortexm0ds_logic.v(1435)
  wire Q09ow6;  // ../RTL/cortexm0ds_logic.v(967)
  wire Q0fiu6;  // ../RTL/cortexm0ds_logic.v(504)
  wire Q0gow6;  // ../RTL/cortexm0ds_logic.v(1061)
  wire Q0miu6;  // ../RTL/cortexm0ds_logic.v(598)
  wire Q0now6;  // ../RTL/cortexm0ds_logic.v(1154)
  wire Q0tiu6;  // ../RTL/cortexm0ds_logic.v(691)
  wire Q0uhu6;  // ../RTL/cortexm0ds_logic.v(223)
  wire Q0uow6;  // ../RTL/cortexm0ds_logic.v(1248)
  wire Q10iu6;  // ../RTL/cortexm0ds_logic.v(304)
  wire Q10pw6;  // ../RTL/cortexm0ds_logic.v(1328)
  wire Q16ju6;  // ../RTL/cortexm0ds_logic.v(866)
  wire Q17iu6;  // ../RTL/cortexm0ds_logic.v(398)
  wire Q17pw6;  // ../RTL/cortexm0ds_logic.v(1422)
  wire Q18ow6;  // ../RTL/cortexm0ds_logic.v(954)
  wire Q1eiu6;  // ../RTL/cortexm0ds_logic.v(491)
  wire Q1epw6;  // ../RTL/cortexm0ds_logic.v(1516)
  wire Q1fow6;  // ../RTL/cortexm0ds_logic.v(1048)
  wire Q1hbx6;  // ../RTL/cortexm0ds_logic.v(1710)
  wire Q1liu6;  // ../RTL/cortexm0ds_logic.v(585)
  wire Q1mow6;  // ../RTL/cortexm0ds_logic.v(1141)
  wire Q1siu6;  // ../RTL/cortexm0ds_logic.v(678)
  wire Q1thu6;  // ../RTL/cortexm0ds_logic.v(210)
  wire Q1tow6;  // ../RTL/cortexm0ds_logic.v(1235)
  wire Q1ziu6;  // ../RTL/cortexm0ds_logic.v(772)
  wire Q25ju6;  // ../RTL/cortexm0ds_logic.v(853)
  wire Q26iu6;  // ../RTL/cortexm0ds_logic.v(385)
  wire Q26pw6;  // ../RTL/cortexm0ds_logic.v(1409)
  wire Q27ow6;  // ../RTL/cortexm0ds_logic.v(941)
  wire Q2diu6;  // ../RTL/cortexm0ds_logic.v(478)
  wire Q2dpw6;  // ../RTL/cortexm0ds_logic.v(1503)
  wire Q2eow6;  // ../RTL/cortexm0ds_logic.v(1035)
  wire Q2gax6;  // ../RTL/cortexm0ds_logic.v(1643)
  wire Q2ibx6;  // ../RTL/cortexm0ds_logic.v(1712)
  wire Q2kiu6;  // ../RTL/cortexm0ds_logic.v(572)
  wire Q2low6;  // ../RTL/cortexm0ds_logic.v(1128)
  wire Q2riu6;  // ../RTL/cortexm0ds_logic.v(665)
  wire Q2shu6;  // ../RTL/cortexm0ds_logic.v(197)
  wire Q2sow6;  // ../RTL/cortexm0ds_logic.v(1222)
  wire Q2yiu6;  // ../RTL/cortexm0ds_logic.v(759)
  wire Q2zhu6;  // ../RTL/cortexm0ds_logic.v(291)
  wire Q2zow6;  // ../RTL/cortexm0ds_logic.v(1315)
  wire Q34ju6;  // ../RTL/cortexm0ds_logic.v(840)
  wire Q35iu6;  // ../RTL/cortexm0ds_logic.v(372)
  wire Q35pw6;  // ../RTL/cortexm0ds_logic.v(1396)
  wire Q3ciu6;  // ../RTL/cortexm0ds_logic.v(465)
  wire Q3cpw6;  // ../RTL/cortexm0ds_logic.v(1490)
  wire Q3dow6;  // ../RTL/cortexm0ds_logic.v(1022)
  wire Q3jiu6;  // ../RTL/cortexm0ds_logic.v(559)
  wire Q3kow6;  // ../RTL/cortexm0ds_logic.v(1115)
  wire Q3qiu6;  // ../RTL/cortexm0ds_logic.v(652)
  wire Q3rhu6;  // ../RTL/cortexm0ds_logic.v(184)
  wire Q3row6;  // ../RTL/cortexm0ds_logic.v(1209)
  wire Q3xiu6;  // ../RTL/cortexm0ds_logic.v(746)
  wire Q3yhu6;  // ../RTL/cortexm0ds_logic.v(278)
  wire Q3yow6;  // ../RTL/cortexm0ds_logic.v(1302)
  wire Q43ju6;  // ../RTL/cortexm0ds_logic.v(827)
  wire Q44iu6;  // ../RTL/cortexm0ds_logic.v(359)
  wire Q44pw6;  // ../RTL/cortexm0ds_logic.v(1383)
  wire Q4aju6;  // ../RTL/cortexm0ds_logic.v(920)
  wire Q4biu6;  // ../RTL/cortexm0ds_logic.v(452)
  wire Q4bpw6;  // ../RTL/cortexm0ds_logic.v(1477)
  wire Q4cow6;  // ../RTL/cortexm0ds_logic.v(1009)
  wire Q4dbx6;  // ../RTL/cortexm0ds_logic.v(1703)
  wire Q4iiu6;  // ../RTL/cortexm0ds_logic.v(546)
  wire Q4jow6;  // ../RTL/cortexm0ds_logic.v(1102)
  wire Q4lhu6;  // ../RTL/cortexm0ds_logic.v(138)
  wire Q4piu6;  // ../RTL/cortexm0ds_logic.v(639)
  wire Q4qhu6;  // ../RTL/cortexm0ds_logic.v(171)
  wire Q4qow6;  // ../RTL/cortexm0ds_logic.v(1196)
  wire Q4wiu6;  // ../RTL/cortexm0ds_logic.v(733)
  wire Q4xhu6;  // ../RTL/cortexm0ds_logic.v(265)
  wire Q4xow6;  // ../RTL/cortexm0ds_logic.v(1289)
  wire Q52ju6;  // ../RTL/cortexm0ds_logic.v(814)
  wire Q53pw6;  // ../RTL/cortexm0ds_logic.v(1370)
  wire Q59ju6;  // ../RTL/cortexm0ds_logic.v(907)
  wire Q5aiu6;  // ../RTL/cortexm0ds_logic.v(439)
  wire Q5apw6;  // ../RTL/cortexm0ds_logic.v(1464)
  wire Q5bow6;  // ../RTL/cortexm0ds_logic.v(996)
  wire Q5hiu6;  // ../RTL/cortexm0ds_logic.v(533)
  wire Q5iow6;  // ../RTL/cortexm0ds_logic.v(1089)
  wire Q5mhu6;  // ../RTL/cortexm0ds_logic.v(141)
  wire Q5oiu6;  // ../RTL/cortexm0ds_logic.v(626)
  wire Q5phu6;  // ../RTL/cortexm0ds_logic.v(158)
  wire Q5pow6;  // ../RTL/cortexm0ds_logic.v(1183)
  wire Q5viu6;  // ../RTL/cortexm0ds_logic.v(720)
  wire Q5whu6;  // ../RTL/cortexm0ds_logic.v(252)
  wire Q5wow6;  // ../RTL/cortexm0ds_logic.v(1276)
  wire Q61ju6;  // ../RTL/cortexm0ds_logic.v(801)
  wire Q62iu6;  // ../RTL/cortexm0ds_logic.v(333)
  wire Q62pw6;  // ../RTL/cortexm0ds_logic.v(1357)
  wire Q68ju6;  // ../RTL/cortexm0ds_logic.v(894)
  wire Q69iu6;  // ../RTL/cortexm0ds_logic.v(426)
  wire Q69pw6;  // ../RTL/cortexm0ds_logic.v(1451)
  wire Q6aow6;  // ../RTL/cortexm0ds_logic.v(983)
  wire Q6fax6;  // ../RTL/cortexm0ds_logic.v(1641)
  wire Q6giu6;  // ../RTL/cortexm0ds_logic.v(520)
  wire Q6how6;  // ../RTL/cortexm0ds_logic.v(1076)
  wire Q6khu6;  // ../RTL/cortexm0ds_logic.v(136)
  wire Q6niu6;  // ../RTL/cortexm0ds_logic.v(613)
  wire Q6oow6;  // ../RTL/cortexm0ds_logic.v(1170)
  wire Q6uiu6;  // ../RTL/cortexm0ds_logic.v(707)
  wire Q6vhu6;  // ../RTL/cortexm0ds_logic.v(239)
  wire Q6vow6;  // ../RTL/cortexm0ds_logic.v(1263)
  wire Q70ju6;  // ../RTL/cortexm0ds_logic.v(788)
  wire Q71iu6;  // ../RTL/cortexm0ds_logic.v(320)
  wire Q71pw6;  // ../RTL/cortexm0ds_logic.v(1344)
  wire Q77ju6;  // ../RTL/cortexm0ds_logic.v(881)
  wire Q78iu6;  // ../RTL/cortexm0ds_logic.v(413)
  wire Q78pw6;  // ../RTL/cortexm0ds_logic.v(1438)
  wire Q79ow6;  // ../RTL/cortexm0ds_logic.v(970)
  wire Q7fiu6;  // ../RTL/cortexm0ds_logic.v(507)
  wire Q7gow6;  // ../RTL/cortexm0ds_logic.v(1063)
  wire Q7miu6;  // ../RTL/cortexm0ds_logic.v(600)
  wire Q7now6;  // ../RTL/cortexm0ds_logic.v(1157)
  wire Q7ohu6;  // ../RTL/cortexm0ds_logic.v(146)
  wire Q7tiu6;  // ../RTL/cortexm0ds_logic.v(694)
  wire Q7uhu6;  // ../RTL/cortexm0ds_logic.v(226)
  wire Q7uow6;  // ../RTL/cortexm0ds_logic.v(1250)
  wire Q80iu6;  // ../RTL/cortexm0ds_logic.v(307)
  wire Q80pw6;  // ../RTL/cortexm0ds_logic.v(1331)
  wire Q86ju6;  // ../RTL/cortexm0ds_logic.v(868)
  wire Q87iu6;  // ../RTL/cortexm0ds_logic.v(400)
  wire Q87pw6;  // ../RTL/cortexm0ds_logic.v(1425)
  wire Q88ow6;  // ../RTL/cortexm0ds_logic.v(957)
  wire Q89bx6;  // ../RTL/cortexm0ds_logic.v(1696)
  wire Q8aax6;  // ../RTL/cortexm0ds_logic.v(1632)
  wire Q8eiu6;  // ../RTL/cortexm0ds_logic.v(494)
  wire Q8fow6;  // ../RTL/cortexm0ds_logic.v(1050)
  wire Q8jhu6;  // ../RTL/cortexm0ds_logic.v(133)
  wire Q8liu6;  // ../RTL/cortexm0ds_logic.v(587)
  wire Q8mow6;  // ../RTL/cortexm0ds_logic.v(1144)
  wire Q8nhu6;  // ../RTL/cortexm0ds_logic.v(144)
  wire Q8siu6;  // ../RTL/cortexm0ds_logic.v(681)
  wire Q8thu6;  // ../RTL/cortexm0ds_logic.v(213)
  wire Q8tow6;  // ../RTL/cortexm0ds_logic.v(1237)
  wire Q8ziu6;  // ../RTL/cortexm0ds_logic.v(775)
  wire Q95ju6;  // ../RTL/cortexm0ds_logic.v(855)
  wire Q96iu6;  // ../RTL/cortexm0ds_logic.v(387)
  wire Q96pw6;  // ../RTL/cortexm0ds_logic.v(1412)
  wire Q97ow6;  // ../RTL/cortexm0ds_logic.v(944)
  wire Q9dax6;  // ../RTL/cortexm0ds_logic.v(1638)
  wire Q9diu6;  // ../RTL/cortexm0ds_logic.v(481)
  wire Q9dpw6;  // ../RTL/cortexm0ds_logic.v(1505)
  wire Q9eow6;  // ../RTL/cortexm0ds_logic.v(1037)
  wire Q9kiu6;  // ../RTL/cortexm0ds_logic.v(574)
  wire Q9low6;  // ../RTL/cortexm0ds_logic.v(1131)
  wire Q9nax6;  // ../RTL/cortexm0ds_logic.v(1656)
  wire Q9riu6;  // ../RTL/cortexm0ds_logic.v(668)
  wire Q9shu6;  // ../RTL/cortexm0ds_logic.v(200)
  wire Q9sow6;  // ../RTL/cortexm0ds_logic.v(1224)
  wire Q9yiu6;  // ../RTL/cortexm0ds_logic.v(762)
  wire Q9zhu6;  // ../RTL/cortexm0ds_logic.v(294)
  wire Q9zow6;  // ../RTL/cortexm0ds_logic.v(1318)
  wire Qa1qw6;  // ../RTL/cortexm0ds_logic.v(1619)
  wire Qa4ju6;  // ../RTL/cortexm0ds_logic.v(842)
  wire Qa5iu6;  // ../RTL/cortexm0ds_logic.v(374)
  wire Qa5pw6;  // ../RTL/cortexm0ds_logic.v(1399)
  wire Qa6ow6;  // ../RTL/cortexm0ds_logic.v(931)
  wire Qaciu6;  // ../RTL/cortexm0ds_logic.v(468)
  wire Qacpw6;  // ../RTL/cortexm0ds_logic.v(1492)
  wire Qadow6;  // ../RTL/cortexm0ds_logic.v(1024)
  wire Qaihu6;  // ../RTL/cortexm0ds_logic.v(130)
  wire Qaipw6;  // ../RTL/cortexm0ds_logic.v(1584)
  wire Qajiu6;  // ../RTL/cortexm0ds_logic.v(561)
  wire Qakbx6;  // ../RTL/cortexm0ds_logic.v(1716)
  wire Qakow6;  // ../RTL/cortexm0ds_logic.v(1118)
  wire Qaqiu6;  // ../RTL/cortexm0ds_logic.v(655)
  wire Qarhu6;  // ../RTL/cortexm0ds_logic.v(187)
  wire Qarow6;  // ../RTL/cortexm0ds_logic.v(1211)
  wire Qaxiu6;  // ../RTL/cortexm0ds_logic.v(749)
  wire Qayhu6;  // ../RTL/cortexm0ds_logic.v(281)
  wire Qayow6;  // ../RTL/cortexm0ds_logic.v(1305)
  wire Qb3ju6;  // ../RTL/cortexm0ds_logic.v(829)
  wire Qb4iu6;  // ../RTL/cortexm0ds_logic.v(361)
  wire Qb4pw6;  // ../RTL/cortexm0ds_logic.v(1386)
  wire Qbaju6;  // ../RTL/cortexm0ds_logic.v(923)
  wire Qbbiu6;  // ../RTL/cortexm0ds_logic.v(455)
  wire Qbbpw6;  // ../RTL/cortexm0ds_logic.v(1479)
  wire Qbcow6;  // ../RTL/cortexm0ds_logic.v(1011)
  wire Qbehu6;  // ../RTL/cortexm0ds_logic.v(121)
  wire Qbiiu6;  // ../RTL/cortexm0ds_logic.v(548)
  wire Qbjow6;  // ../RTL/cortexm0ds_logic.v(1105)
  wire Qbmpw6;  // ../RTL/cortexm0ds_logic.v(1592)
  wire Qbpiu6;  // ../RTL/cortexm0ds_logic.v(642)
  wire Qbqhu6;  // ../RTL/cortexm0ds_logic.v(174)
  wire Qbqow6;  // ../RTL/cortexm0ds_logic.v(1198)
  wire Qbwiu6;  // ../RTL/cortexm0ds_logic.v(736)
  wire Qbxhu6;  // ../RTL/cortexm0ds_logic.v(268)
  wire Qbxow6;  // ../RTL/cortexm0ds_logic.v(1292)
  wire Qc2ju6;  // ../RTL/cortexm0ds_logic.v(816)
  wire Qc3iu6;  // ../RTL/cortexm0ds_logic.v(348)
  wire Qc3pw6;  // ../RTL/cortexm0ds_logic.v(1373)
  wire Qc5bx6;  // ../RTL/cortexm0ds_logic.v(1689)
  wire Qc9ju6;  // ../RTL/cortexm0ds_logic.v(910)
  wire Qcaiu6;  // ../RTL/cortexm0ds_logic.v(442)
  wire Qcapw6;  // ../RTL/cortexm0ds_logic.v(1466)
  wire Qcbow6;  // ../RTL/cortexm0ds_logic.v(998)
  wire Qchiu6;  // ../RTL/cortexm0ds_logic.v(535)
  wire Qciow6;  // ../RTL/cortexm0ds_logic.v(1092)
  wire Qcoiu6;  // ../RTL/cortexm0ds_logic.v(629)
  wire Qcphu6;  // ../RTL/cortexm0ds_logic.v(161)
  wire Qcpow6;  // ../RTL/cortexm0ds_logic.v(1185)
  wire Qcviu6;  // ../RTL/cortexm0ds_logic.v(723)
  wire Qcwhu6;  // ../RTL/cortexm0ds_logic.v(255)
  wire Qcwow6;  // ../RTL/cortexm0ds_logic.v(1279)
  wire Qd1ju6;  // ../RTL/cortexm0ds_logic.v(803)
  wire Qd2iu6;  // ../RTL/cortexm0ds_logic.v(335)
  wire Qd2pw6;  // ../RTL/cortexm0ds_logic.v(1360)
  wire Qd8ju6;  // ../RTL/cortexm0ds_logic.v(897)
  wire Qd9iu6;  // ../RTL/cortexm0ds_logic.v(429)
  wire Qd9pw6;  // ../RTL/cortexm0ds_logic.v(1453)
  wire Qdaow6;  // ../RTL/cortexm0ds_logic.v(985)
  wire Qdgiu6;  // ../RTL/cortexm0ds_logic.v(522)
  wire Qdhow6;  // ../RTL/cortexm0ds_logic.v(1079)
  wire Qdniu6;  // ../RTL/cortexm0ds_logic.v(616)
  wire Qdohu6;  // ../RTL/cortexm0ds_logic.v(148)
  wire Qdoow6;  // ../RTL/cortexm0ds_logic.v(1172)
  wire Qduiu6;  // ../RTL/cortexm0ds_logic.v(710)
  wire Qdvhu6;  // ../RTL/cortexm0ds_logic.v(242)
  wire Qdvow6;  // ../RTL/cortexm0ds_logic.v(1266)
  wire Qe0ju6;  // ../RTL/cortexm0ds_logic.v(790)
  wire Qe1iu6;  // ../RTL/cortexm0ds_logic.v(322)
  wire Qe1pw6;  // ../RTL/cortexm0ds_logic.v(1347)
  wire Qe7ju6;  // ../RTL/cortexm0ds_logic.v(884)
  wire Qe8iu6;  // ../RTL/cortexm0ds_logic.v(416)
  wire Qe8pw6;  // ../RTL/cortexm0ds_logic.v(1440)
  wire Qe9ow6;  // ../RTL/cortexm0ds_logic.v(972)
  wire Qefiu6;  // ../RTL/cortexm0ds_logic.v(509)
  wire Qegow6;  // ../RTL/cortexm0ds_logic.v(1066)
  wire Qehbx6;  // ../RTL/cortexm0ds_logic.v(1711)
  wire Qemiu6;  // ../RTL/cortexm0ds_logic.v(603)
  wire Qenow6;  // ../RTL/cortexm0ds_logic.v(1159)
  wire Qetiu6;  // ../RTL/cortexm0ds_logic.v(697)
  wire Qeuhu6;  // ../RTL/cortexm0ds_logic.v(229)
  wire Qeuow6;  // ../RTL/cortexm0ds_logic.v(1253)
  wire Qf0iu6;  // ../RTL/cortexm0ds_logic.v(309)
  wire Qf0pw6;  // ../RTL/cortexm0ds_logic.v(1334)
  wire Qf4bx6;  // ../RTL/cortexm0ds_logic.v(1687)
  wire Qf6ju6;  // ../RTL/cortexm0ds_logic.v(871)
  wire Qf7iu6;  // ../RTL/cortexm0ds_logic.v(403)
  wire Qf7pw6;  // ../RTL/cortexm0ds_logic.v(1427)
  wire Qf8ow6;  // ../RTL/cortexm0ds_logic.v(959)
  wire Qfeiu6;  // ../RTL/cortexm0ds_logic.v(496)
  wire Qffhu6;  // ../RTL/cortexm0ds_logic.v(124)
  wire Qffow6;  // ../RTL/cortexm0ds_logic.v(1053)
  wire Qfliu6;  // ../RTL/cortexm0ds_logic.v(590)
  wire Qfmow6;  // ../RTL/cortexm0ds_logic.v(1146)
  wire Qfsiu6;  // ../RTL/cortexm0ds_logic.v(684)
  wire Qfthu6;  // ../RTL/cortexm0ds_logic.v(216)
  wire Qftow6;  // ../RTL/cortexm0ds_logic.v(1240)
  wire Qfziu6;  // ../RTL/cortexm0ds_logic.v(777)
  wire Qg5ju6;  // ../RTL/cortexm0ds_logic.v(858)
  wire Qg6iu6;  // ../RTL/cortexm0ds_logic.v(390)
  wire Qg6pw6;  // ../RTL/cortexm0ds_logic.v(1414)
  wire Qg7ow6;  // ../RTL/cortexm0ds_logic.v(946)
  wire Qgdiu6;  // ../RTL/cortexm0ds_logic.v(483)
  wire Qgdpw6;  // ../RTL/cortexm0ds_logic.v(1508)
  wire Qgeow6;  // ../RTL/cortexm0ds_logic.v(1040)
  wire Qgkiu6;  // ../RTL/cortexm0ds_logic.v(577)
  wire Qglow6;  // ../RTL/cortexm0ds_logic.v(1133)
  wire Qgriu6;  // ../RTL/cortexm0ds_logic.v(671)
  wire Qgshu6;  // ../RTL/cortexm0ds_logic.v(203)
  wire Qgsow6;  // ../RTL/cortexm0ds_logic.v(1227)
  wire Qgyiu6;  // ../RTL/cortexm0ds_logic.v(764)
  wire Qgzhu6;  // ../RTL/cortexm0ds_logic.v(296)
  wire Qgzow6;  // ../RTL/cortexm0ds_logic.v(1321)
  wire Qh4ju6;  // ../RTL/cortexm0ds_logic.v(845)
  wire Qh5iu6;  // ../RTL/cortexm0ds_logic.v(377)
  wire Qh5pw6;  // ../RTL/cortexm0ds_logic.v(1401)
  wire Qh6ow6;  // ../RTL/cortexm0ds_logic.v(933)
  wire Qhciu6;  // ../RTL/cortexm0ds_logic.v(470)
  wire Qhcpw6;  // ../RTL/cortexm0ds_logic.v(1495)
  wire Qhdow6;  // ../RTL/cortexm0ds_logic.v(1027)
  wire Qhhhu6;  // ../RTL/cortexm0ds_logic.v(128)
  wire Qhjiu6;  // ../RTL/cortexm0ds_logic.v(564)
  wire Qhkow6;  // ../RTL/cortexm0ds_logic.v(1120)
  wire Qhmpw6;  // ../RTL/cortexm0ds_logic.v(1592)
  wire Qhqiu6;  // ../RTL/cortexm0ds_logic.v(658)
  wire Qhrhu6;  // ../RTL/cortexm0ds_logic.v(190)
  wire Qhrow6;  // ../RTL/cortexm0ds_logic.v(1214)
  wire Qhxiu6;  // ../RTL/cortexm0ds_logic.v(751)
  wire Qhyhu6;  // ../RTL/cortexm0ds_logic.v(283)
  wire Qhyow6;  // ../RTL/cortexm0ds_logic.v(1308)
  wire Qi3ju6;  // ../RTL/cortexm0ds_logic.v(832)
  wire Qi4iu6;  // ../RTL/cortexm0ds_logic.v(364)
  wire Qi4pw6;  // ../RTL/cortexm0ds_logic.v(1388)
  wire Qiaju6;  // ../RTL/cortexm0ds_logic.v(925)
  wire Qibiu6;  // ../RTL/cortexm0ds_logic.v(457)
  wire Qibpw6;  // ../RTL/cortexm0ds_logic.v(1482)
  wire Qicow6;  // ../RTL/cortexm0ds_logic.v(1014)
  wire Qifhu6;  // ../RTL/cortexm0ds_logic.v(124)
  wire Qiiiu6;  // ../RTL/cortexm0ds_logic.v(551)
  wire Qijow6;  // ../RTL/cortexm0ds_logic.v(1107)
  wire Qijpw6;  // ../RTL/cortexm0ds_logic.v(1587)
  wire Qipiu6;  // ../RTL/cortexm0ds_logic.v(645)
  wire Qiqhu6;  // ../RTL/cortexm0ds_logic.v(177)
  wire Qiqow6;  // ../RTL/cortexm0ds_logic.v(1201)
  wire Qirax6;  // ../RTL/cortexm0ds_logic.v(1664)
  wire Qiwiu6;  // ../RTL/cortexm0ds_logic.v(738)
  wire Qixhu6;  // ../RTL/cortexm0ds_logic.v(270)
  wire Qixow6;  // ../RTL/cortexm0ds_logic.v(1295)
  wire Qj1qw6;  // ../RTL/cortexm0ds_logic.v(1620)
  wire Qj2ju6;  // ../RTL/cortexm0ds_logic.v(819)
  wire Qj3iu6;  // ../RTL/cortexm0ds_logic.v(351)
  wire Qj3pw6;  // ../RTL/cortexm0ds_logic.v(1375)
  wire Qj9ju6;  // ../RTL/cortexm0ds_logic.v(912)
  wire Qjaiu6;  // ../RTL/cortexm0ds_logic.v(444)
  wire Qjapw6;  // ../RTL/cortexm0ds_logic.v(1469)
  wire Qjbbx6;  // ../RTL/cortexm0ds_logic.v(1700)
  wire Qjbow6;  // ../RTL/cortexm0ds_logic.v(1001)
  wire Qjcbx6;  // ../RTL/cortexm0ds_logic.v(1702)
  wire Qjhax6;  // ../RTL/cortexm0ds_logic.v(1646)
  wire Qjhiu6;  // ../RTL/cortexm0ds_logic.v(538)
  wire Qjiow6;  // ../RTL/cortexm0ds_logic.v(1094)
  wire Qjoiu6;  // ../RTL/cortexm0ds_logic.v(632)
  wire Qjphu6;  // ../RTL/cortexm0ds_logic.v(164)
  wire Qjpow6;  // ../RTL/cortexm0ds_logic.v(1188)
  wire Qjviu6;  // ../RTL/cortexm0ds_logic.v(725)
  wire Qjwhu6;  // ../RTL/cortexm0ds_logic.v(257)
  wire Qjwow6;  // ../RTL/cortexm0ds_logic.v(1282)
  wire Qjyax6;  // ../RTL/cortexm0ds_logic.v(1677)
  wire Qjypw6;  // ../RTL/cortexm0ds_logic.v(1614)
  wire Qk1ju6;  // ../RTL/cortexm0ds_logic.v(806)
  wire Qk2iu6;  // ../RTL/cortexm0ds_logic.v(338)
  wire Qk2pw6;  // ../RTL/cortexm0ds_logic.v(1362)
  wire Qk8ju6;  // ../RTL/cortexm0ds_logic.v(899)
  wire Qk9iu6;  // ../RTL/cortexm0ds_logic.v(431)
  wire Qk9pw6;  // ../RTL/cortexm0ds_logic.v(1456)
  wire Qkabx6;  // ../RTL/cortexm0ds_logic.v(1698)
  wire Qkaow6;  // ../RTL/cortexm0ds_logic.v(988)
  wire Qkgiu6;  // ../RTL/cortexm0ds_logic.v(525)
  wire Qkhow6;  // ../RTL/cortexm0ds_logic.v(1081)
  wire Qkniu6;  // ../RTL/cortexm0ds_logic.v(619)
  wire Qkohu6;  // ../RTL/cortexm0ds_logic.v(151)
  wire Qkoow6;  // ../RTL/cortexm0ds_logic.v(1175)
  wire Qkrax6;  // ../RTL/cortexm0ds_logic.v(1664)
  wire Qkuiu6;  // ../RTL/cortexm0ds_logic.v(712)
  wire Qkvhu6;  // ../RTL/cortexm0ds_logic.v(244)
  wire Qkvow6;  // ../RTL/cortexm0ds_logic.v(1269)
  wire Ql0ju6;  // ../RTL/cortexm0ds_logic.v(793)
  wire Ql1iu6;  // ../RTL/cortexm0ds_logic.v(325)
  wire Ql1pw6;  // ../RTL/cortexm0ds_logic.v(1349)
  wire Ql7ju6;  // ../RTL/cortexm0ds_logic.v(886)
  wire Ql8iu6;  // ../RTL/cortexm0ds_logic.v(418)
  wire Ql8pw6;  // ../RTL/cortexm0ds_logic.v(1443)
  wire Ql9ow6;  // ../RTL/cortexm0ds_logic.v(975)
  wire Qlfbx6;  // ../RTL/cortexm0ds_logic.v(1707)
  wire Qlfhu6;  // ../RTL/cortexm0ds_logic.v(124)
  wire Qlfiu6;  // ../RTL/cortexm0ds_logic.v(512)
  wire Qlgow6;  // ../RTL/cortexm0ds_logic.v(1068)
  wire Qlmiu6;  // ../RTL/cortexm0ds_logic.v(606)
  wire Qlnow6;  // ../RTL/cortexm0ds_logic.v(1162)
  wire Qlopw6;  // ../RTL/cortexm0ds_logic.v(1596)
  wire Qltiu6;  // ../RTL/cortexm0ds_logic.v(699)
  wire Qluhu6;  // ../RTL/cortexm0ds_logic.v(231)
  wire Qluow6;  // ../RTL/cortexm0ds_logic.v(1256)
  wire Qm0iu6;  // ../RTL/cortexm0ds_logic.v(312)
  wire Qm0pw6;  // ../RTL/cortexm0ds_logic.v(1336)
  wire Qm6ju6;  // ../RTL/cortexm0ds_logic.v(873)
  wire Qm7iu6;  // ../RTL/cortexm0ds_logic.v(405)
  wire Qm7pw6;  // ../RTL/cortexm0ds_logic.v(1430)
  wire Qm8ow6;  // ../RTL/cortexm0ds_logic.v(962)
  wire Qmdax6;  // ../RTL/cortexm0ds_logic.v(1638)
  wire Qmdhu6;  // ../RTL/cortexm0ds_logic.v(120)
  wire Qmeiu6;  // ../RTL/cortexm0ds_logic.v(499)
  wire Qmfow6;  // ../RTL/cortexm0ds_logic.v(1055)
  wire Qmliu6;  // ../RTL/cortexm0ds_logic.v(593)
  wire Qmmow6;  // ../RTL/cortexm0ds_logic.v(1149)
  wire Qmrax6;  // ../RTL/cortexm0ds_logic.v(1664)
  wire Qmsiu6;  // ../RTL/cortexm0ds_logic.v(686)
  wire Qmthu6;  // ../RTL/cortexm0ds_logic.v(218)
  wire Qmtow6;  // ../RTL/cortexm0ds_logic.v(1243)
  wire Qmziu6;  // ../RTL/cortexm0ds_logic.v(780)
  wire Qn5ju6;  // ../RTL/cortexm0ds_logic.v(860)
  wire Qn6iu6;  // ../RTL/cortexm0ds_logic.v(392)
  wire Qn6pw6;  // ../RTL/cortexm0ds_logic.v(1417)
  wire Qn7ow6;  // ../RTL/cortexm0ds_logic.v(949)
  wire Qndiu6;  // ../RTL/cortexm0ds_logic.v(486)
  wire Qndpw6;  // ../RTL/cortexm0ds_logic.v(1510)
  wire Qneow6;  // ../RTL/cortexm0ds_logic.v(1042)
  wire Qnghu6;  // ../RTL/cortexm0ds_logic.v(127)
  wire Qnkhu6;  // ../RTL/cortexm0ds_logic.v(137)
  wire Qnkiu6;  // ../RTL/cortexm0ds_logic.v(580)
  wire Qnlow6;  // ../RTL/cortexm0ds_logic.v(1136)
  wire Qnopw6;  // ../RTL/cortexm0ds_logic.v(1596)
  wire Qnriu6;  // ../RTL/cortexm0ds_logic.v(673)
  wire Qnshu6;  // ../RTL/cortexm0ds_logic.v(205)
  wire Qnsow6;  // ../RTL/cortexm0ds_logic.v(1230)
  wire Qnyiu6;  // ../RTL/cortexm0ds_logic.v(767)
  wire Qnzhu6;  // ../RTL/cortexm0ds_logic.v(299)
  wire Qnzow6;  // ../RTL/cortexm0ds_logic.v(1323)
  wire Qo3bx6;  // ../RTL/cortexm0ds_logic.v(1686)
  wire Qo4ju6;  // ../RTL/cortexm0ds_logic.v(847)
  wire Qo5iu6;  // ../RTL/cortexm0ds_logic.v(379)
  wire Qo5pw6;  // ../RTL/cortexm0ds_logic.v(1404)
  wire Qo6ow6;  // ../RTL/cortexm0ds_logic.v(936)
  wire Qociu6;  // ../RTL/cortexm0ds_logic.v(473)
  wire Qocpw6;  // ../RTL/cortexm0ds_logic.v(1497)
  wire Qodow6;  // ../RTL/cortexm0ds_logic.v(1029)
  wire Qofhu6;  // ../RTL/cortexm0ds_logic.v(125)
  wire Qojiu6;  // ../RTL/cortexm0ds_logic.v(567)
  wire Qokow6;  // ../RTL/cortexm0ds_logic.v(1123)
  wire Qoqiu6;  // ../RTL/cortexm0ds_logic.v(660)
  wire Qorax6;  // ../RTL/cortexm0ds_logic.v(1664)
  wire Qorhu6;  // ../RTL/cortexm0ds_logic.v(192)
  wire Qorow6;  // ../RTL/cortexm0ds_logic.v(1217)
  wire Qoxiu6;  // ../RTL/cortexm0ds_logic.v(754)
  wire Qoyhu6;  // ../RTL/cortexm0ds_logic.v(286)
  wire Qoyow6;  // ../RTL/cortexm0ds_logic.v(1310)
  wire Qp3ju6;  // ../RTL/cortexm0ds_logic.v(834)
  wire Qp4iu6;  // ../RTL/cortexm0ds_logic.v(366)
  wire Qp4pw6;  // ../RTL/cortexm0ds_logic.v(1391)
  wire Qpaju6;  // ../RTL/cortexm0ds_logic.v(928)
  wire Qpbiu6;  // ../RTL/cortexm0ds_logic.v(460)
  wire Qpbpw6;  // ../RTL/cortexm0ds_logic.v(1484)
  wire Qpcow6;  // ../RTL/cortexm0ds_logic.v(1016)
  wire Qpiiu6;  // ../RTL/cortexm0ds_logic.v(554)
  wire Qpjhu6;  // ../RTL/cortexm0ds_logic.v(134)
  wire Qpjow6;  // ../RTL/cortexm0ds_logic.v(1110)
  wire Qpopw6;  // ../RTL/cortexm0ds_logic.v(1596)
  wire Qppiu6;  // ../RTL/cortexm0ds_logic.v(647)
  wire Qpqhu6;  // ../RTL/cortexm0ds_logic.v(179)
  wire Qpqow6;  // ../RTL/cortexm0ds_logic.v(1204)
  wire Qpwiu6;  // ../RTL/cortexm0ds_logic.v(741)
  wire Qpxhu6;  // ../RTL/cortexm0ds_logic.v(273)
  wire Qpxow6;  // ../RTL/cortexm0ds_logic.v(1297)
  wire Qq2ju6;  // ../RTL/cortexm0ds_logic.v(821)
  wire Qq3iu6;  // ../RTL/cortexm0ds_logic.v(353)
  wire Qq3pw6;  // ../RTL/cortexm0ds_logic.v(1378)
  wire Qq9ju6;  // ../RTL/cortexm0ds_logic.v(915)
  wire Qqaiu6;  // ../RTL/cortexm0ds_logic.v(447)
  wire Qqapw6;  // ../RTL/cortexm0ds_logic.v(1471)
  wire Qqbow6;  // ../RTL/cortexm0ds_logic.v(1003)
  wire Qqdhu6;  // ../RTL/cortexm0ds_logic.v(120)
  wire Qqhiu6;  // ../RTL/cortexm0ds_logic.v(541)
  wire Qqiow6;  // ../RTL/cortexm0ds_logic.v(1097)
  wire Qqoiu6;  // ../RTL/cortexm0ds_logic.v(634)
  wire Qqphu6;  // ../RTL/cortexm0ds_logic.v(166)
  wire Qqpow6;  // ../RTL/cortexm0ds_logic.v(1191)
  wire Qqviu6;  // ../RTL/cortexm0ds_logic.v(728)
  wire Qqwhu6;  // ../RTL/cortexm0ds_logic.v(260)
  wire Qqwow6;  // ../RTL/cortexm0ds_logic.v(1284)
  wire Qr1ju6;  // ../RTL/cortexm0ds_logic.v(808)
  wire Qr2iu6;  // ../RTL/cortexm0ds_logic.v(340)
  wire Qr2pw6;  // ../RTL/cortexm0ds_logic.v(1365)
  wire Qr8ju6;  // ../RTL/cortexm0ds_logic.v(902)
  wire Qr9iu6;  // ../RTL/cortexm0ds_logic.v(434)
  wire Qr9pw6;  // ../RTL/cortexm0ds_logic.v(1458)
  wire Qraow6;  // ../RTL/cortexm0ds_logic.v(990)
  wire Qrgiu6;  // ../RTL/cortexm0ds_logic.v(528)
  wire Qrhow6;  // ../RTL/cortexm0ds_logic.v(1084)
  wire Qrihu6;  // ../RTL/cortexm0ds_logic.v(132)
  wire Qrniu6;  // ../RTL/cortexm0ds_logic.v(621)
  wire Qrohu6;  // ../RTL/cortexm0ds_logic.v(153)
  wire Qroow6;  // ../RTL/cortexm0ds_logic.v(1178)
  wire Qruiu6;  // ../RTL/cortexm0ds_logic.v(715)
  wire Qrvhu6;  // ../RTL/cortexm0ds_logic.v(247)
  wire Qrvow6;  // ../RTL/cortexm0ds_logic.v(1271)
  wire Qs0ju6;  // ../RTL/cortexm0ds_logic.v(795)
  wire Qs1iu6;  // ../RTL/cortexm0ds_logic.v(327)
  wire Qs1pw6;  // ../RTL/cortexm0ds_logic.v(1352)
  wire Qs7ju6;  // ../RTL/cortexm0ds_logic.v(889)
  wire Qs8iu6;  // ../RTL/cortexm0ds_logic.v(421)
  wire Qs8pw6;  // ../RTL/cortexm0ds_logic.v(1445)
  wire Qs9ow6;  // ../RTL/cortexm0ds_logic.v(977)
  wire Qsfax6;  // ../RTL/cortexm0ds_logic.v(1642)
  wire Qsfiu6;  // ../RTL/cortexm0ds_logic.v(515)
  wire Qsgow6;  // ../RTL/cortexm0ds_logic.v(1071)
  wire Qsmiu6;  // ../RTL/cortexm0ds_logic.v(608)
  wire Qsnow6;  // ../RTL/cortexm0ds_logic.v(1165)
  wire Qstiu6;  // ../RTL/cortexm0ds_logic.v(702)
  wire Qsuhu6;  // ../RTL/cortexm0ds_logic.v(234)
  wire Qsuow6;  // ../RTL/cortexm0ds_logic.v(1258)
  wire Qt0iu6;  // ../RTL/cortexm0ds_logic.v(314)
  wire Qt0pw6;  // ../RTL/cortexm0ds_logic.v(1339)
  wire Qt6ju6;  // ../RTL/cortexm0ds_logic.v(876)
  wire Qt7iu6;  // ../RTL/cortexm0ds_logic.v(408)
  wire Qt7pw6;  // ../RTL/cortexm0ds_logic.v(1432)
  wire Qt8ow6;  // ../RTL/cortexm0ds_logic.v(964)
  wire Qteiu6;  // ../RTL/cortexm0ds_logic.v(502)
  wire Qtfow6;  // ../RTL/cortexm0ds_logic.v(1058)
  wire Qtliu6;  // ../RTL/cortexm0ds_logic.v(595)
  wire Qtmow6;  // ../RTL/cortexm0ds_logic.v(1152)
  wire Qtsiu6;  // ../RTL/cortexm0ds_logic.v(689)
  wire Qtthu6;  // ../RTL/cortexm0ds_logic.v(221)
  wire Qttow6;  // ../RTL/cortexm0ds_logic.v(1245)
  wire Qtziu6;  // ../RTL/cortexm0ds_logic.v(782)
  wire Qu5ju6;  // ../RTL/cortexm0ds_logic.v(863)
  wire Qu6iu6;  // ../RTL/cortexm0ds_logic.v(395)
  wire Qu6pw6;  // ../RTL/cortexm0ds_logic.v(1419)
  wire Qu7ow6;  // ../RTL/cortexm0ds_logic.v(951)
  wire Qudbx6;  // ../RTL/cortexm0ds_logic.v(1704)
  wire Qudiu6;  // ../RTL/cortexm0ds_logic.v(489)
  wire Qudpw6;  // ../RTL/cortexm0ds_logic.v(1513)
  wire Queow6;  // ../RTL/cortexm0ds_logic.v(1045)
  wire Qufax6;  // ../RTL/cortexm0ds_logic.v(1643)
  wire Qukax6;  // ../RTL/cortexm0ds_logic.v(1652)
  wire Qukiu6;  // ../RTL/cortexm0ds_logic.v(582)
  wire Qulow6;  // ../RTL/cortexm0ds_logic.v(1139)
  wire Quriu6;  // ../RTL/cortexm0ds_logic.v(676)
  wire Qushu6;  // ../RTL/cortexm0ds_logic.v(208)
  wire Qusow6;  // ../RTL/cortexm0ds_logic.v(1232)
  wire Quyiu6;  // ../RTL/cortexm0ds_logic.v(769)
  wire Quzhu6;  // ../RTL/cortexm0ds_logic.v(301)
  wire Quzow6;  // ../RTL/cortexm0ds_logic.v(1326)
  wire Qv4ju6;  // ../RTL/cortexm0ds_logic.v(850)
  wire Qv5iu6;  // ../RTL/cortexm0ds_logic.v(382)
  wire Qv5pw6;  // ../RTL/cortexm0ds_logic.v(1406)
  wire Qv6ow6;  // ../RTL/cortexm0ds_logic.v(938)
  wire Qvciu6;  // ../RTL/cortexm0ds_logic.v(476)
  wire Qvcpw6;  // ../RTL/cortexm0ds_logic.v(1500)
  wire Qvdow6;  // ../RTL/cortexm0ds_logic.v(1032)
  wire Qvehu6;  // ../RTL/cortexm0ds_logic.v(123)
  wire Qvjiu6;  // ../RTL/cortexm0ds_logic.v(569)
  wire Qvkow6;  // ../RTL/cortexm0ds_logic.v(1126)
  wire Qvqiu6;  // ../RTL/cortexm0ds_logic.v(663)
  wire Qvrhu6;  // ../RTL/cortexm0ds_logic.v(195)
  wire Qvrow6;  // ../RTL/cortexm0ds_logic.v(1219)
  wire Qvvax6;  // ../RTL/cortexm0ds_logic.v(1672)
  wire Qvxiu6;  // ../RTL/cortexm0ds_logic.v(756)
  wire Qvyhu6;  // ../RTL/cortexm0ds_logic.v(288)
  wire Qvyow6;  // ../RTL/cortexm0ds_logic.v(1313)
  wire Qw3ju6;  // ../RTL/cortexm0ds_logic.v(837)
  wire Qw4iu6;  // ../RTL/cortexm0ds_logic.v(369)
  wire Qw4pw6;  // ../RTL/cortexm0ds_logic.v(1393)
  wire Qwbiu6;  // ../RTL/cortexm0ds_logic.v(463)
  wire Qwbpw6;  // ../RTL/cortexm0ds_logic.v(1487)
  wire Qwcow6;  // ../RTL/cortexm0ds_logic.v(1019)
  wire Qwdhu6;  // ../RTL/cortexm0ds_logic.v(120)
  wire Qwfax6;  // ../RTL/cortexm0ds_logic.v(1643)
  wire Qwfbx6;  // ../RTL/cortexm0ds_logic.v(1708)
  wire Qwiiu6;  // ../RTL/cortexm0ds_logic.v(556)
  wire Qwjow6;  // ../RTL/cortexm0ds_logic.v(1113)
  wire Qwpiu6;  // ../RTL/cortexm0ds_logic.v(650)
  wire Qwqhu6;  // ../RTL/cortexm0ds_logic.v(182)
  wire Qwqow6;  // ../RTL/cortexm0ds_logic.v(1206)
  wire Qwwiu6;  // ../RTL/cortexm0ds_logic.v(743)
  wire Qwxhu6;  // ../RTL/cortexm0ds_logic.v(275)
  wire Qwxow6;  // ../RTL/cortexm0ds_logic.v(1300)
  wire Qx0bx6;  // ../RTL/cortexm0ds_logic.v(1681)
  wire Qx2ju6;  // ../RTL/cortexm0ds_logic.v(824)
  wire Qx3iu6;  // ../RTL/cortexm0ds_logic.v(356)
  wire Qx3pw6;  // ../RTL/cortexm0ds_logic.v(1380)
  wire Qx9ju6;  // ../RTL/cortexm0ds_logic.v(918)
  wire Qxaiu6;  // ../RTL/cortexm0ds_logic.v(450)
  wire Qxapw6;  // ../RTL/cortexm0ds_logic.v(1474)
  wire Qxbow6;  // ../RTL/cortexm0ds_logic.v(1006)
  wire Qxhiu6;  // ../RTL/cortexm0ds_logic.v(543)
  wire Qxibx6;  // ../RTL/cortexm0ds_logic.v(1714)
  wire Qxiow6;  // ../RTL/cortexm0ds_logic.v(1100)
  wire Qxoiu6;  // ../RTL/cortexm0ds_logic.v(637)
  wire Qxphu6;  // ../RTL/cortexm0ds_logic.v(169)
  wire Qxpow6;  // ../RTL/cortexm0ds_logic.v(1193)
  wire Qxviu6;  // ../RTL/cortexm0ds_logic.v(730)
  wire Qxwhu6;  // ../RTL/cortexm0ds_logic.v(262)
  wire Qxwow6;  // ../RTL/cortexm0ds_logic.v(1287)
  wire Qy1ju6;  // ../RTL/cortexm0ds_logic.v(811)
  wire Qy2iu6;  // ../RTL/cortexm0ds_logic.v(343)
  wire Qy2pw6;  // ../RTL/cortexm0ds_logic.v(1367)
  wire Qy8ju6;  // ../RTL/cortexm0ds_logic.v(905)
  wire Qy9iu6;  // ../RTL/cortexm0ds_logic.v(437)
  wire Qy9pw6;  // ../RTL/cortexm0ds_logic.v(1461)
  wire Qyaow6;  // ../RTL/cortexm0ds_logic.v(993)
  wire Qygiu6;  // ../RTL/cortexm0ds_logic.v(530)
  wire Qyhow6;  // ../RTL/cortexm0ds_logic.v(1087)
  wire Qyjax6;  // ../RTL/cortexm0ds_logic.v(1650)
  wire Qyniu6;  // ../RTL/cortexm0ds_logic.v(624)
  wire Qyohu6;  // ../RTL/cortexm0ds_logic.v(156)
  wire Qyoow6;  // ../RTL/cortexm0ds_logic.v(1180)
  wire Qyuiu6;  // ../RTL/cortexm0ds_logic.v(717)
  wire Qyvhu6;  // ../RTL/cortexm0ds_logic.v(249)
  wire Qyvow6;  // ../RTL/cortexm0ds_logic.v(1274)
  wire Qz0ju6;  // ../RTL/cortexm0ds_logic.v(798)
  wire Qz1iu6;  // ../RTL/cortexm0ds_logic.v(330)
  wire Qz1pw6;  // ../RTL/cortexm0ds_logic.v(1354)
  wire Qz7ju6;  // ../RTL/cortexm0ds_logic.v(892)
  wire Qz8iu6;  // ../RTL/cortexm0ds_logic.v(424)
  wire Qz8pw6;  // ../RTL/cortexm0ds_logic.v(1448)
  wire Qz9ow6;  // ../RTL/cortexm0ds_logic.v(980)
  wire Qzfiu6;  // ../RTL/cortexm0ds_logic.v(517)
  wire Qzgow6;  // ../RTL/cortexm0ds_logic.v(1074)
  wire Qzmiu6;  // ../RTL/cortexm0ds_logic.v(611)
  wire Qznow6;  // ../RTL/cortexm0ds_logic.v(1167)
  wire Qztiu6;  // ../RTL/cortexm0ds_logic.v(704)
  wire Qzuhu6;  // ../RTL/cortexm0ds_logic.v(236)
  wire Qzuow6;  // ../RTL/cortexm0ds_logic.v(1261)
  wire R04ju6;  // ../RTL/cortexm0ds_logic.v(838)
  wire R05iu6;  // ../RTL/cortexm0ds_logic.v(370)
  wire R05pw6;  // ../RTL/cortexm0ds_logic.v(1395)
  wire R0ciu6;  // ../RTL/cortexm0ds_logic.v(464)
  wire R0cpw6;  // ../RTL/cortexm0ds_logic.v(1488)
  wire R0dow6;  // ../RTL/cortexm0ds_logic.v(1020)
  wire R0ghu6;  // ../RTL/cortexm0ds_logic.v(125)
  wire R0jiu6;  // ../RTL/cortexm0ds_logic.v(558)
  wire R0kow6;  // ../RTL/cortexm0ds_logic.v(1114)
  wire R0nhu6;  // ../RTL/cortexm0ds_logic.v(144)
  wire R0qiu6;  // ../RTL/cortexm0ds_logic.v(651)
  wire R0rhu6;  // ../RTL/cortexm0ds_logic.v(183)
  wire R0row6;  // ../RTL/cortexm0ds_logic.v(1208)
  wire R0xiu6;  // ../RTL/cortexm0ds_logic.v(745)
  wire R0yhu6;  // ../RTL/cortexm0ds_logic.v(277)
  wire R0yow6;  // ../RTL/cortexm0ds_logic.v(1301)
  wire R13ju6;  // ../RTL/cortexm0ds_logic.v(825)
  wire R14iu6;  // ../RTL/cortexm0ds_logic.v(357)
  wire R14pw6;  // ../RTL/cortexm0ds_logic.v(1382)
  wire R19ax6;  // ../RTL/cortexm0ds_logic.v(1629)
  wire R1abx6;  // ../RTL/cortexm0ds_logic.v(1697)
  wire R1aju6;  // ../RTL/cortexm0ds_logic.v(919)
  wire R1biu6;  // ../RTL/cortexm0ds_logic.v(451)
  wire R1bpw6;  // ../RTL/cortexm0ds_logic.v(1475)
  wire R1cow6;  // ../RTL/cortexm0ds_logic.v(1007)
  wire R1eax6;  // ../RTL/cortexm0ds_logic.v(1639)
  wire R1iiu6;  // ../RTL/cortexm0ds_logic.v(545)
  wire R1jow6;  // ../RTL/cortexm0ds_logic.v(1101)
  wire R1piu6;  // ../RTL/cortexm0ds_logic.v(638)
  wire R1qhu6;  // ../RTL/cortexm0ds_logic.v(170)
  wire R1qow6;  // ../RTL/cortexm0ds_logic.v(1195)
  wire R1wiu6;  // ../RTL/cortexm0ds_logic.v(732)
  wire R1xhu6;  // ../RTL/cortexm0ds_logic.v(264)
  wire R1xow6;  // ../RTL/cortexm0ds_logic.v(1288)
  wire R22ju6;  // ../RTL/cortexm0ds_logic.v(812)
  wire R23iu6;  // ../RTL/cortexm0ds_logic.v(344)
  wire R23pw6;  // ../RTL/cortexm0ds_logic.v(1369)
  wire R29ju6;  // ../RTL/cortexm0ds_logic.v(906)
  wire R2aiu6;  // ../RTL/cortexm0ds_logic.v(438)
  wire R2apw6;  // ../RTL/cortexm0ds_logic.v(1462)
  wire R2bow6;  // ../RTL/cortexm0ds_logic.v(994)
  wire R2hax6;  // ../RTL/cortexm0ds_logic.v(1645)
  wire R2hiu6;  // ../RTL/cortexm0ds_logic.v(532)
  wire R2iow6;  // ../RTL/cortexm0ds_logic.v(1088)
  wire R2oiu6;  // ../RTL/cortexm0ds_logic.v(625)
  wire R2phu6;  // ../RTL/cortexm0ds_logic.v(157)
  wire R2pow6;  // ../RTL/cortexm0ds_logic.v(1182)
  wire R2viu6;  // ../RTL/cortexm0ds_logic.v(719)
  wire R2whu6;  // ../RTL/cortexm0ds_logic.v(251)
  wire R2wow6;  // ../RTL/cortexm0ds_logic.v(1275)
  wire R31ju6;  // ../RTL/cortexm0ds_logic.v(799)
  wire R32iu6;  // ../RTL/cortexm0ds_logic.v(331)
  wire R32pw6;  // ../RTL/cortexm0ds_logic.v(1356)
  wire R38ju6;  // ../RTL/cortexm0ds_logic.v(893)
  wire R39iu6;  // ../RTL/cortexm0ds_logic.v(425)
  wire R39pw6;  // ../RTL/cortexm0ds_logic.v(1449)
  wire R3aow6;  // ../RTL/cortexm0ds_logic.v(981)
  wire R3giu6;  // ../RTL/cortexm0ds_logic.v(519)
  wire R3how6;  // ../RTL/cortexm0ds_logic.v(1075)
  wire R3niu6;  // ../RTL/cortexm0ds_logic.v(612)
  wire R3oow6;  // ../RTL/cortexm0ds_logic.v(1169)
  wire R3uiu6;  // ../RTL/cortexm0ds_logic.v(706)
  wire R3vhu6;  // ../RTL/cortexm0ds_logic.v(238)
  wire R3vow6;  // ../RTL/cortexm0ds_logic.v(1262)
  wire R3vpw6;  // ../RTL/cortexm0ds_logic.v(1608)
  wire R40ju6;  // ../RTL/cortexm0ds_logic.v(786)
  wire R41iu6;  // ../RTL/cortexm0ds_logic.v(318)
  wire R41pw6;  // ../RTL/cortexm0ds_logic.v(1343)
  wire R47ju6;  // ../RTL/cortexm0ds_logic.v(880)
  wire R48iu6;  // ../RTL/cortexm0ds_logic.v(412)
  wire R48pw6;  // ../RTL/cortexm0ds_logic.v(1436)
  wire R49ow6;  // ../RTL/cortexm0ds_logic.v(968)
  wire R4fiu6;  // ../RTL/cortexm0ds_logic.v(506)
  wire R4gow6;  // ../RTL/cortexm0ds_logic.v(1062)
  wire R4miu6;  // ../RTL/cortexm0ds_logic.v(599)
  wire R4now6;  // ../RTL/cortexm0ds_logic.v(1156)
  wire R4tiu6;  // ../RTL/cortexm0ds_logic.v(693)
  wire R4uhu6;  // ../RTL/cortexm0ds_logic.v(225)
  wire R4uow6;  // ../RTL/cortexm0ds_logic.v(1249)
  wire R50iu6;  // ../RTL/cortexm0ds_logic.v(305)
  wire R50pw6;  // ../RTL/cortexm0ds_logic.v(1330)
  wire R56ju6;  // ../RTL/cortexm0ds_logic.v(867)
  wire R57iu6;  // ../RTL/cortexm0ds_logic.v(399)
  wire R57pw6;  // ../RTL/cortexm0ds_logic.v(1423)
  wire R58ow6;  // ../RTL/cortexm0ds_logic.v(955)
  wire R5eiu6;  // ../RTL/cortexm0ds_logic.v(493)
  wire R5fow6;  // ../RTL/cortexm0ds_logic.v(1049)
  wire R5liu6;  // ../RTL/cortexm0ds_logic.v(586)
  wire R5mow6;  // ../RTL/cortexm0ds_logic.v(1143)
  wire R5siu6;  // ../RTL/cortexm0ds_logic.v(680)
  wire R5thu6;  // ../RTL/cortexm0ds_logic.v(212)
  wire R5tow6;  // ../RTL/cortexm0ds_logic.v(1236)
  wire R5ziu6;  // ../RTL/cortexm0ds_logic.v(773)
  wire R65ju6;  // ../RTL/cortexm0ds_logic.v(854)
  wire R66iu6;  // ../RTL/cortexm0ds_logic.v(386)
  wire R66pw6;  // ../RTL/cortexm0ds_logic.v(1410)
  wire R67ow6;  // ../RTL/cortexm0ds_logic.v(942)
  wire R6diu6;  // ../RTL/cortexm0ds_logic.v(480)
  wire R6dpw6;  // ../RTL/cortexm0ds_logic.v(1504)
  wire R6eow6;  // ../RTL/cortexm0ds_logic.v(1036)
  wire R6hhu6;  // ../RTL/cortexm0ds_logic.v(128)
  wire R6kiu6;  // ../RTL/cortexm0ds_logic.v(573)
  wire R6low6;  // ../RTL/cortexm0ds_logic.v(1130)
  wire R6riu6;  // ../RTL/cortexm0ds_logic.v(667)
  wire R6shu6;  // ../RTL/cortexm0ds_logic.v(199)
  wire R6sow6;  // ../RTL/cortexm0ds_logic.v(1223)
  wire R6yiu6;  // ../RTL/cortexm0ds_logic.v(760)
  wire R6zhu6;  // ../RTL/cortexm0ds_logic.v(292)
  wire R6zow6;  // ../RTL/cortexm0ds_logic.v(1317)
  wire R74ju6;  // ../RTL/cortexm0ds_logic.v(841)
  wire R75iu6;  // ../RTL/cortexm0ds_logic.v(373)
  wire R75pw6;  // ../RTL/cortexm0ds_logic.v(1397)
  wire R76ow6;  // ../RTL/cortexm0ds_logic.v(929)
  wire R7ciu6;  // ../RTL/cortexm0ds_logic.v(467)
  wire R7cpw6;  // ../RTL/cortexm0ds_logic.v(1491)
  wire R7dow6;  // ../RTL/cortexm0ds_logic.v(1023)
  wire R7ibx6;  // ../RTL/cortexm0ds_logic.v(1712)
  wire R7jiu6;  // ../RTL/cortexm0ds_logic.v(560)
  wire R7kow6;  // ../RTL/cortexm0ds_logic.v(1117)
  wire R7kpw6;  // ../RTL/cortexm0ds_logic.v(1588)
  wire R7nax6;  // ../RTL/cortexm0ds_logic.v(1656)
  wire R7qiu6;  // ../RTL/cortexm0ds_logic.v(654)
  wire R7rhu6;  // ../RTL/cortexm0ds_logic.v(186)
  wire R7row6;  // ../RTL/cortexm0ds_logic.v(1210)
  wire R7xiu6;  // ../RTL/cortexm0ds_logic.v(747)
  wire R7yhu6;  // ../RTL/cortexm0ds_logic.v(279)
  wire R7yow6;  // ../RTL/cortexm0ds_logic.v(1304)
  wire R83ju6;  // ../RTL/cortexm0ds_logic.v(828)
  wire R84iu6;  // ../RTL/cortexm0ds_logic.v(360)
  wire R84pw6;  // ../RTL/cortexm0ds_logic.v(1384)
  wire R8aju6;  // ../RTL/cortexm0ds_logic.v(922)
  wire R8biu6;  // ../RTL/cortexm0ds_logic.v(454)
  wire R8bpw6;  // ../RTL/cortexm0ds_logic.v(1478)
  wire R8cow6;  // ../RTL/cortexm0ds_logic.v(1010)
  wire R8iiu6;  // ../RTL/cortexm0ds_logic.v(547)
  wire R8jow6;  // ../RTL/cortexm0ds_logic.v(1104)
  wire R8piu6;  // ../RTL/cortexm0ds_logic.v(641)
  wire R8qhu6;  // ../RTL/cortexm0ds_logic.v(173)
  wire R8qow6;  // ../RTL/cortexm0ds_logic.v(1197)
  wire R8wiu6;  // ../RTL/cortexm0ds_logic.v(734)
  wire R8xhu6;  // ../RTL/cortexm0ds_logic.v(266)
  wire R8xow6;  // ../RTL/cortexm0ds_logic.v(1291)
  wire R92ju6;  // ../RTL/cortexm0ds_logic.v(815)
  wire R93iu6;  // ../RTL/cortexm0ds_logic.v(347)
  wire R93pw6;  // ../RTL/cortexm0ds_logic.v(1371)
  wire R99ju6;  // ../RTL/cortexm0ds_logic.v(909)
  wire R9aiu6;  // ../RTL/cortexm0ds_logic.v(441)
  wire R9apw6;  // ../RTL/cortexm0ds_logic.v(1465)
  wire R9bow6;  // ../RTL/cortexm0ds_logic.v(997)
  wire R9hiu6;  // ../RTL/cortexm0ds_logic.v(534)
  wire R9ibx6;  // ../RTL/cortexm0ds_logic.v(1712)
  wire R9iow6;  // ../RTL/cortexm0ds_logic.v(1091)
  wire R9mpw6;  // ../RTL/cortexm0ds_logic.v(1592)
  wire R9ohu6;  // ../RTL/cortexm0ds_logic.v(146)
  wire R9oiu6;  // ../RTL/cortexm0ds_logic.v(628)
  wire R9phu6;  // ../RTL/cortexm0ds_logic.v(160)
  wire R9pow6;  // ../RTL/cortexm0ds_logic.v(1184)
  wire R9viu6;  // ../RTL/cortexm0ds_logic.v(721)
  wire R9whu6;  // ../RTL/cortexm0ds_logic.v(253)
  wire R9wow6;  // ../RTL/cortexm0ds_logic.v(1278)
  wire R9yax6;  // ../RTL/cortexm0ds_logic.v(1676)
  wire Ra1ju6;  // ../RTL/cortexm0ds_logic.v(802)
  wire Ra2iu6;  // ../RTL/cortexm0ds_logic.v(334)
  wire Ra2pw6;  // ../RTL/cortexm0ds_logic.v(1358)
  wire Ra2qw6;  // ../RTL/cortexm0ds_logic.v(1621)
  wire Ra8ju6;  // ../RTL/cortexm0ds_logic.v(896)
  wire Ra9iu6;  // ../RTL/cortexm0ds_logic.v(428)
  wire Ra9pw6;  // ../RTL/cortexm0ds_logic.v(1452)
  wire Raaow6;  // ../RTL/cortexm0ds_logic.v(984)
  wire Ragiu6;  // ../RTL/cortexm0ds_logic.v(521)
  wire Rahow6;  // ../RTL/cortexm0ds_logic.v(1078)
  wire Raniu6;  // ../RTL/cortexm0ds_logic.v(615)
  wire Raohu6;  // ../RTL/cortexm0ds_logic.v(147)
  wire Raoow6;  // ../RTL/cortexm0ds_logic.v(1171)
  wire Rauiu6;  // ../RTL/cortexm0ds_logic.v(708)
  wire Ravhu6;  // ../RTL/cortexm0ds_logic.v(240)
  wire Ravow6;  // ../RTL/cortexm0ds_logic.v(1265)
  wire Rb0ju6;  // ../RTL/cortexm0ds_logic.v(789)
  wire Rb1iu6;  // ../RTL/cortexm0ds_logic.v(321)
  wire Rb1pw6;  // ../RTL/cortexm0ds_logic.v(1345)
  wire Rb7ju6;  // ../RTL/cortexm0ds_logic.v(883)
  wire Rb8iu6;  // ../RTL/cortexm0ds_logic.v(415)
  wire Rb8pw6;  // ../RTL/cortexm0ds_logic.v(1439)
  wire Rb9ow6;  // ../RTL/cortexm0ds_logic.v(971)
  wire Rbfiu6;  // ../RTL/cortexm0ds_logic.v(508)
  wire Rbgow6;  // ../RTL/cortexm0ds_logic.v(1065)
  wire Rbibx6;  // ../RTL/cortexm0ds_logic.v(1712)
  wire Rbmiu6;  // ../RTL/cortexm0ds_logic.v(602)
  wire Rbnow6;  // ../RTL/cortexm0ds_logic.v(1158)
  wire Rbtiu6;  // ../RTL/cortexm0ds_logic.v(695)
  wire Rbuhu6;  // ../RTL/cortexm0ds_logic.v(227)
  wire Rbuow6;  // ../RTL/cortexm0ds_logic.v(1252)
  wire Rc0iu6;  // ../RTL/cortexm0ds_logic.v(308)
  wire Rc0pw6;  // ../RTL/cortexm0ds_logic.v(1332)
  wire Rc6ju6;  // ../RTL/cortexm0ds_logic.v(870)
  wire Rc7iu6;  // ../RTL/cortexm0ds_logic.v(402)
  wire Rc7pw6;  // ../RTL/cortexm0ds_logic.v(1426)
  wire Rc8ow6;  // ../RTL/cortexm0ds_logic.v(958)
  wire Rceiu6;  // ../RTL/cortexm0ds_logic.v(495)
  wire Rcfow6;  // ../RTL/cortexm0ds_logic.v(1052)
  wire Rcliu6;  // ../RTL/cortexm0ds_logic.v(589)
  wire Rcmow6;  // ../RTL/cortexm0ds_logic.v(1145)
  wire Rcsiu6;  // ../RTL/cortexm0ds_logic.v(682)
  wire Rcthu6;  // ../RTL/cortexm0ds_logic.v(214)
  wire Rctow6;  // ../RTL/cortexm0ds_logic.v(1239)
  wire Rcziu6;  // ../RTL/cortexm0ds_logic.v(776)
  wire Rd5ju6;  // ../RTL/cortexm0ds_logic.v(857)
  wire Rd6iu6;  // ../RTL/cortexm0ds_logic.v(389)
  wire Rd6pw6;  // ../RTL/cortexm0ds_logic.v(1413)
  wire Rd7ow6;  // ../RTL/cortexm0ds_logic.v(945)
  wire Rddiu6;  // ../RTL/cortexm0ds_logic.v(482)
  wire Rddpw6;  // ../RTL/cortexm0ds_logic.v(1507)
  wire Rdeow6;  // ../RTL/cortexm0ds_logic.v(1039)
  wire Rdibx6;  // ../RTL/cortexm0ds_logic.v(1713)
  wire Rdkiu6;  // ../RTL/cortexm0ds_logic.v(576)
  wire Rdkpw6;  // ../RTL/cortexm0ds_logic.v(1588)
  wire Rdlow6;  // ../RTL/cortexm0ds_logic.v(1132)
  wire Rdriu6;  // ../RTL/cortexm0ds_logic.v(669)
  wire Rdshu6;  // ../RTL/cortexm0ds_logic.v(201)
  wire Rdsow6;  // ../RTL/cortexm0ds_logic.v(1226)
  wire Rdyiu6;  // ../RTL/cortexm0ds_logic.v(763)
  wire Rdzhu6;  // ../RTL/cortexm0ds_logic.v(295)
  wire Rdzow6;  // ../RTL/cortexm0ds_logic.v(1319)
  wire Re4ju6;  // ../RTL/cortexm0ds_logic.v(844)
  wire Re5iu6;  // ../RTL/cortexm0ds_logic.v(376)
  wire Re5pw6;  // ../RTL/cortexm0ds_logic.v(1400)
  wire Re6ow6;  // ../RTL/cortexm0ds_logic.v(932)
  wire Reciu6;  // ../RTL/cortexm0ds_logic.v(469)
  wire Recpw6;  // ../RTL/cortexm0ds_logic.v(1494)
  wire Redow6;  // ../RTL/cortexm0ds_logic.v(1026)
  wire Rejiu6;  // ../RTL/cortexm0ds_logic.v(563)
  wire Rekbx6;  // ../RTL/cortexm0ds_logic.v(1716)
  wire Rekow6;  // ../RTL/cortexm0ds_logic.v(1119)
  wire Reqiu6;  // ../RTL/cortexm0ds_logic.v(656)
  wire Rerhu6;  // ../RTL/cortexm0ds_logic.v(188)
  wire Rerow6;  // ../RTL/cortexm0ds_logic.v(1213)
  wire Rexiu6;  // ../RTL/cortexm0ds_logic.v(750)
  wire Reyhu6;  // ../RTL/cortexm0ds_logic.v(282)
  wire Reyow6;  // ../RTL/cortexm0ds_logic.v(1306)
  wire Rezax6;  // ../RTL/cortexm0ds_logic.v(1678)
  wire Rf3ju6;  // ../RTL/cortexm0ds_logic.v(831)
  wire Rf4iu6;  // ../RTL/cortexm0ds_logic.v(363)
  wire Rf4pw6;  // ../RTL/cortexm0ds_logic.v(1387)
  wire Rfaju6;  // ../RTL/cortexm0ds_logic.v(924)
  wire Rfbiu6;  // ../RTL/cortexm0ds_logic.v(456)
  wire Rfbpw6;  // ../RTL/cortexm0ds_logic.v(1481)
  wire Rfcow6;  // ../RTL/cortexm0ds_logic.v(1013)
  wire Rfibx6;  // ../RTL/cortexm0ds_logic.v(1713)
  wire Rfiiu6;  // ../RTL/cortexm0ds_logic.v(550)
  wire Rfjow6;  // ../RTL/cortexm0ds_logic.v(1106)
  wire Rfkpw6;  // ../RTL/cortexm0ds_logic.v(1588)
  wire Rfpiu6;  // ../RTL/cortexm0ds_logic.v(643)
  wire Rfqhu6;  // ../RTL/cortexm0ds_logic.v(175)
  wire Rfqow6;  // ../RTL/cortexm0ds_logic.v(1200)
  wire Rfwiu6;  // ../RTL/cortexm0ds_logic.v(737)
  wire Rfxax6;  // ../RTL/cortexm0ds_logic.v(1675)
  wire Rfxhu6;  // ../RTL/cortexm0ds_logic.v(269)
  wire Rfxow6;  // ../RTL/cortexm0ds_logic.v(1293)
  wire Rg2ju6;  // ../RTL/cortexm0ds_logic.v(818)
  wire Rg3iu6;  // ../RTL/cortexm0ds_logic.v(350)
  wire Rg3pw6;  // ../RTL/cortexm0ds_logic.v(1374)
  wire Rg9ax6;  // ../RTL/cortexm0ds_logic.v(1630)
  wire Rg9ju6;  // ../RTL/cortexm0ds_logic.v(911)
  wire Rgaiu6;  // ../RTL/cortexm0ds_logic.v(443)
  wire Rgapw6;  // ../RTL/cortexm0ds_logic.v(1468)
  wire Rgbow6;  // ../RTL/cortexm0ds_logic.v(1000)
  wire Rghiu6;  // ../RTL/cortexm0ds_logic.v(537)
  wire Rgiow6;  // ../RTL/cortexm0ds_logic.v(1093)
  wire Rgnhu6;  // ../RTL/cortexm0ds_logic.v(145)
  wire Rgoiu6;  // ../RTL/cortexm0ds_logic.v(630)
  wire Rgphu6;  // ../RTL/cortexm0ds_logic.v(162)
  wire Rgpow6;  // ../RTL/cortexm0ds_logic.v(1187)
  wire Rgrax6;  // ../RTL/cortexm0ds_logic.v(1664)
  wire Rgviu6;  // ../RTL/cortexm0ds_logic.v(724)
  wire Rgwhu6;  // ../RTL/cortexm0ds_logic.v(256)
  wire Rgwow6;  // ../RTL/cortexm0ds_logic.v(1280)
  wire Rh1ju6;  // ../RTL/cortexm0ds_logic.v(805)
  wire Rh2iu6;  // ../RTL/cortexm0ds_logic.v(337)
  wire Rh2pw6;  // ../RTL/cortexm0ds_logic.v(1361)
  wire Rh8ju6;  // ../RTL/cortexm0ds_logic.v(898)
  wire Rh9iu6;  // ../RTL/cortexm0ds_logic.v(430)
  wire Rh9pw6;  // ../RTL/cortexm0ds_logic.v(1455)
  wire Rhaow6;  // ../RTL/cortexm0ds_logic.v(987)
  wire Rhgiu6;  // ../RTL/cortexm0ds_logic.v(524)
  wire Rhhow6;  // ../RTL/cortexm0ds_logic.v(1080)
  wire Rhibx6;  // ../RTL/cortexm0ds_logic.v(1713)
  wire Rhkpw6;  // ../RTL/cortexm0ds_logic.v(1588)
  wire Rhniu6;  // ../RTL/cortexm0ds_logic.v(617)
  wire Rhohu6;  // ../RTL/cortexm0ds_logic.v(149)
  wire Rhoow6;  // ../RTL/cortexm0ds_logic.v(1174)
  wire Rhuiu6;  // ../RTL/cortexm0ds_logic.v(711)
  wire Rhvhu6;  // ../RTL/cortexm0ds_logic.v(243)
  wire Rhvow6;  // ../RTL/cortexm0ds_logic.v(1267)
  wire Rhypw6;  // ../RTL/cortexm0ds_logic.v(1614)
  wire Ri0ju6;  // ../RTL/cortexm0ds_logic.v(792)
  wire Ri1iu6;  // ../RTL/cortexm0ds_logic.v(324)
  wire Ri1pw6;  // ../RTL/cortexm0ds_logic.v(1348)
  wire Ri7ju6;  // ../RTL/cortexm0ds_logic.v(885)
  wire Ri8iu6;  // ../RTL/cortexm0ds_logic.v(417)
  wire Ri8pw6;  // ../RTL/cortexm0ds_logic.v(1442)
  wire Ri9ow6;  // ../RTL/cortexm0ds_logic.v(974)
  wire Rifiu6;  // ../RTL/cortexm0ds_logic.v(511)
  wire Righu6;  // ../RTL/cortexm0ds_logic.v(126)
  wire Rigow6;  // ../RTL/cortexm0ds_logic.v(1067)
  wire Rijbx6;  // ../RTL/cortexm0ds_logic.v(1715)
  wire Rilpw6;  // ../RTL/cortexm0ds_logic.v(1590)
  wire Rimiu6;  // ../RTL/cortexm0ds_logic.v(604)
  wire Rinow6;  // ../RTL/cortexm0ds_logic.v(1161)
  wire Ritiu6;  // ../RTL/cortexm0ds_logic.v(698)
  wire Riuhu6;  // ../RTL/cortexm0ds_logic.v(230)
  wire Riuow6;  // ../RTL/cortexm0ds_logic.v(1254)
  wire Rj0iu6;  // ../RTL/cortexm0ds_logic.v(311)
  wire Rj0pw6;  // ../RTL/cortexm0ds_logic.v(1335)
  wire Rj6ju6;  // ../RTL/cortexm0ds_logic.v(872)
  wire Rj7iu6;  // ../RTL/cortexm0ds_logic.v(404)
  wire Rj7pw6;  // ../RTL/cortexm0ds_logic.v(1429)
  wire Rj8ow6;  // ../RTL/cortexm0ds_logic.v(961)
  wire Rjeiu6;  // ../RTL/cortexm0ds_logic.v(498)
  wire Rjfow6;  // ../RTL/cortexm0ds_logic.v(1054)
  wire Rjibx6;  // ../RTL/cortexm0ds_logic.v(1713)
  wire Rjliu6;  // ../RTL/cortexm0ds_logic.v(591)
  wire Rjmow6;  // ../RTL/cortexm0ds_logic.v(1148)
  wire Rjopw6;  // ../RTL/cortexm0ds_logic.v(1596)
  wire Rjsiu6;  // ../RTL/cortexm0ds_logic.v(685)
  wire Rjthu6;  // ../RTL/cortexm0ds_logic.v(217)
  wire Rjtow6;  // ../RTL/cortexm0ds_logic.v(1241)
  wire Rjziu6;  // ../RTL/cortexm0ds_logic.v(779)
  wire Rk1bx6;  // ../RTL/cortexm0ds_logic.v(1682)
  wire Rk5ju6;  // ../RTL/cortexm0ds_logic.v(859)
  wire Rk6iu6;  // ../RTL/cortexm0ds_logic.v(391)
  wire Rk6pw6;  // ../RTL/cortexm0ds_logic.v(1416)
  wire Rk7ow6;  // ../RTL/cortexm0ds_logic.v(948)
  wire Rkbax6;  // ../RTL/cortexm0ds_logic.v(1634)
  wire Rkdiu6;  // ../RTL/cortexm0ds_logic.v(485)
  wire Rkdpw6;  // ../RTL/cortexm0ds_logic.v(1509)
  wire Rkeow6;  // ../RTL/cortexm0ds_logic.v(1041)
  wire Rkkax6;  // ../RTL/cortexm0ds_logic.v(1651)
  wire Rkkiu6;  // ../RTL/cortexm0ds_logic.v(578)
  wire Rklow6;  // ../RTL/cortexm0ds_logic.v(1135)
  wire Rkriu6;  // ../RTL/cortexm0ds_logic.v(672)
  wire Rkshu6;  // ../RTL/cortexm0ds_logic.v(204)
  wire Rksow6;  // ../RTL/cortexm0ds_logic.v(1228)
  wire Rkyiu6;  // ../RTL/cortexm0ds_logic.v(766)
  wire Rkzhu6;  // ../RTL/cortexm0ds_logic.v(298)
  wire Rkzow6;  // ../RTL/cortexm0ds_logic.v(1322)
  wire Rl4ju6;  // ../RTL/cortexm0ds_logic.v(846)
  wire Rl5iu6;  // ../RTL/cortexm0ds_logic.v(378)
  wire Rl5pw6;  // ../RTL/cortexm0ds_logic.v(1403)
  wire Rl6ow6;  // ../RTL/cortexm0ds_logic.v(935)
  wire Rlciu6;  // ../RTL/cortexm0ds_logic.v(472)
  wire Rlcpw6;  // ../RTL/cortexm0ds_logic.v(1496)
  wire Rldow6;  // ../RTL/cortexm0ds_logic.v(1028)
  wire Rlgbx6;  // ../RTL/cortexm0ds_logic.v(1709)
  wire Rlibx6;  // ../RTL/cortexm0ds_logic.v(1713)
  wire Rljiu6;  // ../RTL/cortexm0ds_logic.v(565)
  wire Rlkow6;  // ../RTL/cortexm0ds_logic.v(1122)
  wire Rlqiu6;  // ../RTL/cortexm0ds_logic.v(659)
  wire Rlrhu6;  // ../RTL/cortexm0ds_logic.v(191)
  wire Rlrow6;  // ../RTL/cortexm0ds_logic.v(1215)
  wire Rlxiu6;  // ../RTL/cortexm0ds_logic.v(753)
  wire Rlyhu6;  // ../RTL/cortexm0ds_logic.v(285)
  wire Rlyow6;  // ../RTL/cortexm0ds_logic.v(1309)
  wire Rm2bx6;  // ../RTL/cortexm0ds_logic.v(1684)
  wire Rm3ju6;  // ../RTL/cortexm0ds_logic.v(833)
  wire Rm4iu6;  // ../RTL/cortexm0ds_logic.v(365)
  wire Rm4pw6;  // ../RTL/cortexm0ds_logic.v(1390)
  wire Rmaju6;  // ../RTL/cortexm0ds_logic.v(927)
  wire Rmbiu6;  // ../RTL/cortexm0ds_logic.v(459)
  wire Rmbpw6;  // ../RTL/cortexm0ds_logic.v(1483)
  wire Rmcow6;  // ../RTL/cortexm0ds_logic.v(1015)
  wire Rmiiu6;  // ../RTL/cortexm0ds_logic.v(552)
  wire Rmjow6;  // ../RTL/cortexm0ds_logic.v(1109)
  wire Rmpiu6;  // ../RTL/cortexm0ds_logic.v(646)
  wire Rmqhu6;  // ../RTL/cortexm0ds_logic.v(178)
  wire Rmqow6;  // ../RTL/cortexm0ds_logic.v(1202)
  wire Rmwiu6;  // ../RTL/cortexm0ds_logic.v(740)
  wire Rmxhu6;  // ../RTL/cortexm0ds_logic.v(272)
  wire Rmxow6;  // ../RTL/cortexm0ds_logic.v(1296)
  wire Rn2ju6;  // ../RTL/cortexm0ds_logic.v(820)
  wire Rn3iu6;  // ../RTL/cortexm0ds_logic.v(352)
  wire Rn3pw6;  // ../RTL/cortexm0ds_logic.v(1377)
  wire Rn9ju6;  // ../RTL/cortexm0ds_logic.v(914)
  wire Rnaax6;  // ../RTL/cortexm0ds_logic.v(1632)
  wire Rnaiu6;  // ../RTL/cortexm0ds_logic.v(446)
  wire Rnapw6;  // ../RTL/cortexm0ds_logic.v(1470)
  wire Rnbow6;  // ../RTL/cortexm0ds_logic.v(1002)
  wire Rnhiu6;  // ../RTL/cortexm0ds_logic.v(539)
  wire Rnibx6;  // ../RTL/cortexm0ds_logic.v(1713)
  wire Rniow6;  // ../RTL/cortexm0ds_logic.v(1096)
  wire Rnoiu6;  // ../RTL/cortexm0ds_logic.v(633)
  wire Rnphu6;  // ../RTL/cortexm0ds_logic.v(165)
  wire Rnpow6;  // ../RTL/cortexm0ds_logic.v(1189)
  wire Rnvax6;  // ../RTL/cortexm0ds_logic.v(1672)
  wire Rnviu6;  // ../RTL/cortexm0ds_logic.v(727)
  wire Rnwhu6;  // ../RTL/cortexm0ds_logic.v(259)
  wire Rnwow6;  // ../RTL/cortexm0ds_logic.v(1283)
  wire Ro1ju6;  // ../RTL/cortexm0ds_logic.v(807)
  wire Ro2iu6;  // ../RTL/cortexm0ds_logic.v(339)
  wire Ro2pw6;  // ../RTL/cortexm0ds_logic.v(1364)
  wire Ro8ax6;  // ../RTL/cortexm0ds_logic.v(1629)
  wire Ro8ju6;  // ../RTL/cortexm0ds_logic.v(901)
  wire Ro9iu6;  // ../RTL/cortexm0ds_logic.v(433)
  wire Ro9pw6;  // ../RTL/cortexm0ds_logic.v(1457)
  wire Roaow6;  // ../RTL/cortexm0ds_logic.v(989)
  wire Rogiu6;  // ../RTL/cortexm0ds_logic.v(526)
  wire Rohow6;  // ../RTL/cortexm0ds_logic.v(1083)
  wire Romhu6;  // ../RTL/cortexm0ds_logic.v(143)
  wire Roniu6;  // ../RTL/cortexm0ds_logic.v(620)
  wire Roohu6;  // ../RTL/cortexm0ds_logic.v(152)
  wire Rooow6;  // ../RTL/cortexm0ds_logic.v(1176)
  wire Rouiu6;  // ../RTL/cortexm0ds_logic.v(714)
  wire Rovhu6;  // ../RTL/cortexm0ds_logic.v(246)
  wire Rovow6;  // ../RTL/cortexm0ds_logic.v(1270)
  wire Rp0ju6;  // ../RTL/cortexm0ds_logic.v(794)
  wire Rp1iu6;  // ../RTL/cortexm0ds_logic.v(326)
  wire Rp1pw6;  // ../RTL/cortexm0ds_logic.v(1351)
  wire Rp7ju6;  // ../RTL/cortexm0ds_logic.v(888)
  wire Rp8iu6;  // ../RTL/cortexm0ds_logic.v(420)
  wire Rp8pw6;  // ../RTL/cortexm0ds_logic.v(1444)
  wire Rp9ow6;  // ../RTL/cortexm0ds_logic.v(976)
  wire Rpfiu6;  // ../RTL/cortexm0ds_logic.v(513)
  wire Rpgow6;  // ../RTL/cortexm0ds_logic.v(1070)
  wire Rpibx6;  // ../RTL/cortexm0ds_logic.v(1713)
  wire Rpmiu6;  // ../RTL/cortexm0ds_logic.v(607)
  wire Rpnow6;  // ../RTL/cortexm0ds_logic.v(1163)
  wire Rptiu6;  // ../RTL/cortexm0ds_logic.v(701)
  wire Rpuhu6;  // ../RTL/cortexm0ds_logic.v(233)
  wire Rpuow6;  // ../RTL/cortexm0ds_logic.v(1257)
  wire Rpvax6;  // ../RTL/cortexm0ds_logic.v(1672)
  wire Rq0iu6;  // ../RTL/cortexm0ds_logic.v(313)
  wire Rq0pw6;  // ../RTL/cortexm0ds_logic.v(1338)
  wire Rq0qw6;  // ../RTL/cortexm0ds_logic.v(1618)
  wire Rq6ju6;  // ../RTL/cortexm0ds_logic.v(875)
  wire Rq7iu6;  // ../RTL/cortexm0ds_logic.v(407)
  wire Rq7pw6;  // ../RTL/cortexm0ds_logic.v(1431)
  wire Rq8ow6;  // ../RTL/cortexm0ds_logic.v(963)
  wire Rqeiu6;  // ../RTL/cortexm0ds_logic.v(500)
  wire Rqfow6;  // ../RTL/cortexm0ds_logic.v(1057)
  wire Rqliu6;  // ../RTL/cortexm0ds_logic.v(594)
  wire Rqmow6;  // ../RTL/cortexm0ds_logic.v(1150)
  wire Rqsiu6;  // ../RTL/cortexm0ds_logic.v(688)
  wire Rqthu6;  // ../RTL/cortexm0ds_logic.v(220)
  wire Rqtow6;  // ../RTL/cortexm0ds_logic.v(1244)
  wire Rqziu6;  // ../RTL/cortexm0ds_logic.v(781)
  wire Rr3qw6;  // ../RTL/cortexm0ds_logic.v(1624)
  wire Rr5ju6;  // ../RTL/cortexm0ds_logic.v(862)
  wire Rr6iu6;  // ../RTL/cortexm0ds_logic.v(394)
  wire Rr6pw6;  // ../RTL/cortexm0ds_logic.v(1418)
  wire Rr7ow6;  // ../RTL/cortexm0ds_logic.v(950)
  wire Rrdiu6;  // ../RTL/cortexm0ds_logic.v(487)
  wire Rrdpw6;  // ../RTL/cortexm0ds_logic.v(1512)
  wire Rreow6;  // ../RTL/cortexm0ds_logic.v(1044)
  wire Rribx6;  // ../RTL/cortexm0ds_logic.v(1713)
  wire Rrkiu6;  // ../RTL/cortexm0ds_logic.v(581)
  wire Rrlhu6;  // ../RTL/cortexm0ds_logic.v(140)
  wire Rrlow6;  // ../RTL/cortexm0ds_logic.v(1137)
  wire Rrnhu6;  // ../RTL/cortexm0ds_logic.v(145)
  wire Rrriu6;  // ../RTL/cortexm0ds_logic.v(675)
  wire Rrshu6;  // ../RTL/cortexm0ds_logic.v(207)
  wire Rrsow6;  // ../RTL/cortexm0ds_logic.v(1231)
  wire Rrvax6;  // ../RTL/cortexm0ds_logic.v(1672)
  wire Rryiu6;  // ../RTL/cortexm0ds_logic.v(768)
  wire Rrzhu6;  // ../RTL/cortexm0ds_logic.v(300)
  wire Rrzow6;  // ../RTL/cortexm0ds_logic.v(1325)
  wire Rs4ju6;  // ../RTL/cortexm0ds_logic.v(849)
  wire Rs5iu6;  // ../RTL/cortexm0ds_logic.v(381)
  wire Rs5pw6;  // ../RTL/cortexm0ds_logic.v(1405)
  wire Rs6ow6;  // ../RTL/cortexm0ds_logic.v(937)
  wire Rsciu6;  // ../RTL/cortexm0ds_logic.v(474)
  wire Rscpw6;  // ../RTL/cortexm0ds_logic.v(1499)
  wire Rsdow6;  // ../RTL/cortexm0ds_logic.v(1031)
  wire Rsjiu6;  // ../RTL/cortexm0ds_logic.v(568)
  wire Rskax6;  // ../RTL/cortexm0ds_logic.v(1652)
  wire Rskow6;  // ../RTL/cortexm0ds_logic.v(1124)
  wire Rsqiu6;  // ../RTL/cortexm0ds_logic.v(662)
  wire Rsrhu6;  // ../RTL/cortexm0ds_logic.v(194)
  wire Rsrow6;  // ../RTL/cortexm0ds_logic.v(1218)
  wire Rsxiu6;  // ../RTL/cortexm0ds_logic.v(755)
  wire Rsyhu6;  // ../RTL/cortexm0ds_logic.v(287)
  wire Rsyow6;  // ../RTL/cortexm0ds_logic.v(1312)
  wire Rt3ju6;  // ../RTL/cortexm0ds_logic.v(836)
  wire Rt4iu6;  // ../RTL/cortexm0ds_logic.v(368)
  wire Rt4pw6;  // ../RTL/cortexm0ds_logic.v(1392)
  wire Rtbiu6;  // ../RTL/cortexm0ds_logic.v(461)
  wire Rtbpw6;  // ../RTL/cortexm0ds_logic.v(1486)
  wire Rtcow6;  // ../RTL/cortexm0ds_logic.v(1018)
  wire Rteax6;  // ../RTL/cortexm0ds_logic.v(1641)
  wire Rthhu6;  // ../RTL/cortexm0ds_logic.v(129)
  wire Rtibx6;  // ../RTL/cortexm0ds_logic.v(1713)
  wire Rtiiu6;  // ../RTL/cortexm0ds_logic.v(555)
  wire Rtjow6;  // ../RTL/cortexm0ds_logic.v(1111)
  wire Rtpiu6;  // ../RTL/cortexm0ds_logic.v(649)
  wire Rtqhu6;  // ../RTL/cortexm0ds_logic.v(181)
  wire Rtqow6;  // ../RTL/cortexm0ds_logic.v(1205)
  wire Rtvax6;  // ../RTL/cortexm0ds_logic.v(1672)
  wire Rtwiu6;  // ../RTL/cortexm0ds_logic.v(742)
  wire Rtxhu6;  // ../RTL/cortexm0ds_logic.v(274)
  wire Rtxow6;  // ../RTL/cortexm0ds_logic.v(1299)
  wire Ru2ju6;  // ../RTL/cortexm0ds_logic.v(823)
  wire Ru3iu6;  // ../RTL/cortexm0ds_logic.v(355)
  wire Ru3pw6;  // ../RTL/cortexm0ds_logic.v(1379)
  wire Ru9ju6;  // ../RTL/cortexm0ds_logic.v(916)
  wire Ruaiu6;  // ../RTL/cortexm0ds_logic.v(448)
  wire Ruapw6;  // ../RTL/cortexm0ds_logic.v(1473)
  wire Rubow6;  // ../RTL/cortexm0ds_logic.v(1005)
  wire Rucax6;  // ../RTL/cortexm0ds_logic.v(1637)
  wire Ruhiu6;  // ../RTL/cortexm0ds_logic.v(542)
  wire Ruiow6;  // ../RTL/cortexm0ds_logic.v(1098)
  wire Ruoiu6;  // ../RTL/cortexm0ds_logic.v(636)
  wire Ruphu6;  // ../RTL/cortexm0ds_logic.v(168)
  wire Rupow6;  // ../RTL/cortexm0ds_logic.v(1192)
  wire Ruviu6;  // ../RTL/cortexm0ds_logic.v(729)
  wire Ruwhu6;  // ../RTL/cortexm0ds_logic.v(261)
  wire Ruwow6;  // ../RTL/cortexm0ds_logic.v(1286)
  wire Rv1ju6;  // ../RTL/cortexm0ds_logic.v(810)
  wire Rv2iu6;  // ../RTL/cortexm0ds_logic.v(342)
  wire Rv2pw6;  // ../RTL/cortexm0ds_logic.v(1366)
  wire Rv7ax6;  // ../RTL/cortexm0ds_logic.v(1627)
  wire Rv8ju6;  // ../RTL/cortexm0ds_logic.v(903)
  wire Rv9iu6;  // ../RTL/cortexm0ds_logic.v(435)
  wire Rv9pw6;  // ../RTL/cortexm0ds_logic.v(1460)
  wire Rvaow6;  // ../RTL/cortexm0ds_logic.v(992)
  wire Rvgiu6;  // ../RTL/cortexm0ds_logic.v(529)
  wire Rvhow6;  // ../RTL/cortexm0ds_logic.v(1085)
  wire Rvibx6;  // ../RTL/cortexm0ds_logic.v(1713)
  wire Rvniu6;  // ../RTL/cortexm0ds_logic.v(623)
  wire Rvohu6;  // ../RTL/cortexm0ds_logic.v(155)
  wire Rvoow6;  // ../RTL/cortexm0ds_logic.v(1179)
  wire Rvuiu6;  // ../RTL/cortexm0ds_logic.v(716)
  wire Rvvhu6;  // ../RTL/cortexm0ds_logic.v(248)
  wire Rvvow6;  // ../RTL/cortexm0ds_logic.v(1273)
  wire Rw0ju6;  // ../RTL/cortexm0ds_logic.v(797)
  wire Rw1iu6;  // ../RTL/cortexm0ds_logic.v(329)
  wire Rw1pw6;  // ../RTL/cortexm0ds_logic.v(1353)
  wire Rw7ju6;  // ../RTL/cortexm0ds_logic.v(890)
  wire Rw8iu6;  // ../RTL/cortexm0ds_logic.v(422)
  wire Rw8pw6;  // ../RTL/cortexm0ds_logic.v(1447)
  wire Rw9ow6;  // ../RTL/cortexm0ds_logic.v(979)
  wire Rwfiu6;  // ../RTL/cortexm0ds_logic.v(516)
  wire Rwgow6;  // ../RTL/cortexm0ds_logic.v(1072)
  wire Rwhax6;  // ../RTL/cortexm0ds_logic.v(1647)
  wire Rwjax6;  // ../RTL/cortexm0ds_logic.v(1650)
  wire Rwmiu6;  // ../RTL/cortexm0ds_logic.v(610)
  wire Rwnow6;  // ../RTL/cortexm0ds_logic.v(1166)
  wire Rwtiu6;  // ../RTL/cortexm0ds_logic.v(703)
  wire Rwuhu6;  // ../RTL/cortexm0ds_logic.v(235)
  wire Rwuow6;  // ../RTL/cortexm0ds_logic.v(1260)
  wire Rx0iu6;  // ../RTL/cortexm0ds_logic.v(316)
  wire Rx0pw6;  // ../RTL/cortexm0ds_logic.v(1340)
  wire Rx6ju6;  // ../RTL/cortexm0ds_logic.v(877)
  wire Rx7iu6;  // ../RTL/cortexm0ds_logic.v(409)
  wire Rx7pw6;  // ../RTL/cortexm0ds_logic.v(1434)
  wire Rx8ow6;  // ../RTL/cortexm0ds_logic.v(966)
  wire Rxeiu6;  // ../RTL/cortexm0ds_logic.v(503)
  wire Rxfow6;  // ../RTL/cortexm0ds_logic.v(1059)
  wire Rxliu6;  // ../RTL/cortexm0ds_logic.v(597)
  wire Rxmow6;  // ../RTL/cortexm0ds_logic.v(1153)
  wire Rxsiu6;  // ../RTL/cortexm0ds_logic.v(690)
  wire Rxthu6;  // ../RTL/cortexm0ds_logic.v(222)
  wire Rxtow6;  // ../RTL/cortexm0ds_logic.v(1247)
  wire Rxziu6;  // ../RTL/cortexm0ds_logic.v(784)
  wire Ry0qw6;  // ../RTL/cortexm0ds_logic.v(1619)
  wire Ry2qw6;  // ../RTL/cortexm0ds_logic.v(1622)
  wire Ry5ju6;  // ../RTL/cortexm0ds_logic.v(864)
  wire Ry6iu6;  // ../RTL/cortexm0ds_logic.v(396)
  wire Ry6pw6;  // ../RTL/cortexm0ds_logic.v(1421)
  wire Ry7ow6;  // ../RTL/cortexm0ds_logic.v(953)
  wire Rydiu6;  // ../RTL/cortexm0ds_logic.v(490)
  wire Rydpw6;  // ../RTL/cortexm0ds_logic.v(1514)
  wire Ryeow6;  // ../RTL/cortexm0ds_logic.v(1046)
  wire Ryfax6;  // ../RTL/cortexm0ds_logic.v(1643)
  wire Rykiu6;  // ../RTL/cortexm0ds_logic.v(584)
  wire Rylow6;  // ../RTL/cortexm0ds_logic.v(1140)
  wire Ryriu6;  // ../RTL/cortexm0ds_logic.v(677)
  wire Ryshu6;  // ../RTL/cortexm0ds_logic.v(209)
  wire Rysow6;  // ../RTL/cortexm0ds_logic.v(1234)
  wire Ryyiu6;  // ../RTL/cortexm0ds_logic.v(771)
  wire Ryzhu6;  // ../RTL/cortexm0ds_logic.v(303)
  wire Ryzow6;  // ../RTL/cortexm0ds_logic.v(1327)
  wire Rz0bx6;  // ../RTL/cortexm0ds_logic.v(1681)
  wire Rz4ju6;  // ../RTL/cortexm0ds_logic.v(851)
  wire Rz5iu6;  // ../RTL/cortexm0ds_logic.v(383)
  wire Rz5pw6;  // ../RTL/cortexm0ds_logic.v(1408)
  wire Rz6ow6;  // ../RTL/cortexm0ds_logic.v(940)
  wire Rz8bx6;  // ../RTL/cortexm0ds_logic.v(1695)
  wire Rzciu6;  // ../RTL/cortexm0ds_logic.v(477)
  wire Rzcpw6;  // ../RTL/cortexm0ds_logic.v(1501)
  wire Rzdow6;  // ../RTL/cortexm0ds_logic.v(1033)
  wire Rzjiu6;  // ../RTL/cortexm0ds_logic.v(571)
  wire Rzkow6;  // ../RTL/cortexm0ds_logic.v(1127)
  wire Rzqiu6;  // ../RTL/cortexm0ds_logic.v(664)
  wire Rzrhu6;  // ../RTL/cortexm0ds_logic.v(196)
  wire Rzrow6;  // ../RTL/cortexm0ds_logic.v(1221)
  wire Rzxiu6;  // ../RTL/cortexm0ds_logic.v(758)
  wire Rzyhu6;  // ../RTL/cortexm0ds_logic.v(290)
  wire Rzyow6;  // ../RTL/cortexm0ds_logic.v(1314)
  wire S01ju6;  // ../RTL/cortexm0ds_logic.v(798)
  wire S02iu6;  // ../RTL/cortexm0ds_logic.v(330)
  wire S02pw6;  // ../RTL/cortexm0ds_logic.v(1355)
  wire S08ju6;  // ../RTL/cortexm0ds_logic.v(892)
  wire S09iu6;  // ../RTL/cortexm0ds_logic.v(424)
  wire S09pw6;  // ../RTL/cortexm0ds_logic.v(1448)
  wire S0aow6;  // ../RTL/cortexm0ds_logic.v(980)
  wire S0giu6;  // ../RTL/cortexm0ds_logic.v(518)
  wire S0how6;  // ../RTL/cortexm0ds_logic.v(1074)
  wire S0kbx6;  // ../RTL/cortexm0ds_logic.v(1716)
  wire S0lhu6;  // ../RTL/cortexm0ds_logic.v(138)
  wire S0niu6;  // ../RTL/cortexm0ds_logic.v(611)
  wire S0oow6;  // ../RTL/cortexm0ds_logic.v(1168)
  wire S0uiu6;  // ../RTL/cortexm0ds_logic.v(705)
  wire S0vhu6;  // ../RTL/cortexm0ds_logic.v(237)
  wire S0vow6;  // ../RTL/cortexm0ds_logic.v(1261)
  wire S10ju6;  // ../RTL/cortexm0ds_logic.v(785)
  wire S11bx6;  // ../RTL/cortexm0ds_logic.v(1681)
  wire S11iu6;  // ../RTL/cortexm0ds_logic.v(317)
  wire S11pw6;  // ../RTL/cortexm0ds_logic.v(1342)
  wire S17ju6;  // ../RTL/cortexm0ds_logic.v(879)
  wire S18ax6;  // ../RTL/cortexm0ds_logic.v(1627)
  wire S18iu6;  // ../RTL/cortexm0ds_logic.v(411)
  wire S18pw6;  // ../RTL/cortexm0ds_logic.v(1435)
  wire S19ow6;  // ../RTL/cortexm0ds_logic.v(967)
  wire S1ehu6;  // ../RTL/cortexm0ds_logic.v(121)
  wire S1fiu6;  // ../RTL/cortexm0ds_logic.v(505)
  wire S1gow6;  // ../RTL/cortexm0ds_logic.v(1061)
  wire S1miu6;  // ../RTL/cortexm0ds_logic.v(598)
  wire S1nax6;  // ../RTL/cortexm0ds_logic.v(1656)
  wire S1now6;  // ../RTL/cortexm0ds_logic.v(1155)
  wire S1tiu6;  // ../RTL/cortexm0ds_logic.v(692)
  wire S1uhu6;  // ../RTL/cortexm0ds_logic.v(224)
  wire S1uow6;  // ../RTL/cortexm0ds_logic.v(1248)
  wire S20iu6;  // ../RTL/cortexm0ds_logic.v(304)
  wire S20pw6;  // ../RTL/cortexm0ds_logic.v(1329)
  wire S26ju6;  // ../RTL/cortexm0ds_logic.v(866)
  wire S27iu6;  // ../RTL/cortexm0ds_logic.v(398)
  wire S27pw6;  // ../RTL/cortexm0ds_logic.v(1422)
  wire S28ow6;  // ../RTL/cortexm0ds_logic.v(954)
  wire S2cax6;  // ../RTL/cortexm0ds_logic.v(1635)
  wire S2cbx6;  // ../RTL/cortexm0ds_logic.v(1701)
  wire S2eiu6;  // ../RTL/cortexm0ds_logic.v(492)
  wire S2epw6;  // ../RTL/cortexm0ds_logic.v(1516)
  wire S2fow6;  // ../RTL/cortexm0ds_logic.v(1048)
  wire S2khu6;  // ../RTL/cortexm0ds_logic.v(135)
  wire S2liu6;  // ../RTL/cortexm0ds_logic.v(585)
  wire S2mow6;  // ../RTL/cortexm0ds_logic.v(1142)
  wire S2siu6;  // ../RTL/cortexm0ds_logic.v(679)
  wire S2thu6;  // ../RTL/cortexm0ds_logic.v(211)
  wire S2tow6;  // ../RTL/cortexm0ds_logic.v(1235)
  wire S2ziu6;  // ../RTL/cortexm0ds_logic.v(772)
  wire S32bx6;  // ../RTL/cortexm0ds_logic.v(1683)
  wire S35ju6;  // ../RTL/cortexm0ds_logic.v(853)
  wire S36iu6;  // ../RTL/cortexm0ds_logic.v(385)
  wire S36pw6;  // ../RTL/cortexm0ds_logic.v(1409)
  wire S37ow6;  // ../RTL/cortexm0ds_logic.v(941)
  wire S38ax6;  // ../RTL/cortexm0ds_logic.v(1628)
  wire S3diu6;  // ../RTL/cortexm0ds_logic.v(479)
  wire S3dpw6;  // ../RTL/cortexm0ds_logic.v(1503)
  wire S3eow6;  // ../RTL/cortexm0ds_logic.v(1035)
  wire S3hhu6;  // ../RTL/cortexm0ds_logic.v(127)
  wire S3kiu6;  // ../RTL/cortexm0ds_logic.v(572)
  wire S3low6;  // ../RTL/cortexm0ds_logic.v(1129)
  wire S3mpw6;  // ../RTL/cortexm0ds_logic.v(1592)
  wire S3nax6;  // ../RTL/cortexm0ds_logic.v(1656)
  wire S3ohu6;  // ../RTL/cortexm0ds_logic.v(146)
  wire S3riu6;  // ../RTL/cortexm0ds_logic.v(666)
  wire S3shu6;  // ../RTL/cortexm0ds_logic.v(198)
  wire S3sow6;  // ../RTL/cortexm0ds_logic.v(1222)
  wire S3yiu6;  // ../RTL/cortexm0ds_logic.v(759)
  wire S3zhu6;  // ../RTL/cortexm0ds_logic.v(291)
  wire S3zow6;  // ../RTL/cortexm0ds_logic.v(1316)
  wire S44ju6;  // ../RTL/cortexm0ds_logic.v(840)
  wire S45iu6;  // ../RTL/cortexm0ds_logic.v(372)
  wire S45pw6;  // ../RTL/cortexm0ds_logic.v(1396)
  wire S4ciu6;  // ../RTL/cortexm0ds_logic.v(466)
  wire S4cpw6;  // ../RTL/cortexm0ds_logic.v(1490)
  wire S4dow6;  // ../RTL/cortexm0ds_logic.v(1022)
  wire S4jhu6;  // ../RTL/cortexm0ds_logic.v(133)
  wire S4jiu6;  // ../RTL/cortexm0ds_logic.v(559)
  wire S4kbx6;  // ../RTL/cortexm0ds_logic.v(1716)
  wire S4kow6;  // ../RTL/cortexm0ds_logic.v(1116)
  wire S4qiu6;  // ../RTL/cortexm0ds_logic.v(653)
  wire S4rhu6;  // ../RTL/cortexm0ds_logic.v(185)
  wire S4row6;  // ../RTL/cortexm0ds_logic.v(1209)
  wire S4xiu6;  // ../RTL/cortexm0ds_logic.v(746)
  wire S4yhu6;  // ../RTL/cortexm0ds_logic.v(278)
  wire S4yow6;  // ../RTL/cortexm0ds_logic.v(1303)
  wire S53bx6;  // ../RTL/cortexm0ds_logic.v(1685)
  wire S53ju6;  // ../RTL/cortexm0ds_logic.v(827)
  wire S54iu6;  // ../RTL/cortexm0ds_logic.v(359)
  wire S54pw6;  // ../RTL/cortexm0ds_logic.v(1383)
  wire S58ax6;  // ../RTL/cortexm0ds_logic.v(1628)
  wire S5aju6;  // ../RTL/cortexm0ds_logic.v(921)
  wire S5biu6;  // ../RTL/cortexm0ds_logic.v(453)
  wire S5bpw6;  // ../RTL/cortexm0ds_logic.v(1477)
  wire S5cow6;  // ../RTL/cortexm0ds_logic.v(1009)
  wire S5iiu6;  // ../RTL/cortexm0ds_logic.v(546)
  wire S5jow6;  // ../RTL/cortexm0ds_logic.v(1103)
  wire S5kpw6;  // ../RTL/cortexm0ds_logic.v(1588)
  wire S5nax6;  // ../RTL/cortexm0ds_logic.v(1656)
  wire S5piu6;  // ../RTL/cortexm0ds_logic.v(640)
  wire S5qhu6;  // ../RTL/cortexm0ds_logic.v(172)
  wire S5qow6;  // ../RTL/cortexm0ds_logic.v(1196)
  wire S5wiu6;  // ../RTL/cortexm0ds_logic.v(733)
  wire S5xhu6;  // ../RTL/cortexm0ds_logic.v(265)
  wire S5xow6;  // ../RTL/cortexm0ds_logic.v(1290)
  wire S62ju6;  // ../RTL/cortexm0ds_logic.v(814)
  wire S63iu6;  // ../RTL/cortexm0ds_logic.v(346)
  wire S63pw6;  // ../RTL/cortexm0ds_logic.v(1370)
  wire S69ju6;  // ../RTL/cortexm0ds_logic.v(908)
  wire S6aiu6;  // ../RTL/cortexm0ds_logic.v(440)
  wire S6apw6;  // ../RTL/cortexm0ds_logic.v(1464)
  wire S6bow6;  // ../RTL/cortexm0ds_logic.v(996)
  wire S6hiu6;  // ../RTL/cortexm0ds_logic.v(533)
  wire S6ihu6;  // ../RTL/cortexm0ds_logic.v(130)
  wire S6iow6;  // ../RTL/cortexm0ds_logic.v(1090)
  wire S6oiu6;  // ../RTL/cortexm0ds_logic.v(627)
  wire S6phu6;  // ../RTL/cortexm0ds_logic.v(159)
  wire S6pow6;  // ../RTL/cortexm0ds_logic.v(1183)
  wire S6viu6;  // ../RTL/cortexm0ds_logic.v(720)
  wire S6whu6;  // ../RTL/cortexm0ds_logic.v(252)
  wire S6wow6;  // ../RTL/cortexm0ds_logic.v(1277)
  wire S71ju6;  // ../RTL/cortexm0ds_logic.v(801)
  wire S72iu6;  // ../RTL/cortexm0ds_logic.v(333)
  wire S72pw6;  // ../RTL/cortexm0ds_logic.v(1357)
  wire S78ax6;  // ../RTL/cortexm0ds_logic.v(1628)
  wire S78ju6;  // ../RTL/cortexm0ds_logic.v(895)
  wire S79iu6;  // ../RTL/cortexm0ds_logic.v(427)
  wire S79pw6;  // ../RTL/cortexm0ds_logic.v(1451)
  wire S7aow6;  // ../RTL/cortexm0ds_logic.v(983)
  wire S7giu6;  // ../RTL/cortexm0ds_logic.v(520)
  wire S7how6;  // ../RTL/cortexm0ds_logic.v(1077)
  wire S7mpw6;  // ../RTL/cortexm0ds_logic.v(1592)
  wire S7niu6;  // ../RTL/cortexm0ds_logic.v(614)
  wire S7oow6;  // ../RTL/cortexm0ds_logic.v(1170)
  wire S7uiu6;  // ../RTL/cortexm0ds_logic.v(707)
  wire S7vhu6;  // ../RTL/cortexm0ds_logic.v(239)
  wire S7vow6;  // ../RTL/cortexm0ds_logic.v(1264)
  wire S7yax6;  // ../RTL/cortexm0ds_logic.v(1676)
  wire S80ju6;  // ../RTL/cortexm0ds_logic.v(788)
  wire S81iu6;  // ../RTL/cortexm0ds_logic.v(320)
  wire S81pw6;  // ../RTL/cortexm0ds_logic.v(1344)
  wire S87ju6;  // ../RTL/cortexm0ds_logic.v(882)
  wire S88iu6;  // ../RTL/cortexm0ds_logic.v(414)
  wire S88pw6;  // ../RTL/cortexm0ds_logic.v(1438)
  wire S89ow6;  // ../RTL/cortexm0ds_logic.v(970)
  wire S8fiu6;  // ../RTL/cortexm0ds_logic.v(507)
  wire S8gow6;  // ../RTL/cortexm0ds_logic.v(1064)
  wire S8miu6;  // ../RTL/cortexm0ds_logic.v(601)
  wire S8now6;  // ../RTL/cortexm0ds_logic.v(1157)
  wire S8tiu6;  // ../RTL/cortexm0ds_logic.v(694)
  wire S8uhu6;  // ../RTL/cortexm0ds_logic.v(226)
  wire S8uow6;  // ../RTL/cortexm0ds_logic.v(1251)
  wire S90iu6;  // ../RTL/cortexm0ds_logic.v(307)
  wire S90pw6;  // ../RTL/cortexm0ds_logic.v(1331)
  wire S96ju6;  // ../RTL/cortexm0ds_logic.v(869)
  wire S97iu6;  // ../RTL/cortexm0ds_logic.v(401)
  wire S97pw6;  // ../RTL/cortexm0ds_logic.v(1425)
  wire S98ax6;  // ../RTL/cortexm0ds_logic.v(1628)
  wire S98ow6;  // ../RTL/cortexm0ds_logic.v(957)
  wire S9eiu6;  // ../RTL/cortexm0ds_logic.v(494)
  wire S9fow6;  // ../RTL/cortexm0ds_logic.v(1051)
  wire S9liu6;  // ../RTL/cortexm0ds_logic.v(588)
  wire S9mow6;  // ../RTL/cortexm0ds_logic.v(1144)
  wire S9siu6;  // ../RTL/cortexm0ds_logic.v(681)
  wire S9thu6;  // ../RTL/cortexm0ds_logic.v(213)
  wire S9tow6;  // ../RTL/cortexm0ds_logic.v(1238)
  wire S9ziu6;  // ../RTL/cortexm0ds_logic.v(775)
  wire Sa5ju6;  // ../RTL/cortexm0ds_logic.v(856)
  wire Sa6iu6;  // ../RTL/cortexm0ds_logic.v(388)
  wire Sa6pw6;  // ../RTL/cortexm0ds_logic.v(1412)
  wire Sa7ow6;  // ../RTL/cortexm0ds_logic.v(944)
  wire Sadiu6;  // ../RTL/cortexm0ds_logic.v(481)
  wire Sadpw6;  // ../RTL/cortexm0ds_logic.v(1506)
  wire Saeow6;  // ../RTL/cortexm0ds_logic.v(1038)
  wire Sakiu6;  // ../RTL/cortexm0ds_logic.v(575)
  wire Salow6;  // ../RTL/cortexm0ds_logic.v(1131)
  wire Samhu6;  // ../RTL/cortexm0ds_logic.v(142)
  wire Sariu6;  // ../RTL/cortexm0ds_logic.v(668)
  wire Sashu6;  // ../RTL/cortexm0ds_logic.v(200)
  wire Sasow6;  // ../RTL/cortexm0ds_logic.v(1225)
  wire Sayiu6;  // ../RTL/cortexm0ds_logic.v(762)
  wire Sazhu6;  // ../RTL/cortexm0ds_logic.v(294)
  wire Sazow6;  // ../RTL/cortexm0ds_logic.v(1318)
  wire Sb4ju6;  // ../RTL/cortexm0ds_logic.v(843)
  wire Sb5iu6;  // ../RTL/cortexm0ds_logic.v(375)
  wire Sb5pw6;  // ../RTL/cortexm0ds_logic.v(1399)
  wire Sb6ow6;  // ../RTL/cortexm0ds_logic.v(931)
  wire Sb8ax6;  // ../RTL/cortexm0ds_logic.v(1628)
  wire Sbciu6;  // ../RTL/cortexm0ds_logic.v(468)
  wire Sbcpw6;  // ../RTL/cortexm0ds_logic.v(1493)
  wire Sbdow6;  // ../RTL/cortexm0ds_logic.v(1025)
  wire Sbfax6;  // ../RTL/cortexm0ds_logic.v(1642)
  wire Sbghu6;  // ../RTL/cortexm0ds_logic.v(126)
  wire Sbjiu6;  // ../RTL/cortexm0ds_logic.v(562)
  wire Sbkow6;  // ../RTL/cortexm0ds_logic.v(1118)
  wire Sbqiu6;  // ../RTL/cortexm0ds_logic.v(655)
  wire Sbrhu6;  // ../RTL/cortexm0ds_logic.v(187)
  wire Sbrow6;  // ../RTL/cortexm0ds_logic.v(1212)
  wire Sbxiu6;  // ../RTL/cortexm0ds_logic.v(749)
  wire Sbyax6;  // ../RTL/cortexm0ds_logic.v(1676)
  wire Sbyhu6;  // ../RTL/cortexm0ds_logic.v(281)
  wire Sbyow6;  // ../RTL/cortexm0ds_logic.v(1305)
  wire Sc3ju6;  // ../RTL/cortexm0ds_logic.v(830)
  wire Sc4iu6;  // ../RTL/cortexm0ds_logic.v(362)
  wire Sc4pw6;  // ../RTL/cortexm0ds_logic.v(1386)
  wire Scaju6;  // ../RTL/cortexm0ds_logic.v(923)
  wire Scbiu6;  // ../RTL/cortexm0ds_logic.v(455)
  wire Scbpw6;  // ../RTL/cortexm0ds_logic.v(1480)
  wire Sccow6;  // ../RTL/cortexm0ds_logic.v(1012)
  wire Sciiu6;  // ../RTL/cortexm0ds_logic.v(549)
  wire Scjow6;  // ../RTL/cortexm0ds_logic.v(1105)
  wire Scpiu6;  // ../RTL/cortexm0ds_logic.v(642)
  wire Scqhu6;  // ../RTL/cortexm0ds_logic.v(174)
  wire Scqow6;  // ../RTL/cortexm0ds_logic.v(1199)
  wire Scwiu6;  // ../RTL/cortexm0ds_logic.v(736)
  wire Scxhu6;  // ../RTL/cortexm0ds_logic.v(268)
  wire Scxow6;  // ../RTL/cortexm0ds_logic.v(1292)
  wire Sd2ju6;  // ../RTL/cortexm0ds_logic.v(817)
  wire Sd3iu6;  // ../RTL/cortexm0ds_logic.v(349)
  wire Sd3pw6;  // ../RTL/cortexm0ds_logic.v(1373)
  wire Sd8ax6;  // ../RTL/cortexm0ds_logic.v(1628)
  wire Sd9ju6;  // ../RTL/cortexm0ds_logic.v(910)
  wire Sdaiu6;  // ../RTL/cortexm0ds_logic.v(442)
  wire Sdapw6;  // ../RTL/cortexm0ds_logic.v(1467)
  wire Sdbow6;  // ../RTL/cortexm0ds_logic.v(999)
  wire Sddbx6;  // ../RTL/cortexm0ds_logic.v(1703)
  wire Sdhiu6;  // ../RTL/cortexm0ds_logic.v(536)
  wire Sdiow6;  // ../RTL/cortexm0ds_logic.v(1092)
  wire Sdlhu6;  // ../RTL/cortexm0ds_logic.v(139)
  wire Sdlpw6;  // ../RTL/cortexm0ds_logic.v(1590)
  wire Sdoiu6;  // ../RTL/cortexm0ds_logic.v(629)
  wire Sdphu6;  // ../RTL/cortexm0ds_logic.v(161)
  wire Sdpow6;  // ../RTL/cortexm0ds_logic.v(1186)
  wire Sdviu6;  // ../RTL/cortexm0ds_logic.v(723)
  wire Sdwhu6;  // ../RTL/cortexm0ds_logic.v(255)
  wire Sdwow6;  // ../RTL/cortexm0ds_logic.v(1279)
  wire Se1ju6;  // ../RTL/cortexm0ds_logic.v(804)
  wire Se2iu6;  // ../RTL/cortexm0ds_logic.v(336)
  wire Se2pw6;  // ../RTL/cortexm0ds_logic.v(1360)
  wire Se8ju6;  // ../RTL/cortexm0ds_logic.v(897)
  wire Se9iu6;  // ../RTL/cortexm0ds_logic.v(429)
  wire Se9pw6;  // ../RTL/cortexm0ds_logic.v(1454)
  wire Seaow6;  // ../RTL/cortexm0ds_logic.v(986)
  wire Seehu6;  // ../RTL/cortexm0ds_logic.v(122)
  wire Segiu6;  // ../RTL/cortexm0ds_logic.v(523)
  wire Sehow6;  // ../RTL/cortexm0ds_logic.v(1079)
  wire Sejax6;  // ../RTL/cortexm0ds_logic.v(1649)
  wire Seniu6;  // ../RTL/cortexm0ds_logic.v(616)
  wire Seohu6;  // ../RTL/cortexm0ds_logic.v(148)
  wire Seoow6;  // ../RTL/cortexm0ds_logic.v(1173)
  wire Serax6;  // ../RTL/cortexm0ds_logic.v(1664)
  wire Seuiu6;  // ../RTL/cortexm0ds_logic.v(710)
  wire Sevhu6;  // ../RTL/cortexm0ds_logic.v(242)
  wire Sevow6;  // ../RTL/cortexm0ds_logic.v(1266)
  wire Sf0ju6;  // ../RTL/cortexm0ds_logic.v(791)
  wire Sf1iu6;  // ../RTL/cortexm0ds_logic.v(323)
  wire Sf1pw6;  // ../RTL/cortexm0ds_logic.v(1347)
  wire Sf7ju6;  // ../RTL/cortexm0ds_logic.v(884)
  wire Sf8iu6;  // ../RTL/cortexm0ds_logic.v(416)
  wire Sf8pw6;  // ../RTL/cortexm0ds_logic.v(1441)
  wire Sf9ow6;  // ../RTL/cortexm0ds_logic.v(973)
  wire Sffiu6;  // ../RTL/cortexm0ds_logic.v(510)
  wire Sfmiu6;  // ../RTL/cortexm0ds_logic.v(603)
  wire Sfnow6;  // ../RTL/cortexm0ds_logic.v(1160)
  wire Sftiu6;  // ../RTL/cortexm0ds_logic.v(697)
  wire Sfuhu6;  // ../RTL/cortexm0ds_logic.v(229)
  wire Sfuow6;  // ../RTL/cortexm0ds_logic.v(1253)
  wire Sfypw6;  // ../RTL/cortexm0ds_logic.v(1614)
  wire Sg0iu6;  // ../RTL/cortexm0ds_logic.v(310)
  wire Sg0pw6;  // ../RTL/cortexm0ds_logic.v(1334)
  wire Sg6ju6;  // ../RTL/cortexm0ds_logic.v(871)
  wire Sg7iu6;  // ../RTL/cortexm0ds_logic.v(403)
  wire Sg7pw6;  // ../RTL/cortexm0ds_logic.v(1428)
  wire Sg8ow6;  // ../RTL/cortexm0ds_logic.v(960)
  wire Sgeiu6;  // ../RTL/cortexm0ds_logic.v(497)
  wire Sgfow6;  // ../RTL/cortexm0ds_logic.v(1053)
  wire Sgjax6;  // ../RTL/cortexm0ds_logic.v(1649)
  wire Sgliu6;  // ../RTL/cortexm0ds_logic.v(590)
  wire Sgmow6;  // ../RTL/cortexm0ds_logic.v(1147)
  wire Sgsiu6;  // ../RTL/cortexm0ds_logic.v(684)
  wire Sgthu6;  // ../RTL/cortexm0ds_logic.v(216)
  wire Sgtow6;  // ../RTL/cortexm0ds_logic.v(1240)
  wire Sgziu6;  // ../RTL/cortexm0ds_logic.v(778)
  wire Sh4bx6;  // ../RTL/cortexm0ds_logic.v(1687)
  wire Sh5ju6;  // ../RTL/cortexm0ds_logic.v(858)
  wire Sh6iu6;  // ../RTL/cortexm0ds_logic.v(390)
  wire Sh6pw6;  // ../RTL/cortexm0ds_logic.v(1415)
  wire Sh7ow6;  // ../RTL/cortexm0ds_logic.v(947)
  wire Shdiu6;  // ../RTL/cortexm0ds_logic.v(484)
  wire Shdpw6;  // ../RTL/cortexm0ds_logic.v(1508)
  wire Sheow6;  // ../RTL/cortexm0ds_logic.v(1040)
  wire Shkiu6;  // ../RTL/cortexm0ds_logic.v(577)
  wire Shlow6;  // ../RTL/cortexm0ds_logic.v(1134)
  wire Shopw6;  // ../RTL/cortexm0ds_logic.v(1596)
  wire Shriu6;  // ../RTL/cortexm0ds_logic.v(671)
  wire Shshu6;  // ../RTL/cortexm0ds_logic.v(203)
  wire Shsow6;  // ../RTL/cortexm0ds_logic.v(1227)
  wire Shyiu6;  // ../RTL/cortexm0ds_logic.v(765)
  wire Shzhu6;  // ../RTL/cortexm0ds_logic.v(297)
  wire Shzow6;  // ../RTL/cortexm0ds_logic.v(1321)
  wire Si4ju6;  // ../RTL/cortexm0ds_logic.v(845)
  wire Si5iu6;  // ../RTL/cortexm0ds_logic.v(377)
  wire Si5pw6;  // ../RTL/cortexm0ds_logic.v(1402)
  wire Si6ow6;  // ../RTL/cortexm0ds_logic.v(934)
  wire Siciu6;  // ../RTL/cortexm0ds_logic.v(471)
  wire Sicpw6;  // ../RTL/cortexm0ds_logic.v(1495)
  wire Sidow6;  // ../RTL/cortexm0ds_logic.v(1027)
  wire Sijax6;  // ../RTL/cortexm0ds_logic.v(1650)
  wire Sijiu6;  // ../RTL/cortexm0ds_logic.v(564)
  wire Sikow6;  // ../RTL/cortexm0ds_logic.v(1121)
  wire Siqiu6;  // ../RTL/cortexm0ds_logic.v(658)
  wire Sirhu6;  // ../RTL/cortexm0ds_logic.v(190)
  wire Sirow6;  // ../RTL/cortexm0ds_logic.v(1214)
  wire Sixiu6;  // ../RTL/cortexm0ds_logic.v(752)
  wire Siyhu6;  // ../RTL/cortexm0ds_logic.v(284)
  wire Siyow6;  // ../RTL/cortexm0ds_logic.v(1308)
  wire Sj3ju6;  // ../RTL/cortexm0ds_logic.v(832)
  wire Sj4iu6;  // ../RTL/cortexm0ds_logic.v(364)
  wire Sj4pw6;  // ../RTL/cortexm0ds_logic.v(1389)
  wire Sjaju6;  // ../RTL/cortexm0ds_logic.v(926)
  wire Sjbiu6;  // ../RTL/cortexm0ds_logic.v(458)
  wire Sjbpw6;  // ../RTL/cortexm0ds_logic.v(1482)
  wire Sjcow6;  // ../RTL/cortexm0ds_logic.v(1014)
  wire Sjiiu6;  // ../RTL/cortexm0ds_logic.v(551)
  wire Sjjow6;  // ../RTL/cortexm0ds_logic.v(1108)
  wire Sjkhu6;  // ../RTL/cortexm0ds_logic.v(137)
  wire Sjpiu6;  // ../RTL/cortexm0ds_logic.v(645)
  wire Sjqhu6;  // ../RTL/cortexm0ds_logic.v(177)
  wire Sjqow6;  // ../RTL/cortexm0ds_logic.v(1201)
  wire Sjwiu6;  // ../RTL/cortexm0ds_logic.v(739)
  wire Sjxhu6;  // ../RTL/cortexm0ds_logic.v(271)
  wire Sjxow6;  // ../RTL/cortexm0ds_logic.v(1295)
  wire Sk2ju6;  // ../RTL/cortexm0ds_logic.v(819)
  wire Sk3iu6;  // ../RTL/cortexm0ds_logic.v(351)
  wire Sk3pw6;  // ../RTL/cortexm0ds_logic.v(1376)
  wire Sk9ju6;  // ../RTL/cortexm0ds_logic.v(913)
  wire Skaiu6;  // ../RTL/cortexm0ds_logic.v(445)
  wire Skapw6;  // ../RTL/cortexm0ds_logic.v(1469)
  wire Skbow6;  // ../RTL/cortexm0ds_logic.v(1001)
  wire Skhiu6;  // ../RTL/cortexm0ds_logic.v(538)
  wire Skiow6;  // ../RTL/cortexm0ds_logic.v(1095)
  wire Skjax6;  // ../RTL/cortexm0ds_logic.v(1650)
  wire Skoiu6;  // ../RTL/cortexm0ds_logic.v(632)
  wire Skphu6;  // ../RTL/cortexm0ds_logic.v(164)
  wire Skpow6;  // ../RTL/cortexm0ds_logic.v(1188)
  wire Skviu6;  // ../RTL/cortexm0ds_logic.v(726)
  wire Skwhu6;  // ../RTL/cortexm0ds_logic.v(258)
  wire Skwow6;  // ../RTL/cortexm0ds_logic.v(1282)
  wire Sl1ju6;  // ../RTL/cortexm0ds_logic.v(806)
  wire Sl2iu6;  // ../RTL/cortexm0ds_logic.v(338)
  wire Sl2pw6;  // ../RTL/cortexm0ds_logic.v(1363)
  wire Sl8ju6;  // ../RTL/cortexm0ds_logic.v(900)
  wire Sl9iu6;  // ../RTL/cortexm0ds_logic.v(432)
  wire Sl9pw6;  // ../RTL/cortexm0ds_logic.v(1456)
  wire Slaow6;  // ../RTL/cortexm0ds_logic.v(988)
  wire Slgiu6;  // ../RTL/cortexm0ds_logic.v(525)
  wire Slhow6;  // ../RTL/cortexm0ds_logic.v(1082)
  wire Sljhu6;  // ../RTL/cortexm0ds_logic.v(134)
  wire Slniu6;  // ../RTL/cortexm0ds_logic.v(619)
  wire Slohu6;  // ../RTL/cortexm0ds_logic.v(151)
  wire Sloow6;  // ../RTL/cortexm0ds_logic.v(1175)
  wire Sluiu6;  // ../RTL/cortexm0ds_logic.v(713)
  wire Slvax6;  // ../RTL/cortexm0ds_logic.v(1671)
  wire Slvhu6;  // ../RTL/cortexm0ds_logic.v(245)
  wire Slvow6;  // ../RTL/cortexm0ds_logic.v(1269)
  wire Slyax6;  // ../RTL/cortexm0ds_logic.v(1677)
  wire Sm0ju6;  // ../RTL/cortexm0ds_logic.v(793)
  wire Sm1iu6;  // ../RTL/cortexm0ds_logic.v(325)
  wire Sm1pw6;  // ../RTL/cortexm0ds_logic.v(1350)
  wire Sm7ju6;  // ../RTL/cortexm0ds_logic.v(887)
  wire Sm8iu6;  // ../RTL/cortexm0ds_logic.v(419)
  wire Sm8pw6;  // ../RTL/cortexm0ds_logic.v(1443)
  wire Sm9ow6;  // ../RTL/cortexm0ds_logic.v(975)
  wire Smfiu6;  // ../RTL/cortexm0ds_logic.v(512)
  wire Smgow6;  // ../RTL/cortexm0ds_logic.v(1069)
  wire Smhhu6;  // ../RTL/cortexm0ds_logic.v(129)
  wire Smjax6;  // ../RTL/cortexm0ds_logic.v(1650)
  wire Smmiu6;  // ../RTL/cortexm0ds_logic.v(606)
  wire Smnow6;  // ../RTL/cortexm0ds_logic.v(1162)
  wire Smtiu6;  // ../RTL/cortexm0ds_logic.v(700)
  wire Smuhu6;  // ../RTL/cortexm0ds_logic.v(232)
  wire Smuow6;  // ../RTL/cortexm0ds_logic.v(1256)
  wire Sn0iu6;  // ../RTL/cortexm0ds_logic.v(312)
  wire Sn0pw6;  // ../RTL/cortexm0ds_logic.v(1337)
  wire Sn4bx6;  // ../RTL/cortexm0ds_logic.v(1687)
  wire Sn6ju6;  // ../RTL/cortexm0ds_logic.v(874)
  wire Sn7iu6;  // ../RTL/cortexm0ds_logic.v(406)
  wire Sn7pw6;  // ../RTL/cortexm0ds_logic.v(1430)
  wire Sn8ow6;  // ../RTL/cortexm0ds_logic.v(962)
  wire Sneiu6;  // ../RTL/cortexm0ds_logic.v(499)
  wire Snfow6;  // ../RTL/cortexm0ds_logic.v(1056)
  wire Snihu6;  // ../RTL/cortexm0ds_logic.v(131)
  wire Snliu6;  // ../RTL/cortexm0ds_logic.v(593)
  wire Snmow6;  // ../RTL/cortexm0ds_logic.v(1149)
  wire Snsiu6;  // ../RTL/cortexm0ds_logic.v(687)
  wire Snthu6;  // ../RTL/cortexm0ds_logic.v(219)
  wire Sntow6;  // ../RTL/cortexm0ds_logic.v(1243)
  wire Snziu6;  // ../RTL/cortexm0ds_logic.v(780)
  wire So0qw6;  // ../RTL/cortexm0ds_logic.v(1618)
  wire So5ju6;  // ../RTL/cortexm0ds_logic.v(861)
  wire So6iu6;  // ../RTL/cortexm0ds_logic.v(393)
  wire So6pw6;  // ../RTL/cortexm0ds_logic.v(1417)
  wire So7ow6;  // ../RTL/cortexm0ds_logic.v(949)
  wire Sodiu6;  // ../RTL/cortexm0ds_logic.v(486)
  wire Sodpw6;  // ../RTL/cortexm0ds_logic.v(1511)
  wire Soeow6;  // ../RTL/cortexm0ds_logic.v(1043)
  wire Sojax6;  // ../RTL/cortexm0ds_logic.v(1650)
  wire Sokiu6;  // ../RTL/cortexm0ds_logic.v(580)
  wire Solow6;  // ../RTL/cortexm0ds_logic.v(1136)
  wire Soriu6;  // ../RTL/cortexm0ds_logic.v(674)
  wire Soshu6;  // ../RTL/cortexm0ds_logic.v(206)
  wire Sosow6;  // ../RTL/cortexm0ds_logic.v(1230)
  wire Soyiu6;  // ../RTL/cortexm0ds_logic.v(767)
  wire Sozhu6;  // ../RTL/cortexm0ds_logic.v(299)
  wire Sozow6;  // ../RTL/cortexm0ds_logic.v(1324)
  wire Sp4ju6;  // ../RTL/cortexm0ds_logic.v(848)
  wire Sp5iu6;  // ../RTL/cortexm0ds_logic.v(380)
  wire Sp5pw6;  // ../RTL/cortexm0ds_logic.v(1404)
  wire Sp6ow6;  // ../RTL/cortexm0ds_logic.v(936)
  wire Spciu6;  // ../RTL/cortexm0ds_logic.v(473)
  wire Spcpw6;  // ../RTL/cortexm0ds_logic.v(1498)
  wire Spdow6;  // ../RTL/cortexm0ds_logic.v(1030)
  wire Spjiu6;  // ../RTL/cortexm0ds_logic.v(567)
  wire Spkow6;  // ../RTL/cortexm0ds_logic.v(1123)
  wire Spqiu6;  // ../RTL/cortexm0ds_logic.v(661)
  wire Sprhu6;  // ../RTL/cortexm0ds_logic.v(193)
  wire Sprow6;  // ../RTL/cortexm0ds_logic.v(1217)
  wire Spxiu6;  // ../RTL/cortexm0ds_logic.v(754)
  wire Spyhu6;  // ../RTL/cortexm0ds_logic.v(286)
  wire Spyow6;  // ../RTL/cortexm0ds_logic.v(1311)
  wire Sq3bx6;  // ../RTL/cortexm0ds_logic.v(1686)
  wire Sq3ju6;  // ../RTL/cortexm0ds_logic.v(835)
  wire Sq4iu6;  // ../RTL/cortexm0ds_logic.v(367)
  wire Sq4pw6;  // ../RTL/cortexm0ds_logic.v(1391)
  wire Sqaju6;  // ../RTL/cortexm0ds_logic.v(928)
  wire Sqbiu6;  // ../RTL/cortexm0ds_logic.v(460)
  wire Sqbpw6;  // ../RTL/cortexm0ds_logic.v(1485)
  wire Sqcow6;  // ../RTL/cortexm0ds_logic.v(1017)
  wire Sqfax6;  // ../RTL/cortexm0ds_logic.v(1642)
  wire Sqiiu6;  // ../RTL/cortexm0ds_logic.v(554)
  wire Sqjax6;  // ../RTL/cortexm0ds_logic.v(1650)
  wire Sqjow6;  // ../RTL/cortexm0ds_logic.v(1110)
  wire Sqkax6;  // ../RTL/cortexm0ds_logic.v(1652)
  wire Sqpiu6;  // ../RTL/cortexm0ds_logic.v(648)
  wire Sqqhu6;  // ../RTL/cortexm0ds_logic.v(180)
  wire Sqqow6;  // ../RTL/cortexm0ds_logic.v(1204)
  wire Sqwiu6;  // ../RTL/cortexm0ds_logic.v(741)
  wire Sqwpw6;  // ../RTL/cortexm0ds_logic.v(1611)
  wire Sqxhu6;  // ../RTL/cortexm0ds_logic.v(273)
  wire Sqxow6;  // ../RTL/cortexm0ds_logic.v(1298)
  wire Sr2ju6;  // ../RTL/cortexm0ds_logic.v(822)
  wire Sr3iu6;  // ../RTL/cortexm0ds_logic.v(354)
  wire Sr3pw6;  // ../RTL/cortexm0ds_logic.v(1378)
  wire Sr9ju6;  // ../RTL/cortexm0ds_logic.v(915)
  wire Sraiu6;  // ../RTL/cortexm0ds_logic.v(447)
  wire Srapw6;  // ../RTL/cortexm0ds_logic.v(1472)
  wire Srbow6;  // ../RTL/cortexm0ds_logic.v(1004)
  wire Srhiu6;  // ../RTL/cortexm0ds_logic.v(541)
  wire Sriow6;  // ../RTL/cortexm0ds_logic.v(1097)
  wire Sroiu6;  // ../RTL/cortexm0ds_logic.v(635)
  wire Srphu6;  // ../RTL/cortexm0ds_logic.v(167)
  wire Srpow6;  // ../RTL/cortexm0ds_logic.v(1191)
  wire Srviu6;  // ../RTL/cortexm0ds_logic.v(728)
  wire Srwhu6;  // ../RTL/cortexm0ds_logic.v(260)
  wire Srwow6;  // ../RTL/cortexm0ds_logic.v(1285)
  wire Ss0qw6;  // ../RTL/cortexm0ds_logic.v(1618)
  wire Ss1ju6;  // ../RTL/cortexm0ds_logic.v(809)
  wire Ss2iu6;  // ../RTL/cortexm0ds_logic.v(341)
  wire Ss2pw6;  // ../RTL/cortexm0ds_logic.v(1365)
  wire Ss8ju6;  // ../RTL/cortexm0ds_logic.v(902)
  wire Ss9iu6;  // ../RTL/cortexm0ds_logic.v(434)
  wire Ss9pw6;  // ../RTL/cortexm0ds_logic.v(1459)
  wire Ssaow6;  // ../RTL/cortexm0ds_logic.v(991)
  wire Ssgiu6;  // ../RTL/cortexm0ds_logic.v(528)
  wire Sshow6;  // ../RTL/cortexm0ds_logic.v(1084)
  wire Ssjax6;  // ../RTL/cortexm0ds_logic.v(1650)
  wire Ssniu6;  // ../RTL/cortexm0ds_logic.v(622)
  wire Ssohu6;  // ../RTL/cortexm0ds_logic.v(154)
  wire Ssoow6;  // ../RTL/cortexm0ds_logic.v(1178)
  wire Ssuiu6;  // ../RTL/cortexm0ds_logic.v(715)
  wire Ssvhu6;  // ../RTL/cortexm0ds_logic.v(247)
  wire Ssvow6;  // ../RTL/cortexm0ds_logic.v(1272)
  wire St0ju6;  // ../RTL/cortexm0ds_logic.v(796)
  wire St1iu6;  // ../RTL/cortexm0ds_logic.v(328)
  wire St1pw6;  // ../RTL/cortexm0ds_logic.v(1352)
  wire St7ju6;  // ../RTL/cortexm0ds_logic.v(889)
  wire St8iu6;  // ../RTL/cortexm0ds_logic.v(421)
  wire St8pw6;  // ../RTL/cortexm0ds_logic.v(1446)
  wire St9ow6;  // ../RTL/cortexm0ds_logic.v(978)
  wire Stdhu6;  // ../RTL/cortexm0ds_logic.v(120)
  wire Stfiu6;  // ../RTL/cortexm0ds_logic.v(515)
  wire Stgow6;  // ../RTL/cortexm0ds_logic.v(1071)
  wire Stkpw6;  // ../RTL/cortexm0ds_logic.v(1589)
  wire Stmiu6;  // ../RTL/cortexm0ds_logic.v(609)
  wire Stnow6;  // ../RTL/cortexm0ds_logic.v(1165)
  wire Sttiu6;  // ../RTL/cortexm0ds_logic.v(702)
  wire Stuhu6;  // ../RTL/cortexm0ds_logic.v(234)
  wire Stuow6;  // ../RTL/cortexm0ds_logic.v(1259)
  wire Su0iu6;  // ../RTL/cortexm0ds_logic.v(315)
  wire Su0pw6;  // ../RTL/cortexm0ds_logic.v(1339)
  wire Su6ju6;  // ../RTL/cortexm0ds_logic.v(876)
  wire Su7iu6;  // ../RTL/cortexm0ds_logic.v(408)
  wire Su7pw6;  // ../RTL/cortexm0ds_logic.v(1433)
  wire Su8ax6;  // ../RTL/cortexm0ds_logic.v(1629)
  wire Su8ow6;  // ../RTL/cortexm0ds_logic.v(965)
  wire Sueiu6;  // ../RTL/cortexm0ds_logic.v(502)
  wire Sufow6;  // ../RTL/cortexm0ds_logic.v(1058)
  wire Sujax6;  // ../RTL/cortexm0ds_logic.v(1650)
  wire Suliu6;  // ../RTL/cortexm0ds_logic.v(596)
  wire Sumow6;  // ../RTL/cortexm0ds_logic.v(1152)
  wire Susiu6;  // ../RTL/cortexm0ds_logic.v(689)
  wire Suthu6;  // ../RTL/cortexm0ds_logic.v(221)
  wire Sutow6;  // ../RTL/cortexm0ds_logic.v(1246)
  wire Suziu6;  // ../RTL/cortexm0ds_logic.v(783)
  wire Sv5ju6;  // ../RTL/cortexm0ds_logic.v(863)
  wire Sv6iu6;  // ../RTL/cortexm0ds_logic.v(395)
  wire Sv6pw6;  // ../RTL/cortexm0ds_logic.v(1420)
  wire Sv7ow6;  // ../RTL/cortexm0ds_logic.v(952)
  wire Svdiu6;  // ../RTL/cortexm0ds_logic.v(489)
  wire Svdpw6;  // ../RTL/cortexm0ds_logic.v(1513)
  wire Sveow6;  // ../RTL/cortexm0ds_logic.v(1045)
  wire Svkiu6;  // ../RTL/cortexm0ds_logic.v(583)
  wire Svlow6;  // ../RTL/cortexm0ds_logic.v(1139)
  wire Svriu6;  // ../RTL/cortexm0ds_logic.v(676)
  wire Svshu6;  // ../RTL/cortexm0ds_logic.v(208)
  wire Svsow6;  // ../RTL/cortexm0ds_logic.v(1233)
  wire Svyiu6;  // ../RTL/cortexm0ds_logic.v(770)
  wire Svzhu6;  // ../RTL/cortexm0ds_logic.v(302)
  wire Svzow6;  // ../RTL/cortexm0ds_logic.v(1326)
  wire Sw0qw6;  // ../RTL/cortexm0ds_logic.v(1619)
  wire Sw4ju6;  // ../RTL/cortexm0ds_logic.v(850)
  wire Sw5iu6;  // ../RTL/cortexm0ds_logic.v(382)
  wire Sw5pw6;  // ../RTL/cortexm0ds_logic.v(1407)
  wire Sw6ow6;  // ../RTL/cortexm0ds_logic.v(939)
  wire Swciu6;  // ../RTL/cortexm0ds_logic.v(476)
  wire Swcpw6;  // ../RTL/cortexm0ds_logic.v(1500)
  wire Swdow6;  // ../RTL/cortexm0ds_logic.v(1032)
  wire Swjbx6;  // ../RTL/cortexm0ds_logic.v(1715)
  wire Swjiu6;  // ../RTL/cortexm0ds_logic.v(570)
  wire Swkow6;  // ../RTL/cortexm0ds_logic.v(1126)
  wire Swqiu6;  // ../RTL/cortexm0ds_logic.v(663)
  wire Swrhu6;  // ../RTL/cortexm0ds_logic.v(195)
  wire Swrow6;  // ../RTL/cortexm0ds_logic.v(1220)
  wire Swxiu6;  // ../RTL/cortexm0ds_logic.v(757)
  wire Swyhu6;  // ../RTL/cortexm0ds_logic.v(289)
  wire Swyow6;  // ../RTL/cortexm0ds_logic.v(1313)
  wire Sx3ju6;  // ../RTL/cortexm0ds_logic.v(837)
  wire Sx3qw6;  // ../RTL/cortexm0ds_logic.v(1624)
  wire Sx4iu6;  // ../RTL/cortexm0ds_logic.v(369)
  wire Sx4pw6;  // ../RTL/cortexm0ds_logic.v(1394)
  wire Sx7ax6;  // ../RTL/cortexm0ds_logic.v(1627)
  wire Sxbiu6;  // ../RTL/cortexm0ds_logic.v(463)
  wire Sxbpw6;  // ../RTL/cortexm0ds_logic.v(1487)
  wire Sxcow6;  // ../RTL/cortexm0ds_logic.v(1019)
  wire Sxiiu6;  // ../RTL/cortexm0ds_logic.v(557)
  wire Sxjow6;  // ../RTL/cortexm0ds_logic.v(1113)
  wire Sxpiu6;  // ../RTL/cortexm0ds_logic.v(650)
  wire Sxqhu6;  // ../RTL/cortexm0ds_logic.v(182)
  wire Sxqow6;  // ../RTL/cortexm0ds_logic.v(1207)
  wire Sxwiu6;  // ../RTL/cortexm0ds_logic.v(744)
  wire Sxxhu6;  // ../RTL/cortexm0ds_logic.v(276)
  wire Sxxow6;  // ../RTL/cortexm0ds_logic.v(1300)
  wire Sy2ju6;  // ../RTL/cortexm0ds_logic.v(824)
  wire Sy3iu6;  // ../RTL/cortexm0ds_logic.v(356)
  wire Sy3pw6;  // ../RTL/cortexm0ds_logic.v(1381)
  wire Sy9ju6;  // ../RTL/cortexm0ds_logic.v(918)
  wire Syaiu6;  // ../RTL/cortexm0ds_logic.v(450)
  wire Syapw6;  // ../RTL/cortexm0ds_logic.v(1474)
  wire Sybow6;  // ../RTL/cortexm0ds_logic.v(1006)
  wire Syehu6;  // ../RTL/cortexm0ds_logic.v(123)
  wire Syhiu6;  // ../RTL/cortexm0ds_logic.v(544)
  wire Syiow6;  // ../RTL/cortexm0ds_logic.v(1100)
  wire Syjbx6;  // ../RTL/cortexm0ds_logic.v(1715)
  wire Syoiu6;  // ../RTL/cortexm0ds_logic.v(637)
  wire Syphu6;  // ../RTL/cortexm0ds_logic.v(169)
  wire Sypow6;  // ../RTL/cortexm0ds_logic.v(1194)
  wire Syviu6;  // ../RTL/cortexm0ds_logic.v(731)
  wire Sywhu6;  // ../RTL/cortexm0ds_logic.v(263)
  wire Sywow6;  // ../RTL/cortexm0ds_logic.v(1287)
  wire Sz1ju6;  // ../RTL/cortexm0ds_logic.v(811)
  wire Sz2iu6;  // ../RTL/cortexm0ds_logic.v(343)
  wire Sz2pw6;  // ../RTL/cortexm0ds_logic.v(1368)
  wire Sz3qw6;  // ../RTL/cortexm0ds_logic.v(1625)
  wire Sz7ax6;  // ../RTL/cortexm0ds_logic.v(1627)
  wire Sz8ju6;  // ../RTL/cortexm0ds_logic.v(905)
  wire Sz9iu6;  // ../RTL/cortexm0ds_logic.v(437)
  wire Sz9pw6;  // ../RTL/cortexm0ds_logic.v(1461)
  wire Szaow6;  // ../RTL/cortexm0ds_logic.v(993)
  wire Szgiu6;  // ../RTL/cortexm0ds_logic.v(531)
  wire Szhow6;  // ../RTL/cortexm0ds_logic.v(1087)
  wire Szmax6;  // ../RTL/cortexm0ds_logic.v(1656)
  wire Szniu6;  // ../RTL/cortexm0ds_logic.v(624)
  wire Szohu6;  // ../RTL/cortexm0ds_logic.v(156)
  wire Szoow6;  // ../RTL/cortexm0ds_logic.v(1181)
  wire Szuiu6;  // ../RTL/cortexm0ds_logic.v(718)
  wire Szvhu6;  // ../RTL/cortexm0ds_logic.v(250)
  wire Szvow6;  // ../RTL/cortexm0ds_logic.v(1274)
  wire T00qw6;  // ../RTL/cortexm0ds_logic.v(1617)
  wire T05ju6;  // ../RTL/cortexm0ds_logic.v(852)
  wire T06iu6;  // ../RTL/cortexm0ds_logic.v(384)
  wire T06pw6;  // ../RTL/cortexm0ds_logic.v(1408)
  wire T07ow6;  // ../RTL/cortexm0ds_logic.v(940)
  wire T0diu6;  // ../RTL/cortexm0ds_logic.v(477)
  wire T0dpw6;  // ../RTL/cortexm0ds_logic.v(1502)
  wire T0eow6;  // ../RTL/cortexm0ds_logic.v(1034)
  wire T0hhu6;  // ../RTL/cortexm0ds_logic.v(127)
  wire T0ipw6;  // ../RTL/cortexm0ds_logic.v(1584)
  wire T0kiu6;  // ../RTL/cortexm0ds_logic.v(571)
  wire T0low6;  // ../RTL/cortexm0ds_logic.v(1127)
  wire T0riu6;  // ../RTL/cortexm0ds_logic.v(665)
  wire T0shu6;  // ../RTL/cortexm0ds_logic.v(197)
  wire T0sow6;  // ../RTL/cortexm0ds_logic.v(1221)
  wire T0yiu6;  // ../RTL/cortexm0ds_logic.v(758)
  wire T0zhu6;  // ../RTL/cortexm0ds_logic.v(290)
  wire T0zow6;  // ../RTL/cortexm0ds_logic.v(1315)
  wire T14ju6;  // ../RTL/cortexm0ds_logic.v(839)
  wire T15iu6;  // ../RTL/cortexm0ds_logic.v(371)
  wire T15pw6;  // ../RTL/cortexm0ds_logic.v(1395)
  wire T1ciu6;  // ../RTL/cortexm0ds_logic.v(464)
  wire T1cpw6;  // ../RTL/cortexm0ds_logic.v(1489)
  wire T1dow6;  // ../RTL/cortexm0ds_logic.v(1021)
  wire T1fbx6;  // ../RTL/cortexm0ds_logic.v(1706)
  wire T1jiu6;  // ../RTL/cortexm0ds_logic.v(558)
  wire T1kow6;  // ../RTL/cortexm0ds_logic.v(1114)
  wire T1qiu6;  // ../RTL/cortexm0ds_logic.v(652)
  wire T1rhu6;  // ../RTL/cortexm0ds_logic.v(184)
  wire T1row6;  // ../RTL/cortexm0ds_logic.v(1208)
  wire T1vpw6;  // ../RTL/cortexm0ds_logic.v(1608)
  wire T1xiu6;  // ../RTL/cortexm0ds_logic.v(745)
  wire T1yhu6;  // ../RTL/cortexm0ds_logic.v(277)
  wire T1yow6;  // ../RTL/cortexm0ds_logic.v(1302)
  wire T20qw6;  // ../RTL/cortexm0ds_logic.v(1617)
  wire T23ju6;  // ../RTL/cortexm0ds_logic.v(826)
  wire T24iu6;  // ../RTL/cortexm0ds_logic.v(358)
  wire T24pw6;  // ../RTL/cortexm0ds_logic.v(1382)
  wire T2aju6;  // ../RTL/cortexm0ds_logic.v(919)
  wire T2biu6;  // ../RTL/cortexm0ds_logic.v(451)
  wire T2bpw6;  // ../RTL/cortexm0ds_logic.v(1476)
  wire T2cow6;  // ../RTL/cortexm0ds_logic.v(1008)
  wire T2dbx6;  // ../RTL/cortexm0ds_logic.v(1703)
  wire T2iiu6;  // ../RTL/cortexm0ds_logic.v(545)
  wire T2jow6;  // ../RTL/cortexm0ds_logic.v(1101)
  wire T2kbx6;  // ../RTL/cortexm0ds_logic.v(1716)
  wire T2piu6;  // ../RTL/cortexm0ds_logic.v(639)
  wire T2qhu6;  // ../RTL/cortexm0ds_logic.v(171)
  wire T2qow6;  // ../RTL/cortexm0ds_logic.v(1195)
  wire T2wiu6;  // ../RTL/cortexm0ds_logic.v(732)
  wire T2xhu6;  // ../RTL/cortexm0ds_logic.v(264)
  wire T2xow6;  // ../RTL/cortexm0ds_logic.v(1289)
  wire T32ju6;  // ../RTL/cortexm0ds_logic.v(813)
  wire T33iu6;  // ../RTL/cortexm0ds_logic.v(345)
  wire T33pw6;  // ../RTL/cortexm0ds_logic.v(1369)
  wire T39ju6;  // ../RTL/cortexm0ds_logic.v(906)
  wire T3abx6;  // ../RTL/cortexm0ds_logic.v(1697)
  wire T3aiu6;  // ../RTL/cortexm0ds_logic.v(438)
  wire T3apw6;  // ../RTL/cortexm0ds_logic.v(1463)
  wire T3bow6;  // ../RTL/cortexm0ds_logic.v(995)
  wire T3fbx6;  // ../RTL/cortexm0ds_logic.v(1707)
  wire T3hiu6;  // ../RTL/cortexm0ds_logic.v(532)
  wire T3iow6;  // ../RTL/cortexm0ds_logic.v(1088)
  wire T3kpw6;  // ../RTL/cortexm0ds_logic.v(1588)
  wire T3oiu6;  // ../RTL/cortexm0ds_logic.v(626)
  wire T3opw6;  // ../RTL/cortexm0ds_logic.v(1595)
  wire T3phu6;  // ../RTL/cortexm0ds_logic.v(158)
  wire T3pow6;  // ../RTL/cortexm0ds_logic.v(1182)
  wire T3viu6;  // ../RTL/cortexm0ds_logic.v(719)
  wire T3whu6;  // ../RTL/cortexm0ds_logic.v(251)
  wire T3wow6;  // ../RTL/cortexm0ds_logic.v(1276)
  wire T40qw6;  // ../RTL/cortexm0ds_logic.v(1617)
  wire T41ju6;  // ../RTL/cortexm0ds_logic.v(800)
  wire T42iu6;  // ../RTL/cortexm0ds_logic.v(332)
  wire T42pw6;  // ../RTL/cortexm0ds_logic.v(1356)
  wire T48ju6;  // ../RTL/cortexm0ds_logic.v(893)
  wire T49iu6;  // ../RTL/cortexm0ds_logic.v(425)
  wire T49pw6;  // ../RTL/cortexm0ds_logic.v(1450)
  wire T4aow6;  // ../RTL/cortexm0ds_logic.v(982)
  wire T4giu6;  // ../RTL/cortexm0ds_logic.v(519)
  wire T4how6;  // ../RTL/cortexm0ds_logic.v(1075)
  wire T4niu6;  // ../RTL/cortexm0ds_logic.v(613)
  wire T4oow6;  // ../RTL/cortexm0ds_logic.v(1169)
  wire T4uiu6;  // ../RTL/cortexm0ds_logic.v(706)
  wire T4vhu6;  // ../RTL/cortexm0ds_logic.v(238)
  wire T4vow6;  // ../RTL/cortexm0ds_logic.v(1263)
  wire T50ju6;  // ../RTL/cortexm0ds_logic.v(787)
  wire T51iu6;  // ../RTL/cortexm0ds_logic.v(319)
  wire T51pw6;  // ../RTL/cortexm0ds_logic.v(1343)
  wire T57ju6;  // ../RTL/cortexm0ds_logic.v(880)
  wire T58iu6;  // ../RTL/cortexm0ds_logic.v(412)
  wire T58pw6;  // ../RTL/cortexm0ds_logic.v(1437)
  wire T59ow6;  // ../RTL/cortexm0ds_logic.v(969)
  wire T5fbx6;  // ../RTL/cortexm0ds_logic.v(1707)
  wire T5fiu6;  // ../RTL/cortexm0ds_logic.v(506)
  wire T5gow6;  // ../RTL/cortexm0ds_logic.v(1062)
  wire T5miu6;  // ../RTL/cortexm0ds_logic.v(600)
  wire T5mpw6;  // ../RTL/cortexm0ds_logic.v(1592)
  wire T5now6;  // ../RTL/cortexm0ds_logic.v(1156)
  wire T5tiu6;  // ../RTL/cortexm0ds_logic.v(693)
  wire T5uhu6;  // ../RTL/cortexm0ds_logic.v(225)
  wire T5uow6;  // ../RTL/cortexm0ds_logic.v(1250)
  wire T5yax6;  // ../RTL/cortexm0ds_logic.v(1676)
  wire T60iu6;  // ../RTL/cortexm0ds_logic.v(306)
  wire T60pw6;  // ../RTL/cortexm0ds_logic.v(1330)
  wire T60qw6;  // ../RTL/cortexm0ds_logic.v(1617)
  wire T66ju6;  // ../RTL/cortexm0ds_logic.v(867)
  wire T67iu6;  // ../RTL/cortexm0ds_logic.v(399)
  wire T67pw6;  // ../RTL/cortexm0ds_logic.v(1424)
  wire T68ow6;  // ../RTL/cortexm0ds_logic.v(956)
  wire T6aax6;  // ../RTL/cortexm0ds_logic.v(1632)
  wire T6ehu6;  // ../RTL/cortexm0ds_logic.v(121)
  wire T6eiu6;  // ../RTL/cortexm0ds_logic.v(493)
  wire T6fow6;  // ../RTL/cortexm0ds_logic.v(1049)
  wire T6kbx6;  // ../RTL/cortexm0ds_logic.v(1716)
  wire T6liu6;  // ../RTL/cortexm0ds_logic.v(587)
  wire T6mow6;  // ../RTL/cortexm0ds_logic.v(1143)
  wire T6siu6;  // ../RTL/cortexm0ds_logic.v(680)
  wire T6thu6;  // ../RTL/cortexm0ds_logic.v(212)
  wire T6tow6;  // ../RTL/cortexm0ds_logic.v(1237)
  wire T6ziu6;  // ../RTL/cortexm0ds_logic.v(774)
  wire T75ju6;  // ../RTL/cortexm0ds_logic.v(854)
  wire T76iu6;  // ../RTL/cortexm0ds_logic.v(386)
  wire T76pw6;  // ../RTL/cortexm0ds_logic.v(1411)
  wire T77ow6;  // ../RTL/cortexm0ds_logic.v(943)
  wire T7bax6;  // ../RTL/cortexm0ds_logic.v(1634)
  wire T7diu6;  // ../RTL/cortexm0ds_logic.v(480)
  wire T7dpw6;  // ../RTL/cortexm0ds_logic.v(1504)
  wire T7eow6;  // ../RTL/cortexm0ds_logic.v(1036)
  wire T7fbx6;  // ../RTL/cortexm0ds_logic.v(1707)
  wire T7kiu6;  // ../RTL/cortexm0ds_logic.v(574)
  wire T7low6;  // ../RTL/cortexm0ds_logic.v(1130)
  wire T7riu6;  // ../RTL/cortexm0ds_logic.v(667)
  wire T7shu6;  // ../RTL/cortexm0ds_logic.v(199)
  wire T7sow6;  // ../RTL/cortexm0ds_logic.v(1224)
  wire T7yiu6;  // ../RTL/cortexm0ds_logic.v(761)
  wire T7zhu6;  // ../RTL/cortexm0ds_logic.v(293)
  wire T7zow6;  // ../RTL/cortexm0ds_logic.v(1317)
  wire T80qw6;  // ../RTL/cortexm0ds_logic.v(1617)
  wire T82qw6;  // ../RTL/cortexm0ds_logic.v(1621)
  wire T84ju6;  // ../RTL/cortexm0ds_logic.v(841)
  wire T85iu6;  // ../RTL/cortexm0ds_logic.v(373)
  wire T85pw6;  // ../RTL/cortexm0ds_logic.v(1398)
  wire T86ow6;  // ../RTL/cortexm0ds_logic.v(930)
  wire T8ciu6;  // ../RTL/cortexm0ds_logic.v(467)
  wire T8cpw6;  // ../RTL/cortexm0ds_logic.v(1491)
  wire T8dow6;  // ../RTL/cortexm0ds_logic.v(1023)
  wire T8jiu6;  // ../RTL/cortexm0ds_logic.v(561)
  wire T8kbx6;  // ../RTL/cortexm0ds_logic.v(1716)
  wire T8kow6;  // ../RTL/cortexm0ds_logic.v(1117)
  wire T8qiu6;  // ../RTL/cortexm0ds_logic.v(654)
  wire T8rhu6;  // ../RTL/cortexm0ds_logic.v(186)
  wire T8row6;  // ../RTL/cortexm0ds_logic.v(1211)
  wire T8xiu6;  // ../RTL/cortexm0ds_logic.v(748)
  wire T8yhu6;  // ../RTL/cortexm0ds_logic.v(280)
  wire T8yow6;  // ../RTL/cortexm0ds_logic.v(1304)
  wire T93ju6;  // ../RTL/cortexm0ds_logic.v(828)
  wire T94iu6;  // ../RTL/cortexm0ds_logic.v(360)
  wire T94pw6;  // ../RTL/cortexm0ds_logic.v(1385)
  wire T9aju6;  // ../RTL/cortexm0ds_logic.v(922)
  wire T9biu6;  // ../RTL/cortexm0ds_logic.v(454)
  wire T9bpw6;  // ../RTL/cortexm0ds_logic.v(1478)
  wire T9cow6;  // ../RTL/cortexm0ds_logic.v(1010)
  wire T9fbx6;  // ../RTL/cortexm0ds_logic.v(1707)
  wire T9iiu6;  // ../RTL/cortexm0ds_logic.v(548)
  wire T9jow6;  // ../RTL/cortexm0ds_logic.v(1104)
  wire T9kpw6;  // ../RTL/cortexm0ds_logic.v(1588)
  wire T9piu6;  // ../RTL/cortexm0ds_logic.v(641)
  wire T9qhu6;  // ../RTL/cortexm0ds_logic.v(173)
  wire T9qow6;  // ../RTL/cortexm0ds_logic.v(1198)
  wire T9wiu6;  // ../RTL/cortexm0ds_logic.v(735)
  wire T9xhu6;  // ../RTL/cortexm0ds_logic.v(267)
  wire T9xow6;  // ../RTL/cortexm0ds_logic.v(1291)
  wire Ta0qw6;  // ../RTL/cortexm0ds_logic.v(1617)
  wire Ta2ju6;  // ../RTL/cortexm0ds_logic.v(815)
  wire Ta3iu6;  // ../RTL/cortexm0ds_logic.v(347)
  wire Ta3pw6;  // ../RTL/cortexm0ds_logic.v(1372)
  wire Ta9ju6;  // ../RTL/cortexm0ds_logic.v(909)
  wire Taaiu6;  // ../RTL/cortexm0ds_logic.v(441)
  wire Taapw6;  // ../RTL/cortexm0ds_logic.v(1465)
  wire Tabow6;  // ../RTL/cortexm0ds_logic.v(997)
  wire Tahiu6;  // ../RTL/cortexm0ds_logic.v(535)
  wire Taiow6;  // ../RTL/cortexm0ds_logic.v(1091)
  wire Tajax6;  // ../RTL/cortexm0ds_logic.v(1649)
  wire Taoiu6;  // ../RTL/cortexm0ds_logic.v(628)
  wire Taphu6;  // ../RTL/cortexm0ds_logic.v(160)
  wire Tapow6;  // ../RTL/cortexm0ds_logic.v(1185)
  wire Taviu6;  // ../RTL/cortexm0ds_logic.v(722)
  wire Tawhu6;  // ../RTL/cortexm0ds_logic.v(254)
  wire Tawow6;  // ../RTL/cortexm0ds_logic.v(1278)
  wire Tb1ju6;  // ../RTL/cortexm0ds_logic.v(802)
  wire Tb2iu6;  // ../RTL/cortexm0ds_logic.v(334)
  wire Tb2pw6;  // ../RTL/cortexm0ds_logic.v(1359)
  wire Tb3qw6;  // ../RTL/cortexm0ds_logic.v(1623)
  wire Tb8ju6;  // ../RTL/cortexm0ds_logic.v(896)
  wire Tb9iu6;  // ../RTL/cortexm0ds_logic.v(428)
  wire Tb9pw6;  // ../RTL/cortexm0ds_logic.v(1452)
  wire Tbaow6;  // ../RTL/cortexm0ds_logic.v(984)
  wire Tbfbx6;  // ../RTL/cortexm0ds_logic.v(1707)
  wire Tbgiu6;  // ../RTL/cortexm0ds_logic.v(522)
  wire Tbhow6;  // ../RTL/cortexm0ds_logic.v(1078)
  wire Tbniu6;  // ../RTL/cortexm0ds_logic.v(615)
  wire Tbohu6;  // ../RTL/cortexm0ds_logic.v(147)
  wire Tboow6;  // ../RTL/cortexm0ds_logic.v(1172)
  wire Tbuiu6;  // ../RTL/cortexm0ds_logic.v(709)
  wire Tbvhu6;  // ../RTL/cortexm0ds_logic.v(241)
  wire Tbvow6;  // ../RTL/cortexm0ds_logic.v(1265)
  wire Tc0ju6;  // ../RTL/cortexm0ds_logic.v(789)
  wire Tc0qw6;  // ../RTL/cortexm0ds_logic.v(1618)
  wire Tc1iu6;  // ../RTL/cortexm0ds_logic.v(321)
  wire Tc1pw6;  // ../RTL/cortexm0ds_logic.v(1346)
  wire Tc7ju6;  // ../RTL/cortexm0ds_logic.v(883)
  wire Tc8iu6;  // ../RTL/cortexm0ds_logic.v(415)
  wire Tc8pw6;  // ../RTL/cortexm0ds_logic.v(1439)
  wire Tc9bx6;  // ../RTL/cortexm0ds_logic.v(1696)
  wire Tc9ow6;  // ../RTL/cortexm0ds_logic.v(971)
  wire Tceax6;  // ../RTL/cortexm0ds_logic.v(1640)
  wire Tcfiu6;  // ../RTL/cortexm0ds_logic.v(509)
  wire Tcgow6;  // ../RTL/cortexm0ds_logic.v(1065)
  wire Tchbx6;  // ../RTL/cortexm0ds_logic.v(1711)
  wire Tcipw6;  // ../RTL/cortexm0ds_logic.v(1585)
  wire Tcjax6;  // ../RTL/cortexm0ds_logic.v(1649)
  wire Tcjbx6;  // ../RTL/cortexm0ds_logic.v(1714)
  wire Tcmiu6;  // ../RTL/cortexm0ds_logic.v(602)
  wire Tcnow6;  // ../RTL/cortexm0ds_logic.v(1159)
  wire Tcrax6;  // ../RTL/cortexm0ds_logic.v(1664)
  wire Tctiu6;  // ../RTL/cortexm0ds_logic.v(696)
  wire Tcuhu6;  // ../RTL/cortexm0ds_logic.v(228)
  wire Tcuow6;  // ../RTL/cortexm0ds_logic.v(1252)
  wire Td0iu6;  // ../RTL/cortexm0ds_logic.v(308)
  wire Td0pw6;  // ../RTL/cortexm0ds_logic.v(1333)
  wire Td6ju6;  // ../RTL/cortexm0ds_logic.v(870)
  wire Td7iu6;  // ../RTL/cortexm0ds_logic.v(402)
  wire Td7pw6;  // ../RTL/cortexm0ds_logic.v(1426)
  wire Td8ow6;  // ../RTL/cortexm0ds_logic.v(958)
  wire Tdeiu6;  // ../RTL/cortexm0ds_logic.v(496)
  wire Tdfbx6;  // ../RTL/cortexm0ds_logic.v(1707)
  wire Tdfow6;  // ../RTL/cortexm0ds_logic.v(1052)
  wire Tdliu6;  // ../RTL/cortexm0ds_logic.v(589)
  wire Tdmow6;  // ../RTL/cortexm0ds_logic.v(1146)
  wire Tdsiu6;  // ../RTL/cortexm0ds_logic.v(683)
  wire Tdthu6;  // ../RTL/cortexm0ds_logic.v(215)
  wire Tdtow6;  // ../RTL/cortexm0ds_logic.v(1239)
  wire Tdypw6;  // ../RTL/cortexm0ds_logic.v(1614)
  wire Tdziu6;  // ../RTL/cortexm0ds_logic.v(776)
  wire Te0qw6;  // ../RTL/cortexm0ds_logic.v(1618)
  wire Te5ju6;  // ../RTL/cortexm0ds_logic.v(857)
  wire Te6iu6;  // ../RTL/cortexm0ds_logic.v(389)
  wire Te6pw6;  // ../RTL/cortexm0ds_logic.v(1413)
  wire Te7ow6;  // ../RTL/cortexm0ds_logic.v(945)
  wire Tediu6;  // ../RTL/cortexm0ds_logic.v(483)
  wire Tedpw6;  // ../RTL/cortexm0ds_logic.v(1507)
  wire Teeow6;  // ../RTL/cortexm0ds_logic.v(1039)
  wire Tekiu6;  // ../RTL/cortexm0ds_logic.v(576)
  wire Telow6;  // ../RTL/cortexm0ds_logic.v(1133)
  wire Teriu6;  // ../RTL/cortexm0ds_logic.v(670)
  wire Teshu6;  // ../RTL/cortexm0ds_logic.v(202)
  wire Tesow6;  // ../RTL/cortexm0ds_logic.v(1226)
  wire Teyiu6;  // ../RTL/cortexm0ds_logic.v(763)
  wire Tezhu6;  // ../RTL/cortexm0ds_logic.v(295)
  wire Tezow6;  // ../RTL/cortexm0ds_logic.v(1320)
  wire Tf4ju6;  // ../RTL/cortexm0ds_logic.v(844)
  wire Tf5iu6;  // ../RTL/cortexm0ds_logic.v(376)
  wire Tf5pw6;  // ../RTL/cortexm0ds_logic.v(1400)
  wire Tf6ow6;  // ../RTL/cortexm0ds_logic.v(932)
  wire Tfcax6;  // ../RTL/cortexm0ds_logic.v(1636)
  wire Tfciu6;  // ../RTL/cortexm0ds_logic.v(470)
  wire Tfcpw6;  // ../RTL/cortexm0ds_logic.v(1494)
  wire Tfdow6;  // ../RTL/cortexm0ds_logic.v(1026)
  wire Tffbx6;  // ../RTL/cortexm0ds_logic.v(1707)
  wire Tfjiu6;  // ../RTL/cortexm0ds_logic.v(563)
  wire Tfkow6;  // ../RTL/cortexm0ds_logic.v(1120)
  wire Tfqiu6;  // ../RTL/cortexm0ds_logic.v(657)
  wire Tfrhu6;  // ../RTL/cortexm0ds_logic.v(189)
  wire Tfrow6;  // ../RTL/cortexm0ds_logic.v(1213)
  wire Tfxiu6;  // ../RTL/cortexm0ds_logic.v(750)
  wire Tfyhu6;  // ../RTL/cortexm0ds_logic.v(282)
  wire Tfyow6;  // ../RTL/cortexm0ds_logic.v(1307)
  wire Tg0qw6;  // ../RTL/cortexm0ds_logic.v(1618)
  wire Tg3ju6;  // ../RTL/cortexm0ds_logic.v(831)
  wire Tg4iu6;  // ../RTL/cortexm0ds_logic.v(363)
  wire Tg4pw6;  // ../RTL/cortexm0ds_logic.v(1387)
  wire Tgaju6;  // ../RTL/cortexm0ds_logic.v(925)
  wire Tgbiu6;  // ../RTL/cortexm0ds_logic.v(457)
  wire Tgbpw6;  // ../RTL/cortexm0ds_logic.v(1481)
  wire Tgcow6;  // ../RTL/cortexm0ds_logic.v(1013)
  wire Tgiiu6;  // ../RTL/cortexm0ds_logic.v(550)
  wire Tgjow6;  // ../RTL/cortexm0ds_logic.v(1107)
  wire Tgkbx6;  // ../RTL/cortexm0ds_logic.v(1716)
  wire Tgpiu6;  // ../RTL/cortexm0ds_logic.v(644)
  wire Tgqhu6;  // ../RTL/cortexm0ds_logic.v(176)
  wire Tgqow6;  // ../RTL/cortexm0ds_logic.v(1200)
  wire Tgwiu6;  // ../RTL/cortexm0ds_logic.v(737)
  wire Tgxhu6;  // ../RTL/cortexm0ds_logic.v(269)
  wire Tgxow6;  // ../RTL/cortexm0ds_logic.v(1294)
  wire Tgzax6;  // ../RTL/cortexm0ds_logic.v(1678)
  wire Th2ju6;  // ../RTL/cortexm0ds_logic.v(818)
  wire Th3iu6;  // ../RTL/cortexm0ds_logic.v(350)
  wire Th3pw6;  // ../RTL/cortexm0ds_logic.v(1374)
  wire Th9ju6;  // ../RTL/cortexm0ds_logic.v(912)
  wire Thaiu6;  // ../RTL/cortexm0ds_logic.v(444)
  wire Thapw6;  // ../RTL/cortexm0ds_logic.v(1468)
  wire Thbow6;  // ../RTL/cortexm0ds_logic.v(1000)
  wire Thcbx6;  // ../RTL/cortexm0ds_logic.v(1702)
  wire Thfbx6;  // ../RTL/cortexm0ds_logic.v(1707)
  wire Thhax6;  // ../RTL/cortexm0ds_logic.v(1646)
  wire Thhiu6;  // ../RTL/cortexm0ds_logic.v(537)
  wire Thiax6;  // ../RTL/cortexm0ds_logic.v(1648)
  wire Thiow6;  // ../RTL/cortexm0ds_logic.v(1094)
  wire Thoiu6;  // ../RTL/cortexm0ds_logic.v(631)
  wire Thphu6;  // ../RTL/cortexm0ds_logic.v(163)
  wire Thpow6;  // ../RTL/cortexm0ds_logic.v(1187)
  wire Thviu6;  // ../RTL/cortexm0ds_logic.v(724)
  wire Thwhu6;  // ../RTL/cortexm0ds_logic.v(256)
  wire Thwow6;  // ../RTL/cortexm0ds_logic.v(1281)
  wire Thxax6;  // ../RTL/cortexm0ds_logic.v(1675)
  wire Ti0qw6;  // ../RTL/cortexm0ds_logic.v(1618)
  wire Ti1ju6;  // ../RTL/cortexm0ds_logic.v(805)
  wire Ti2iu6;  // ../RTL/cortexm0ds_logic.v(337)
  wire Ti2pw6;  // ../RTL/cortexm0ds_logic.v(1361)
  wire Ti8ju6;  // ../RTL/cortexm0ds_logic.v(899)
  wire Ti9iu6;  // ../RTL/cortexm0ds_logic.v(431)
  wire Ti9pw6;  // ../RTL/cortexm0ds_logic.v(1455)
  wire Tiaow6;  // ../RTL/cortexm0ds_logic.v(987)
  wire Tigiu6;  // ../RTL/cortexm0ds_logic.v(524)
  wire Tihow6;  // ../RTL/cortexm0ds_logic.v(1081)
  wire Tikbx6;  // ../RTL/cortexm0ds_logic.v(1716)
  wire Tiniu6;  // ../RTL/cortexm0ds_logic.v(618)
  wire Tiohu6;  // ../RTL/cortexm0ds_logic.v(150)
  wire Tioow6;  // ../RTL/cortexm0ds_logic.v(1174)
  wire Tiuiu6;  // ../RTL/cortexm0ds_logic.v(711)
  wire Tivhu6;  // ../RTL/cortexm0ds_logic.v(243)
  wire Tivow6;  // ../RTL/cortexm0ds_logic.v(1268)
  wire Tj0ju6;  // ../RTL/cortexm0ds_logic.v(792)
  wire Tj1iu6;  // ../RTL/cortexm0ds_logic.v(324)
  wire Tj1pw6;  // ../RTL/cortexm0ds_logic.v(1348)
  wire Tj7ju6;  // ../RTL/cortexm0ds_logic.v(886)
  wire Tj8iu6;  // ../RTL/cortexm0ds_logic.v(418)
  wire Tj8pw6;  // ../RTL/cortexm0ds_logic.v(1442)
  wire Tj9ow6;  // ../RTL/cortexm0ds_logic.v(974)
  wire Tjfbx6;  // ../RTL/cortexm0ds_logic.v(1707)
  wire Tjfiu6;  // ../RTL/cortexm0ds_logic.v(511)
  wire Tjgow6;  // ../RTL/cortexm0ds_logic.v(1068)
  wire Tjkpw6;  // ../RTL/cortexm0ds_logic.v(1589)
  wire Tjmiu6;  // ../RTL/cortexm0ds_logic.v(605)
  wire Tjnow6;  // ../RTL/cortexm0ds_logic.v(1161)
  wire Tjtiu6;  // ../RTL/cortexm0ds_logic.v(698)
  wire Tjuhu6;  // ../RTL/cortexm0ds_logic.v(230)
  wire Tjuow6;  // ../RTL/cortexm0ds_logic.v(1255)
  wire Tjvax6;  // ../RTL/cortexm0ds_logic.v(1671)
  wire Tk0iu6;  // ../RTL/cortexm0ds_logic.v(311)
  wire Tk0pw6;  // ../RTL/cortexm0ds_logic.v(1335)
  wire Tk0qw6;  // ../RTL/cortexm0ds_logic.v(1618)
  wire Tk6ju6;  // ../RTL/cortexm0ds_logic.v(873)
  wire Tk7iu6;  // ../RTL/cortexm0ds_logic.v(405)
  wire Tk7pw6;  // ../RTL/cortexm0ds_logic.v(1429)
  wire Tk8ow6;  // ../RTL/cortexm0ds_logic.v(961)
  wire Tkdax6;  // ../RTL/cortexm0ds_logic.v(1638)
  wire Tkeiu6;  // ../RTL/cortexm0ds_logic.v(498)
  wire Tkfow6;  // ../RTL/cortexm0ds_logic.v(1055)
  wire Tkjbx6;  // ../RTL/cortexm0ds_logic.v(1715)
  wire Tkliu6;  // ../RTL/cortexm0ds_logic.v(592)
  wire Tkmow6;  // ../RTL/cortexm0ds_logic.v(1148)
  wire Tksiu6;  // ../RTL/cortexm0ds_logic.v(685)
  wire Tkthu6;  // ../RTL/cortexm0ds_logic.v(217)
  wire Tktow6;  // ../RTL/cortexm0ds_logic.v(1242)
  wire Tkziu6;  // ../RTL/cortexm0ds_logic.v(779)
  wire Tl4bx6;  // ../RTL/cortexm0ds_logic.v(1687)
  wire Tl5ju6;  // ../RTL/cortexm0ds_logic.v(860)
  wire Tl6iu6;  // ../RTL/cortexm0ds_logic.v(392)
  wire Tl6pw6;  // ../RTL/cortexm0ds_logic.v(1416)
  wire Tl7ow6;  // ../RTL/cortexm0ds_logic.v(948)
  wire Tldiu6;  // ../RTL/cortexm0ds_logic.v(485)
  wire Tldpw6;  // ../RTL/cortexm0ds_logic.v(1510)
  wire Tlebx6;  // ../RTL/cortexm0ds_logic.v(1706)
  wire Tleow6;  // ../RTL/cortexm0ds_logic.v(1042)
  wire Tlkiu6;  // ../RTL/cortexm0ds_logic.v(579)
  wire Tllow6;  // ../RTL/cortexm0ds_logic.v(1135)
  wire Tlriu6;  // ../RTL/cortexm0ds_logic.v(672)
  wire Tlshu6;  // ../RTL/cortexm0ds_logic.v(204)
  wire Tlsow6;  // ../RTL/cortexm0ds_logic.v(1229)
  wire Tlyiu6;  // ../RTL/cortexm0ds_logic.v(766)
  wire Tlzhu6;  // ../RTL/cortexm0ds_logic.v(298)
  wire Tlzow6;  // ../RTL/cortexm0ds_logic.v(1322)
  wire Tm0qw6;  // ../RTL/cortexm0ds_logic.v(1618)
  wire Tm4ju6;  // ../RTL/cortexm0ds_logic.v(847)
  wire Tm5iu6;  // ../RTL/cortexm0ds_logic.v(379)
  wire Tm5pw6;  // ../RTL/cortexm0ds_logic.v(1403)
  wire Tm6ow6;  // ../RTL/cortexm0ds_logic.v(935)
  wire Tmciu6;  // ../RTL/cortexm0ds_logic.v(472)
  wire Tmcpw6;  // ../RTL/cortexm0ds_logic.v(1497)
  wire Tmdow6;  // ../RTL/cortexm0ds_logic.v(1029)
  wire Tmjbx6;  // ../RTL/cortexm0ds_logic.v(1715)
  wire Tmjiu6;  // ../RTL/cortexm0ds_logic.v(566)
  wire Tmkow6;  // ../RTL/cortexm0ds_logic.v(1122)
  wire Tmqiu6;  // ../RTL/cortexm0ds_logic.v(659)
  wire Tmrhu6;  // ../RTL/cortexm0ds_logic.v(191)
  wire Tmrow6;  // ../RTL/cortexm0ds_logic.v(1216)
  wire Tmxiu6;  // ../RTL/cortexm0ds_logic.v(753)
  wire Tmyhu6;  // ../RTL/cortexm0ds_logic.v(285)
  wire Tmyow6;  // ../RTL/cortexm0ds_logic.v(1309)
  wire Tn3ju6;  // ../RTL/cortexm0ds_logic.v(834)
  wire Tn4iu6;  // ../RTL/cortexm0ds_logic.v(366)
  wire Tn4pw6;  // ../RTL/cortexm0ds_logic.v(1390)
  wire Tnaju6;  // ../RTL/cortexm0ds_logic.v(927)
  wire Tnbiu6;  // ../RTL/cortexm0ds_logic.v(459)
  wire Tnbpw6;  // ../RTL/cortexm0ds_logic.v(1484)
  wire Tncow6;  // ../RTL/cortexm0ds_logic.v(1016)
  wire Tnebx6;  // ../RTL/cortexm0ds_logic.v(1706)
  wire Tngbx6;  // ../RTL/cortexm0ds_logic.v(1709)
  wire Tniiu6;  // ../RTL/cortexm0ds_logic.v(553)
  wire Tnjow6;  // ../RTL/cortexm0ds_logic.v(1109)
  wire Tnpiu6;  // ../RTL/cortexm0ds_logic.v(646)
  wire Tnqhu6;  // ../RTL/cortexm0ds_logic.v(178)
  wire Tnqow6;  // ../RTL/cortexm0ds_logic.v(1203)
  wire Tnwiu6;  // ../RTL/cortexm0ds_logic.v(740)
  wire Tnxhu6;  // ../RTL/cortexm0ds_logic.v(272)
  wire Tnxow6;  // ../RTL/cortexm0ds_logic.v(1296)
  wire To2ju6;  // ../RTL/cortexm0ds_logic.v(821)
  wire To3iu6;  // ../RTL/cortexm0ds_logic.v(353)
  wire To3pw6;  // ../RTL/cortexm0ds_logic.v(1377)
  wire To9ju6;  // ../RTL/cortexm0ds_logic.v(914)
  wire Toaiu6;  // ../RTL/cortexm0ds_logic.v(446)
  wire Toapw6;  // ../RTL/cortexm0ds_logic.v(1471)
  wire Tobow6;  // ../RTL/cortexm0ds_logic.v(1003)
  wire Tohiu6;  // ../RTL/cortexm0ds_logic.v(540)
  wire Toiow6;  // ../RTL/cortexm0ds_logic.v(1096)
  wire Tokax6;  // ../RTL/cortexm0ds_logic.v(1652)
  wire Tonhu6;  // ../RTL/cortexm0ds_logic.v(145)
  wire Tooiu6;  // ../RTL/cortexm0ds_logic.v(633)
  wire Tophu6;  // ../RTL/cortexm0ds_logic.v(165)
  wire Topow6;  // ../RTL/cortexm0ds_logic.v(1190)
  wire Toviu6;  // ../RTL/cortexm0ds_logic.v(727)
  wire Towhu6;  // ../RTL/cortexm0ds_logic.v(259)
  wire Towow6;  // ../RTL/cortexm0ds_logic.v(1283)
  wire Tp1ju6;  // ../RTL/cortexm0ds_logic.v(808)
  wire Tp2iu6;  // ../RTL/cortexm0ds_logic.v(340)
  wire Tp2pw6;  // ../RTL/cortexm0ds_logic.v(1364)
  wire Tp8ju6;  // ../RTL/cortexm0ds_logic.v(901)
  wire Tp9iu6;  // ../RTL/cortexm0ds_logic.v(433)
  wire Tp9pw6;  // ../RTL/cortexm0ds_logic.v(1458)
  wire Tpaow6;  // ../RTL/cortexm0ds_logic.v(990)
  wire Tpebx6;  // ../RTL/cortexm0ds_logic.v(1706)
  wire Tpgiu6;  // ../RTL/cortexm0ds_logic.v(527)
  wire Tphow6;  // ../RTL/cortexm0ds_logic.v(1083)
  wire Tpniu6;  // ../RTL/cortexm0ds_logic.v(620)
  wire Tpohu6;  // ../RTL/cortexm0ds_logic.v(152)
  wire Tpoow6;  // ../RTL/cortexm0ds_logic.v(1177)
  wire Tptpw6;  // ../RTL/cortexm0ds_logic.v(1605)
  wire Tpuiu6;  // ../RTL/cortexm0ds_logic.v(714)
  wire Tpvhu6;  // ../RTL/cortexm0ds_logic.v(246)
  wire Tpvow6;  // ../RTL/cortexm0ds_logic.v(1270)
  wire Tq0ju6;  // ../RTL/cortexm0ds_logic.v(795)
  wire Tq1iu6;  // ../RTL/cortexm0ds_logic.v(327)
  wire Tq1pw6;  // ../RTL/cortexm0ds_logic.v(1351)
  wire Tq7ju6;  // ../RTL/cortexm0ds_logic.v(888)
  wire Tq8iu6;  // ../RTL/cortexm0ds_logic.v(420)
  wire Tq8pw6;  // ../RTL/cortexm0ds_logic.v(1445)
  wire Tq9ow6;  // ../RTL/cortexm0ds_logic.v(977)
  wire Tqfiu6;  // ../RTL/cortexm0ds_logic.v(514)
  wire Tqgow6;  // ../RTL/cortexm0ds_logic.v(1070)
  wire Tqmiu6;  // ../RTL/cortexm0ds_logic.v(607)
  wire Tqnow6;  // ../RTL/cortexm0ds_logic.v(1164)
  wire Tqtiu6;  // ../RTL/cortexm0ds_logic.v(701)
  wire Tquhu6;  // ../RTL/cortexm0ds_logic.v(233)
  wire Tquow6;  // ../RTL/cortexm0ds_logic.v(1257)
  wire Tr0iu6;  // ../RTL/cortexm0ds_logic.v(314)
  wire Tr0pw6;  // ../RTL/cortexm0ds_logic.v(1338)
  wire Tr6ju6;  // ../RTL/cortexm0ds_logic.v(875)
  wire Tr7iu6;  // ../RTL/cortexm0ds_logic.v(407)
  wire Tr7pw6;  // ../RTL/cortexm0ds_logic.v(1432)
  wire Tr8ow6;  // ../RTL/cortexm0ds_logic.v(964)
  wire Trebx6;  // ../RTL/cortexm0ds_logic.v(1706)
  wire Treiu6;  // ../RTL/cortexm0ds_logic.v(501)
  wire Trfow6;  // ../RTL/cortexm0ds_logic.v(1057)
  wire Trliu6;  // ../RTL/cortexm0ds_logic.v(594)
  wire Trmow6;  // ../RTL/cortexm0ds_logic.v(1151)
  wire Trsiu6;  // ../RTL/cortexm0ds_logic.v(688)
  wire Trthu6;  // ../RTL/cortexm0ds_logic.v(220)
  wire Trtow6;  // ../RTL/cortexm0ds_logic.v(1244)
  wire Trziu6;  // ../RTL/cortexm0ds_logic.v(782)
  wire Ts5ju6;  // ../RTL/cortexm0ds_logic.v(862)
  wire Ts6iu6;  // ../RTL/cortexm0ds_logic.v(394)
  wire Ts6pw6;  // ../RTL/cortexm0ds_logic.v(1419)
  wire Ts7ow6;  // ../RTL/cortexm0ds_logic.v(951)
  wire Tsdbx6;  // ../RTL/cortexm0ds_logic.v(1704)
  wire Tsdiu6;  // ../RTL/cortexm0ds_logic.v(488)
  wire Tsdpw6;  // ../RTL/cortexm0ds_logic.v(1512)
  wire Tseow6;  // ../RTL/cortexm0ds_logic.v(1044)
  wire Tskiu6;  // ../RTL/cortexm0ds_logic.v(581)
  wire Tslow6;  // ../RTL/cortexm0ds_logic.v(1138)
  wire Tsriu6;  // ../RTL/cortexm0ds_logic.v(675)
  wire Tsshu6;  // ../RTL/cortexm0ds_logic.v(207)
  wire Tssow6;  // ../RTL/cortexm0ds_logic.v(1231)
  wire Tsyiu6;  // ../RTL/cortexm0ds_logic.v(769)
  wire Tszhu6;  // ../RTL/cortexm0ds_logic.v(301)
  wire Tszow6;  // ../RTL/cortexm0ds_logic.v(1325)
  wire Tt4ju6;  // ../RTL/cortexm0ds_logic.v(849)
  wire Tt5iu6;  // ../RTL/cortexm0ds_logic.v(381)
  wire Tt5pw6;  // ../RTL/cortexm0ds_logic.v(1406)
  wire Tt6ow6;  // ../RTL/cortexm0ds_logic.v(938)
  wire Tt9ax6;  // ../RTL/cortexm0ds_logic.v(1631)
  wire Ttciu6;  // ../RTL/cortexm0ds_logic.v(475)
  wire Ttcpw6;  // ../RTL/cortexm0ds_logic.v(1499)
  wire Ttdow6;  // ../RTL/cortexm0ds_logic.v(1031)
  wire Ttebx6;  // ../RTL/cortexm0ds_logic.v(1706)
  wire Ttjiu6;  // ../RTL/cortexm0ds_logic.v(568)
  wire Ttkow6;  // ../RTL/cortexm0ds_logic.v(1125)
  wire Ttmhu6;  // ../RTL/cortexm0ds_logic.v(143)
  wire Ttqiu6;  // ../RTL/cortexm0ds_logic.v(662)
  wire Ttrhu6;  // ../RTL/cortexm0ds_logic.v(194)
  wire Ttrow6;  // ../RTL/cortexm0ds_logic.v(1218)
  wire Ttxiu6;  // ../RTL/cortexm0ds_logic.v(756)
  wire Ttyhu6;  // ../RTL/cortexm0ds_logic.v(288)
  wire Ttyow6;  // ../RTL/cortexm0ds_logic.v(1312)
  wire Tu0qw6;  // ../RTL/cortexm0ds_logic.v(1618)
  wire Tu3ju6;  // ../RTL/cortexm0ds_logic.v(836)
  wire Tu4iu6;  // ../RTL/cortexm0ds_logic.v(368)
  wire Tu4pw6;  // ../RTL/cortexm0ds_logic.v(1393)
  wire Tubiu6;  // ../RTL/cortexm0ds_logic.v(462)
  wire Tubpw6;  // ../RTL/cortexm0ds_logic.v(1486)
  wire Tucow6;  // ../RTL/cortexm0ds_logic.v(1018)
  wire Tuiiu6;  // ../RTL/cortexm0ds_logic.v(555)
  wire Tujbx6;  // ../RTL/cortexm0ds_logic.v(1715)
  wire Tujow6;  // ../RTL/cortexm0ds_logic.v(1112)
  wire Tupiu6;  // ../RTL/cortexm0ds_logic.v(649)
  wire Tuqhu6;  // ../RTL/cortexm0ds_logic.v(181)
  wire Tuqow6;  // ../RTL/cortexm0ds_logic.v(1205)
  wire Tuwiu6;  // ../RTL/cortexm0ds_logic.v(743)
  wire Tuxhu6;  // ../RTL/cortexm0ds_logic.v(275)
  wire Tuxow6;  // ../RTL/cortexm0ds_logic.v(1299)
  wire Tv2ju6;  // ../RTL/cortexm0ds_logic.v(823)
  wire Tv3iu6;  // ../RTL/cortexm0ds_logic.v(355)
  wire Tv3pw6;  // ../RTL/cortexm0ds_logic.v(1380)
  wire Tv9ju6;  // ../RTL/cortexm0ds_logic.v(917)
  wire Tvaiu6;  // ../RTL/cortexm0ds_logic.v(449)
  wire Tvapw6;  // ../RTL/cortexm0ds_logic.v(1473)
  wire Tvbow6;  // ../RTL/cortexm0ds_logic.v(1005)
  wire Tvebx6;  // ../RTL/cortexm0ds_logic.v(1706)
  wire Tvhiu6;  // ../RTL/cortexm0ds_logic.v(542)
  wire Tviow6;  // ../RTL/cortexm0ds_logic.v(1099)
  wire Tvoiu6;  // ../RTL/cortexm0ds_logic.v(636)
  wire Tvphu6;  // ../RTL/cortexm0ds_logic.v(168)
  wire Tvpow6;  // ../RTL/cortexm0ds_logic.v(1192)
  wire Tvviu6;  // ../RTL/cortexm0ds_logic.v(730)
  wire Tvwhu6;  // ../RTL/cortexm0ds_logic.v(262)
  wire Tvwow6;  // ../RTL/cortexm0ds_logic.v(1286)
  wire Tw1ju6;  // ../RTL/cortexm0ds_logic.v(810)
  wire Tw2iu6;  // ../RTL/cortexm0ds_logic.v(342)
  wire Tw2pw6;  // ../RTL/cortexm0ds_logic.v(1367)
  wire Tw8ju6;  // ../RTL/cortexm0ds_logic.v(904)
  wire Tw9iu6;  // ../RTL/cortexm0ds_logic.v(436)
  wire Tw9pw6;  // ../RTL/cortexm0ds_logic.v(1460)
  wire Twaow6;  // ../RTL/cortexm0ds_logic.v(992)
  wire Twgiu6;  // ../RTL/cortexm0ds_logic.v(529)
  wire Twhow6;  // ../RTL/cortexm0ds_logic.v(1086)
  wire Twlhu6;  // ../RTL/cortexm0ds_logic.v(140)
  wire Twniu6;  // ../RTL/cortexm0ds_logic.v(623)
  wire Twohu6;  // ../RTL/cortexm0ds_logic.v(155)
  wire Twoow6;  // ../RTL/cortexm0ds_logic.v(1179)
  wire Twuiu6;  // ../RTL/cortexm0ds_logic.v(717)
  wire Twvhu6;  // ../RTL/cortexm0ds_logic.v(249)
  wire Twvow6;  // ../RTL/cortexm0ds_logic.v(1273)
  wire Twzpw6;  // ../RTL/cortexm0ds_logic.v(1617)
  wire Tx0ju6;  // ../RTL/cortexm0ds_logic.v(797)
  wire Tx1iu6;  // ../RTL/cortexm0ds_logic.v(329)
  wire Tx1pw6;  // ../RTL/cortexm0ds_logic.v(1354)
  wire Tx7ju6;  // ../RTL/cortexm0ds_logic.v(891)
  wire Tx8iu6;  // ../RTL/cortexm0ds_logic.v(423)
  wire Tx8pw6;  // ../RTL/cortexm0ds_logic.v(1447)
  wire Tx9ow6;  // ../RTL/cortexm0ds_logic.v(979)
  wire Txebx6;  // ../RTL/cortexm0ds_logic.v(1706)
  wire Txfiu6;  // ../RTL/cortexm0ds_logic.v(516)
  wire Txgow6;  // ../RTL/cortexm0ds_logic.v(1073)
  wire Txmax6;  // ../RTL/cortexm0ds_logic.v(1656)
  wire Txmiu6;  // ../RTL/cortexm0ds_logic.v(610)
  wire Txnow6;  // ../RTL/cortexm0ds_logic.v(1166)
  wire Txtiu6;  // ../RTL/cortexm0ds_logic.v(704)
  wire Txuhu6;  // ../RTL/cortexm0ds_logic.v(236)
  wire Txuow6;  // ../RTL/cortexm0ds_logic.v(1260)
  wire Ty0iu6;  // ../RTL/cortexm0ds_logic.v(316)
  wire Ty0pw6;  // ../RTL/cortexm0ds_logic.v(1341)
  wire Ty6ju6;  // ../RTL/cortexm0ds_logic.v(878)
  wire Ty7iu6;  // ../RTL/cortexm0ds_logic.v(410)
  wire Ty7pw6;  // ../RTL/cortexm0ds_logic.v(1434)
  wire Ty8ow6;  // ../RTL/cortexm0ds_logic.v(966)
  wire Tyaax6;  // ../RTL/cortexm0ds_logic.v(1633)
  wire Tyeiu6;  // ../RTL/cortexm0ds_logic.v(503)
  wire Tyfow6;  // ../RTL/cortexm0ds_logic.v(1060)
  wire Tyipw6;  // ../RTL/cortexm0ds_logic.v(1586)
  wire Tyliu6;  // ../RTL/cortexm0ds_logic.v(597)
  wire Tymow6;  // ../RTL/cortexm0ds_logic.v(1153)
  wire Tysiu6;  // ../RTL/cortexm0ds_logic.v(691)
  wire Tythu6;  // ../RTL/cortexm0ds_logic.v(223)
  wire Tytow6;  // ../RTL/cortexm0ds_logic.v(1247)
  wire Tyziu6;  // ../RTL/cortexm0ds_logic.v(784)
  wire Tyzpw6;  // ../RTL/cortexm0ds_logic.v(1617)
  wire Tz5ju6;  // ../RTL/cortexm0ds_logic.v(865)
  wire Tz6iu6;  // ../RTL/cortexm0ds_logic.v(397)
  wire Tz6pw6;  // ../RTL/cortexm0ds_logic.v(1421)
  wire Tz7ow6;  // ../RTL/cortexm0ds_logic.v(953)
  wire Tzdiu6;  // ../RTL/cortexm0ds_logic.v(490)
  wire Tzdpw6;  // ../RTL/cortexm0ds_logic.v(1515)
  wire Tzebx6;  // ../RTL/cortexm0ds_logic.v(1706)
  wire Tzeow6;  // ../RTL/cortexm0ds_logic.v(1047)
  wire Tzgbx6;  // ../RTL/cortexm0ds_logic.v(1710)
  wire Tzkiu6;  // ../RTL/cortexm0ds_logic.v(584)
  wire Tzlow6;  // ../RTL/cortexm0ds_logic.v(1140)
  wire Tzriu6;  // ../RTL/cortexm0ds_logic.v(678)
  wire Tzshu6;  // ../RTL/cortexm0ds_logic.v(210)
  wire Tzsow6;  // ../RTL/cortexm0ds_logic.v(1234)
  wire Tzyiu6;  // ../RTL/cortexm0ds_logic.v(771)
  wire Tzzhu6;  // ../RTL/cortexm0ds_logic.v(303)
  wire Tzzow6;  // ../RTL/cortexm0ds_logic.v(1328)
  wire U02ju6;  // ../RTL/cortexm0ds_logic.v(812)
  wire U03iu6;  // ../RTL/cortexm0ds_logic.v(344)
  wire U03pw6;  // ../RTL/cortexm0ds_logic.v(1368)
  wire U09ju6;  // ../RTL/cortexm0ds_logic.v(905)
  wire U0aiu6;  // ../RTL/cortexm0ds_logic.v(437)
  wire U0apw6;  // ../RTL/cortexm0ds_logic.v(1462)
  wire U0bow6;  // ../RTL/cortexm0ds_logic.v(994)
  wire U0hax6;  // ../RTL/cortexm0ds_logic.v(1645)
  wire U0hiu6;  // ../RTL/cortexm0ds_logic.v(531)
  wire U0iow6;  // ../RTL/cortexm0ds_logic.v(1087)
  wire U0jhu6;  // ../RTL/cortexm0ds_logic.v(132)
  wire U0oiu6;  // ../RTL/cortexm0ds_logic.v(625)
  wire U0phu6;  // ../RTL/cortexm0ds_logic.v(157)
  wire U0pow6;  // ../RTL/cortexm0ds_logic.v(1181)
  wire U0rax6;  // ../RTL/cortexm0ds_logic.v(1663)
  wire U0viu6;  // ../RTL/cortexm0ds_logic.v(718)
  wire U0whu6;  // ../RTL/cortexm0ds_logic.v(250)
  wire U0wow6;  // ../RTL/cortexm0ds_logic.v(1275)
  wire U11ju6;  // ../RTL/cortexm0ds_logic.v(799)
  wire U12iu6;  // ../RTL/cortexm0ds_logic.v(331)
  wire U12pw6;  // ../RTL/cortexm0ds_logic.v(1355)
  wire U18ju6;  // ../RTL/cortexm0ds_logic.v(892)
  wire U19iu6;  // ../RTL/cortexm0ds_logic.v(424)
  wire U19pw6;  // ../RTL/cortexm0ds_logic.v(1449)
  wire U1aow6;  // ../RTL/cortexm0ds_logic.v(981)
  wire U1fhu6;  // ../RTL/cortexm0ds_logic.v(123)
  wire U1giu6;  // ../RTL/cortexm0ds_logic.v(518)
  wire U1how6;  // ../RTL/cortexm0ds_logic.v(1074)
  wire U1kpw6;  // ../RTL/cortexm0ds_logic.v(1588)
  wire U1niu6;  // ../RTL/cortexm0ds_logic.v(612)
  wire U1oow6;  // ../RTL/cortexm0ds_logic.v(1168)
  wire U1uiu6;  // ../RTL/cortexm0ds_logic.v(705)
  wire U1vhu6;  // ../RTL/cortexm0ds_logic.v(237)
  wire U1vow6;  // ../RTL/cortexm0ds_logic.v(1262)
  wire U20ju6;  // ../RTL/cortexm0ds_logic.v(786)
  wire U21iu6;  // ../RTL/cortexm0ds_logic.v(318)
  wire U21pw6;  // ../RTL/cortexm0ds_logic.v(1342)
  wire U27ju6;  // ../RTL/cortexm0ds_logic.v(879)
  wire U28iu6;  // ../RTL/cortexm0ds_logic.v(411)
  wire U28pw6;  // ../RTL/cortexm0ds_logic.v(1436)
  wire U29ow6;  // ../RTL/cortexm0ds_logic.v(968)
  wire U2fiu6;  // ../RTL/cortexm0ds_logic.v(505)
  wire U2gow6;  // ../RTL/cortexm0ds_logic.v(1061)
  wire U2ihu6;  // ../RTL/cortexm0ds_logic.v(130)
  wire U2miu6;  // ../RTL/cortexm0ds_logic.v(599)
  wire U2now6;  // ../RTL/cortexm0ds_logic.v(1155)
  wire U2rax6;  // ../RTL/cortexm0ds_logic.v(1663)
  wire U2tiu6;  // ../RTL/cortexm0ds_logic.v(692)
  wire U2uhu6;  // ../RTL/cortexm0ds_logic.v(224)
  wire U2uow6;  // ../RTL/cortexm0ds_logic.v(1249)
  wire U30iu6;  // ../RTL/cortexm0ds_logic.v(305)
  wire U30pw6;  // ../RTL/cortexm0ds_logic.v(1329)
  wire U31bx6;  // ../RTL/cortexm0ds_logic.v(1681)
  wire U36ju6;  // ../RTL/cortexm0ds_logic.v(866)
  wire U37iu6;  // ../RTL/cortexm0ds_logic.v(398)
  wire U37pw6;  // ../RTL/cortexm0ds_logic.v(1423)
  wire U38ow6;  // ../RTL/cortexm0ds_logic.v(955)
  wire U3eiu6;  // ../RTL/cortexm0ds_logic.v(492)
  wire U3epw6;  // ../RTL/cortexm0ds_logic.v(1516)
  wire U3fow6;  // ../RTL/cortexm0ds_logic.v(1048)
  wire U3liu6;  // ../RTL/cortexm0ds_logic.v(586)
  wire U3mow6;  // ../RTL/cortexm0ds_logic.v(1142)
  wire U3siu6;  // ../RTL/cortexm0ds_logic.v(679)
  wire U3thu6;  // ../RTL/cortexm0ds_logic.v(211)
  wire U3tow6;  // ../RTL/cortexm0ds_logic.v(1236)
  wire U3yax6;  // ../RTL/cortexm0ds_logic.v(1676)
  wire U3ziu6;  // ../RTL/cortexm0ds_logic.v(773)
  wire U45ju6;  // ../RTL/cortexm0ds_logic.v(853)
  wire U46iu6;  // ../RTL/cortexm0ds_logic.v(385)
  wire U46pw6;  // ../RTL/cortexm0ds_logic.v(1410)
  wire U47ow6;  // ../RTL/cortexm0ds_logic.v(942)
  wire U4diu6;  // ../RTL/cortexm0ds_logic.v(479)
  wire U4dpw6;  // ../RTL/cortexm0ds_logic.v(1503)
  wire U4eow6;  // ../RTL/cortexm0ds_logic.v(1035)
  wire U4fax6;  // ../RTL/cortexm0ds_logic.v(1641)
  wire U4kiu6;  // ../RTL/cortexm0ds_logic.v(573)
  wire U4low6;  // ../RTL/cortexm0ds_logic.v(1129)
  wire U4rax6;  // ../RTL/cortexm0ds_logic.v(1663)
  wire U4riu6;  // ../RTL/cortexm0ds_logic.v(666)
  wire U4shu6;  // ../RTL/cortexm0ds_logic.v(198)
  wire U4sow6;  // ../RTL/cortexm0ds_logic.v(1223)
  wire U4yiu6;  // ../RTL/cortexm0ds_logic.v(760)
  wire U4zhu6;  // ../RTL/cortexm0ds_logic.v(292)
  wire U4zow6;  // ../RTL/cortexm0ds_logic.v(1316)
  wire U54ju6;  // ../RTL/cortexm0ds_logic.v(840)
  wire U55iu6;  // ../RTL/cortexm0ds_logic.v(372)
  wire U55pw6;  // ../RTL/cortexm0ds_logic.v(1397)
  wire U5ciu6;  // ../RTL/cortexm0ds_logic.v(466)
  wire U5cpw6;  // ../RTL/cortexm0ds_logic.v(1490)
  wire U5dow6;  // ../RTL/cortexm0ds_logic.v(1022)
  wire U5jiu6;  // ../RTL/cortexm0ds_logic.v(560)
  wire U5kow6;  // ../RTL/cortexm0ds_logic.v(1116)
  wire U5qiu6;  // ../RTL/cortexm0ds_logic.v(653)
  wire U5rhu6;  // ../RTL/cortexm0ds_logic.v(185)
  wire U5row6;  // ../RTL/cortexm0ds_logic.v(1210)
  wire U5xiu6;  // ../RTL/cortexm0ds_logic.v(747)
  wire U5yhu6;  // ../RTL/cortexm0ds_logic.v(279)
  wire U5yow6;  // ../RTL/cortexm0ds_logic.v(1303)
  wire U63ju6;  // ../RTL/cortexm0ds_logic.v(827)
  wire U64iu6;  // ../RTL/cortexm0ds_logic.v(359)
  wire U64pw6;  // ../RTL/cortexm0ds_logic.v(1384)
  wire U6aju6;  // ../RTL/cortexm0ds_logic.v(921)
  wire U6biu6;  // ../RTL/cortexm0ds_logic.v(453)
  wire U6bpw6;  // ../RTL/cortexm0ds_logic.v(1477)
  wire U6cow6;  // ../RTL/cortexm0ds_logic.v(1009)
  wire U6iiu6;  // ../RTL/cortexm0ds_logic.v(547)
  wire U6jow6;  // ../RTL/cortexm0ds_logic.v(1103)
  wire U6piu6;  // ../RTL/cortexm0ds_logic.v(640)
  wire U6qhu6;  // ../RTL/cortexm0ds_logic.v(172)
  wire U6qow6;  // ../RTL/cortexm0ds_logic.v(1197)
  wire U6rax6;  // ../RTL/cortexm0ds_logic.v(1663)
  wire U6wiu6;  // ../RTL/cortexm0ds_logic.v(734)
  wire U6xhu6;  // ../RTL/cortexm0ds_logic.v(266)
  wire U6xow6;  // ../RTL/cortexm0ds_logic.v(1290)
  wire U72ju6;  // ../RTL/cortexm0ds_logic.v(814)
  wire U73iu6;  // ../RTL/cortexm0ds_logic.v(346)
  wire U73pw6;  // ../RTL/cortexm0ds_logic.v(1371)
  wire U79ju6;  // ../RTL/cortexm0ds_logic.v(908)
  wire U7aiu6;  // ../RTL/cortexm0ds_logic.v(440)
  wire U7apw6;  // ../RTL/cortexm0ds_logic.v(1464)
  wire U7bow6;  // ../RTL/cortexm0ds_logic.v(996)
  wire U7dax6;  // ../RTL/cortexm0ds_logic.v(1637)
  wire U7hiu6;  // ../RTL/cortexm0ds_logic.v(534)
  wire U7iow6;  // ../RTL/cortexm0ds_logic.v(1090)
  wire U7oiu6;  // ../RTL/cortexm0ds_logic.v(627)
  wire U7phu6;  // ../RTL/cortexm0ds_logic.v(159)
  wire U7pow6;  // ../RTL/cortexm0ds_logic.v(1184)
  wire U7viu6;  // ../RTL/cortexm0ds_logic.v(721)
  wire U7whu6;  // ../RTL/cortexm0ds_logic.v(253)
  wire U7wow6;  // ../RTL/cortexm0ds_logic.v(1277)
  wire U81ju6;  // ../RTL/cortexm0ds_logic.v(801)
  wire U82iu6;  // ../RTL/cortexm0ds_logic.v(333)
  wire U82pw6;  // ../RTL/cortexm0ds_logic.v(1358)
  wire U88ju6;  // ../RTL/cortexm0ds_logic.v(895)
  wire U89iu6;  // ../RTL/cortexm0ds_logic.v(427)
  wire U89pw6;  // ../RTL/cortexm0ds_logic.v(1451)
  wire U8aow6;  // ../RTL/cortexm0ds_logic.v(983)
  wire U8giu6;  // ../RTL/cortexm0ds_logic.v(521)
  wire U8how6;  // ../RTL/cortexm0ds_logic.v(1077)
  wire U8jax6;  // ../RTL/cortexm0ds_logic.v(1649)
  wire U8niu6;  // ../RTL/cortexm0ds_logic.v(614)
  wire U8oow6;  // ../RTL/cortexm0ds_logic.v(1171)
  wire U8rax6;  // ../RTL/cortexm0ds_logic.v(1664)
  wire U8uiu6;  // ../RTL/cortexm0ds_logic.v(708)
  wire U8vhu6;  // ../RTL/cortexm0ds_logic.v(240)
  wire U8vow6;  // ../RTL/cortexm0ds_logic.v(1264)
  wire U90ju6;  // ../RTL/cortexm0ds_logic.v(788)
  wire U91iu6;  // ../RTL/cortexm0ds_logic.v(320)
  wire U91pw6;  // ../RTL/cortexm0ds_logic.v(1345)
  wire U97ju6;  // ../RTL/cortexm0ds_logic.v(882)
  wire U98iu6;  // ../RTL/cortexm0ds_logic.v(414)
  wire U98pw6;  // ../RTL/cortexm0ds_logic.v(1438)
  wire U99ow6;  // ../RTL/cortexm0ds_logic.v(970)
  wire U9fiu6;  // ../RTL/cortexm0ds_logic.v(508)
  wire U9gow6;  // ../RTL/cortexm0ds_logic.v(1064)
  wire U9miu6;  // ../RTL/cortexm0ds_logic.v(601)
  wire U9now6;  // ../RTL/cortexm0ds_logic.v(1158)
  wire U9tiu6;  // ../RTL/cortexm0ds_logic.v(695)
  wire U9uhu6;  // ../RTL/cortexm0ds_logic.v(227)
  wire U9uow6;  // ../RTL/cortexm0ds_logic.v(1251)
  wire U9ypw6;  // ../RTL/cortexm0ds_logic.v(1614)
  wire Ua0iu6;  // ../RTL/cortexm0ds_logic.v(307)
  wire Ua0pw6;  // ../RTL/cortexm0ds_logic.v(1332)
  wire Ua6ju6;  // ../RTL/cortexm0ds_logic.v(869)
  wire Ua7iu6;  // ../RTL/cortexm0ds_logic.v(401)
  wire Ua7pw6;  // ../RTL/cortexm0ds_logic.v(1425)
  wire Ua8ow6;  // ../RTL/cortexm0ds_logic.v(957)
  wire Ua9bx6;  // ../RTL/cortexm0ds_logic.v(1696)
  wire Uaeiu6;  // ../RTL/cortexm0ds_logic.v(495)
  wire Uafow6;  // ../RTL/cortexm0ds_logic.v(1051)
  wire Ualiu6;  // ../RTL/cortexm0ds_logic.v(588)
  wire Uamow6;  // ../RTL/cortexm0ds_logic.v(1145)
  wire Uarax6;  // ../RTL/cortexm0ds_logic.v(1664)
  wire Uasiu6;  // ../RTL/cortexm0ds_logic.v(682)
  wire Uathu6;  // ../RTL/cortexm0ds_logic.v(214)
  wire Uatow6;  // ../RTL/cortexm0ds_logic.v(1238)
  wire Uaziu6;  // ../RTL/cortexm0ds_logic.v(775)
  wire Ub5ju6;  // ../RTL/cortexm0ds_logic.v(856)
  wire Ub6iu6;  // ../RTL/cortexm0ds_logic.v(388)
  wire Ub6pw6;  // ../RTL/cortexm0ds_logic.v(1412)
  wire Ub7ow6;  // ../RTL/cortexm0ds_logic.v(944)
  wire Ubdiu6;  // ../RTL/cortexm0ds_logic.v(482)
  wire Ubdpw6;  // ../RTL/cortexm0ds_logic.v(1506)
  wire Ubeow6;  // ../RTL/cortexm0ds_logic.v(1038)
  wire Ubkiu6;  // ../RTL/cortexm0ds_logic.v(575)
  wire Ublow6;  // ../RTL/cortexm0ds_logic.v(1132)
  wire Ubnhu6;  // ../RTL/cortexm0ds_logic.v(144)
  wire Ubriu6;  // ../RTL/cortexm0ds_logic.v(669)
  wire Ubshu6;  // ../RTL/cortexm0ds_logic.v(201)
  wire Ubsow6;  // ../RTL/cortexm0ds_logic.v(1225)
  wire Ubyiu6;  // ../RTL/cortexm0ds_logic.v(762)
  wire Ubypw6;  // ../RTL/cortexm0ds_logic.v(1614)
  wire Ubzhu6;  // ../RTL/cortexm0ds_logic.v(294)
  wire Ubzow6;  // ../RTL/cortexm0ds_logic.v(1319)
  wire Uc4ju6;  // ../RTL/cortexm0ds_logic.v(843)
  wire Uc5iu6;  // ../RTL/cortexm0ds_logic.v(375)
  wire Uc5pw6;  // ../RTL/cortexm0ds_logic.v(1399)
  wire Uc6ow6;  // ../RTL/cortexm0ds_logic.v(931)
  wire Ucciu6;  // ../RTL/cortexm0ds_logic.v(469)
  wire Uccpw6;  // ../RTL/cortexm0ds_logic.v(1493)
  wire Ucdow6;  // ../RTL/cortexm0ds_logic.v(1025)
  wire Ucjiu6;  // ../RTL/cortexm0ds_logic.v(562)
  wire Uckow6;  // ../RTL/cortexm0ds_logic.v(1119)
  wire Ucqiu6;  // ../RTL/cortexm0ds_logic.v(656)
  wire Ucrhu6;  // ../RTL/cortexm0ds_logic.v(188)
  wire Ucrow6;  // ../RTL/cortexm0ds_logic.v(1212)
  wire Ucxiu6;  // ../RTL/cortexm0ds_logic.v(749)
  wire Ucyhu6;  // ../RTL/cortexm0ds_logic.v(281)
  wire Ucyow6;  // ../RTL/cortexm0ds_logic.v(1306)
  wire Ud3ju6;  // ../RTL/cortexm0ds_logic.v(830)
  wire Ud4iu6;  // ../RTL/cortexm0ds_logic.v(362)
  wire Ud4pw6;  // ../RTL/cortexm0ds_logic.v(1386)
  wire Udaju6;  // ../RTL/cortexm0ds_logic.v(924)
  wire Udbiu6;  // ../RTL/cortexm0ds_logic.v(456)
  wire Udbpw6;  // ../RTL/cortexm0ds_logic.v(1480)
  wire Udcow6;  // ../RTL/cortexm0ds_logic.v(1012)
  wire Udiiu6;  // ../RTL/cortexm0ds_logic.v(549)
  wire Udjow6;  // ../RTL/cortexm0ds_logic.v(1106)
  wire Udpiu6;  // ../RTL/cortexm0ds_logic.v(643)
  wire Udqhu6;  // ../RTL/cortexm0ds_logic.v(175)
  wire Udqow6;  // ../RTL/cortexm0ds_logic.v(1199)
  wire Udwiu6;  // ../RTL/cortexm0ds_logic.v(736)
  wire Udxhu6;  // ../RTL/cortexm0ds_logic.v(268)
  wire Udxow6;  // ../RTL/cortexm0ds_logic.v(1293)
  wire Ue2ju6;  // ../RTL/cortexm0ds_logic.v(817)
  wire Ue3iu6;  // ../RTL/cortexm0ds_logic.v(349)
  wire Ue3pw6;  // ../RTL/cortexm0ds_logic.v(1373)
  wire Ue9ax6;  // ../RTL/cortexm0ds_logic.v(1630)
  wire Ue9ju6;  // ../RTL/cortexm0ds_logic.v(911)
  wire Ueaiu6;  // ../RTL/cortexm0ds_logic.v(443)
  wire Ueapw6;  // ../RTL/cortexm0ds_logic.v(1467)
  wire Uebow6;  // ../RTL/cortexm0ds_logic.v(999)
  wire Uehiu6;  // ../RTL/cortexm0ds_logic.v(536)
  wire Ueiow6;  // ../RTL/cortexm0ds_logic.v(1093)
  wire Ueoiu6;  // ../RTL/cortexm0ds_logic.v(630)
  wire Uephu6;  // ../RTL/cortexm0ds_logic.v(162)
  wire Uepow6;  // ../RTL/cortexm0ds_logic.v(1186)
  wire Ueviu6;  // ../RTL/cortexm0ds_logic.v(723)
  wire Uewhu6;  // ../RTL/cortexm0ds_logic.v(255)
  wire Uewow6;  // ../RTL/cortexm0ds_logic.v(1280)
  wire Uf1ju6;  // ../RTL/cortexm0ds_logic.v(804)
  wire Uf2iu6;  // ../RTL/cortexm0ds_logic.v(336)
  wire Uf2pw6;  // ../RTL/cortexm0ds_logic.v(1360)
  wire Uf8ju6;  // ../RTL/cortexm0ds_logic.v(898)
  wire Uf9iu6;  // ../RTL/cortexm0ds_logic.v(430)
  wire Uf9pw6;  // ../RTL/cortexm0ds_logic.v(1454)
  wire Ufaow6;  // ../RTL/cortexm0ds_logic.v(986)
  wire Ufbbx6;  // ../RTL/cortexm0ds_logic.v(1700)
  wire Ufebx6;  // ../RTL/cortexm0ds_logic.v(1705)
  wire Ufgiu6;  // ../RTL/cortexm0ds_logic.v(523)
  wire Ufhow6;  // ../RTL/cortexm0ds_logic.v(1080)
  wire Ufkhu6;  // ../RTL/cortexm0ds_logic.v(136)
  wire Ufmhu6;  // ../RTL/cortexm0ds_logic.v(142)
  wire Ufniu6;  // ../RTL/cortexm0ds_logic.v(617)
  wire Ufohu6;  // ../RTL/cortexm0ds_logic.v(149)
  wire Ufoow6;  // ../RTL/cortexm0ds_logic.v(1173)
  wire Ufopw6;  // ../RTL/cortexm0ds_logic.v(1596)
  wire Ufuiu6;  // ../RTL/cortexm0ds_logic.v(710)
  wire Ufvhu6;  // ../RTL/cortexm0ds_logic.v(242)
  wire Ufvow6;  // ../RTL/cortexm0ds_logic.v(1267)
  wire Ug0ju6;  // ../RTL/cortexm0ds_logic.v(791)
  wire Ug1iu6;  // ../RTL/cortexm0ds_logic.v(323)
  wire Ug1pw6;  // ../RTL/cortexm0ds_logic.v(1347)
  wire Ug7ju6;  // ../RTL/cortexm0ds_logic.v(885)
  wire Ug8iu6;  // ../RTL/cortexm0ds_logic.v(417)
  wire Ug8pw6;  // ../RTL/cortexm0ds_logic.v(1441)
  wire Ug9ow6;  // ../RTL/cortexm0ds_logic.v(973)
  wire Ugfiu6;  // ../RTL/cortexm0ds_logic.v(510)
  wire Uggow6;  // ../RTL/cortexm0ds_logic.v(1067)
  wire Ugmiu6;  // ../RTL/cortexm0ds_logic.v(604)
  wire Ugnow6;  // ../RTL/cortexm0ds_logic.v(1160)
  wire Ugtiu6;  // ../RTL/cortexm0ds_logic.v(697)
  wire Uguhu6;  // ../RTL/cortexm0ds_logic.v(229)
  wire Uguow6;  // ../RTL/cortexm0ds_logic.v(1254)
  wire Uh0iu6;  // ../RTL/cortexm0ds_logic.v(310)
  wire Uh0pw6;  // ../RTL/cortexm0ds_logic.v(1334)
  wire Uh2qw6;  // ../RTL/cortexm0ds_logic.v(1622)
  wire Uh6ju6;  // ../RTL/cortexm0ds_logic.v(872)
  wire Uh7iu6;  // ../RTL/cortexm0ds_logic.v(404)
  wire Uh7pw6;  // ../RTL/cortexm0ds_logic.v(1428)
  wire Uh8ow6;  // ../RTL/cortexm0ds_logic.v(960)
  wire Uhehu6;  // ../RTL/cortexm0ds_logic.v(122)
  wire Uheiu6;  // ../RTL/cortexm0ds_logic.v(497)
  wire Uhfow6;  // ../RTL/cortexm0ds_logic.v(1054)
  wire Uhjhu6;  // ../RTL/cortexm0ds_logic.v(134)
  wire Uhliu6;  // ../RTL/cortexm0ds_logic.v(591)
  wire Uhmow6;  // ../RTL/cortexm0ds_logic.v(1147)
  wire Uhsiu6;  // ../RTL/cortexm0ds_logic.v(684)
  wire Uhthu6;  // ../RTL/cortexm0ds_logic.v(216)
  wire Uhtow6;  // ../RTL/cortexm0ds_logic.v(1241)
  wire Uhvax6;  // ../RTL/cortexm0ds_logic.v(1671)
  wire Uhziu6;  // ../RTL/cortexm0ds_logic.v(778)
  wire Ui5ju6;  // ../RTL/cortexm0ds_logic.v(859)
  wire Ui6iu6;  // ../RTL/cortexm0ds_logic.v(391)
  wire Ui6pw6;  // ../RTL/cortexm0ds_logic.v(1415)
  wire Ui7ow6;  // ../RTL/cortexm0ds_logic.v(947)
  wire Uidiu6;  // ../RTL/cortexm0ds_logic.v(484)
  wire Uidpw6;  // ../RTL/cortexm0ds_logic.v(1509)
  wire Uieow6;  // ../RTL/cortexm0ds_logic.v(1041)
  wire Uikiu6;  // ../RTL/cortexm0ds_logic.v(578)
  wire Uilhu6;  // ../RTL/cortexm0ds_logic.v(139)
  wire Uilow6;  // ../RTL/cortexm0ds_logic.v(1134)
  wire Uiriu6;  // ../RTL/cortexm0ds_logic.v(671)
  wire Uishu6;  // ../RTL/cortexm0ds_logic.v(203)
  wire Uisow6;  // ../RTL/cortexm0ds_logic.v(1228)
  wire Uiyiu6;  // ../RTL/cortexm0ds_logic.v(765)
  wire Uizax6;  // ../RTL/cortexm0ds_logic.v(1678)
  wire Uizhu6;  // ../RTL/cortexm0ds_logic.v(297)
  wire Uizow6;  // ../RTL/cortexm0ds_logic.v(1321)
  wire Uj4bx6;  // ../RTL/cortexm0ds_logic.v(1687)
  wire Uj4ju6;  // ../RTL/cortexm0ds_logic.v(846)
  wire Uj5iu6;  // ../RTL/cortexm0ds_logic.v(378)
  wire Uj5pw6;  // ../RTL/cortexm0ds_logic.v(1402)
  wire Uj6ow6;  // ../RTL/cortexm0ds_logic.v(934)
  wire Ujciu6;  // ../RTL/cortexm0ds_logic.v(471)
  wire Ujcpw6;  // ../RTL/cortexm0ds_logic.v(1496)
  wire Ujdow6;  // ../RTL/cortexm0ds_logic.v(1028)
  wire Ujihu6;  // ../RTL/cortexm0ds_logic.v(131)
  wire Ujjiu6;  // ../RTL/cortexm0ds_logic.v(565)
  wire Ujkow6;  // ../RTL/cortexm0ds_logic.v(1121)
  wire Ujqiu6;  // ../RTL/cortexm0ds_logic.v(658)
  wire Ujrhu6;  // ../RTL/cortexm0ds_logic.v(190)
  wire Ujrow6;  // ../RTL/cortexm0ds_logic.v(1215)
  wire Ujspw6;  // ../RTL/cortexm0ds_logic.v(1603)
  wire Ujxax6;  // ../RTL/cortexm0ds_logic.v(1675)
  wire Ujxiu6;  // ../RTL/cortexm0ds_logic.v(752)
  wire Ujyhu6;  // ../RTL/cortexm0ds_logic.v(284)
  wire Ujyow6;  // ../RTL/cortexm0ds_logic.v(1308)
  wire Uk3ju6;  // ../RTL/cortexm0ds_logic.v(833)
  wire Uk4iu6;  // ../RTL/cortexm0ds_logic.v(365)
  wire Uk4pw6;  // ../RTL/cortexm0ds_logic.v(1389)
  wire Ukaju6;  // ../RTL/cortexm0ds_logic.v(926)
  wire Ukbiu6;  // ../RTL/cortexm0ds_logic.v(458)
  wire Ukbpw6;  // ../RTL/cortexm0ds_logic.v(1483)
  wire Ukcow6;  // ../RTL/cortexm0ds_logic.v(1015)
  wire Ukiiu6;  // ../RTL/cortexm0ds_logic.v(552)
  wire Ukjow6;  // ../RTL/cortexm0ds_logic.v(1108)
  wire Ukpiu6;  // ../RTL/cortexm0ds_logic.v(645)
  wire Ukqhu6;  // ../RTL/cortexm0ds_logic.v(177)
  wire Ukqow6;  // ../RTL/cortexm0ds_logic.v(1202)
  wire Ukwiu6;  // ../RTL/cortexm0ds_logic.v(739)
  wire Ukxhu6;  // ../RTL/cortexm0ds_logic.v(271)
  wire Ukxow6;  // ../RTL/cortexm0ds_logic.v(1295)
  wire Ul2ju6;  // ../RTL/cortexm0ds_logic.v(820)
  wire Ul3iu6;  // ../RTL/cortexm0ds_logic.v(352)
  wire Ul3pw6;  // ../RTL/cortexm0ds_logic.v(1376)
  wire Ul9ju6;  // ../RTL/cortexm0ds_logic.v(913)
  wire Ulaiu6;  // ../RTL/cortexm0ds_logic.v(445)
  wire Ulapw6;  // ../RTL/cortexm0ds_logic.v(1470)
  wire Ulbow6;  // ../RTL/cortexm0ds_logic.v(1002)
  wire Ulhiu6;  // ../RTL/cortexm0ds_logic.v(539)
  wire Uliow6;  // ../RTL/cortexm0ds_logic.v(1095)
  wire Ulnhu6;  // ../RTL/cortexm0ds_logic.v(145)
  wire Uloiu6;  // ../RTL/cortexm0ds_logic.v(632)
  wire Ulphu6;  // ../RTL/cortexm0ds_logic.v(164)
  wire Ulpow6;  // ../RTL/cortexm0ds_logic.v(1189)
  wire Ulviu6;  // ../RTL/cortexm0ds_logic.v(726)
  wire Ulwhu6;  // ../RTL/cortexm0ds_logic.v(258)
  wire Ulwow6;  // ../RTL/cortexm0ds_logic.v(1282)
  wire Um1bx6;  // ../RTL/cortexm0ds_logic.v(1682)
  wire Um1ju6;  // ../RTL/cortexm0ds_logic.v(807)
  wire Um2iu6;  // ../RTL/cortexm0ds_logic.v(339)
  wire Um2pw6;  // ../RTL/cortexm0ds_logic.v(1363)
  wire Um8ju6;  // ../RTL/cortexm0ds_logic.v(900)
  wire Um9iu6;  // ../RTL/cortexm0ds_logic.v(432)
  wire Um9pw6;  // ../RTL/cortexm0ds_logic.v(1457)
  wire Umaow6;  // ../RTL/cortexm0ds_logic.v(989)
  wire Umgiu6;  // ../RTL/cortexm0ds_logic.v(526)
  wire Umhow6;  // ../RTL/cortexm0ds_logic.v(1082)
  wire Umkax6;  // ../RTL/cortexm0ds_logic.v(1652)
  wire Umniu6;  // ../RTL/cortexm0ds_logic.v(619)
  wire Umohu6;  // ../RTL/cortexm0ds_logic.v(151)
  wire Umoow6;  // ../RTL/cortexm0ds_logic.v(1176)
  wire Umuiu6;  // ../RTL/cortexm0ds_logic.v(713)
  wire Umvhu6;  // ../RTL/cortexm0ds_logic.v(245)
  wire Umvow6;  // ../RTL/cortexm0ds_logic.v(1269)
  wire Un0ju6;  // ../RTL/cortexm0ds_logic.v(794)
  wire Un1iu6;  // ../RTL/cortexm0ds_logic.v(326)
  wire Un1pw6;  // ../RTL/cortexm0ds_logic.v(1350)
  wire Un7ju6;  // ../RTL/cortexm0ds_logic.v(887)
  wire Un8iu6;  // ../RTL/cortexm0ds_logic.v(419)
  wire Un8pw6;  // ../RTL/cortexm0ds_logic.v(1444)
  wire Un9ow6;  // ../RTL/cortexm0ds_logic.v(976)
  wire Unfiu6;  // ../RTL/cortexm0ds_logic.v(513)
  wire Ungow6;  // ../RTL/cortexm0ds_logic.v(1069)
  wire Unmiu6;  // ../RTL/cortexm0ds_logic.v(606)
  wire Unnow6;  // ../RTL/cortexm0ds_logic.v(1163)
  wire Untiu6;  // ../RTL/cortexm0ds_logic.v(700)
  wire Untpw6;  // ../RTL/cortexm0ds_logic.v(1605)
  wire Unuhu6;  // ../RTL/cortexm0ds_logic.v(232)
  wire Unuow6;  // ../RTL/cortexm0ds_logic.v(1256)
  wire Unyax6;  // ../RTL/cortexm0ds_logic.v(1677)
  wire Uo0iu6;  // ../RTL/cortexm0ds_logic.v(313)
  wire Uo0pw6;  // ../RTL/cortexm0ds_logic.v(1337)
  wire Uo2bx6;  // ../RTL/cortexm0ds_logic.v(1684)
  wire Uo6ju6;  // ../RTL/cortexm0ds_logic.v(874)
  wire Uo7iu6;  // ../RTL/cortexm0ds_logic.v(406)
  wire Uo7pw6;  // ../RTL/cortexm0ds_logic.v(1431)
  wire Uo8ow6;  // ../RTL/cortexm0ds_logic.v(963)
  wire Uoeiu6;  // ../RTL/cortexm0ds_logic.v(500)
  wire Uofax6;  // ../RTL/cortexm0ds_logic.v(1642)
  wire Uofow6;  // ../RTL/cortexm0ds_logic.v(1056)
  wire Uoipw6;  // ../RTL/cortexm0ds_logic.v(1585)
  wire Uojbx6;  // ../RTL/cortexm0ds_logic.v(1715)
  wire Uoliu6;  // ../RTL/cortexm0ds_logic.v(593)
  wire Uomow6;  // ../RTL/cortexm0ds_logic.v(1150)
  wire Uoqax6;  // ../RTL/cortexm0ds_logic.v(1663)
  wire Uosiu6;  // ../RTL/cortexm0ds_logic.v(687)
  wire Uothu6;  // ../RTL/cortexm0ds_logic.v(219)
  wire Uotow6;  // ../RTL/cortexm0ds_logic.v(1243)
  wire Uoziu6;  // ../RTL/cortexm0ds_logic.v(781)
  wire Up4bx6;  // ../RTL/cortexm0ds_logic.v(1687)
  wire Up5ju6;  // ../RTL/cortexm0ds_logic.v(861)
  wire Up6iu6;  // ../RTL/cortexm0ds_logic.v(393)
  wire Up6pw6;  // ../RTL/cortexm0ds_logic.v(1418)
  wire Up7ow6;  // ../RTL/cortexm0ds_logic.v(950)
  wire Updiu6;  // ../RTL/cortexm0ds_logic.v(487)
  wire Updpw6;  // ../RTL/cortexm0ds_logic.v(1511)
  wire Upeow6;  // ../RTL/cortexm0ds_logic.v(1043)
  wire Upkiu6;  // ../RTL/cortexm0ds_logic.v(580)
  wire Uplow6;  // ../RTL/cortexm0ds_logic.v(1137)
  wire Upriu6;  // ../RTL/cortexm0ds_logic.v(674)
  wire Upshu6;  // ../RTL/cortexm0ds_logic.v(206)
  wire Upsow6;  // ../RTL/cortexm0ds_logic.v(1230)
  wire Upyiu6;  // ../RTL/cortexm0ds_logic.v(768)
  wire Upzhu6;  // ../RTL/cortexm0ds_logic.v(300)
  wire Upzow6;  // ../RTL/cortexm0ds_logic.v(1324)
  wire Uq4ju6;  // ../RTL/cortexm0ds_logic.v(848)
  wire Uq5iu6;  // ../RTL/cortexm0ds_logic.v(380)
  wire Uq5pw6;  // ../RTL/cortexm0ds_logic.v(1405)
  wire Uq6ow6;  // ../RTL/cortexm0ds_logic.v(937)
  wire Uqciu6;  // ../RTL/cortexm0ds_logic.v(474)
  wire Uqcpw6;  // ../RTL/cortexm0ds_logic.v(1498)
  wire Uqdow6;  // ../RTL/cortexm0ds_logic.v(1030)
  wire Uqipw6;  // ../RTL/cortexm0ds_logic.v(1585)
  wire Uqjiu6;  // ../RTL/cortexm0ds_logic.v(567)
  wire Uqkow6;  // ../RTL/cortexm0ds_logic.v(1124)
  wire Uqqax6;  // ../RTL/cortexm0ds_logic.v(1663)
  wire Uqqiu6;  // ../RTL/cortexm0ds_logic.v(661)
  wire Uqrhu6;  // ../RTL/cortexm0ds_logic.v(193)
  wire Uqrow6;  // ../RTL/cortexm0ds_logic.v(1217)
  wire Uqxiu6;  // ../RTL/cortexm0ds_logic.v(755)
  wire Uqyhu6;  // ../RTL/cortexm0ds_logic.v(287)
  wire Uqyow6;  // ../RTL/cortexm0ds_logic.v(1311)
  wire Ur3ju6;  // ../RTL/cortexm0ds_logic.v(835)
  wire Ur4iu6;  // ../RTL/cortexm0ds_logic.v(367)
  wire Ur4pw6;  // ../RTL/cortexm0ds_logic.v(1392)
  wire Uraju6;  // ../RTL/cortexm0ds_logic.v(929)
  wire Urbiu6;  // ../RTL/cortexm0ds_logic.v(461)
  wire Urbpw6;  // ../RTL/cortexm0ds_logic.v(1485)
  wire Urcow6;  // ../RTL/cortexm0ds_logic.v(1017)
  wire Ureax6;  // ../RTL/cortexm0ds_logic.v(1640)
  wire Urgbx6;  // ../RTL/cortexm0ds_logic.v(1710)
  wire Uriiu6;  // ../RTL/cortexm0ds_logic.v(554)
  wire Urjow6;  // ../RTL/cortexm0ds_logic.v(1111)
  wire Urpiu6;  // ../RTL/cortexm0ds_logic.v(648)
  wire Urqhu6;  // ../RTL/cortexm0ds_logic.v(180)
  wire Urqow6;  // ../RTL/cortexm0ds_logic.v(1204)
  wire Urwiu6;  // ../RTL/cortexm0ds_logic.v(742)
  wire Urxhu6;  // ../RTL/cortexm0ds_logic.v(274)
  wire Urxow6;  // ../RTL/cortexm0ds_logic.v(1298)
  wire Us2ju6;  // ../RTL/cortexm0ds_logic.v(822)
  wire Us3bx6;  // ../RTL/cortexm0ds_logic.v(1686)
  wire Us3iu6;  // ../RTL/cortexm0ds_logic.v(354)
  wire Us3pw6;  // ../RTL/cortexm0ds_logic.v(1379)
  wire Us9ju6;  // ../RTL/cortexm0ds_logic.v(916)
  wire Usaiu6;  // ../RTL/cortexm0ds_logic.v(448)
  wire Usapw6;  // ../RTL/cortexm0ds_logic.v(1472)
  wire Usbow6;  // ../RTL/cortexm0ds_logic.v(1004)
  wire Uscax6;  // ../RTL/cortexm0ds_logic.v(1637)
  wire Ushiu6;  // ../RTL/cortexm0ds_logic.v(541)
  wire Usiow6;  // ../RTL/cortexm0ds_logic.v(1098)
  wire Usipw6;  // ../RTL/cortexm0ds_logic.v(1585)
  wire Usjbx6;  // ../RTL/cortexm0ds_logic.v(1715)
  wire Usnpw6;  // ../RTL/cortexm0ds_logic.v(1595)
  wire Usoiu6;  // ../RTL/cortexm0ds_logic.v(635)
  wire Usphu6;  // ../RTL/cortexm0ds_logic.v(167)
  wire Uspow6;  // ../RTL/cortexm0ds_logic.v(1191)
  wire Usqax6;  // ../RTL/cortexm0ds_logic.v(1663)
  wire Usviu6;  // ../RTL/cortexm0ds_logic.v(729)
  wire Uswhu6;  // ../RTL/cortexm0ds_logic.v(261)
  wire Uswow6;  // ../RTL/cortexm0ds_logic.v(1285)
  wire Ut1ju6;  // ../RTL/cortexm0ds_logic.v(809)
  wire Ut2iu6;  // ../RTL/cortexm0ds_logic.v(341)
  wire Ut2pw6;  // ../RTL/cortexm0ds_logic.v(1366)
  wire Ut8ju6;  // ../RTL/cortexm0ds_logic.v(903)
  wire Ut9iu6;  // ../RTL/cortexm0ds_logic.v(435)
  wire Ut9pw6;  // ../RTL/cortexm0ds_logic.v(1459)
  wire Utaow6;  // ../RTL/cortexm0ds_logic.v(991)
  wire Utgiu6;  // ../RTL/cortexm0ds_logic.v(528)
  wire Uthow6;  // ../RTL/cortexm0ds_logic.v(1085)
  wire Utniu6;  // ../RTL/cortexm0ds_logic.v(622)
  wire Utohu6;  // ../RTL/cortexm0ds_logic.v(154)
  wire Utoow6;  // ../RTL/cortexm0ds_logic.v(1178)
  wire Utqpw6;  // ../RTL/cortexm0ds_logic.v(1600)
  wire Utuiu6;  // ../RTL/cortexm0ds_logic.v(716)
  wire Utvhu6;  // ../RTL/cortexm0ds_logic.v(248)
  wire Utvow6;  // ../RTL/cortexm0ds_logic.v(1272)
  wire Uu0ju6;  // ../RTL/cortexm0ds_logic.v(796)
  wire Uu1iu6;  // ../RTL/cortexm0ds_logic.v(328)
  wire Uu1pw6;  // ../RTL/cortexm0ds_logic.v(1353)
  wire Uu7ju6;  // ../RTL/cortexm0ds_logic.v(890)
  wire Uu8iu6;  // ../RTL/cortexm0ds_logic.v(422)
  wire Uu8pw6;  // ../RTL/cortexm0ds_logic.v(1446)
  wire Uu9ow6;  // ../RTL/cortexm0ds_logic.v(978)
  wire Uufiu6;  // ../RTL/cortexm0ds_logic.v(515)
  wire Uugow6;  // ../RTL/cortexm0ds_logic.v(1072)
  wire Uumiu6;  // ../RTL/cortexm0ds_logic.v(609)
  wire Uunow6;  // ../RTL/cortexm0ds_logic.v(1165)
  wire Uunpw6;  // ../RTL/cortexm0ds_logic.v(1595)
  wire Uuqax6;  // ../RTL/cortexm0ds_logic.v(1663)
  wire Uutiu6;  // ../RTL/cortexm0ds_logic.v(703)
  wire Uuuhu6;  // ../RTL/cortexm0ds_logic.v(235)
  wire Uuuow6;  // ../RTL/cortexm0ds_logic.v(1259)
  wire Uuzpw6;  // ../RTL/cortexm0ds_logic.v(1617)
  wire Uv0iu6;  // ../RTL/cortexm0ds_logic.v(315)
  wire Uv0pw6;  // ../RTL/cortexm0ds_logic.v(1340)
  wire Uv6ju6;  // ../RTL/cortexm0ds_logic.v(877)
  wire Uv7iu6;  // ../RTL/cortexm0ds_logic.v(409)
  wire Uv7pw6;  // ../RTL/cortexm0ds_logic.v(1433)
  wire Uv8ow6;  // ../RTL/cortexm0ds_logic.v(965)
  wire Uveiu6;  // ../RTL/cortexm0ds_logic.v(502)
  wire Uvfow6;  // ../RTL/cortexm0ds_logic.v(1059)
  wire Uvliu6;  // ../RTL/cortexm0ds_logic.v(596)
  wire Uvmax6;  // ../RTL/cortexm0ds_logic.v(1656)
  wire Uvmow6;  // ../RTL/cortexm0ds_logic.v(1152)
  wire Uvsiu6;  // ../RTL/cortexm0ds_logic.v(690)
  wire Uvthu6;  // ../RTL/cortexm0ds_logic.v(222)
  wire Uvtow6;  // ../RTL/cortexm0ds_logic.v(1246)
  wire Uvziu6;  // ../RTL/cortexm0ds_logic.v(783)
  wire Uw5ju6;  // ../RTL/cortexm0ds_logic.v(864)
  wire Uw6iu6;  // ../RTL/cortexm0ds_logic.v(396)
  wire Uw6pw6;  // ../RTL/cortexm0ds_logic.v(1420)
  wire Uw7ow6;  // ../RTL/cortexm0ds_logic.v(952)
  wire Uwdiu6;  // ../RTL/cortexm0ds_logic.v(489)
  wire Uwdpw6;  // ../RTL/cortexm0ds_logic.v(1514)
  wire Uweow6;  // ../RTL/cortexm0ds_logic.v(1046)
  wire Uwipw6;  // ../RTL/cortexm0ds_logic.v(1586)
  wire Uwkhu6;  // ../RTL/cortexm0ds_logic.v(138)
  wire Uwkiu6;  // ../RTL/cortexm0ds_logic.v(583)
  wire Uwlow6;  // ../RTL/cortexm0ds_logic.v(1139)
  wire Uwqax6;  // ../RTL/cortexm0ds_logic.v(1663)
  wire Uwriu6;  // ../RTL/cortexm0ds_logic.v(677)
  wire Uwshu6;  // ../RTL/cortexm0ds_logic.v(209)
  wire Uwsow6;  // ../RTL/cortexm0ds_logic.v(1233)
  wire Uwyiu6;  // ../RTL/cortexm0ds_logic.v(770)
  wire Uwzhu6;  // ../RTL/cortexm0ds_logic.v(302)
  wire Uwzow6;  // ../RTL/cortexm0ds_logic.v(1327)
  wire Ux4ju6;  // ../RTL/cortexm0ds_logic.v(851)
  wire Ux5iu6;  // ../RTL/cortexm0ds_logic.v(383)
  wire Ux5pw6;  // ../RTL/cortexm0ds_logic.v(1407)
  wire Ux6ow6;  // ../RTL/cortexm0ds_logic.v(939)
  wire Ux8bx6;  // ../RTL/cortexm0ds_logic.v(1695)
  wire Uxciu6;  // ../RTL/cortexm0ds_logic.v(476)
  wire Uxcpw6;  // ../RTL/cortexm0ds_logic.v(1501)
  wire Uxdow6;  // ../RTL/cortexm0ds_logic.v(1033)
  wire Uxjiu6;  // ../RTL/cortexm0ds_logic.v(570)
  wire Uxkow6;  // ../RTL/cortexm0ds_logic.v(1126)
  wire Uxqiu6;  // ../RTL/cortexm0ds_logic.v(664)
  wire Uxrhu6;  // ../RTL/cortexm0ds_logic.v(196)
  wire Uxrow6;  // ../RTL/cortexm0ds_logic.v(1220)
  wire Uxxiu6;  // ../RTL/cortexm0ds_logic.v(757)
  wire Uxyhu6;  // ../RTL/cortexm0ds_logic.v(289)
  wire Uxyow6;  // ../RTL/cortexm0ds_logic.v(1314)
  wire Uy3ju6;  // ../RTL/cortexm0ds_logic.v(838)
  wire Uy4iu6;  // ../RTL/cortexm0ds_logic.v(370)
  wire Uy4pw6;  // ../RTL/cortexm0ds_logic.v(1394)
  wire Uybiu6;  // ../RTL/cortexm0ds_logic.v(463)
  wire Uybpw6;  // ../RTL/cortexm0ds_logic.v(1488)
  wire Uycow6;  // ../RTL/cortexm0ds_logic.v(1020)
  wire Uyiiu6;  // ../RTL/cortexm0ds_logic.v(557)
  wire Uyjhu6;  // ../RTL/cortexm0ds_logic.v(135)
  wire Uyjow6;  // ../RTL/cortexm0ds_logic.v(1113)
  wire Uypiu6;  // ../RTL/cortexm0ds_logic.v(651)
  wire Uyqax6;  // ../RTL/cortexm0ds_logic.v(1663)
  wire Uyqhu6;  // ../RTL/cortexm0ds_logic.v(183)
  wire Uyqow6;  // ../RTL/cortexm0ds_logic.v(1207)
  wire Uywiu6;  // ../RTL/cortexm0ds_logic.v(744)
  wire Uyxhu6;  // ../RTL/cortexm0ds_logic.v(276)
  wire Uyxow6;  // ../RTL/cortexm0ds_logic.v(1301)
  wire Uz2ju6;  // ../RTL/cortexm0ds_logic.v(825)
  wire Uz3iu6;  // ../RTL/cortexm0ds_logic.v(357)
  wire Uz3pw6;  // ../RTL/cortexm0ds_logic.v(1381)
  wire Uz9ju6;  // ../RTL/cortexm0ds_logic.v(918)
  wire Uzaiu6;  // ../RTL/cortexm0ds_logic.v(450)
  wire Uzapw6;  // ../RTL/cortexm0ds_logic.v(1475)
  wire Uzbow6;  // ../RTL/cortexm0ds_logic.v(1007)
  wire Uzhiu6;  // ../RTL/cortexm0ds_logic.v(544)
  wire Uziow6;  // ../RTL/cortexm0ds_logic.v(1100)
  wire Uzoiu6;  // ../RTL/cortexm0ds_logic.v(638)
  wire Uzphu6;  // ../RTL/cortexm0ds_logic.v(170)
  wire Uzpow6;  // ../RTL/cortexm0ds_logic.v(1194)
  wire Uzviu6;  // ../RTL/cortexm0ds_logic.v(731)
  wire Uzwhu6;  // ../RTL/cortexm0ds_logic.v(263)
  wire Uzwow6;  // ../RTL/cortexm0ds_logic.v(1288)
  wire V00iu6;  // ../RTL/cortexm0ds_logic.v(304)
  wire V00pw6;  // ../RTL/cortexm0ds_logic.v(1328)
  wire V06ju6;  // ../RTL/cortexm0ds_logic.v(865)
  wire V07iu6;  // ../RTL/cortexm0ds_logic.v(397)
  wire V07pw6;  // ../RTL/cortexm0ds_logic.v(1422)
  wire V08ow6;  // ../RTL/cortexm0ds_logic.v(954)
  wire V0cax6;  // ../RTL/cortexm0ds_logic.v(1635)
  wire V0eiu6;  // ../RTL/cortexm0ds_logic.v(491)
  wire V0epw6;  // ../RTL/cortexm0ds_logic.v(1515)
  wire V0fow6;  // ../RTL/cortexm0ds_logic.v(1047)
  wire V0jpw6;  // ../RTL/cortexm0ds_logic.v(1586)
  wire V0liu6;  // ../RTL/cortexm0ds_logic.v(584)
  wire V0mow6;  // ../RTL/cortexm0ds_logic.v(1141)
  wire V0siu6;  // ../RTL/cortexm0ds_logic.v(678)
  wire V0thu6;  // ../RTL/cortexm0ds_logic.v(210)
  wire V0tow6;  // ../RTL/cortexm0ds_logic.v(1234)
  wire V0ziu6;  // ../RTL/cortexm0ds_logic.v(772)
  wire V15ju6;  // ../RTL/cortexm0ds_logic.v(852)
  wire V16iu6;  // ../RTL/cortexm0ds_logic.v(384)
  wire V16pw6;  // ../RTL/cortexm0ds_logic.v(1409)
  wire V17ow6;  // ../RTL/cortexm0ds_logic.v(941)
  wire V1diu6;  // ../RTL/cortexm0ds_logic.v(478)
  wire V1dpw6;  // ../RTL/cortexm0ds_logic.v(1502)
  wire V1eow6;  // ../RTL/cortexm0ds_logic.v(1034)
  wire V1kiu6;  // ../RTL/cortexm0ds_logic.v(571)
  wire V1low6;  // ../RTL/cortexm0ds_logic.v(1128)
  wire V1mhu6;  // ../RTL/cortexm0ds_logic.v(141)
  wire V1riu6;  // ../RTL/cortexm0ds_logic.v(665)
  wire V1shu6;  // ../RTL/cortexm0ds_logic.v(197)
  wire V1sow6;  // ../RTL/cortexm0ds_logic.v(1221)
  wire V1vax6;  // ../RTL/cortexm0ds_logic.v(1670)
  wire V1yax6;  // ../RTL/cortexm0ds_logic.v(1676)
  wire V1yiu6;  // ../RTL/cortexm0ds_logic.v(759)
  wire V1zhu6;  // ../RTL/cortexm0ds_logic.v(291)
  wire V1zow6;  // ../RTL/cortexm0ds_logic.v(1315)
  wire V24ju6;  // ../RTL/cortexm0ds_logic.v(839)
  wire V25iu6;  // ../RTL/cortexm0ds_logic.v(371)
  wire V25pw6;  // ../RTL/cortexm0ds_logic.v(1396)
  wire V2ciu6;  // ../RTL/cortexm0ds_logic.v(465)
  wire V2cpw6;  // ../RTL/cortexm0ds_logic.v(1489)
  wire V2dow6;  // ../RTL/cortexm0ds_logic.v(1021)
  wire V2jiu6;  // ../RTL/cortexm0ds_logic.v(558)
  wire V2kow6;  // ../RTL/cortexm0ds_logic.v(1115)
  wire V2qiu6;  // ../RTL/cortexm0ds_logic.v(652)
  wire V2rhu6;  // ../RTL/cortexm0ds_logic.v(184)
  wire V2row6;  // ../RTL/cortexm0ds_logic.v(1208)
  wire V2xiu6;  // ../RTL/cortexm0ds_logic.v(746)
  wire V2yhu6;  // ../RTL/cortexm0ds_logic.v(278)
  wire V2yow6;  // ../RTL/cortexm0ds_logic.v(1302)
  wire V33ju6;  // ../RTL/cortexm0ds_logic.v(826)
  wire V34iu6;  // ../RTL/cortexm0ds_logic.v(358)
  wire V34pw6;  // ../RTL/cortexm0ds_logic.v(1383)
  wire V3aju6;  // ../RTL/cortexm0ds_logic.v(920)
  wire V3biu6;  // ../RTL/cortexm0ds_logic.v(452)
  wire V3bpw6;  // ../RTL/cortexm0ds_logic.v(1476)
  wire V3cow6;  // ../RTL/cortexm0ds_logic.v(1008)
  wire V3iiu6;  // ../RTL/cortexm0ds_logic.v(545)
  wire V3jow6;  // ../RTL/cortexm0ds_logic.v(1102)
  wire V3piu6;  // ../RTL/cortexm0ds_logic.v(639)
  wire V3qhu6;  // ../RTL/cortexm0ds_logic.v(171)
  wire V3qow6;  // ../RTL/cortexm0ds_logic.v(1195)
  wire V3vax6;  // ../RTL/cortexm0ds_logic.v(1671)
  wire V3wiu6;  // ../RTL/cortexm0ds_logic.v(733)
  wire V3xhu6;  // ../RTL/cortexm0ds_logic.v(265)
  wire V3xow6;  // ../RTL/cortexm0ds_logic.v(1289)
  wire V42ju6;  // ../RTL/cortexm0ds_logic.v(813)
  wire V43pw6;  // ../RTL/cortexm0ds_logic.v(1370)
  wire V49ju6;  // ../RTL/cortexm0ds_logic.v(907)
  wire V4aiu6;  // ../RTL/cortexm0ds_logic.v(439)
  wire V4apw6;  // ../RTL/cortexm0ds_logic.v(1463)
  wire V4bow6;  // ../RTL/cortexm0ds_logic.v(995)
  wire V4hiu6;  // ../RTL/cortexm0ds_logic.v(532)
  wire V4iow6;  // ../RTL/cortexm0ds_logic.v(1089)
  wire V4oiu6;  // ../RTL/cortexm0ds_logic.v(626)
  wire V4phu6;  // ../RTL/cortexm0ds_logic.v(158)
  wire V4pow6;  // ../RTL/cortexm0ds_logic.v(1182)
  wire V4viu6;  // ../RTL/cortexm0ds_logic.v(720)
  wire V4whu6;  // ../RTL/cortexm0ds_logic.v(252)
  wire V4wow6;  // ../RTL/cortexm0ds_logic.v(1276)
  wire V51ju6;  // ../RTL/cortexm0ds_logic.v(800)
  wire V52bx6;  // ../RTL/cortexm0ds_logic.v(1683)
  wire V52iu6;  // ../RTL/cortexm0ds_logic.v(332)
  wire V52pw6;  // ../RTL/cortexm0ds_logic.v(1357)
  wire V53qw6;  // ../RTL/cortexm0ds_logic.v(1623)
  wire V58ju6;  // ../RTL/cortexm0ds_logic.v(894)
  wire V59iu6;  // ../RTL/cortexm0ds_logic.v(426)
  wire V59pw6;  // ../RTL/cortexm0ds_logic.v(1450)
  wire V5abx6;  // ../RTL/cortexm0ds_logic.v(1697)
  wire V5aow6;  // ../RTL/cortexm0ds_logic.v(982)
  wire V5giu6;  // ../RTL/cortexm0ds_logic.v(519)
  wire V5how6;  // ../RTL/cortexm0ds_logic.v(1076)
  wire V5niu6;  // ../RTL/cortexm0ds_logic.v(613)
  wire V5oow6;  // ../RTL/cortexm0ds_logic.v(1169)
  wire V5uiu6;  // ../RTL/cortexm0ds_logic.v(707)
  wire V5vax6;  // ../RTL/cortexm0ds_logic.v(1671)
  wire V5vhu6;  // ../RTL/cortexm0ds_logic.v(239)
  wire V5vow6;  // ../RTL/cortexm0ds_logic.v(1263)
  wire V60ju6;  // ../RTL/cortexm0ds_logic.v(787)
  wire V61iu6;  // ../RTL/cortexm0ds_logic.v(319)
  wire V61pw6;  // ../RTL/cortexm0ds_logic.v(1344)
  wire V67ju6;  // ../RTL/cortexm0ds_logic.v(881)
  wire V68iu6;  // ../RTL/cortexm0ds_logic.v(413)
  wire V68pw6;  // ../RTL/cortexm0ds_logic.v(1437)
  wire V69ow6;  // ../RTL/cortexm0ds_logic.v(969)
  wire V6fiu6;  // ../RTL/cortexm0ds_logic.v(506)
  wire V6gow6;  // ../RTL/cortexm0ds_logic.v(1063)
  wire V6jax6;  // ../RTL/cortexm0ds_logic.v(1649)
  wire V6miu6;  // ../RTL/cortexm0ds_logic.v(600)
  wire V6now6;  // ../RTL/cortexm0ds_logic.v(1156)
  wire V6tiu6;  // ../RTL/cortexm0ds_logic.v(694)
  wire V6uhu6;  // ../RTL/cortexm0ds_logic.v(226)
  wire V6uow6;  // ../RTL/cortexm0ds_logic.v(1250)
  wire V70iu6;  // ../RTL/cortexm0ds_logic.v(306)
  wire V70pw6;  // ../RTL/cortexm0ds_logic.v(1331)
  wire V73bx6;  // ../RTL/cortexm0ds_logic.v(1685)
  wire V76ju6;  // ../RTL/cortexm0ds_logic.v(868)
  wire V77iu6;  // ../RTL/cortexm0ds_logic.v(400)
  wire V77pw6;  // ../RTL/cortexm0ds_logic.v(1424)
  wire V78ow6;  // ../RTL/cortexm0ds_logic.v(956)
  wire V7eiu6;  // ../RTL/cortexm0ds_logic.v(493)
  wire V7fow6;  // ../RTL/cortexm0ds_logic.v(1050)
  wire V7liu6;  // ../RTL/cortexm0ds_logic.v(587)
  wire V7mow6;  // ../RTL/cortexm0ds_logic.v(1143)
  wire V7siu6;  // ../RTL/cortexm0ds_logic.v(681)
  wire V7thu6;  // ../RTL/cortexm0ds_logic.v(213)
  wire V7tow6;  // ../RTL/cortexm0ds_logic.v(1237)
  wire V7vax6;  // ../RTL/cortexm0ds_logic.v(1671)
  wire V7ziu6;  // ../RTL/cortexm0ds_logic.v(774)
  wire V85ju6;  // ../RTL/cortexm0ds_logic.v(855)
  wire V86iu6;  // ../RTL/cortexm0ds_logic.v(387)
  wire V86pw6;  // ../RTL/cortexm0ds_logic.v(1411)
  wire V87ow6;  // ../RTL/cortexm0ds_logic.v(943)
  wire V8diu6;  // ../RTL/cortexm0ds_logic.v(480)
  wire V8dpw6;  // ../RTL/cortexm0ds_logic.v(1505)
  wire V8eow6;  // ../RTL/cortexm0ds_logic.v(1037)
  wire V8kiu6;  // ../RTL/cortexm0ds_logic.v(574)
  wire V8low6;  // ../RTL/cortexm0ds_logic.v(1130)
  wire V8riu6;  // ../RTL/cortexm0ds_logic.v(668)
  wire V8shu6;  // ../RTL/cortexm0ds_logic.v(200)
  wire V8sow6;  // ../RTL/cortexm0ds_logic.v(1224)
  wire V8yiu6;  // ../RTL/cortexm0ds_logic.v(761)
  wire V8zhu6;  // ../RTL/cortexm0ds_logic.v(293)
  wire V8zow6;  // ../RTL/cortexm0ds_logic.v(1318)
  wire V94ju6;  // ../RTL/cortexm0ds_logic.v(842)
  wire V95iu6;  // ../RTL/cortexm0ds_logic.v(374)
  wire V95pw6;  // ../RTL/cortexm0ds_logic.v(1398)
  wire V96ow6;  // ../RTL/cortexm0ds_logic.v(930)
  wire V9ciu6;  // ../RTL/cortexm0ds_logic.v(467)
  wire V9cpw6;  // ../RTL/cortexm0ds_logic.v(1492)
  wire V9dow6;  // ../RTL/cortexm0ds_logic.v(1024)
  wire V9ghu6;  // ../RTL/cortexm0ds_logic.v(126)
  wire V9jiu6;  // ../RTL/cortexm0ds_logic.v(561)
  wire V9kow6;  // ../RTL/cortexm0ds_logic.v(1117)
  wire V9qiu6;  // ../RTL/cortexm0ds_logic.v(655)
  wire V9rhu6;  // ../RTL/cortexm0ds_logic.v(187)
  wire V9row6;  // ../RTL/cortexm0ds_logic.v(1211)
  wire V9vax6;  // ../RTL/cortexm0ds_logic.v(1671)
  wire V9xiu6;  // ../RTL/cortexm0ds_logic.v(748)
  wire V9yhu6;  // ../RTL/cortexm0ds_logic.v(280)
  wire V9yow6;  // ../RTL/cortexm0ds_logic.v(1305)
  wire Va3ju6;  // ../RTL/cortexm0ds_logic.v(829)
  wire Va4iu6;  // ../RTL/cortexm0ds_logic.v(361)
  wire Va4pw6;  // ../RTL/cortexm0ds_logic.v(1385)
  wire Va7ax6;  // ../RTL/cortexm0ds_logic.v(1626)
  wire Vaaju6;  // ../RTL/cortexm0ds_logic.v(922)
  wire Vabiu6;  // ../RTL/cortexm0ds_logic.v(454)
  wire Vabpw6;  // ../RTL/cortexm0ds_logic.v(1479)
  wire Vacow6;  // ../RTL/cortexm0ds_logic.v(1011)
  wire Vaiiu6;  // ../RTL/cortexm0ds_logic.v(548)
  wire Vajow6;  // ../RTL/cortexm0ds_logic.v(1104)
  wire Vapiu6;  // ../RTL/cortexm0ds_logic.v(642)
  wire Vaqhu6;  // ../RTL/cortexm0ds_logic.v(174)
  wire Vaqow6;  // ../RTL/cortexm0ds_logic.v(1198)
  wire Vawiu6;  // ../RTL/cortexm0ds_logic.v(735)
  wire Vaxhu6;  // ../RTL/cortexm0ds_logic.v(267)
  wire Vaxow6;  // ../RTL/cortexm0ds_logic.v(1292)
  wire Vb2ju6;  // ../RTL/cortexm0ds_logic.v(816)
  wire Vb3iu6;  // ../RTL/cortexm0ds_logic.v(348)
  wire Vb3pw6;  // ../RTL/cortexm0ds_logic.v(1372)
  wire Vb9ju6;  // ../RTL/cortexm0ds_logic.v(909)
  wire Vbaiu6;  // ../RTL/cortexm0ds_logic.v(441)
  wire Vbapw6;  // ../RTL/cortexm0ds_logic.v(1466)
  wire Vbbow6;  // ../RTL/cortexm0ds_logic.v(998)
  wire Vbhiu6;  // ../RTL/cortexm0ds_logic.v(535)
  wire Vbiow6;  // ../RTL/cortexm0ds_logic.v(1091)
  wire Vbkpw6;  // ../RTL/cortexm0ds_logic.v(1588)
  wire Vboiu6;  // ../RTL/cortexm0ds_logic.v(629)
  wire Vbphu6;  // ../RTL/cortexm0ds_logic.v(161)
  wire Vbpow6;  // ../RTL/cortexm0ds_logic.v(1185)
  wire Vbspw6;  // ../RTL/cortexm0ds_logic.v(1603)
  wire Vbvax6;  // ../RTL/cortexm0ds_logic.v(1671)
  wire Vbviu6;  // ../RTL/cortexm0ds_logic.v(722)
  wire Vbwhu6;  // ../RTL/cortexm0ds_logic.v(254)
  wire Vbwow6;  // ../RTL/cortexm0ds_logic.v(1279)
  wire Vc1ju6;  // ../RTL/cortexm0ds_logic.v(803)
  wire Vc2iu6;  // ../RTL/cortexm0ds_logic.v(335)
  wire Vc2pw6;  // ../RTL/cortexm0ds_logic.v(1359)
  wire Vc8ju6;  // ../RTL/cortexm0ds_logic.v(896)
  wire Vc9iu6;  // ../RTL/cortexm0ds_logic.v(428)
  wire Vc9pw6;  // ../RTL/cortexm0ds_logic.v(1453)
  wire Vcaow6;  // ../RTL/cortexm0ds_logic.v(985)
  wire Vcgiu6;  // ../RTL/cortexm0ds_logic.v(522)
  wire Vchhu6;  // ../RTL/cortexm0ds_logic.v(128)
  wire Vchow6;  // ../RTL/cortexm0ds_logic.v(1078)
  wire Vcniu6;  // ../RTL/cortexm0ds_logic.v(616)
  wire Vcohu6;  // ../RTL/cortexm0ds_logic.v(148)
  wire Vcoow6;  // ../RTL/cortexm0ds_logic.v(1172)
  wire Vcuiu6;  // ../RTL/cortexm0ds_logic.v(709)
  wire Vcvhu6;  // ../RTL/cortexm0ds_logic.v(241)
  wire Vcvow6;  // ../RTL/cortexm0ds_logic.v(1266)
  wire Vd0ju6;  // ../RTL/cortexm0ds_logic.v(790)
  wire Vd1iu6;  // ../RTL/cortexm0ds_logic.v(322)
  wire Vd1pw6;  // ../RTL/cortexm0ds_logic.v(1346)
  wire Vd7ju6;  // ../RTL/cortexm0ds_logic.v(883)
  wire Vd8iu6;  // ../RTL/cortexm0ds_logic.v(415)
  wire Vd8pw6;  // ../RTL/cortexm0ds_logic.v(1440)
  wire Vd9ow6;  // ../RTL/cortexm0ds_logic.v(972)
  wire Vdfiu6;  // ../RTL/cortexm0ds_logic.v(509)
  wire Vdgow6;  // ../RTL/cortexm0ds_logic.v(1065)
  wire Vdmiu6;  // ../RTL/cortexm0ds_logic.v(603)
  wire Vdnow6;  // ../RTL/cortexm0ds_logic.v(1159)
  wire Vdtiu6;  // ../RTL/cortexm0ds_logic.v(696)
  wire Vduhu6;  // ../RTL/cortexm0ds_logic.v(228)
  wire Vduow6;  // ../RTL/cortexm0ds_logic.v(1253)
  wire Vdvax6;  // ../RTL/cortexm0ds_logic.v(1671)
  wire Ve0iu6;  // ../RTL/cortexm0ds_logic.v(309)
  wire Ve0pw6;  // ../RTL/cortexm0ds_logic.v(1333)
  wire Ve6ju6;  // ../RTL/cortexm0ds_logic.v(870)
  wire Ve7iu6;  // ../RTL/cortexm0ds_logic.v(402)
  wire Ve7pw6;  // ../RTL/cortexm0ds_logic.v(1427)
  wire Ve8ow6;  // ../RTL/cortexm0ds_logic.v(959)
  wire Veeiu6;  // ../RTL/cortexm0ds_logic.v(496)
  wire Vefax6;  // ../RTL/cortexm0ds_logic.v(1642)
  wire Vefow6;  // ../RTL/cortexm0ds_logic.v(1052)
  wire Veliu6;  // ../RTL/cortexm0ds_logic.v(590)
  wire Vemow6;  // ../RTL/cortexm0ds_logic.v(1146)
  wire Veqax6;  // ../RTL/cortexm0ds_logic.v(1662)
  wire Vesiu6;  // ../RTL/cortexm0ds_logic.v(683)
  wire Vethu6;  // ../RTL/cortexm0ds_logic.v(215)
  wire Vetow6;  // ../RTL/cortexm0ds_logic.v(1240)
  wire Veziu6;  // ../RTL/cortexm0ds_logic.v(777)
  wire Vf5ju6;  // ../RTL/cortexm0ds_logic.v(857)
  wire Vf6iu6;  // ../RTL/cortexm0ds_logic.v(389)
  wire Vf6pw6;  // ../RTL/cortexm0ds_logic.v(1414)
  wire Vf7ow6;  // ../RTL/cortexm0ds_logic.v(946)
  wire Vfdiu6;  // ../RTL/cortexm0ds_logic.v(483)
  wire Vfdpw6;  // ../RTL/cortexm0ds_logic.v(1507)
  wire Vfeow6;  // ../RTL/cortexm0ds_logic.v(1039)
  wire Vfkiu6;  // ../RTL/cortexm0ds_logic.v(577)
  wire Vflow6;  // ../RTL/cortexm0ds_logic.v(1133)
  wire Vfriu6;  // ../RTL/cortexm0ds_logic.v(670)
  wire Vfshu6;  // ../RTL/cortexm0ds_logic.v(202)
  wire Vfsow6;  // ../RTL/cortexm0ds_logic.v(1227)
  wire Vfvax6;  // ../RTL/cortexm0ds_logic.v(1671)
  wire Vfyiu6;  // ../RTL/cortexm0ds_logic.v(764)
  wire Vfzhu6;  // ../RTL/cortexm0ds_logic.v(296)
  wire Vfzow6;  // ../RTL/cortexm0ds_logic.v(1320)
  wire Vg4ju6;  // ../RTL/cortexm0ds_logic.v(844)
  wire Vg5iu6;  // ../RTL/cortexm0ds_logic.v(376)
  wire Vg5pw6;  // ../RTL/cortexm0ds_logic.v(1401)
  wire Vg6ow6;  // ../RTL/cortexm0ds_logic.v(933)
  wire Vgciu6;  // ../RTL/cortexm0ds_logic.v(470)
  wire Vgcpw6;  // ../RTL/cortexm0ds_logic.v(1494)
  wire Vgdow6;  // ../RTL/cortexm0ds_logic.v(1026)
  wire Vgjiu6;  // ../RTL/cortexm0ds_logic.v(564)
  wire Vgjpw6;  // ../RTL/cortexm0ds_logic.v(1587)
  wire Vgkow6;  // ../RTL/cortexm0ds_logic.v(1120)
  wire Vgqax6;  // ../RTL/cortexm0ds_logic.v(1662)
  wire Vgqiu6;  // ../RTL/cortexm0ds_logic.v(657)
  wire Vgrhu6;  // ../RTL/cortexm0ds_logic.v(189)
  wire Vgrow6;  // ../RTL/cortexm0ds_logic.v(1214)
  wire Vgxiu6;  // ../RTL/cortexm0ds_logic.v(751)
  wire Vgyhu6;  // ../RTL/cortexm0ds_logic.v(283)
  wire Vgyow6;  // ../RTL/cortexm0ds_logic.v(1307)
  wire Vh3ju6;  // ../RTL/cortexm0ds_logic.v(831)
  wire Vh4iu6;  // ../RTL/cortexm0ds_logic.v(363)
  wire Vh4pw6;  // ../RTL/cortexm0ds_logic.v(1388)
  wire Vhaju6;  // ../RTL/cortexm0ds_logic.v(925)
  wire Vhbiu6;  // ../RTL/cortexm0ds_logic.v(457)
  wire Vhbpw6;  // ../RTL/cortexm0ds_logic.v(1481)
  wire Vhcow6;  // ../RTL/cortexm0ds_logic.v(1013)
  wire Vhiiu6;  // ../RTL/cortexm0ds_logic.v(551)
  wire Vhjow6;  // ../RTL/cortexm0ds_logic.v(1107)
  wire Vhpiu6;  // ../RTL/cortexm0ds_logic.v(644)
  wire Vhqhu6;  // ../RTL/cortexm0ds_logic.v(176)
  wire Vhqow6;  // ../RTL/cortexm0ds_logic.v(1201)
  wire Vhspw6;  // ../RTL/cortexm0ds_logic.v(1603)
  wire Vhwiu6;  // ../RTL/cortexm0ds_logic.v(738)
  wire Vhxhu6;  // ../RTL/cortexm0ds_logic.v(270)
  wire Vhxow6;  // ../RTL/cortexm0ds_logic.v(1294)
  wire Vi2ju6;  // ../RTL/cortexm0ds_logic.v(818)
  wire Vi3iu6;  // ../RTL/cortexm0ds_logic.v(350)
  wire Vi3pw6;  // ../RTL/cortexm0ds_logic.v(1375)
  wire Vi9ju6;  // ../RTL/cortexm0ds_logic.v(912)
  wire Viaiu6;  // ../RTL/cortexm0ds_logic.v(444)
  wire Viapw6;  // ../RTL/cortexm0ds_logic.v(1468)
  wire Vibax6;  // ../RTL/cortexm0ds_logic.v(1634)
  wire Vibow6;  // ../RTL/cortexm0ds_logic.v(1000)
  wire Vihiu6;  // ../RTL/cortexm0ds_logic.v(538)
  wire Viiow6;  // ../RTL/cortexm0ds_logic.v(1094)
  wire Vioiu6;  // ../RTL/cortexm0ds_logic.v(631)
  wire Viphu6;  // ../RTL/cortexm0ds_logic.v(163)
  wire Vipow6;  // ../RTL/cortexm0ds_logic.v(1188)
  wire Viqax6;  // ../RTL/cortexm0ds_logic.v(1662)
  wire Viviu6;  // ../RTL/cortexm0ds_logic.v(725)
  wire Viwhu6;  // ../RTL/cortexm0ds_logic.v(257)
  wire Viwow6;  // ../RTL/cortexm0ds_logic.v(1281)
  wire Vj1ju6;  // ../RTL/cortexm0ds_logic.v(805)
  wire Vj2iu6;  // ../RTL/cortexm0ds_logic.v(337)
  wire Vj2pw6;  // ../RTL/cortexm0ds_logic.v(1362)
  wire Vj3qw6;  // ../RTL/cortexm0ds_logic.v(1624)
  wire Vj8ju6;  // ../RTL/cortexm0ds_logic.v(899)
  wire Vj9iu6;  // ../RTL/cortexm0ds_logic.v(431)
  wire Vj9pw6;  // ../RTL/cortexm0ds_logic.v(1455)
  wire Vjaow6;  // ../RTL/cortexm0ds_logic.v(987)
  wire Vjgiu6;  // ../RTL/cortexm0ds_logic.v(525)
  wire Vjhow6;  // ../RTL/cortexm0ds_logic.v(1081)
  wire Vjniu6;  // ../RTL/cortexm0ds_logic.v(618)
  wire Vjohu6;  // ../RTL/cortexm0ds_logic.v(150)
  wire Vjoow6;  // ../RTL/cortexm0ds_logic.v(1175)
  wire Vjuiu6;  // ../RTL/cortexm0ds_logic.v(712)
  wire Vjvhu6;  // ../RTL/cortexm0ds_logic.v(244)
  wire Vjvow6;  // ../RTL/cortexm0ds_logic.v(1268)
  wire Vk0ju6;  // ../RTL/cortexm0ds_logic.v(792)
  wire Vk1iu6;  // ../RTL/cortexm0ds_logic.v(324)
  wire Vk1pw6;  // ../RTL/cortexm0ds_logic.v(1349)
  wire Vk7ju6;  // ../RTL/cortexm0ds_logic.v(886)
  wire Vk8iu6;  // ../RTL/cortexm0ds_logic.v(418)
  wire Vk8pw6;  // ../RTL/cortexm0ds_logic.v(1442)
  wire Vk9ow6;  // ../RTL/cortexm0ds_logic.v(974)
  wire Vkfiu6;  // ../RTL/cortexm0ds_logic.v(512)
  wire Vkgow6;  // ../RTL/cortexm0ds_logic.v(1068)
  wire Vkmiu6;  // ../RTL/cortexm0ds_logic.v(605)
  wire Vknow6;  // ../RTL/cortexm0ds_logic.v(1162)
  wire Vkqax6;  // ../RTL/cortexm0ds_logic.v(1662)
  wire Vktiu6;  // ../RTL/cortexm0ds_logic.v(699)
  wire Vkuhu6;  // ../RTL/cortexm0ds_logic.v(231)
  wire Vkuow6;  // ../RTL/cortexm0ds_logic.v(1255)
  wire Vkzax6;  // ../RTL/cortexm0ds_logic.v(1679)
  wire Vl0iu6;  // ../RTL/cortexm0ds_logic.v(311)
  wire Vl0pw6;  // ../RTL/cortexm0ds_logic.v(1336)
  wire Vl6ju6;  // ../RTL/cortexm0ds_logic.v(873)
  wire Vl7iu6;  // ../RTL/cortexm0ds_logic.v(405)
  wire Vl7pw6;  // ../RTL/cortexm0ds_logic.v(1429)
  wire Vl8ow6;  // ../RTL/cortexm0ds_logic.v(961)
  wire Vlaax6;  // ../RTL/cortexm0ds_logic.v(1632)
  wire Vleiu6;  // ../RTL/cortexm0ds_logic.v(499)
  wire Vlfow6;  // ../RTL/cortexm0ds_logic.v(1055)
  wire Vlkpw6;  // ../RTL/cortexm0ds_logic.v(1589)
  wire Vlliu6;  // ../RTL/cortexm0ds_logic.v(592)
  wire Vlmow6;  // ../RTL/cortexm0ds_logic.v(1149)
  wire Vlsiu6;  // ../RTL/cortexm0ds_logic.v(686)
  wire Vlthu6;  // ../RTL/cortexm0ds_logic.v(218)
  wire Vltow6;  // ../RTL/cortexm0ds_logic.v(1242)
  wire Vltpw6;  // ../RTL/cortexm0ds_logic.v(1605)
  wire Vlxax6;  // ../RTL/cortexm0ds_logic.v(1675)
  wire Vlziu6;  // ../RTL/cortexm0ds_logic.v(779)
  wire Vm5ju6;  // ../RTL/cortexm0ds_logic.v(860)
  wire Vm6iu6;  // ../RTL/cortexm0ds_logic.v(392)
  wire Vm6pw6;  // ../RTL/cortexm0ds_logic.v(1416)
  wire Vm7ow6;  // ../RTL/cortexm0ds_logic.v(948)
  wire Vmdiu6;  // ../RTL/cortexm0ds_logic.v(486)
  wire Vmdpw6;  // ../RTL/cortexm0ds_logic.v(1510)
  wire Vmeow6;  // ../RTL/cortexm0ds_logic.v(1042)
  wire Vmipw6;  // ../RTL/cortexm0ds_logic.v(1585)
  wire Vmkiu6;  // ../RTL/cortexm0ds_logic.v(579)
  wire Vmlow6;  // ../RTL/cortexm0ds_logic.v(1136)
  wire Vmqax6;  // ../RTL/cortexm0ds_logic.v(1662)
  wire Vmriu6;  // ../RTL/cortexm0ds_logic.v(673)
  wire Vmshu6;  // ../RTL/cortexm0ds_logic.v(205)
  wire Vmsow6;  // ../RTL/cortexm0ds_logic.v(1229)
  wire Vmyiu6;  // ../RTL/cortexm0ds_logic.v(766)
  wire Vmzhu6;  // ../RTL/cortexm0ds_logic.v(298)
  wire Vmzow6;  // ../RTL/cortexm0ds_logic.v(1323)
  wire Vn4ju6;  // ../RTL/cortexm0ds_logic.v(847)
  wire Vn5iu6;  // ../RTL/cortexm0ds_logic.v(379)
  wire Vn5pw6;  // ../RTL/cortexm0ds_logic.v(1403)
  wire Vn6ow6;  // ../RTL/cortexm0ds_logic.v(935)
  wire Vn9bx6;  // ../RTL/cortexm0ds_logic.v(1696)
  wire Vnciu6;  // ../RTL/cortexm0ds_logic.v(473)
  wire Vncpw6;  // ../RTL/cortexm0ds_logic.v(1497)
  wire Vndow6;  // ../RTL/cortexm0ds_logic.v(1029)
  wire Vnjiu6;  // ../RTL/cortexm0ds_logic.v(566)
  wire Vnkow6;  // ../RTL/cortexm0ds_logic.v(1123)
  wire Vnkpw6;  // ../RTL/cortexm0ds_logic.v(1589)
  wire Vnqiu6;  // ../RTL/cortexm0ds_logic.v(660)
  wire Vnrhu6;  // ../RTL/cortexm0ds_logic.v(192)
  wire Vnrow6;  // ../RTL/cortexm0ds_logic.v(1216)
  wire Vnxiu6;  // ../RTL/cortexm0ds_logic.v(753)
  wire Vnyhu6;  // ../RTL/cortexm0ds_logic.v(285)
  wire Vnyow6;  // ../RTL/cortexm0ds_logic.v(1310)
  wire Vo3ju6;  // ../RTL/cortexm0ds_logic.v(834)
  wire Vo4iu6;  // ../RTL/cortexm0ds_logic.v(366)
  wire Vo4pw6;  // ../RTL/cortexm0ds_logic.v(1390)
  wire Voaju6;  // ../RTL/cortexm0ds_logic.v(928)
  wire Vobiu6;  // ../RTL/cortexm0ds_logic.v(460)
  wire Vobpw6;  // ../RTL/cortexm0ds_logic.v(1484)
  wire Vocow6;  // ../RTL/cortexm0ds_logic.v(1016)
  wire Voiiu6;  // ../RTL/cortexm0ds_logic.v(553)
  wire Vojow6;  // ../RTL/cortexm0ds_logic.v(1110)
  wire Vopiu6;  // ../RTL/cortexm0ds_logic.v(647)
  wire Voqhu6;  // ../RTL/cortexm0ds_logic.v(179)
  wire Voqow6;  // ../RTL/cortexm0ds_logic.v(1203)
  wire Vowiu6;  // ../RTL/cortexm0ds_logic.v(740)
  wire Voxhu6;  // ../RTL/cortexm0ds_logic.v(272)
  wire Voxow6;  // ../RTL/cortexm0ds_logic.v(1297)
  wire Vp2ju6;  // ../RTL/cortexm0ds_logic.v(821)
  wire Vp3iu6;  // ../RTL/cortexm0ds_logic.v(353)
  wire Vp3pw6;  // ../RTL/cortexm0ds_logic.v(1377)
  wire Vp9ju6;  // ../RTL/cortexm0ds_logic.v(915)
  wire Vpaiu6;  // ../RTL/cortexm0ds_logic.v(447)
  wire Vpapw6;  // ../RTL/cortexm0ds_logic.v(1471)
  wire Vpbow6;  // ../RTL/cortexm0ds_logic.v(1003)
  wire Vpgbx6;  // ../RTL/cortexm0ds_logic.v(1709)
  wire Vphiu6;  // ../RTL/cortexm0ds_logic.v(540)
  wire Vpiow6;  // ../RTL/cortexm0ds_logic.v(1097)
  wire Vpkpw6;  // ../RTL/cortexm0ds_logic.v(1589)
  wire Vplpw6;  // ../RTL/cortexm0ds_logic.v(1591)
  wire Vpoiu6;  // ../RTL/cortexm0ds_logic.v(634)
  wire Vpphu6;  // ../RTL/cortexm0ds_logic.v(166)
  wire Vppow6;  // ../RTL/cortexm0ds_logic.v(1190)
  wire Vpviu6;  // ../RTL/cortexm0ds_logic.v(727)
  wire Vpwhu6;  // ../RTL/cortexm0ds_logic.v(259)
  wire Vpwow6;  // ../RTL/cortexm0ds_logic.v(1284)
  wire Vq1ju6;  // ../RTL/cortexm0ds_logic.v(808)
  wire Vq2iu6;  // ../RTL/cortexm0ds_logic.v(340)
  wire Vq2pw6;  // ../RTL/cortexm0ds_logic.v(1364)
  wire Vq8ju6;  // ../RTL/cortexm0ds_logic.v(902)
  wire Vq9iu6;  // ../RTL/cortexm0ds_logic.v(434)
  wire Vq9pw6;  // ../RTL/cortexm0ds_logic.v(1458)
  wire Vqaow6;  // ../RTL/cortexm0ds_logic.v(990)
  wire Vqgax6;  // ../RTL/cortexm0ds_logic.v(1644)
  wire Vqgiu6;  // ../RTL/cortexm0ds_logic.v(527)
  wire Vqhow6;  // ../RTL/cortexm0ds_logic.v(1084)
  wire Vqjbx6;  // ../RTL/cortexm0ds_logic.v(1715)
  wire Vqniu6;  // ../RTL/cortexm0ds_logic.v(621)
  wire Vqohu6;  // ../RTL/cortexm0ds_logic.v(153)
  wire Vqoow6;  // ../RTL/cortexm0ds_logic.v(1177)
  wire Vquiu6;  // ../RTL/cortexm0ds_logic.v(714)
  wire Vqvhu6;  // ../RTL/cortexm0ds_logic.v(246)
  wire Vqvow6;  // ../RTL/cortexm0ds_logic.v(1271)
  wire Vr0ju6;  // ../RTL/cortexm0ds_logic.v(795)
  wire Vr1iu6;  // ../RTL/cortexm0ds_logic.v(327)
  wire Vr1pw6;  // ../RTL/cortexm0ds_logic.v(1351)
  wire Vr7ju6;  // ../RTL/cortexm0ds_logic.v(889)
  wire Vr8iu6;  // ../RTL/cortexm0ds_logic.v(421)
  wire Vr8pw6;  // ../RTL/cortexm0ds_logic.v(1445)
  wire Vr9ow6;  // ../RTL/cortexm0ds_logic.v(977)
  wire Vrfhu6;  // ../RTL/cortexm0ds_logic.v(125)
  wire Vrfiu6;  // ../RTL/cortexm0ds_logic.v(514)
  wire Vrgow6;  // ../RTL/cortexm0ds_logic.v(1071)
  wire Vrmiu6;  // ../RTL/cortexm0ds_logic.v(608)
  wire Vrnow6;  // ../RTL/cortexm0ds_logic.v(1164)
  wire Vrtiu6;  // ../RTL/cortexm0ds_logic.v(701)
  wire Vrtpw6;  // ../RTL/cortexm0ds_logic.v(1606)
  wire Vruhu6;  // ../RTL/cortexm0ds_logic.v(233)
  wire Vruow6;  // ../RTL/cortexm0ds_logic.v(1258)
  wire Vs0iu6;  // ../RTL/cortexm0ds_logic.v(314)
  wire Vs0pw6;  // ../RTL/cortexm0ds_logic.v(1338)
  wire Vs6ju6;  // ../RTL/cortexm0ds_logic.v(876)
  wire Vs7iu6;  // ../RTL/cortexm0ds_logic.v(408)
  wire Vs7pw6;  // ../RTL/cortexm0ds_logic.v(1432)
  wire Vs8ow6;  // ../RTL/cortexm0ds_logic.v(964)
  wire Vseiu6;  // ../RTL/cortexm0ds_logic.v(501)
  wire Vsfow6;  // ../RTL/cortexm0ds_logic.v(1058)
  wire Vsliu6;  // ../RTL/cortexm0ds_logic.v(595)
  wire Vsmow6;  // ../RTL/cortexm0ds_logic.v(1151)
  wire Vssiu6;  // ../RTL/cortexm0ds_logic.v(688)
  wire Vsthu6;  // ../RTL/cortexm0ds_logic.v(220)
  wire Vstow6;  // ../RTL/cortexm0ds_logic.v(1245)
  wire Vsziu6;  // ../RTL/cortexm0ds_logic.v(782)
  wire Vszpw6;  // ../RTL/cortexm0ds_logic.v(1617)
  wire Vt5ju6;  // ../RTL/cortexm0ds_logic.v(863)
  wire Vt6iu6;  // ../RTL/cortexm0ds_logic.v(395)
  wire Vt6pw6;  // ../RTL/cortexm0ds_logic.v(1419)
  wire Vt7ow6;  // ../RTL/cortexm0ds_logic.v(951)
  wire Vtdiu6;  // ../RTL/cortexm0ds_logic.v(488)
  wire Vtdpw6;  // ../RTL/cortexm0ds_logic.v(1513)
  wire Vteow6;  // ../RTL/cortexm0ds_logic.v(1045)
  wire Vtkiu6;  // ../RTL/cortexm0ds_logic.v(582)
  wire Vtlow6;  // ../RTL/cortexm0ds_logic.v(1138)
  wire Vtmax6;  // ../RTL/cortexm0ds_logic.v(1656)
  wire Vtriu6;  // ../RTL/cortexm0ds_logic.v(675)
  wire Vtshu6;  // ../RTL/cortexm0ds_logic.v(207)
  wire Vtsow6;  // ../RTL/cortexm0ds_logic.v(1232)
  wire Vtuax6;  // ../RTL/cortexm0ds_logic.v(1670)
  wire Vtyiu6;  // ../RTL/cortexm0ds_logic.v(769)
  wire Vtzhu6;  // ../RTL/cortexm0ds_logic.v(301)
  wire Vtzow6;  // ../RTL/cortexm0ds_logic.v(1325)
  wire Vu4ju6;  // ../RTL/cortexm0ds_logic.v(850)
  wire Vu5iu6;  // ../RTL/cortexm0ds_logic.v(382)
  wire Vu5pw6;  // ../RTL/cortexm0ds_logic.v(1406)
  wire Vu6ow6;  // ../RTL/cortexm0ds_logic.v(938)
  wire Vuciu6;  // ../RTL/cortexm0ds_logic.v(475)
  wire Vucpw6;  // ../RTL/cortexm0ds_logic.v(1500)
  wire Vudow6;  // ../RTL/cortexm0ds_logic.v(1032)
  wire Vuhax6;  // ../RTL/cortexm0ds_logic.v(1646)
  wire Vuipw6;  // ../RTL/cortexm0ds_logic.v(1585)
  wire Vujiu6;  // ../RTL/cortexm0ds_logic.v(569)
  wire Vukow6;  // ../RTL/cortexm0ds_logic.v(1125)
  wire Vuqiu6;  // ../RTL/cortexm0ds_logic.v(662)
  wire Vurhu6;  // ../RTL/cortexm0ds_logic.v(194)
  wire Vurow6;  // ../RTL/cortexm0ds_logic.v(1219)
  wire Vuxiu6;  // ../RTL/cortexm0ds_logic.v(756)
  wire Vuyhu6;  // ../RTL/cortexm0ds_logic.v(288)
  wire Vuyow6;  // ../RTL/cortexm0ds_logic.v(1312)
  wire Vv3ju6;  // ../RTL/cortexm0ds_logic.v(837)
  wire Vv4iu6;  // ../RTL/cortexm0ds_logic.v(369)
  wire Vv4pw6;  // ../RTL/cortexm0ds_logic.v(1393)
  wire Vvbiu6;  // ../RTL/cortexm0ds_logic.v(462)
  wire Vvbpw6;  // ../RTL/cortexm0ds_logic.v(1487)
  wire Vvcow6;  // ../RTL/cortexm0ds_logic.v(1019)
  wire Vviiu6;  // ../RTL/cortexm0ds_logic.v(556)
  wire Vvjow6;  // ../RTL/cortexm0ds_logic.v(1112)
  wire Vvpiu6;  // ../RTL/cortexm0ds_logic.v(649)
  wire Vvqhu6;  // ../RTL/cortexm0ds_logic.v(181)
  wire Vvqow6;  // ../RTL/cortexm0ds_logic.v(1206)
  wire Vvuax6;  // ../RTL/cortexm0ds_logic.v(1670)
  wire Vvwiu6;  // ../RTL/cortexm0ds_logic.v(743)
  wire Vvxax6;  // ../RTL/cortexm0ds_logic.v(1676)
  wire Vvxhu6;  // ../RTL/cortexm0ds_logic.v(275)
  wire Vvxow6;  // ../RTL/cortexm0ds_logic.v(1299)
  wire Vw2ju6;  // ../RTL/cortexm0ds_logic.v(824)
  wire Vw3iu6;  // ../RTL/cortexm0ds_logic.v(356)
  wire Vw3pw6;  // ../RTL/cortexm0ds_logic.v(1380)
  wire Vw9ju6;  // ../RTL/cortexm0ds_logic.v(917)
  wire Vwaiu6;  // ../RTL/cortexm0ds_logic.v(449)
  wire Vwapw6;  // ../RTL/cortexm0ds_logic.v(1474)
  wire Vwbow6;  // ../RTL/cortexm0ds_logic.v(1006)
  wire Vwhiu6;  // ../RTL/cortexm0ds_logic.v(543)
  wire Vwiow6;  // ../RTL/cortexm0ds_logic.v(1099)
  wire Vwoiu6;  // ../RTL/cortexm0ds_logic.v(636)
  wire Vwphu6;  // ../RTL/cortexm0ds_logic.v(168)
  wire Vwpow6;  // ../RTL/cortexm0ds_logic.v(1193)
  wire Vwviu6;  // ../RTL/cortexm0ds_logic.v(730)
  wire Vwwhu6;  // ../RTL/cortexm0ds_logic.v(262)
  wire Vwwow6;  // ../RTL/cortexm0ds_logic.v(1286)
  wire Vx1ju6;  // ../RTL/cortexm0ds_logic.v(811)
  wire Vx2iu6;  // ../RTL/cortexm0ds_logic.v(343)
  wire Vx2pw6;  // ../RTL/cortexm0ds_logic.v(1367)
  wire Vx8ju6;  // ../RTL/cortexm0ds_logic.v(904)
  wire Vx9iu6;  // ../RTL/cortexm0ds_logic.v(436)
  wire Vx9pw6;  // ../RTL/cortexm0ds_logic.v(1461)
  wire Vxaow6;  // ../RTL/cortexm0ds_logic.v(993)
  wire Vxgiu6;  // ../RTL/cortexm0ds_logic.v(530)
  wire Vxhow6;  // ../RTL/cortexm0ds_logic.v(1086)
  wire Vxmhu6;  // ../RTL/cortexm0ds_logic.v(143)
  wire Vxniu6;  // ../RTL/cortexm0ds_logic.v(623)
  wire Vxohu6;  // ../RTL/cortexm0ds_logic.v(155)
  wire Vxoow6;  // ../RTL/cortexm0ds_logic.v(1180)
  wire Vxuax6;  // ../RTL/cortexm0ds_logic.v(1670)
  wire Vxuiu6;  // ../RTL/cortexm0ds_logic.v(717)
  wire Vxvhu6;  // ../RTL/cortexm0ds_logic.v(249)
  wire Vxvow6;  // ../RTL/cortexm0ds_logic.v(1273)
  wire Vxxax6;  // ../RTL/cortexm0ds_logic.v(1676)
  wire Vy0ju6;  // ../RTL/cortexm0ds_logic.v(798)
  wire Vy1iu6;  // ../RTL/cortexm0ds_logic.v(330)
  wire Vy1pw6;  // ../RTL/cortexm0ds_logic.v(1354)
  wire Vy7ju6;  // ../RTL/cortexm0ds_logic.v(891)
  wire Vy8pw6;  // ../RTL/cortexm0ds_logic.v(1448)
  wire Vy9ow6;  // ../RTL/cortexm0ds_logic.v(980)
  wire Vyfbx6;  // ../RTL/cortexm0ds_logic.v(1708)
  wire Vyfiu6;  // ../RTL/cortexm0ds_logic.v(517)
  wire Vygax6;  // ../RTL/cortexm0ds_logic.v(1645)
  wire Vygow6;  // ../RTL/cortexm0ds_logic.v(1073)
  wire Vymiu6;  // ../RTL/cortexm0ds_logic.v(610)
  wire Vynow6;  // ../RTL/cortexm0ds_logic.v(1167)
  wire Vytiu6;  // ../RTL/cortexm0ds_logic.v(704)
  wire Vyuhu6;  // ../RTL/cortexm0ds_logic.v(236)
  wire Vyuow6;  // ../RTL/cortexm0ds_logic.v(1260)
  wire Vz0iu6;  // ../RTL/cortexm0ds_logic.v(317)
  wire Vz0pw6;  // ../RTL/cortexm0ds_logic.v(1341)
  wire Vz6ju6;  // ../RTL/cortexm0ds_logic.v(878)
  wire Vz7iu6;  // ../RTL/cortexm0ds_logic.v(410)
  wire Vz7pw6;  // ../RTL/cortexm0ds_logic.v(1435)
  wire Vz8ax6;  // ../RTL/cortexm0ds_logic.v(1629)
  wire Vz8ow6;  // ../RTL/cortexm0ds_logic.v(967)
  wire Vzdax6;  // ../RTL/cortexm0ds_logic.v(1639)
  wire Vzeiu6;  // ../RTL/cortexm0ds_logic.v(504)
  wire Vzfow6;  // ../RTL/cortexm0ds_logic.v(1060)
  wire Vzjpw6;  // ../RTL/cortexm0ds_logic.v(1588)
  wire Vzliu6;  // ../RTL/cortexm0ds_logic.v(597)
  wire Vzmow6;  // ../RTL/cortexm0ds_logic.v(1154)
  wire Vzsiu6;  // ../RTL/cortexm0ds_logic.v(691)
  wire Vzthu6;  // ../RTL/cortexm0ds_logic.v(223)
  wire Vztow6;  // ../RTL/cortexm0ds_logic.v(1247)
  wire Vzuax6;  // ../RTL/cortexm0ds_logic.v(1670)
  wire Vzupw6;  // ../RTL/cortexm0ds_logic.v(1608)
  wire Vzxax6;  // ../RTL/cortexm0ds_logic.v(1676)
  wire Vzziu6;  // ../RTL/cortexm0ds_logic.v(785)
  wire W03ju6;  // ../RTL/cortexm0ds_logic.v(825)
  wire W04iu6;  // ../RTL/cortexm0ds_logic.v(357)
  wire W04pw6;  // ../RTL/cortexm0ds_logic.v(1382)
  wire W0aju6;  // ../RTL/cortexm0ds_logic.v(919)
  wire W0biu6;  // ../RTL/cortexm0ds_logic.v(451)
  wire W0bpw6;  // ../RTL/cortexm0ds_logic.v(1475)
  wire W0cow6;  // ../RTL/cortexm0ds_logic.v(1007)
  wire W0dbx6;  // ../RTL/cortexm0ds_logic.v(1703)
  wire W0iiu6;  // ../RTL/cortexm0ds_logic.v(544)
  wire W0jax6;  // ../RTL/cortexm0ds_logic.v(1649)
  wire W0jow6;  // ../RTL/cortexm0ds_logic.v(1101)
  wire W0piu6;  // ../RTL/cortexm0ds_logic.v(638)
  wire W0qhu6;  // ../RTL/cortexm0ds_logic.v(170)
  wire W0qow6;  // ../RTL/cortexm0ds_logic.v(1194)
  wire W0wiu6;  // ../RTL/cortexm0ds_logic.v(732)
  wire W0xhu6;  // ../RTL/cortexm0ds_logic.v(264)
  wire W0xow6;  // ../RTL/cortexm0ds_logic.v(1288)
  wire W12ju6;  // ../RTL/cortexm0ds_logic.v(812)
  wire W13iu6;  // ../RTL/cortexm0ds_logic.v(344)
  wire W13pw6;  // ../RTL/cortexm0ds_logic.v(1369)
  wire W19ju6;  // ../RTL/cortexm0ds_logic.v(906)
  wire W1aiu6;  // ../RTL/cortexm0ds_logic.v(438)
  wire W1apw6;  // ../RTL/cortexm0ds_logic.v(1462)
  wire W1bow6;  // ../RTL/cortexm0ds_logic.v(994)
  wire W1hiu6;  // ../RTL/cortexm0ds_logic.v(531)
  wire W1iow6;  // ../RTL/cortexm0ds_logic.v(1088)
  wire W1oiu6;  // ../RTL/cortexm0ds_logic.v(625)
  wire W1phu6;  // ../RTL/cortexm0ds_logic.v(157)
  wire W1pow6;  // ../RTL/cortexm0ds_logic.v(1181)
  wire W1viu6;  // ../RTL/cortexm0ds_logic.v(719)
  wire W1whu6;  // ../RTL/cortexm0ds_logic.v(251)
  wire W1wow6;  // ../RTL/cortexm0ds_logic.v(1275)
  wire W21ju6;  // ../RTL/cortexm0ds_logic.v(799)
  wire W22iu6;  // ../RTL/cortexm0ds_logic.v(331)
  wire W22pw6;  // ../RTL/cortexm0ds_logic.v(1356)
  wire W28ju6;  // ../RTL/cortexm0ds_logic.v(893)
  wire W29iu6;  // ../RTL/cortexm0ds_logic.v(425)
  wire W29pw6;  // ../RTL/cortexm0ds_logic.v(1449)
  wire W2aow6;  // ../RTL/cortexm0ds_logic.v(981)
  wire W2giu6;  // ../RTL/cortexm0ds_logic.v(518)
  wire W2how6;  // ../RTL/cortexm0ds_logic.v(1075)
  wire W2jax6;  // ../RTL/cortexm0ds_logic.v(1649)
  wire W2niu6;  // ../RTL/cortexm0ds_logic.v(612)
  wire W2oow6;  // ../RTL/cortexm0ds_logic.v(1168)
  wire W2uiu6;  // ../RTL/cortexm0ds_logic.v(706)
  wire W2vhu6;  // ../RTL/cortexm0ds_logic.v(238)
  wire W2vow6;  // ../RTL/cortexm0ds_logic.v(1262)
  wire W30ju6;  // ../RTL/cortexm0ds_logic.v(786)
  wire W31iu6;  // ../RTL/cortexm0ds_logic.v(318)
  wire W31pw6;  // ../RTL/cortexm0ds_logic.v(1343)
  wire W37ju6;  // ../RTL/cortexm0ds_logic.v(880)
  wire W38iu6;  // ../RTL/cortexm0ds_logic.v(412)
  wire W38pw6;  // ../RTL/cortexm0ds_logic.v(1436)
  wire W39ow6;  // ../RTL/cortexm0ds_logic.v(968)
  wire W3fiu6;  // ../RTL/cortexm0ds_logic.v(505)
  wire W3gow6;  // ../RTL/cortexm0ds_logic.v(1062)
  wire W3miu6;  // ../RTL/cortexm0ds_logic.v(599)
  wire W3now6;  // ../RTL/cortexm0ds_logic.v(1155)
  wire W3tiu6;  // ../RTL/cortexm0ds_logic.v(693)
  wire W3uhu6;  // ../RTL/cortexm0ds_logic.v(225)
  wire W3uow6;  // ../RTL/cortexm0ds_logic.v(1249)
  wire W40iu6;  // ../RTL/cortexm0ds_logic.v(305)
  wire W40pw6;  // ../RTL/cortexm0ds_logic.v(1330)
  wire W46ju6;  // ../RTL/cortexm0ds_logic.v(867)
  wire W47iu6;  // ../RTL/cortexm0ds_logic.v(399)
  wire W47pw6;  // ../RTL/cortexm0ds_logic.v(1423)
  wire W48ow6;  // ../RTL/cortexm0ds_logic.v(955)
  wire W4aax6;  // ../RTL/cortexm0ds_logic.v(1631)
  wire W4eiu6;  // ../RTL/cortexm0ds_logic.v(492)
  wire W4epw6;  // ../RTL/cortexm0ds_logic.v(1517)
  wire W4fhu6;  // ../RTL/cortexm0ds_logic.v(123)
  wire W4fow6;  // ../RTL/cortexm0ds_logic.v(1049)
  wire W4jax6;  // ../RTL/cortexm0ds_logic.v(1649)
  wire W4liu6;  // ../RTL/cortexm0ds_logic.v(586)
  wire W4mow6;  // ../RTL/cortexm0ds_logic.v(1142)
  wire W4siu6;  // ../RTL/cortexm0ds_logic.v(680)
  wire W4thu6;  // ../RTL/cortexm0ds_logic.v(212)
  wire W4tow6;  // ../RTL/cortexm0ds_logic.v(1236)
  wire W4ziu6;  // ../RTL/cortexm0ds_logic.v(773)
  wire W51bx6;  // ../RTL/cortexm0ds_logic.v(1681)
  wire W55ju6;  // ../RTL/cortexm0ds_logic.v(854)
  wire W56iu6;  // ../RTL/cortexm0ds_logic.v(386)
  wire W56pw6;  // ../RTL/cortexm0ds_logic.v(1410)
  wire W57ow6;  // ../RTL/cortexm0ds_logic.v(942)
  wire W5diu6;  // ../RTL/cortexm0ds_logic.v(479)
  wire W5dpw6;  // ../RTL/cortexm0ds_logic.v(1504)
  wire W5eow6;  // ../RTL/cortexm0ds_logic.v(1036)
  wire W5kiu6;  // ../RTL/cortexm0ds_logic.v(573)
  wire W5low6;  // ../RTL/cortexm0ds_logic.v(1129)
  wire W5max6;  // ../RTL/cortexm0ds_logic.v(1654)
  wire W5riu6;  // ../RTL/cortexm0ds_logic.v(667)
  wire W5shu6;  // ../RTL/cortexm0ds_logic.v(199)
  wire W5sow6;  // ../RTL/cortexm0ds_logic.v(1223)
  wire W5yiu6;  // ../RTL/cortexm0ds_logic.v(760)
  wire W5ypw6;  // ../RTL/cortexm0ds_logic.v(1614)
  wire W5zhu6;  // ../RTL/cortexm0ds_logic.v(292)
  wire W5zow6;  // ../RTL/cortexm0ds_logic.v(1317)
  wire W64ju6;  // ../RTL/cortexm0ds_logic.v(841)
  wire W65iu6;  // ../RTL/cortexm0ds_logic.v(373)
  wire W65pw6;  // ../RTL/cortexm0ds_logic.v(1397)
  wire W6ciu6;  // ../RTL/cortexm0ds_logic.v(466)
  wire W6cpw6;  // ../RTL/cortexm0ds_logic.v(1491)
  wire W6dow6;  // ../RTL/cortexm0ds_logic.v(1023)
  wire W6ipw6;  // ../RTL/cortexm0ds_logic.v(1584)
  wire W6jiu6;  // ../RTL/cortexm0ds_logic.v(560)
  wire W6kow6;  // ../RTL/cortexm0ds_logic.v(1116)
  wire W6qiu6;  // ../RTL/cortexm0ds_logic.v(654)
  wire W6rhu6;  // ../RTL/cortexm0ds_logic.v(186)
  wire W6row6;  // ../RTL/cortexm0ds_logic.v(1210)
  wire W6xiu6;  // ../RTL/cortexm0ds_logic.v(747)
  wire W6yhu6;  // ../RTL/cortexm0ds_logic.v(279)
  wire W6yow6;  // ../RTL/cortexm0ds_logic.v(1304)
  wire W73ju6;  // ../RTL/cortexm0ds_logic.v(828)
  wire W74iu6;  // ../RTL/cortexm0ds_logic.v(360)
  wire W74pw6;  // ../RTL/cortexm0ds_logic.v(1384)
  wire W7aju6;  // ../RTL/cortexm0ds_logic.v(921)
  wire W7biu6;  // ../RTL/cortexm0ds_logic.v(453)
  wire W7bpw6;  // ../RTL/cortexm0ds_logic.v(1478)
  wire W7cow6;  // ../RTL/cortexm0ds_logic.v(1010)
  wire W7iiu6;  // ../RTL/cortexm0ds_logic.v(547)
  wire W7jow6;  // ../RTL/cortexm0ds_logic.v(1103)
  wire W7max6;  // ../RTL/cortexm0ds_logic.v(1654)
  wire W7piu6;  // ../RTL/cortexm0ds_logic.v(641)
  wire W7qhu6;  // ../RTL/cortexm0ds_logic.v(173)
  wire W7qow6;  // ../RTL/cortexm0ds_logic.v(1197)
  wire W7wiu6;  // ../RTL/cortexm0ds_logic.v(734)
  wire W7xhu6;  // ../RTL/cortexm0ds_logic.v(266)
  wire W7xow6;  // ../RTL/cortexm0ds_logic.v(1291)
  wire W82ju6;  // ../RTL/cortexm0ds_logic.v(815)
  wire W83iu6;  // ../RTL/cortexm0ds_logic.v(347)
  wire W83pw6;  // ../RTL/cortexm0ds_logic.v(1371)
  wire W89ju6;  // ../RTL/cortexm0ds_logic.v(908)
  wire W8aiu6;  // ../RTL/cortexm0ds_logic.v(440)
  wire W8apw6;  // ../RTL/cortexm0ds_logic.v(1465)
  wire W8bow6;  // ../RTL/cortexm0ds_logic.v(997)
  wire W8hbx6;  // ../RTL/cortexm0ds_logic.v(1710)
  wire W8hiu6;  // ../RTL/cortexm0ds_logic.v(534)
  wire W8iow6;  // ../RTL/cortexm0ds_logic.v(1090)
  wire W8oiu6;  // ../RTL/cortexm0ds_logic.v(628)
  wire W8phu6;  // ../RTL/cortexm0ds_logic.v(160)
  wire W8pow6;  // ../RTL/cortexm0ds_logic.v(1184)
  wire W8viu6;  // ../RTL/cortexm0ds_logic.v(721)
  wire W8whu6;  // ../RTL/cortexm0ds_logic.v(253)
  wire W8wow6;  // ../RTL/cortexm0ds_logic.v(1278)
  wire W91ju6;  // ../RTL/cortexm0ds_logic.v(802)
  wire W92iu6;  // ../RTL/cortexm0ds_logic.v(334)
  wire W92pw6;  // ../RTL/cortexm0ds_logic.v(1358)
  wire W98ju6;  // ../RTL/cortexm0ds_logic.v(895)
  wire W99iu6;  // ../RTL/cortexm0ds_logic.v(427)
  wire W99pw6;  // ../RTL/cortexm0ds_logic.v(1452)
  wire W9aow6;  // ../RTL/cortexm0ds_logic.v(984)
  wire W9giu6;  // ../RTL/cortexm0ds_logic.v(521)
  wire W9how6;  // ../RTL/cortexm0ds_logic.v(1077)
  wire W9lhu6;  // ../RTL/cortexm0ds_logic.v(139)
  wire W9max6;  // ../RTL/cortexm0ds_logic.v(1655)
  wire W9niu6;  // ../RTL/cortexm0ds_logic.v(615)
  wire W9ohu6;  // ../RTL/cortexm0ds_logic.v(147)
  wire W9oow6;  // ../RTL/cortexm0ds_logic.v(1171)
  wire W9spw6;  // ../RTL/cortexm0ds_logic.v(1603)
  wire W9uiu6;  // ../RTL/cortexm0ds_logic.v(708)
  wire W9vhu6;  // ../RTL/cortexm0ds_logic.v(240)
  wire W9vow6;  // ../RTL/cortexm0ds_logic.v(1265)
  wire Wa0ju6;  // ../RTL/cortexm0ds_logic.v(789)
  wire Wa1iu6;  // ../RTL/cortexm0ds_logic.v(321)
  wire Wa1pw6;  // ../RTL/cortexm0ds_logic.v(1345)
  wire Wa7ju6;  // ../RTL/cortexm0ds_logic.v(882)
  wire Wa8iu6;  // ../RTL/cortexm0ds_logic.v(414)
  wire Wa8pw6;  // ../RTL/cortexm0ds_logic.v(1439)
  wire Wa9ow6;  // ../RTL/cortexm0ds_logic.v(971)
  wire Wafiu6;  // ../RTL/cortexm0ds_logic.v(508)
  wire Wagow6;  // ../RTL/cortexm0ds_logic.v(1064)
  wire Wahbx6;  // ../RTL/cortexm0ds_logic.v(1711)
  wire Wamiu6;  // ../RTL/cortexm0ds_logic.v(602)
  wire Wanow6;  // ../RTL/cortexm0ds_logic.v(1158)
  wire Watiu6;  // ../RTL/cortexm0ds_logic.v(695)
  wire Wauhu6;  // ../RTL/cortexm0ds_logic.v(227)
  wire Wauow6;  // ../RTL/cortexm0ds_logic.v(1252)
  wire Wb0iu6;  // ../RTL/cortexm0ds_logic.v(308)
  wire Wb0pw6;  // ../RTL/cortexm0ds_logic.v(1332)
  wire Wb6ju6;  // ../RTL/cortexm0ds_logic.v(869)
  wire Wb7iu6;  // ../RTL/cortexm0ds_logic.v(401)
  wire Wb7pw6;  // ../RTL/cortexm0ds_logic.v(1426)
  wire Wb8ow6;  // ../RTL/cortexm0ds_logic.v(958)
  wire Wbeiu6;  // ../RTL/cortexm0ds_logic.v(495)
  wire Wbfow6;  // ../RTL/cortexm0ds_logic.v(1051)
  wire Wbkhu6;  // ../RTL/cortexm0ds_logic.v(136)
  wire Wbliu6;  // ../RTL/cortexm0ds_logic.v(589)
  wire Wbmax6;  // ../RTL/cortexm0ds_logic.v(1655)
  wire Wbmow6;  // ../RTL/cortexm0ds_logic.v(1145)
  wire Wbsiu6;  // ../RTL/cortexm0ds_logic.v(682)
  wire Wbthu6;  // ../RTL/cortexm0ds_logic.v(214)
  wire Wbtow6;  // ../RTL/cortexm0ds_logic.v(1239)
  wire Wbziu6;  // ../RTL/cortexm0ds_logic.v(776)
  wire Wc2qw6;  // ../RTL/cortexm0ds_logic.v(1621)
  wire Wc5ju6;  // ../RTL/cortexm0ds_logic.v(856)
  wire Wc6iu6;  // ../RTL/cortexm0ds_logic.v(388)
  wire Wc6pw6;  // ../RTL/cortexm0ds_logic.v(1413)
  wire Wc7ow6;  // ../RTL/cortexm0ds_logic.v(945)
  wire Wcdiu6;  // ../RTL/cortexm0ds_logic.v(482)
  wire Wcdpw6;  // ../RTL/cortexm0ds_logic.v(1506)
  wire Wceow6;  // ../RTL/cortexm0ds_logic.v(1038)
  wire Wckiu6;  // ../RTL/cortexm0ds_logic.v(576)
  wire Wclow6;  // ../RTL/cortexm0ds_logic.v(1132)
  wire Wcqax6;  // ../RTL/cortexm0ds_logic.v(1662)
  wire Wcriu6;  // ../RTL/cortexm0ds_logic.v(669)
  wire Wcshu6;  // ../RTL/cortexm0ds_logic.v(201)
  wire Wcsow6;  // ../RTL/cortexm0ds_logic.v(1226)
  wire Wcyiu6;  // ../RTL/cortexm0ds_logic.v(763)
  wire Wczhu6;  // ../RTL/cortexm0ds_logic.v(295)
  wire Wczow6;  // ../RTL/cortexm0ds_logic.v(1319)
  wire Wd4ju6;  // ../RTL/cortexm0ds_logic.v(843)
  wire Wd5iu6;  // ../RTL/cortexm0ds_logic.v(375)
  wire Wd5pw6;  // ../RTL/cortexm0ds_logic.v(1400)
  wire Wd6ow6;  // ../RTL/cortexm0ds_logic.v(932)
  wire Wdciu6;  // ../RTL/cortexm0ds_logic.v(469)
  wire Wdcpw6;  // ../RTL/cortexm0ds_logic.v(1493)
  wire Wddow6;  // ../RTL/cortexm0ds_logic.v(1025)
  wire Wdjhu6;  // ../RTL/cortexm0ds_logic.v(133)
  wire Wdjiu6;  // ../RTL/cortexm0ds_logic.v(563)
  wire Wdkow6;  // ../RTL/cortexm0ds_logic.v(1119)
  wire Wdmax6;  // ../RTL/cortexm0ds_logic.v(1655)
  wire Wdqiu6;  // ../RTL/cortexm0ds_logic.v(656)
  wire Wdrhu6;  // ../RTL/cortexm0ds_logic.v(188)
  wire Wdrow6;  // ../RTL/cortexm0ds_logic.v(1213)
  wire Wdxiu6;  // ../RTL/cortexm0ds_logic.v(750)
  wire Wdyhu6;  // ../RTL/cortexm0ds_logic.v(282)
  wire Wdyow6;  // ../RTL/cortexm0ds_logic.v(1306)
  wire We3ju6;  // ../RTL/cortexm0ds_logic.v(830)
  wire We4iu6;  // ../RTL/cortexm0ds_logic.v(362)
  wire We4pw6;  // ../RTL/cortexm0ds_logic.v(1387)
  wire Weaju6;  // ../RTL/cortexm0ds_logic.v(924)
  wire Webiu6;  // ../RTL/cortexm0ds_logic.v(456)
  wire Webpw6;  // ../RTL/cortexm0ds_logic.v(1480)
  wire Wecow6;  // ../RTL/cortexm0ds_logic.v(1012)
  wire Weiiu6;  // ../RTL/cortexm0ds_logic.v(550)
  wire Weipw6;  // ../RTL/cortexm0ds_logic.v(1585)
  wire Wejow6;  // ../RTL/cortexm0ds_logic.v(1106)
  wire Wepiu6;  // ../RTL/cortexm0ds_logic.v(643)
  wire Weqhu6;  // ../RTL/cortexm0ds_logic.v(175)
  wire Weqow6;  // ../RTL/cortexm0ds_logic.v(1200)
  wire Wewiu6;  // ../RTL/cortexm0ds_logic.v(737)
  wire Wexhu6;  // ../RTL/cortexm0ds_logic.v(269)
  wire Wexow6;  // ../RTL/cortexm0ds_logic.v(1293)
  wire Wf2ju6;  // ../RTL/cortexm0ds_logic.v(817)
  wire Wf3iu6;  // ../RTL/cortexm0ds_logic.v(349)
  wire Wf3pw6;  // ../RTL/cortexm0ds_logic.v(1374)
  wire Wf9ju6;  // ../RTL/cortexm0ds_logic.v(911)
  wire Wfaiu6;  // ../RTL/cortexm0ds_logic.v(443)
  wire Wfapw6;  // ../RTL/cortexm0ds_logic.v(1467)
  wire Wfbow6;  // ../RTL/cortexm0ds_logic.v(999)
  wire Wfcbx6;  // ../RTL/cortexm0ds_logic.v(1702)
  wire Wfhax6;  // ../RTL/cortexm0ds_logic.v(1646)
  wire Wfhiu6;  // ../RTL/cortexm0ds_logic.v(537)
  wire Wfihu6;  // ../RTL/cortexm0ds_logic.v(131)
  wire Wfiow6;  // ../RTL/cortexm0ds_logic.v(1093)
  wire Wfmax6;  // ../RTL/cortexm0ds_logic.v(1655)
  wire Wfoiu6;  // ../RTL/cortexm0ds_logic.v(630)
  wire Wfphu6;  // ../RTL/cortexm0ds_logic.v(162)
  wire Wfpow6;  // ../RTL/cortexm0ds_logic.v(1187)
  wire Wfspw6;  // ../RTL/cortexm0ds_logic.v(1603)
  wire Wfviu6;  // ../RTL/cortexm0ds_logic.v(724)
  wire Wfwhu6;  // ../RTL/cortexm0ds_logic.v(256)
  wire Wfwow6;  // ../RTL/cortexm0ds_logic.v(1280)
  wire Wg1ju6;  // ../RTL/cortexm0ds_logic.v(804)
  wire Wg2iu6;  // ../RTL/cortexm0ds_logic.v(336)
  wire Wg2pw6;  // ../RTL/cortexm0ds_logic.v(1361)
  wire Wg8ju6;  // ../RTL/cortexm0ds_logic.v(898)
  wire Wg9iu6;  // ../RTL/cortexm0ds_logic.v(430)
  wire Wg9pw6;  // ../RTL/cortexm0ds_logic.v(1454)
  wire Wgaow6;  // ../RTL/cortexm0ds_logic.v(986)
  wire Wggiu6;  // ../RTL/cortexm0ds_logic.v(524)
  wire Wghow6;  // ../RTL/cortexm0ds_logic.v(1080)
  wire Wgipw6;  // ../RTL/cortexm0ds_logic.v(1585)
  wire Wgniu6;  // ../RTL/cortexm0ds_logic.v(617)
  wire Wgohu6;  // ../RTL/cortexm0ds_logic.v(149)
  wire Wgoow6;  // ../RTL/cortexm0ds_logic.v(1174)
  wire Wguiu6;  // ../RTL/cortexm0ds_logic.v(711)
  wire Wgvhu6;  // ../RTL/cortexm0ds_logic.v(243)
  wire Wgvow6;  // ../RTL/cortexm0ds_logic.v(1267)
  wire Wh0ju6;  // ../RTL/cortexm0ds_logic.v(791)
  wire Wh1iu6;  // ../RTL/cortexm0ds_logic.v(323)
  wire Wh1pw6;  // ../RTL/cortexm0ds_logic.v(1348)
  wire Wh7ju6;  // ../RTL/cortexm0ds_logic.v(885)
  wire Wh8iu6;  // ../RTL/cortexm0ds_logic.v(417)
  wire Wh8pw6;  // ../RTL/cortexm0ds_logic.v(1441)
  wire Wh9ow6;  // ../RTL/cortexm0ds_logic.v(973)
  wire Whfiu6;  // ../RTL/cortexm0ds_logic.v(511)
  wire Whgow6;  // ../RTL/cortexm0ds_logic.v(1067)
  wire Whmax6;  // ../RTL/cortexm0ds_logic.v(1655)
  wire Whmiu6;  // ../RTL/cortexm0ds_logic.v(604)
  wire Whnow6;  // ../RTL/cortexm0ds_logic.v(1161)
  wire Whtiu6;  // ../RTL/cortexm0ds_logic.v(698)
  wire Whuhu6;  // ../RTL/cortexm0ds_logic.v(230)
  wire Whuow6;  // ../RTL/cortexm0ds_logic.v(1254)
  wire Wi0iu6;  // ../RTL/cortexm0ds_logic.v(310)
  wire Wi0pw6;  // ../RTL/cortexm0ds_logic.v(1335)
  wire Wi6ju6;  // ../RTL/cortexm0ds_logic.v(872)
  wire Wi7iu6;  // ../RTL/cortexm0ds_logic.v(404)
  wire Wi7pw6;  // ../RTL/cortexm0ds_logic.v(1428)
  wire Wi8ow6;  // ../RTL/cortexm0ds_logic.v(960)
  wire Widax6;  // ../RTL/cortexm0ds_logic.v(1638)
  wire Wieiu6;  // ../RTL/cortexm0ds_logic.v(498)
  wire Wifow6;  // ../RTL/cortexm0ds_logic.v(1054)
  wire Wiliu6;  // ../RTL/cortexm0ds_logic.v(591)
  wire Wimow6;  // ../RTL/cortexm0ds_logic.v(1148)
  wire Wisiu6;  // ../RTL/cortexm0ds_logic.v(685)
  wire Withu6;  // ../RTL/cortexm0ds_logic.v(217)
  wire Witow6;  // ../RTL/cortexm0ds_logic.v(1241)
  wire Wiziu6;  // ../RTL/cortexm0ds_logic.v(778)
  wire Wj5ju6;  // ../RTL/cortexm0ds_logic.v(859)
  wire Wj6iu6;  // ../RTL/cortexm0ds_logic.v(391)
  wire Wj6pw6;  // ../RTL/cortexm0ds_logic.v(1415)
  wire Wj7ow6;  // ../RTL/cortexm0ds_logic.v(947)
  wire Wjdiu6;  // ../RTL/cortexm0ds_logic.v(485)
  wire Wjdpw6;  // ../RTL/cortexm0ds_logic.v(1509)
  wire Wjeow6;  // ../RTL/cortexm0ds_logic.v(1041)
  wire Wjkiu6;  // ../RTL/cortexm0ds_logic.v(578)
  wire Wjlow6;  // ../RTL/cortexm0ds_logic.v(1135)
  wire Wjmax6;  // ../RTL/cortexm0ds_logic.v(1655)
  wire Wjriu6;  // ../RTL/cortexm0ds_logic.v(672)
  wire Wjshu6;  // ../RTL/cortexm0ds_logic.v(204)
  wire Wjsow6;  // ../RTL/cortexm0ds_logic.v(1228)
  wire Wjtpw6;  // ../RTL/cortexm0ds_logic.v(1605)
  wire Wjuax6;  // ../RTL/cortexm0ds_logic.v(1670)
  wire Wjyiu6;  // ../RTL/cortexm0ds_logic.v(765)
  wire Wjzhu6;  // ../RTL/cortexm0ds_logic.v(297)
  wire Wjzow6;  // ../RTL/cortexm0ds_logic.v(1322)
  wire Wk4ju6;  // ../RTL/cortexm0ds_logic.v(846)
  wire Wk5iu6;  // ../RTL/cortexm0ds_logic.v(378)
  wire Wk5pw6;  // ../RTL/cortexm0ds_logic.v(1402)
  wire Wk6ow6;  // ../RTL/cortexm0ds_logic.v(934)
  wire Wkciu6;  // ../RTL/cortexm0ds_logic.v(472)
  wire Wkcpw6;  // ../RTL/cortexm0ds_logic.v(1496)
  wire Wkdow6;  // ../RTL/cortexm0ds_logic.v(1028)
  wire Wkehu6;  // ../RTL/cortexm0ds_logic.v(122)
  wire Wkipw6;  // ../RTL/cortexm0ds_logic.v(1585)
  wire Wkjiu6;  // ../RTL/cortexm0ds_logic.v(565)
  wire Wkkow6;  // ../RTL/cortexm0ds_logic.v(1122)
  wire Wkmhu6;  // ../RTL/cortexm0ds_logic.v(142)
  wire Wkqiu6;  // ../RTL/cortexm0ds_logic.v(659)
  wire Wkrhu6;  // ../RTL/cortexm0ds_logic.v(191)
  wire Wkrow6;  // ../RTL/cortexm0ds_logic.v(1215)
  wire Wkxiu6;  // ../RTL/cortexm0ds_logic.v(752)
  wire Wkyhu6;  // ../RTL/cortexm0ds_logic.v(284)
  wire Wkyow6;  // ../RTL/cortexm0ds_logic.v(1309)
  wire Wl3ju6;  // ../RTL/cortexm0ds_logic.v(833)
  wire Wl4iu6;  // ../RTL/cortexm0ds_logic.v(365)
  wire Wl4pw6;  // ../RTL/cortexm0ds_logic.v(1389)
  wire Wlaju6;  // ../RTL/cortexm0ds_logic.v(927)
  wire Wlbiu6;  // ../RTL/cortexm0ds_logic.v(459)
  wire Wlbpw6;  // ../RTL/cortexm0ds_logic.v(1483)
  wire Wlcow6;  // ../RTL/cortexm0ds_logic.v(1015)
  wire Wliiu6;  // ../RTL/cortexm0ds_logic.v(552)
  wire Wljow6;  // ../RTL/cortexm0ds_logic.v(1109)
  wire Wlmax6;  // ../RTL/cortexm0ds_logic.v(1655)
  wire Wlpiu6;  // ../RTL/cortexm0ds_logic.v(646)
  wire Wlqhu6;  // ../RTL/cortexm0ds_logic.v(178)
  wire Wlqow6;  // ../RTL/cortexm0ds_logic.v(1202)
  wire Wlspw6;  // ../RTL/cortexm0ds_logic.v(1603)
  wire Wluax6;  // ../RTL/cortexm0ds_logic.v(1670)
  wire Wlwiu6;  // ../RTL/cortexm0ds_logic.v(739)
  wire Wlxhu6;  // ../RTL/cortexm0ds_logic.v(271)
  wire Wlxow6;  // ../RTL/cortexm0ds_logic.v(1296)
  wire Wm2ju6;  // ../RTL/cortexm0ds_logic.v(820)
  wire Wm3iu6;  // ../RTL/cortexm0ds_logic.v(352)
  wire Wm3pw6;  // ../RTL/cortexm0ds_logic.v(1376)
  wire Wm9ju6;  // ../RTL/cortexm0ds_logic.v(914)
  wire Wmaiu6;  // ../RTL/cortexm0ds_logic.v(446)
  wire Wmapw6;  // ../RTL/cortexm0ds_logic.v(1470)
  wire Wmbow6;  // ../RTL/cortexm0ds_logic.v(1002)
  wire Wmhiu6;  // ../RTL/cortexm0ds_logic.v(539)
  wire Wmiow6;  // ../RTL/cortexm0ds_logic.v(1096)
  wire Wmoiu6;  // ../RTL/cortexm0ds_logic.v(633)
  wire Wmphu6;  // ../RTL/cortexm0ds_logic.v(165)
  wire Wmpow6;  // ../RTL/cortexm0ds_logic.v(1189)
  wire Wmviu6;  // ../RTL/cortexm0ds_logic.v(726)
  wire Wmwhu6;  // ../RTL/cortexm0ds_logic.v(258)
  wire Wmwow6;  // ../RTL/cortexm0ds_logic.v(1283)
  wire Wmzax6;  // ../RTL/cortexm0ds_logic.v(1679)
  wire Wn1ju6;  // ../RTL/cortexm0ds_logic.v(807)
  wire Wn2iu6;  // ../RTL/cortexm0ds_logic.v(339)
  wire Wn2pw6;  // ../RTL/cortexm0ds_logic.v(1363)
  wire Wn8ju6;  // ../RTL/cortexm0ds_logic.v(901)
  wire Wn9iu6;  // ../RTL/cortexm0ds_logic.v(433)
  wire Wn9pw6;  // ../RTL/cortexm0ds_logic.v(1457)
  wire Wnaow6;  // ../RTL/cortexm0ds_logic.v(989)
  wire Wngiu6;  // ../RTL/cortexm0ds_logic.v(526)
  wire Wnhow6;  // ../RTL/cortexm0ds_logic.v(1083)
  wire Wnlhu6;  // ../RTL/cortexm0ds_logic.v(140)
  wire Wnmax6;  // ../RTL/cortexm0ds_logic.v(1655)
  wire Wnniu6;  // ../RTL/cortexm0ds_logic.v(620)
  wire Wnohu6;  // ../RTL/cortexm0ds_logic.v(152)
  wire Wnoow6;  // ../RTL/cortexm0ds_logic.v(1176)
  wire Wnuax6;  // ../RTL/cortexm0ds_logic.v(1670)
  wire Wnuiu6;  // ../RTL/cortexm0ds_logic.v(713)
  wire Wnvhu6;  // ../RTL/cortexm0ds_logic.v(245)
  wire Wnvow6;  // ../RTL/cortexm0ds_logic.v(1270)
  wire Wnxax6;  // ../RTL/cortexm0ds_logic.v(1675)
  wire Wo0ju6;  // ../RTL/cortexm0ds_logic.v(794)
  wire Wo1iu6;  // ../RTL/cortexm0ds_logic.v(326)
  wire Wo1pw6;  // ../RTL/cortexm0ds_logic.v(1350)
  wire Wo7ju6;  // ../RTL/cortexm0ds_logic.v(888)
  wire Wo8iu6;  // ../RTL/cortexm0ds_logic.v(420)
  wire Wo8pw6;  // ../RTL/cortexm0ds_logic.v(1444)
  wire Wo9ow6;  // ../RTL/cortexm0ds_logic.v(976)
  wire Wofiu6;  // ../RTL/cortexm0ds_logic.v(513)
  wire Wogow6;  // ../RTL/cortexm0ds_logic.v(1070)
  wire Woiax6;  // ../RTL/cortexm0ds_logic.v(1648)
  wire Womiu6;  // ../RTL/cortexm0ds_logic.v(607)
  wire Wonow6;  // ../RTL/cortexm0ds_logic.v(1163)
  wire Wotiu6;  // ../RTL/cortexm0ds_logic.v(700)
  wire Wouhu6;  // ../RTL/cortexm0ds_logic.v(232)
  wire Wouow6;  // ../RTL/cortexm0ds_logic.v(1257)
  wire Wp0iu6;  // ../RTL/cortexm0ds_logic.v(313)
  wire Wp0pw6;  // ../RTL/cortexm0ds_logic.v(1337)
  wire Wp6ju6;  // ../RTL/cortexm0ds_logic.v(875)
  wire Wp7iu6;  // ../RTL/cortexm0ds_logic.v(407)
  wire Wp7pw6;  // ../RTL/cortexm0ds_logic.v(1431)
  wire Wp8ow6;  // ../RTL/cortexm0ds_logic.v(963)
  wire Wpeiu6;  // ../RTL/cortexm0ds_logic.v(500)
  wire Wpfow6;  // ../RTL/cortexm0ds_logic.v(1057)
  wire Wphhu6;  // ../RTL/cortexm0ds_logic.v(129)
  wire Wpliu6;  // ../RTL/cortexm0ds_logic.v(594)
  wire Wpmax6;  // ../RTL/cortexm0ds_logic.v(1655)
  wire Wpmow6;  // ../RTL/cortexm0ds_logic.v(1150)
  wire Wpsiu6;  // ../RTL/cortexm0ds_logic.v(687)
  wire Wpthu6;  // ../RTL/cortexm0ds_logic.v(219)
  wire Wptow6;  // ../RTL/cortexm0ds_logic.v(1244)
  wire Wpuax6;  // ../RTL/cortexm0ds_logic.v(1670)
  wire Wpyax6;  // ../RTL/cortexm0ds_logic.v(1677)
  wire Wpziu6;  // ../RTL/cortexm0ds_logic.v(781)
  wire Wq5ju6;  // ../RTL/cortexm0ds_logic.v(862)
  wire Wq6iu6;  // ../RTL/cortexm0ds_logic.v(394)
  wire Wq6pw6;  // ../RTL/cortexm0ds_logic.v(1418)
  wire Wq7ow6;  // ../RTL/cortexm0ds_logic.v(950)
  wire Wq8ax6;  // ../RTL/cortexm0ds_logic.v(1629)
  wire Wqdbx6;  // ../RTL/cortexm0ds_logic.v(1704)
  wire Wqdiu6;  // ../RTL/cortexm0ds_logic.v(487)
  wire Wqdpw6;  // ../RTL/cortexm0ds_logic.v(1512)
  wire Wqeow6;  // ../RTL/cortexm0ds_logic.v(1044)
  wire Wqkiu6;  // ../RTL/cortexm0ds_logic.v(581)
  wire Wqlow6;  // ../RTL/cortexm0ds_logic.v(1137)
  wire Wqriu6;  // ../RTL/cortexm0ds_logic.v(674)
  wire Wqshu6;  // ../RTL/cortexm0ds_logic.v(206)
  wire Wqsow6;  // ../RTL/cortexm0ds_logic.v(1231)
  wire Wqyiu6;  // ../RTL/cortexm0ds_logic.v(768)
  wire Wqzhu6;  // ../RTL/cortexm0ds_logic.v(300)
  wire Wqzow6;  // ../RTL/cortexm0ds_logic.v(1324)
  wire Wqzpw6;  // ../RTL/cortexm0ds_logic.v(1616)
  wire Wr4bx6;  // ../RTL/cortexm0ds_logic.v(1688)
  wire Wr4ju6;  // ../RTL/cortexm0ds_logic.v(849)
  wire Wr5iu6;  // ../RTL/cortexm0ds_logic.v(381)
  wire Wr5pw6;  // ../RTL/cortexm0ds_logic.v(1405)
  wire Wr6ow6;  // ../RTL/cortexm0ds_logic.v(937)
  wire Wrciu6;  // ../RTL/cortexm0ds_logic.v(474)
  wire Wrcpw6;  // ../RTL/cortexm0ds_logic.v(1499)
  wire Wrdow6;  // ../RTL/cortexm0ds_logic.v(1031)
  wire Wrjiu6;  // ../RTL/cortexm0ds_logic.v(568)
  wire Wrkow6;  // ../RTL/cortexm0ds_logic.v(1124)
  wire Wrmax6;  // ../RTL/cortexm0ds_logic.v(1655)
  wire Wrqiu6;  // ../RTL/cortexm0ds_logic.v(661)
  wire Wrrhu6;  // ../RTL/cortexm0ds_logic.v(193)
  wire Wrrow6;  // ../RTL/cortexm0ds_logic.v(1218)
  wire Wruax6;  // ../RTL/cortexm0ds_logic.v(1670)
  wire Wrxiu6;  // ../RTL/cortexm0ds_logic.v(755)
  wire Wryhu6;  // ../RTL/cortexm0ds_logic.v(287)
  wire Wryow6;  // ../RTL/cortexm0ds_logic.v(1311)
  wire Ws3ju6;  // ../RTL/cortexm0ds_logic.v(836)
  wire Ws4iu6;  // ../RTL/cortexm0ds_logic.v(368)
  wire Ws4pw6;  // ../RTL/cortexm0ds_logic.v(1392)
  wire Wsaju6;  // ../RTL/cortexm0ds_logic.v(929)
  wire Wsbiu6;  // ../RTL/cortexm0ds_logic.v(461)
  wire Wsbpw6;  // ../RTL/cortexm0ds_logic.v(1486)
  wire Wscow6;  // ../RTL/cortexm0ds_logic.v(1018)
  wire Wsiiu6;  // ../RTL/cortexm0ds_logic.v(555)
  wire Wsjow6;  // ../RTL/cortexm0ds_logic.v(1111)
  wire Wskhu6;  // ../RTL/cortexm0ds_logic.v(137)
  wire Wspiu6;  // ../RTL/cortexm0ds_logic.v(648)
  wire Wsqhu6;  // ../RTL/cortexm0ds_logic.v(180)
  wire Wsqow6;  // ../RTL/cortexm0ds_logic.v(1205)
  wire Wswiu6;  // ../RTL/cortexm0ds_logic.v(742)
  wire Wsxhu6;  // ../RTL/cortexm0ds_logic.v(274)
  wire Wsxow6;  // ../RTL/cortexm0ds_logic.v(1298)
  wire Wt2ju6;  // ../RTL/cortexm0ds_logic.v(823)
  wire Wt3iu6;  // ../RTL/cortexm0ds_logic.v(355)
  wire Wt3pw6;  // ../RTL/cortexm0ds_logic.v(1379)
  wire Wt3qw6;  // ../RTL/cortexm0ds_logic.v(1624)
  wire Wt9ju6;  // ../RTL/cortexm0ds_logic.v(916)
  wire Wtaiu6;  // ../RTL/cortexm0ds_logic.v(448)
  wire Wtapw6;  // ../RTL/cortexm0ds_logic.v(1473)
  wire Wtbow6;  // ../RTL/cortexm0ds_logic.v(1005)
  wire Wthiu6;  // ../RTL/cortexm0ds_logic.v(542)
  wire Wtiow6;  // ../RTL/cortexm0ds_logic.v(1098)
  wire Wtoiu6;  // ../RTL/cortexm0ds_logic.v(635)
  wire Wtphu6;  // ../RTL/cortexm0ds_logic.v(167)
  wire Wtpow6;  // ../RTL/cortexm0ds_logic.v(1192)
  wire Wtviu6;  // ../RTL/cortexm0ds_logic.v(729)
  wire Wtwhu6;  // ../RTL/cortexm0ds_logic.v(261)
  wire Wtwow6;  // ../RTL/cortexm0ds_logic.v(1285)
  wire Wtxax6;  // ../RTL/cortexm0ds_logic.v(1675)
  wire Wu1ju6;  // ../RTL/cortexm0ds_logic.v(810)
  wire Wu2iu6;  // ../RTL/cortexm0ds_logic.v(342)
  wire Wu2pw6;  // ../RTL/cortexm0ds_logic.v(1366)
  wire Wu3bx6;  // ../RTL/cortexm0ds_logic.v(1686)
  wire Wu8ju6;  // ../RTL/cortexm0ds_logic.v(903)
  wire Wu9iu6;  // ../RTL/cortexm0ds_logic.v(435)
  wire Wu9pw6;  // ../RTL/cortexm0ds_logic.v(1460)
  wire Wuaow6;  // ../RTL/cortexm0ds_logic.v(992)
  wire Wugiu6;  // ../RTL/cortexm0ds_logic.v(529)
  wire Wuhow6;  // ../RTL/cortexm0ds_logic.v(1085)
  wire Wujhu6;  // ../RTL/cortexm0ds_logic.v(135)
  wire Wuniu6;  // ../RTL/cortexm0ds_logic.v(622)
  wire Wuohu6;  // ../RTL/cortexm0ds_logic.v(154)
  wire Wuoow6;  // ../RTL/cortexm0ds_logic.v(1179)
  wire Wuuiu6;  // ../RTL/cortexm0ds_logic.v(716)
  wire Wuvhu6;  // ../RTL/cortexm0ds_logic.v(248)
  wire Wuvow6;  // ../RTL/cortexm0ds_logic.v(1272)
  wire Wv0ju6;  // ../RTL/cortexm0ds_logic.v(797)
  wire Wv1iu6;  // ../RTL/cortexm0ds_logic.v(329)
  wire Wv1pw6;  // ../RTL/cortexm0ds_logic.v(1353)
  wire Wv7ju6;  // ../RTL/cortexm0ds_logic.v(890)
  wire Wv8iu6;  // ../RTL/cortexm0ds_logic.v(422)
  wire Wv8pw6;  // ../RTL/cortexm0ds_logic.v(1447)
  wire Wv9ow6;  // ../RTL/cortexm0ds_logic.v(979)
  wire Wvfiu6;  // ../RTL/cortexm0ds_logic.v(516)
  wire Wvgax6;  // ../RTL/cortexm0ds_logic.v(1645)
  wire Wvgow6;  // ../RTL/cortexm0ds_logic.v(1072)
  wire Wvmiu6;  // ../RTL/cortexm0ds_logic.v(609)
  wire Wvnow6;  // ../RTL/cortexm0ds_logic.v(1166)
  wire Wvtiu6;  // ../RTL/cortexm0ds_logic.v(703)
  wire Wvuhu6;  // ../RTL/cortexm0ds_logic.v(235)
  wire Wvuow6;  // ../RTL/cortexm0ds_logic.v(1259)
  wire Ww0iu6;  // ../RTL/cortexm0ds_logic.v(316)
  wire Ww0pw6;  // ../RTL/cortexm0ds_logic.v(1340)
  wire Ww6ju6;  // ../RTL/cortexm0ds_logic.v(877)
  wire Ww7iu6;  // ../RTL/cortexm0ds_logic.v(409)
  wire Ww7pw6;  // ../RTL/cortexm0ds_logic.v(1434)
  wire Ww8ow6;  // ../RTL/cortexm0ds_logic.v(966)
  wire Wweiu6;  // ../RTL/cortexm0ds_logic.v(503)
  wire Wwfow6;  // ../RTL/cortexm0ds_logic.v(1059)
  wire Wwiax6;  // ../RTL/cortexm0ds_logic.v(1648)
  wire Wwihu6;  // ../RTL/cortexm0ds_logic.v(132)
  wire Wwliu6;  // ../RTL/cortexm0ds_logic.v(596)
  wire Wwmow6;  // ../RTL/cortexm0ds_logic.v(1153)
  wire Wwsiu6;  // ../RTL/cortexm0ds_logic.v(690)
  wire Wwthu6;  // ../RTL/cortexm0ds_logic.v(222)
  wire Wwtow6;  // ../RTL/cortexm0ds_logic.v(1246)
  wire Wwziu6;  // ../RTL/cortexm0ds_logic.v(784)
  wire Wx5ju6;  // ../RTL/cortexm0ds_logic.v(864)
  wire Wx6iu6;  // ../RTL/cortexm0ds_logic.v(396)
  wire Wx6pw6;  // ../RTL/cortexm0ds_logic.v(1421)
  wire Wx7ow6;  // ../RTL/cortexm0ds_logic.v(953)
  wire Wxdiu6;  // ../RTL/cortexm0ds_logic.v(490)
  wire Wxdpw6;  // ../RTL/cortexm0ds_logic.v(1514)
  wire Wxeow6;  // ../RTL/cortexm0ds_logic.v(1046)
  wire Wxgbx6;  // ../RTL/cortexm0ds_logic.v(1710)
  wire Wxjpw6;  // ../RTL/cortexm0ds_logic.v(1587)
  wire Wxkiu6;  // ../RTL/cortexm0ds_logic.v(583)
  wire Wxlow6;  // ../RTL/cortexm0ds_logic.v(1140)
  wire Wxriu6;  // ../RTL/cortexm0ds_logic.v(677)
  wire Wxshu6;  // ../RTL/cortexm0ds_logic.v(209)
  wire Wxsow6;  // ../RTL/cortexm0ds_logic.v(1233)
  wire Wxyiu6;  // ../RTL/cortexm0ds_logic.v(771)
  wire Wxzhu6;  // ../RTL/cortexm0ds_logic.v(303)
  wire Wxzow6;  // ../RTL/cortexm0ds_logic.v(1327)
  wire Wy4ju6;  // ../RTL/cortexm0ds_logic.v(851)
  wire Wy5iu6;  // ../RTL/cortexm0ds_logic.v(383)
  wire Wy5pw6;  // ../RTL/cortexm0ds_logic.v(1408)
  wire Wy6ow6;  // ../RTL/cortexm0ds_logic.v(940)
  wire Wyciu6;  // ../RTL/cortexm0ds_logic.v(477)
  wire Wycpw6;  // ../RTL/cortexm0ds_logic.v(1501)
  wire Wydow6;  // ../RTL/cortexm0ds_logic.v(1033)
  wire Wyhhu6;  // ../RTL/cortexm0ds_logic.v(130)
  wire Wyiax6;  // ../RTL/cortexm0ds_logic.v(1649)
  wire Wyjiu6;  // ../RTL/cortexm0ds_logic.v(570)
  wire Wykow6;  // ../RTL/cortexm0ds_logic.v(1127)
  wire Wyqiu6;  // ../RTL/cortexm0ds_logic.v(664)
  wire Wyrhu6;  // ../RTL/cortexm0ds_logic.v(196)
  wire Wyrow6;  // ../RTL/cortexm0ds_logic.v(1220)
  wire Wyxiu6;  // ../RTL/cortexm0ds_logic.v(758)
  wire Wyyhu6;  // ../RTL/cortexm0ds_logic.v(290)
  wire Wyyow6;  // ../RTL/cortexm0ds_logic.v(1314)
  wire Wz3ju6;  // ../RTL/cortexm0ds_logic.v(838)
  wire Wz4iu6;  // ../RTL/cortexm0ds_logic.v(370)
  wire Wz4pw6;  // ../RTL/cortexm0ds_logic.v(1395)
  wire Wzbiu6;  // ../RTL/cortexm0ds_logic.v(464)
  wire Wzbpw6;  // ../RTL/cortexm0ds_logic.v(1488)
  wire Wzcow6;  // ../RTL/cortexm0ds_logic.v(1020)
  wire Wziiu6;  // ../RTL/cortexm0ds_logic.v(557)
  wire Wzjow6;  // ../RTL/cortexm0ds_logic.v(1114)
  wire Wzpiu6;  // ../RTL/cortexm0ds_logic.v(651)
  wire Wzqhu6;  // ../RTL/cortexm0ds_logic.v(183)
  wire Wzqow6;  // ../RTL/cortexm0ds_logic.v(1207)
  wire Wzwiu6;  // ../RTL/cortexm0ds_logic.v(745)
  wire Wzxhu6;  // ../RTL/cortexm0ds_logic.v(277)
  wire Wzxow6;  // ../RTL/cortexm0ds_logic.v(1301)
  wire X00ju6;  // ../RTL/cortexm0ds_logic.v(785)
  wire X01iu6;  // ../RTL/cortexm0ds_logic.v(317)
  wire X01pw6;  // ../RTL/cortexm0ds_logic.v(1341)
  wire X07ju6;  // ../RTL/cortexm0ds_logic.v(879)
  wire X08iu6;  // ../RTL/cortexm0ds_logic.v(411)
  wire X08pw6;  // ../RTL/cortexm0ds_logic.v(1435)
  wire X09ow6;  // ../RTL/cortexm0ds_logic.v(967)
  wire X0fiu6;  // ../RTL/cortexm0ds_logic.v(504)
  wire X0gow6;  // ../RTL/cortexm0ds_logic.v(1061)
  wire X0miu6;  // ../RTL/cortexm0ds_logic.v(598)
  wire X0now6;  // ../RTL/cortexm0ds_logic.v(1154)
  wire X0ohu6;  // ../RTL/cortexm0ds_logic.v(146)
  wire X0tiu6;  // ../RTL/cortexm0ds_logic.v(691)
  wire X0uhu6;  // ../RTL/cortexm0ds_logic.v(223)
  wire X0uow6;  // ../RTL/cortexm0ds_logic.v(1248)
  wire X10iu6;  // ../RTL/cortexm0ds_logic.v(304)
  wire X10pw6;  // ../RTL/cortexm0ds_logic.v(1328)
  wire X16ju6;  // ../RTL/cortexm0ds_logic.v(866)
  wire X17iu6;  // ../RTL/cortexm0ds_logic.v(398)
  wire X17pw6;  // ../RTL/cortexm0ds_logic.v(1422)
  wire X18ow6;  // ../RTL/cortexm0ds_logic.v(954)
  wire X1eiu6;  // ../RTL/cortexm0ds_logic.v(491)
  wire X1epw6;  // ../RTL/cortexm0ds_logic.v(1516)
  wire X1fow6;  // ../RTL/cortexm0ds_logic.v(1048)
  wire X1liu6;  // ../RTL/cortexm0ds_logic.v(585)
  wire X1max6;  // ../RTL/cortexm0ds_logic.v(1654)
  wire X1mow6;  // ../RTL/cortexm0ds_logic.v(1141)
  wire X1siu6;  // ../RTL/cortexm0ds_logic.v(678)
  wire X1thu6;  // ../RTL/cortexm0ds_logic.v(210)
  wire X1tow6;  // ../RTL/cortexm0ds_logic.v(1235)
  wire X1upw6;  // ../RTL/cortexm0ds_logic.v(1606)
  wire X1ziu6;  // ../RTL/cortexm0ds_logic.v(772)
  wire X25ju6;  // ../RTL/cortexm0ds_logic.v(853)
  wire X26iu6;  // ../RTL/cortexm0ds_logic.v(385)
  wire X26pw6;  // ../RTL/cortexm0ds_logic.v(1409)
  wire X27ow6;  // ../RTL/cortexm0ds_logic.v(941)
  wire X2diu6;  // ../RTL/cortexm0ds_logic.v(478)
  wire X2dpw6;  // ../RTL/cortexm0ds_logic.v(1503)
  wire X2eow6;  // ../RTL/cortexm0ds_logic.v(1035)
  wire X2jpw6;  // ../RTL/cortexm0ds_logic.v(1586)
  wire X2kiu6;  // ../RTL/cortexm0ds_logic.v(572)
  wire X2low6;  // ../RTL/cortexm0ds_logic.v(1128)
  wire X2riu6;  // ../RTL/cortexm0ds_logic.v(665)
  wire X2shu6;  // ../RTL/cortexm0ds_logic.v(197)
  wire X2sow6;  // ../RTL/cortexm0ds_logic.v(1222)
  wire X2yiu6;  // ../RTL/cortexm0ds_logic.v(759)
  wire X2zhu6;  // ../RTL/cortexm0ds_logic.v(291)
  wire X2zow6;  // ../RTL/cortexm0ds_logic.v(1315)
  wire X34ju6;  // ../RTL/cortexm0ds_logic.v(840)
  wire X35iu6;  // ../RTL/cortexm0ds_logic.v(372)
  wire X35pw6;  // ../RTL/cortexm0ds_logic.v(1396)
  wire X3ciu6;  // ../RTL/cortexm0ds_logic.v(465)
  wire X3cpw6;  // ../RTL/cortexm0ds_logic.v(1490)
  wire X3dow6;  // ../RTL/cortexm0ds_logic.v(1022)
  wire X3jiu6;  // ../RTL/cortexm0ds_logic.v(559)
  wire X3kow6;  // ../RTL/cortexm0ds_logic.v(1115)
  wire X3max6;  // ../RTL/cortexm0ds_logic.v(1654)
  wire X3qiu6;  // ../RTL/cortexm0ds_logic.v(652)
  wire X3rhu6;  // ../RTL/cortexm0ds_logic.v(184)
  wire X3row6;  // ../RTL/cortexm0ds_logic.v(1209)
  wire X3upw6;  // ../RTL/cortexm0ds_logic.v(1606)
  wire X3xiu6;  // ../RTL/cortexm0ds_logic.v(746)
  wire X3yhu6;  // ../RTL/cortexm0ds_logic.v(278)
  wire X3yow6;  // ../RTL/cortexm0ds_logic.v(1302)
  wire X42qw6;  // ../RTL/cortexm0ds_logic.v(1621)
  wire X43ju6;  // ../RTL/cortexm0ds_logic.v(827)
  wire X44iu6;  // ../RTL/cortexm0ds_logic.v(359)
  wire X44pw6;  // ../RTL/cortexm0ds_logic.v(1383)
  wire X4aju6;  // ../RTL/cortexm0ds_logic.v(920)
  wire X4biu6;  // ../RTL/cortexm0ds_logic.v(452)
  wire X4bpw6;  // ../RTL/cortexm0ds_logic.v(1477)
  wire X4cow6;  // ../RTL/cortexm0ds_logic.v(1009)
  wire X4iiu6;  // ../RTL/cortexm0ds_logic.v(546)
  wire X4jow6;  // ../RTL/cortexm0ds_logic.v(1102)
  wire X4jpw6;  // ../RTL/cortexm0ds_logic.v(1586)
  wire X4piu6;  // ../RTL/cortexm0ds_logic.v(639)
  wire X4qhu6;  // ../RTL/cortexm0ds_logic.v(171)
  wire X4qow6;  // ../RTL/cortexm0ds_logic.v(1196)
  wire X4wiu6;  // ../RTL/cortexm0ds_logic.v(733)
  wire X4xhu6;  // ../RTL/cortexm0ds_logic.v(265)
  wire X4xow6;  // ../RTL/cortexm0ds_logic.v(1289)
  wire X52ju6;  // ../RTL/cortexm0ds_logic.v(814)
  wire X53iu6;  // ../RTL/cortexm0ds_logic.v(346)
  wire X53pw6;  // ../RTL/cortexm0ds_logic.v(1370)
  wire X59ju6;  // ../RTL/cortexm0ds_logic.v(907)
  wire X5aiu6;  // ../RTL/cortexm0ds_logic.v(439)
  wire X5apw6;  // ../RTL/cortexm0ds_logic.v(1464)
  wire X5bax6;  // ../RTL/cortexm0ds_logic.v(1633)
  wire X5bow6;  // ../RTL/cortexm0ds_logic.v(996)
  wire X5hiu6;  // ../RTL/cortexm0ds_logic.v(533)
  wire X5ibx6;  // ../RTL/cortexm0ds_logic.v(1712)
  wire X5iow6;  // ../RTL/cortexm0ds_logic.v(1089)
  wire X5oiu6;  // ../RTL/cortexm0ds_logic.v(626)
  wire X5opw6;  // ../RTL/cortexm0ds_logic.v(1595)
  wire X5phu6;  // ../RTL/cortexm0ds_logic.v(158)
  wire X5pow6;  // ../RTL/cortexm0ds_logic.v(1183)
  wire X5upw6;  // ../RTL/cortexm0ds_logic.v(1606)
  wire X5viu6;  // ../RTL/cortexm0ds_logic.v(720)
  wire X5whu6;  // ../RTL/cortexm0ds_logic.v(252)
  wire X5wow6;  // ../RTL/cortexm0ds_logic.v(1276)
  wire X61ju6;  // ../RTL/cortexm0ds_logic.v(801)
  wire X62iu6;  // ../RTL/cortexm0ds_logic.v(333)
  wire X62pw6;  // ../RTL/cortexm0ds_logic.v(1357)
  wire X68ju6;  // ../RTL/cortexm0ds_logic.v(894)
  wire X69iu6;  // ../RTL/cortexm0ds_logic.v(426)
  wire X69pw6;  // ../RTL/cortexm0ds_logic.v(1451)
  wire X6aow6;  // ../RTL/cortexm0ds_logic.v(983)
  wire X6giu6;  // ../RTL/cortexm0ds_logic.v(520)
  wire X6how6;  // ../RTL/cortexm0ds_logic.v(1076)
  wire X6jpw6;  // ../RTL/cortexm0ds_logic.v(1586)
  wire X6mhu6;  // ../RTL/cortexm0ds_logic.v(141)
  wire X6niu6;  // ../RTL/cortexm0ds_logic.v(613)
  wire X6oow6;  // ../RTL/cortexm0ds_logic.v(1170)
  wire X6uiu6;  // ../RTL/cortexm0ds_logic.v(707)
  wire X6vhu6;  // ../RTL/cortexm0ds_logic.v(239)
  wire X6vow6;  // ../RTL/cortexm0ds_logic.v(1263)
  wire X70ju6;  // ../RTL/cortexm0ds_logic.v(788)
  wire X71iu6;  // ../RTL/cortexm0ds_logic.v(320)
  wire X71pw6;  // ../RTL/cortexm0ds_logic.v(1344)
  wire X77ju6;  // ../RTL/cortexm0ds_logic.v(881)
  wire X78iu6;  // ../RTL/cortexm0ds_logic.v(413)
  wire X78pw6;  // ../RTL/cortexm0ds_logic.v(1438)
  wire X79ow6;  // ../RTL/cortexm0ds_logic.v(970)
  wire X7abx6;  // ../RTL/cortexm0ds_logic.v(1697)
  wire X7fiu6;  // ../RTL/cortexm0ds_logic.v(507)
  wire X7gow6;  // ../RTL/cortexm0ds_logic.v(1063)
  wire X7miu6;  // ../RTL/cortexm0ds_logic.v(600)
  wire X7now6;  // ../RTL/cortexm0ds_logic.v(1157)
  wire X7spw6;  // ../RTL/cortexm0ds_logic.v(1603)
  wire X7tiu6;  // ../RTL/cortexm0ds_logic.v(694)
  wire X7uhu6;  // ../RTL/cortexm0ds_logic.v(226)
  wire X7uow6;  // ../RTL/cortexm0ds_logic.v(1250)
  wire X7ypw6;  // ../RTL/cortexm0ds_logic.v(1614)
  wire X80iu6;  // ../RTL/cortexm0ds_logic.v(307)
  wire X80pw6;  // ../RTL/cortexm0ds_logic.v(1331)
  wire X86ju6;  // ../RTL/cortexm0ds_logic.v(868)
  wire X87iu6;  // ../RTL/cortexm0ds_logic.v(400)
  wire X87pw6;  // ../RTL/cortexm0ds_logic.v(1425)
  wire X88ow6;  // ../RTL/cortexm0ds_logic.v(957)
  wire X8eiu6;  // ../RTL/cortexm0ds_logic.v(494)
  wire X8fow6;  // ../RTL/cortexm0ds_logic.v(1050)
  wire X8liu6;  // ../RTL/cortexm0ds_logic.v(587)
  wire X8mow6;  // ../RTL/cortexm0ds_logic.v(1144)
  wire X8siu6;  // ../RTL/cortexm0ds_logic.v(681)
  wire X8thu6;  // ../RTL/cortexm0ds_logic.v(213)
  wire X8tow6;  // ../RTL/cortexm0ds_logic.v(1237)
  wire X8ziu6;  // ../RTL/cortexm0ds_logic.v(775)
  wire X95ju6;  // ../RTL/cortexm0ds_logic.v(855)
  wire X96iu6;  // ../RTL/cortexm0ds_logic.v(387)
  wire X96pw6;  // ../RTL/cortexm0ds_logic.v(1412)
  wire X97ow6;  // ../RTL/cortexm0ds_logic.v(944)
  wire X9diu6;  // ../RTL/cortexm0ds_logic.v(481)
  wire X9dpw6;  // ../RTL/cortexm0ds_logic.v(1505)
  wire X9eow6;  // ../RTL/cortexm0ds_logic.v(1037)
  wire X9kiu6;  // ../RTL/cortexm0ds_logic.v(574)
  wire X9low6;  // ../RTL/cortexm0ds_logic.v(1131)
  wire X9riu6;  // ../RTL/cortexm0ds_logic.v(668)
  wire X9shu6;  // ../RTL/cortexm0ds_logic.v(200)
  wire X9sow6;  // ../RTL/cortexm0ds_logic.v(1224)
  wire X9yiu6;  // ../RTL/cortexm0ds_logic.v(762)
  wire X9zhu6;  // ../RTL/cortexm0ds_logic.v(294)
  wire X9zow6;  // ../RTL/cortexm0ds_logic.v(1318)
  wire Xa4ju6;  // ../RTL/cortexm0ds_logic.v(842)
  wire Xa5iu6;  // ../RTL/cortexm0ds_logic.v(374)
  wire Xa5pw6;  // ../RTL/cortexm0ds_logic.v(1399)
  wire Xa6ow6;  // ../RTL/cortexm0ds_logic.v(931)
  wire Xaciu6;  // ../RTL/cortexm0ds_logic.v(468)
  wire Xacpw6;  // ../RTL/cortexm0ds_logic.v(1492)
  wire Xadow6;  // ../RTL/cortexm0ds_logic.v(1024)
  wire Xaeax6;  // ../RTL/cortexm0ds_logic.v(1640)
  wire Xajbx6;  // ../RTL/cortexm0ds_logic.v(1714)
  wire Xajiu6;  // ../RTL/cortexm0ds_logic.v(561)
  wire Xakow6;  // ../RTL/cortexm0ds_logic.v(1118)
  wire Xaqax6;  // ../RTL/cortexm0ds_logic.v(1662)
  wire Xaqiu6;  // ../RTL/cortexm0ds_logic.v(655)
  wire Xarhu6;  // ../RTL/cortexm0ds_logic.v(187)
  wire Xarow6;  // ../RTL/cortexm0ds_logic.v(1211)
  wire Xaxiu6;  // ../RTL/cortexm0ds_logic.v(749)
  wire Xayhu6;  // ../RTL/cortexm0ds_logic.v(281)
  wire Xayow6;  // ../RTL/cortexm0ds_logic.v(1305)
  wire Xb3ju6;  // ../RTL/cortexm0ds_logic.v(829)
  wire Xb4iu6;  // ../RTL/cortexm0ds_logic.v(361)
  wire Xb4pw6;  // ../RTL/cortexm0ds_logic.v(1386)
  wire Xbaju6;  // ../RTL/cortexm0ds_logic.v(923)
  wire Xbbiu6;  // ../RTL/cortexm0ds_logic.v(455)
  wire Xbbpw6;  // ../RTL/cortexm0ds_logic.v(1479)
  wire Xbcow6;  // ../RTL/cortexm0ds_logic.v(1011)
  wire Xbiiu6;  // ../RTL/cortexm0ds_logic.v(548)
  wire Xbjow6;  // ../RTL/cortexm0ds_logic.v(1105)
  wire Xbopw6;  // ../RTL/cortexm0ds_logic.v(1596)
  wire Xbpiu6;  // ../RTL/cortexm0ds_logic.v(642)
  wire Xbqhu6;  // ../RTL/cortexm0ds_logic.v(174)
  wire Xbqow6;  // ../RTL/cortexm0ds_logic.v(1198)
  wire Xbwiu6;  // ../RTL/cortexm0ds_logic.v(736)
  wire Xbxhu6;  // ../RTL/cortexm0ds_logic.v(268)
  wire Xbxow6;  // ../RTL/cortexm0ds_logic.v(1292)
  wire Xc2ju6;  // ../RTL/cortexm0ds_logic.v(816)
  wire Xc3iu6;  // ../RTL/cortexm0ds_logic.v(348)
  wire Xc3pw6;  // ../RTL/cortexm0ds_logic.v(1373)
  wire Xc9ax6;  // ../RTL/cortexm0ds_logic.v(1630)
  wire Xc9ju6;  // ../RTL/cortexm0ds_logic.v(910)
  wire Xcaiu6;  // ../RTL/cortexm0ds_logic.v(442)
  wire Xcapw6;  // ../RTL/cortexm0ds_logic.v(1466)
  wire Xcbow6;  // ../RTL/cortexm0ds_logic.v(998)
  wire Xchiu6;  // ../RTL/cortexm0ds_logic.v(535)
  wire Xciow6;  // ../RTL/cortexm0ds_logic.v(1092)
  wire Xcoiu6;  // ../RTL/cortexm0ds_logic.v(629)
  wire Xcphu6;  // ../RTL/cortexm0ds_logic.v(161)
  wire Xcpow6;  // ../RTL/cortexm0ds_logic.v(1185)
  wire Xcviu6;  // ../RTL/cortexm0ds_logic.v(723)
  wire Xcwhu6;  // ../RTL/cortexm0ds_logic.v(255)
  wire Xcwow6;  // ../RTL/cortexm0ds_logic.v(1279)
  wire Xd1ju6;  // ../RTL/cortexm0ds_logic.v(803)
  wire Xd2iu6;  // ../RTL/cortexm0ds_logic.v(335)
  wire Xd2pw6;  // ../RTL/cortexm0ds_logic.v(1360)
  wire Xd8ju6;  // ../RTL/cortexm0ds_logic.v(897)
  wire Xd9iu6;  // ../RTL/cortexm0ds_logic.v(429)
  wire Xd9pw6;  // ../RTL/cortexm0ds_logic.v(1453)
  wire Xdaow6;  // ../RTL/cortexm0ds_logic.v(985)
  wire Xdcax6;  // ../RTL/cortexm0ds_logic.v(1636)
  wire Xdebx6;  // ../RTL/cortexm0ds_logic.v(1705)
  wire Xdgiu6;  // ../RTL/cortexm0ds_logic.v(522)
  wire Xdhow6;  // ../RTL/cortexm0ds_logic.v(1079)
  wire Xdniu6;  // ../RTL/cortexm0ds_logic.v(616)
  wire Xdohu6;  // ../RTL/cortexm0ds_logic.v(148)
  wire Xdoow6;  // ../RTL/cortexm0ds_logic.v(1172)
  wire Xdspw6;  // ../RTL/cortexm0ds_logic.v(1603)
  wire Xduiu6;  // ../RTL/cortexm0ds_logic.v(710)
  wire Xdvhu6;  // ../RTL/cortexm0ds_logic.v(242)
  wire Xdvow6;  // ../RTL/cortexm0ds_logic.v(1266)
  wire Xe0ju6;  // ../RTL/cortexm0ds_logic.v(790)
  wire Xe1iu6;  // ../RTL/cortexm0ds_logic.v(322)
  wire Xe1pw6;  // ../RTL/cortexm0ds_logic.v(1347)
  wire Xe7ju6;  // ../RTL/cortexm0ds_logic.v(884)
  wire Xe8iu6;  // ../RTL/cortexm0ds_logic.v(416)
  wire Xe8pw6;  // ../RTL/cortexm0ds_logic.v(1440)
  wire Xe9ow6;  // ../RTL/cortexm0ds_logic.v(972)
  wire Xefiu6;  // ../RTL/cortexm0ds_logic.v(509)
  wire Xegow6;  // ../RTL/cortexm0ds_logic.v(1066)
  wire Xemiu6;  // ../RTL/cortexm0ds_logic.v(603)
  wire Xenow6;  // ../RTL/cortexm0ds_logic.v(1159)
  wire Xetiu6;  // ../RTL/cortexm0ds_logic.v(697)
  wire Xeuhu6;  // ../RTL/cortexm0ds_logic.v(229)
  wire Xeuow6;  // ../RTL/cortexm0ds_logic.v(1253)
  wire Xf0iu6;  // ../RTL/cortexm0ds_logic.v(309)
  wire Xf0pw6;  // ../RTL/cortexm0ds_logic.v(1334)
  wire Xf6ju6;  // ../RTL/cortexm0ds_logic.v(871)
  wire Xf7iu6;  // ../RTL/cortexm0ds_logic.v(403)
  wire Xf7pw6;  // ../RTL/cortexm0ds_logic.v(1427)
  wire Xf8ax6;  // ../RTL/cortexm0ds_logic.v(1628)
  wire Xf8ow6;  // ../RTL/cortexm0ds_logic.v(959)
  wire Xfeiu6;  // ../RTL/cortexm0ds_logic.v(496)
  wire Xffow6;  // ../RTL/cortexm0ds_logic.v(1053)
  wire Xfiax6;  // ../RTL/cortexm0ds_logic.v(1648)
  wire Xfliu6;  // ../RTL/cortexm0ds_logic.v(590)
  wire Xfmow6;  // ../RTL/cortexm0ds_logic.v(1146)
  wire Xfsiu6;  // ../RTL/cortexm0ds_logic.v(684)
  wire Xfthu6;  // ../RTL/cortexm0ds_logic.v(216)
  wire Xftow6;  // ../RTL/cortexm0ds_logic.v(1240)
  wire Xfziu6;  // ../RTL/cortexm0ds_logic.v(777)
  wire Xg5ju6;  // ../RTL/cortexm0ds_logic.v(858)
  wire Xg6iu6;  // ../RTL/cortexm0ds_logic.v(390)
  wire Xg6pw6;  // ../RTL/cortexm0ds_logic.v(1414)
  wire Xg7ow6;  // ../RTL/cortexm0ds_logic.v(946)
  wire Xgdiu6;  // ../RTL/cortexm0ds_logic.v(483)
  wire Xgdpw6;  // ../RTL/cortexm0ds_logic.v(1508)
  wire Xgeow6;  // ../RTL/cortexm0ds_logic.v(1040)
  wire Xgkiu6;  // ../RTL/cortexm0ds_logic.v(577)
  wire Xglow6;  // ../RTL/cortexm0ds_logic.v(1133)
  wire Xgriu6;  // ../RTL/cortexm0ds_logic.v(671)
  wire Xgshu6;  // ../RTL/cortexm0ds_logic.v(203)
  wire Xgsow6;  // ../RTL/cortexm0ds_logic.v(1227)
  wire Xgyiu6;  // ../RTL/cortexm0ds_logic.v(764)
  wire Xgzhu6;  // ../RTL/cortexm0ds_logic.v(296)
  wire Xgzow6;  // ../RTL/cortexm0ds_logic.v(1321)
  wire Xh4ju6;  // ../RTL/cortexm0ds_logic.v(845)
  wire Xh5iu6;  // ../RTL/cortexm0ds_logic.v(377)
  wire Xh5pw6;  // ../RTL/cortexm0ds_logic.v(1401)
  wire Xh6ow6;  // ../RTL/cortexm0ds_logic.v(933)
  wire Xhciu6;  // ../RTL/cortexm0ds_logic.v(470)
  wire Xhcpw6;  // ../RTL/cortexm0ds_logic.v(1495)
  wire Xhdow6;  // ../RTL/cortexm0ds_logic.v(1027)
  wire Xhjiu6;  // ../RTL/cortexm0ds_logic.v(564)
  wire Xhkow6;  // ../RTL/cortexm0ds_logic.v(1120)
  wire Xhqiu6;  // ../RTL/cortexm0ds_logic.v(658)
  wire Xhrhu6;  // ../RTL/cortexm0ds_logic.v(190)
  wire Xhrow6;  // ../RTL/cortexm0ds_logic.v(1214)
  wire Xhtpw6;  // ../RTL/cortexm0ds_logic.v(1605)
  wire Xhuax6;  // ../RTL/cortexm0ds_logic.v(1669)
  wire Xhxiu6;  // ../RTL/cortexm0ds_logic.v(751)
  wire Xhyhu6;  // ../RTL/cortexm0ds_logic.v(283)
  wire Xhyow6;  // ../RTL/cortexm0ds_logic.v(1308)
  wire Xi3ju6;  // ../RTL/cortexm0ds_logic.v(832)
  wire Xi4iu6;  // ../RTL/cortexm0ds_logic.v(364)
  wire Xi4pw6;  // ../RTL/cortexm0ds_logic.v(1388)
  wire Xiaju6;  // ../RTL/cortexm0ds_logic.v(925)
  wire Xibiu6;  // ../RTL/cortexm0ds_logic.v(457)
  wire Xibpw6;  // ../RTL/cortexm0ds_logic.v(1482)
  wire Xicow6;  // ../RTL/cortexm0ds_logic.v(1014)
  wire Xiiiu6;  // ../RTL/cortexm0ds_logic.v(551)
  wire Xiipw6;  // ../RTL/cortexm0ds_logic.v(1585)
  wire Xijow6;  // ../RTL/cortexm0ds_logic.v(1107)
  wire Xipiu6;  // ../RTL/cortexm0ds_logic.v(645)
  wire Xiqhu6;  // ../RTL/cortexm0ds_logic.v(177)
  wire Xiqow6;  // ../RTL/cortexm0ds_logic.v(1201)
  wire Xiwiu6;  // ../RTL/cortexm0ds_logic.v(738)
  wire Xixhu6;  // ../RTL/cortexm0ds_logic.v(270)
  wire Xixow6;  // ../RTL/cortexm0ds_logic.v(1295)
  wire Xj2ju6;  // ../RTL/cortexm0ds_logic.v(819)
  wire Xj3iu6;  // ../RTL/cortexm0ds_logic.v(351)
  wire Xj3pw6;  // ../RTL/cortexm0ds_logic.v(1375)
  wire Xj9ju6;  // ../RTL/cortexm0ds_logic.v(912)
  wire Xjaiu6;  // ../RTL/cortexm0ds_logic.v(444)
  wire Xjapw6;  // ../RTL/cortexm0ds_logic.v(1469)
  wire Xjbow6;  // ../RTL/cortexm0ds_logic.v(1001)
  wire Xjhiu6;  // ../RTL/cortexm0ds_logic.v(538)
  wire Xjiow6;  // ../RTL/cortexm0ds_logic.v(1094)
  wire Xjoiu6;  // ../RTL/cortexm0ds_logic.v(632)
  wire Xjphu6;  // ../RTL/cortexm0ds_logic.v(164)
  wire Xjpow6;  // ../RTL/cortexm0ds_logic.v(1188)
  wire Xjviu6;  // ../RTL/cortexm0ds_logic.v(725)
  wire Xjwhu6;  // ../RTL/cortexm0ds_logic.v(257)
  wire Xjwow6;  // ../RTL/cortexm0ds_logic.v(1282)
  wire Xk1ju6;  // ../RTL/cortexm0ds_logic.v(806)
  wire Xk2iu6;  // ../RTL/cortexm0ds_logic.v(338)
  wire Xk2pw6;  // ../RTL/cortexm0ds_logic.v(1362)
  wire Xk8ju6;  // ../RTL/cortexm0ds_logic.v(899)
  wire Xk9iu6;  // ../RTL/cortexm0ds_logic.v(431)
  wire Xk9pw6;  // ../RTL/cortexm0ds_logic.v(1456)
  wire Xkaow6;  // ../RTL/cortexm0ds_logic.v(988)
  wire Xkgiu6;  // ../RTL/cortexm0ds_logic.v(525)
  wire Xkhow6;  // ../RTL/cortexm0ds_logic.v(1081)
  wire Xkniu6;  // ../RTL/cortexm0ds_logic.v(619)
  wire Xkohu6;  // ../RTL/cortexm0ds_logic.v(151)
  wire Xkoow6;  // ../RTL/cortexm0ds_logic.v(1175)
  wire Xkqpw6;  // ../RTL/cortexm0ds_logic.v(1600)
  wire Xkuiu6;  // ../RTL/cortexm0ds_logic.v(712)
  wire Xkvhu6;  // ../RTL/cortexm0ds_logic.v(244)
  wire Xkvow6;  // ../RTL/cortexm0ds_logic.v(1269)
  wire Xl0ju6;  // ../RTL/cortexm0ds_logic.v(793)
  wire Xl1iu6;  // ../RTL/cortexm0ds_logic.v(325)
  wire Xl1pw6;  // ../RTL/cortexm0ds_logic.v(1349)
  wire Xl7ju6;  // ../RTL/cortexm0ds_logic.v(886)
  wire Xl8iu6;  // ../RTL/cortexm0ds_logic.v(418)
  wire Xl8pw6;  // ../RTL/cortexm0ds_logic.v(1443)
  wire Xl9ow6;  // ../RTL/cortexm0ds_logic.v(975)
  wire Xlfiu6;  // ../RTL/cortexm0ds_logic.v(512)
  wire Xlgow6;  // ../RTL/cortexm0ds_logic.v(1068)
  wire Xlmiu6;  // ../RTL/cortexm0ds_logic.v(606)
  wire Xlnow6;  // ../RTL/cortexm0ds_logic.v(1162)
  wire Xltiu6;  // ../RTL/cortexm0ds_logic.v(699)
  wire Xluhu6;  // ../RTL/cortexm0ds_logic.v(231)
  wire Xluow6;  // ../RTL/cortexm0ds_logic.v(1256)
  wire Xm0iu6;  // ../RTL/cortexm0ds_logic.v(312)
  wire Xm0pw6;  // ../RTL/cortexm0ds_logic.v(1336)
  wire Xm6ju6;  // ../RTL/cortexm0ds_logic.v(873)
  wire Xm7iu6;  // ../RTL/cortexm0ds_logic.v(405)
  wire Xm7pw6;  // ../RTL/cortexm0ds_logic.v(1430)
  wire Xm8ow6;  // ../RTL/cortexm0ds_logic.v(962)
  wire Xmeiu6;  // ../RTL/cortexm0ds_logic.v(499)
  wire Xmfow6;  // ../RTL/cortexm0ds_logic.v(1055)
  wire Xmliu6;  // ../RTL/cortexm0ds_logic.v(593)
  wire Xmmow6;  // ../RTL/cortexm0ds_logic.v(1149)
  wire Xmsiu6;  // ../RTL/cortexm0ds_logic.v(686)
  wire Xmthu6;  // ../RTL/cortexm0ds_logic.v(218)
  wire Xmtow6;  // ../RTL/cortexm0ds_logic.v(1243)
  wire Xmziu6;  // ../RTL/cortexm0ds_logic.v(780)
  wire Xn5ju6;  // ../RTL/cortexm0ds_logic.v(860)
  wire Xn6iu6;  // ../RTL/cortexm0ds_logic.v(392)
  wire Xn6pw6;  // ../RTL/cortexm0ds_logic.v(1417)
  wire Xn7ax6;  // ../RTL/cortexm0ds_logic.v(1627)
  wire Xn7ow6;  // ../RTL/cortexm0ds_logic.v(949)
  wire Xnbax6;  // ../RTL/cortexm0ds_logic.v(1634)
  wire Xndiu6;  // ../RTL/cortexm0ds_logic.v(486)
  wire Xndpw6;  // ../RTL/cortexm0ds_logic.v(1510)
  wire Xneow6;  // ../RTL/cortexm0ds_logic.v(1042)
  wire Xnkiu6;  // ../RTL/cortexm0ds_logic.v(580)
  wire Xnlow6;  // ../RTL/cortexm0ds_logic.v(1136)
  wire Xnriu6;  // ../RTL/cortexm0ds_logic.v(673)
  wire Xnshu6;  // ../RTL/cortexm0ds_logic.v(205)
  wire Xnsow6;  // ../RTL/cortexm0ds_logic.v(1230)
  wire Xnyiu6;  // ../RTL/cortexm0ds_logic.v(767)
  wire Xnzhu6;  // ../RTL/cortexm0ds_logic.v(299)
  wire Xnzow6;  // ../RTL/cortexm0ds_logic.v(1323)
  wire Xo1bx6;  // ../RTL/cortexm0ds_logic.v(1682)
  wire Xo4ju6;  // ../RTL/cortexm0ds_logic.v(847)
  wire Xo5iu6;  // ../RTL/cortexm0ds_logic.v(379)
  wire Xo5pw6;  // ../RTL/cortexm0ds_logic.v(1404)
  wire Xo6ow6;  // ../RTL/cortexm0ds_logic.v(936)
  wire Xociu6;  // ../RTL/cortexm0ds_logic.v(473)
  wire Xocpw6;  // ../RTL/cortexm0ds_logic.v(1497)
  wire Xodow6;  // ../RTL/cortexm0ds_logic.v(1029)
  wire Xojiu6;  // ../RTL/cortexm0ds_logic.v(567)
  wire Xokow6;  // ../RTL/cortexm0ds_logic.v(1123)
  wire Xoqiu6;  // ../RTL/cortexm0ds_logic.v(660)
  wire Xorhu6;  // ../RTL/cortexm0ds_logic.v(192)
  wire Xorow6;  // ../RTL/cortexm0ds_logic.v(1217)
  wire Xoxiu6;  // ../RTL/cortexm0ds_logic.v(754)
  wire Xoyhu6;  // ../RTL/cortexm0ds_logic.v(286)
  wire Xoyow6;  // ../RTL/cortexm0ds_logic.v(1310)
  wire Xozax6;  // ../RTL/cortexm0ds_logic.v(1679)
  wire Xozpw6;  // ../RTL/cortexm0ds_logic.v(1616)
  wire Xp3ju6;  // ../RTL/cortexm0ds_logic.v(834)
  wire Xp4iu6;  // ../RTL/cortexm0ds_logic.v(366)
  wire Xp4pw6;  // ../RTL/cortexm0ds_logic.v(1391)
  wire Xpaju6;  // ../RTL/cortexm0ds_logic.v(928)
  wire Xpbiu6;  // ../RTL/cortexm0ds_logic.v(460)
  wire Xpbpw6;  // ../RTL/cortexm0ds_logic.v(1484)
  wire Xpcow6;  // ../RTL/cortexm0ds_logic.v(1016)
  wire Xpeax6;  // ../RTL/cortexm0ds_logic.v(1640)
  wire Xpiiu6;  // ../RTL/cortexm0ds_logic.v(554)
  wire Xpjow6;  // ../RTL/cortexm0ds_logic.v(1110)
  wire Xppiu6;  // ../RTL/cortexm0ds_logic.v(647)
  wire Xpqhu6;  // ../RTL/cortexm0ds_logic.v(179)
  wire Xpqow6;  // ../RTL/cortexm0ds_logic.v(1204)
  wire Xpwiu6;  // ../RTL/cortexm0ds_logic.v(741)
  wire Xpxax6;  // ../RTL/cortexm0ds_logic.v(1675)
  wire Xpxhu6;  // ../RTL/cortexm0ds_logic.v(273)
  wire Xpxow6;  // ../RTL/cortexm0ds_logic.v(1297)
  wire Xq2bx6;  // ../RTL/cortexm0ds_logic.v(1684)
  wire Xq2ju6;  // ../RTL/cortexm0ds_logic.v(821)
  wire Xq3iu6;  // ../RTL/cortexm0ds_logic.v(353)
  wire Xq3pw6;  // ../RTL/cortexm0ds_logic.v(1378)
  wire Xq9ju6;  // ../RTL/cortexm0ds_logic.v(915)
  wire Xqaiu6;  // ../RTL/cortexm0ds_logic.v(447)
  wire Xqapw6;  // ../RTL/cortexm0ds_logic.v(1471)
  wire Xqbow6;  // ../RTL/cortexm0ds_logic.v(1003)
  wire Xqcax6;  // ../RTL/cortexm0ds_logic.v(1637)
  wire Xqhiu6;  // ../RTL/cortexm0ds_logic.v(541)
  wire Xqiow6;  // ../RTL/cortexm0ds_logic.v(1097)
  wire Xqoiu6;  // ../RTL/cortexm0ds_logic.v(634)
  wire Xqphu6;  // ../RTL/cortexm0ds_logic.v(166)
  wire Xqpow6;  // ../RTL/cortexm0ds_logic.v(1191)
  wire Xqviu6;  // ../RTL/cortexm0ds_logic.v(728)
  wire Xqwhu6;  // ../RTL/cortexm0ds_logic.v(260)
  wire Xqwow6;  // ../RTL/cortexm0ds_logic.v(1284)
  wire Xr1ju6;  // ../RTL/cortexm0ds_logic.v(808)
  wire Xr2iu6;  // ../RTL/cortexm0ds_logic.v(340)
  wire Xr2pw6;  // ../RTL/cortexm0ds_logic.v(1365)
  wire Xr8ju6;  // ../RTL/cortexm0ds_logic.v(902)
  wire Xr9ax6;  // ../RTL/cortexm0ds_logic.v(1631)
  wire Xr9iu6;  // ../RTL/cortexm0ds_logic.v(434)
  wire Xr9pw6;  // ../RTL/cortexm0ds_logic.v(1458)
  wire Xraow6;  // ../RTL/cortexm0ds_logic.v(990)
  wire Xrgiu6;  // ../RTL/cortexm0ds_logic.v(528)
  wire Xrhow6;  // ../RTL/cortexm0ds_logic.v(1084)
  wire Xrniu6;  // ../RTL/cortexm0ds_logic.v(621)
  wire Xrohu6;  // ../RTL/cortexm0ds_logic.v(153)
  wire Xroow6;  // ../RTL/cortexm0ds_logic.v(1178)
  wire Xruiu6;  // ../RTL/cortexm0ds_logic.v(715)
  wire Xrvhu6;  // ../RTL/cortexm0ds_logic.v(247)
  wire Xrvow6;  // ../RTL/cortexm0ds_logic.v(1271)
  wire Xrxax6;  // ../RTL/cortexm0ds_logic.v(1675)
  wire Xs0ju6;  // ../RTL/cortexm0ds_logic.v(795)
  wire Xs1iu6;  // ../RTL/cortexm0ds_logic.v(327)
  wire Xs1pw6;  // ../RTL/cortexm0ds_logic.v(1352)
  wire Xs7ju6;  // ../RTL/cortexm0ds_logic.v(889)
  wire Xs8iu6;  // ../RTL/cortexm0ds_logic.v(421)
  wire Xs8pw6;  // ../RTL/cortexm0ds_logic.v(1445)
  wire Xs9ow6;  // ../RTL/cortexm0ds_logic.v(977)
  wire Xsfiu6;  // ../RTL/cortexm0ds_logic.v(515)
  wire Xsgow6;  // ../RTL/cortexm0ds_logic.v(1071)
  wire Xsmiu6;  // ../RTL/cortexm0ds_logic.v(608)
  wire Xsnow6;  // ../RTL/cortexm0ds_logic.v(1165)
  wire Xstiu6;  // ../RTL/cortexm0ds_logic.v(702)
  wire Xsuhu6;  // ../RTL/cortexm0ds_logic.v(234)
  wire Xsuow6;  // ../RTL/cortexm0ds_logic.v(1258)
  wire Xt0iu6;  // ../RTL/cortexm0ds_logic.v(314)
  wire Xt0pw6;  // ../RTL/cortexm0ds_logic.v(1339)
  wire Xt6ju6;  // ../RTL/cortexm0ds_logic.v(876)
  wire Xt7iu6;  // ../RTL/cortexm0ds_logic.v(408)
  wire Xt7pw6;  // ../RTL/cortexm0ds_logic.v(1432)
  wire Xt8ow6;  // ../RTL/cortexm0ds_logic.v(964)
  wire Xteiu6;  // ../RTL/cortexm0ds_logic.v(502)
  wire Xtfow6;  // ../RTL/cortexm0ds_logic.v(1058)
  wire Xtliu6;  // ../RTL/cortexm0ds_logic.v(595)
  wire Xtmow6;  // ../RTL/cortexm0ds_logic.v(1152)
  wire Xtsiu6;  // ../RTL/cortexm0ds_logic.v(689)
  wire Xtthu6;  // ../RTL/cortexm0ds_logic.v(221)
  wire Xttow6;  // ../RTL/cortexm0ds_logic.v(1245)
  wire Xttpw6;  // ../RTL/cortexm0ds_logic.v(1606)
  wire Xtziu6;  // ../RTL/cortexm0ds_logic.v(782)
  wire Xu2qw6;  // ../RTL/cortexm0ds_logic.v(1622)
  wire Xu5ju6;  // ../RTL/cortexm0ds_logic.v(863)
  wire Xu6iu6;  // ../RTL/cortexm0ds_logic.v(395)
  wire Xu6pw6;  // ../RTL/cortexm0ds_logic.v(1419)
  wire Xu7ow6;  // ../RTL/cortexm0ds_logic.v(951)
  wire Xudiu6;  // ../RTL/cortexm0ds_logic.v(489)
  wire Xudpw6;  // ../RTL/cortexm0ds_logic.v(1513)
  wire Xueow6;  // ../RTL/cortexm0ds_logic.v(1045)
  wire Xuiax6;  // ../RTL/cortexm0ds_logic.v(1648)
  wire Xukiu6;  // ../RTL/cortexm0ds_logic.v(582)
  wire Xulow6;  // ../RTL/cortexm0ds_logic.v(1139)
  wire Xuriu6;  // ../RTL/cortexm0ds_logic.v(676)
  wire Xushu6;  // ../RTL/cortexm0ds_logic.v(208)
  wire Xusow6;  // ../RTL/cortexm0ds_logic.v(1232)
  wire Xuyiu6;  // ../RTL/cortexm0ds_logic.v(769)
  wire Xuzhu6;  // ../RTL/cortexm0ds_logic.v(301)
  wire Xuzow6;  // ../RTL/cortexm0ds_logic.v(1326)
  wire Xv4ju6;  // ../RTL/cortexm0ds_logic.v(850)
  wire Xv5iu6;  // ../RTL/cortexm0ds_logic.v(382)
  wire Xv5pw6;  // ../RTL/cortexm0ds_logic.v(1406)
  wire Xv6ow6;  // ../RTL/cortexm0ds_logic.v(938)
  wire Xv8bx6;  // ../RTL/cortexm0ds_logic.v(1695)
  wire Xvciu6;  // ../RTL/cortexm0ds_logic.v(476)
  wire Xvcpw6;  // ../RTL/cortexm0ds_logic.v(1500)
  wire Xvdow6;  // ../RTL/cortexm0ds_logic.v(1032)
  wire Xvjiu6;  // ../RTL/cortexm0ds_logic.v(569)
  wire Xvkow6;  // ../RTL/cortexm0ds_logic.v(1126)
  wire Xvlax6;  // ../RTL/cortexm0ds_logic.v(1654)
  wire Xvqiu6;  // ../RTL/cortexm0ds_logic.v(663)
  wire Xvqpw6;  // ../RTL/cortexm0ds_logic.v(1600)
  wire Xvrhu6;  // ../RTL/cortexm0ds_logic.v(195)
  wire Xvrow6;  // ../RTL/cortexm0ds_logic.v(1219)
  wire Xvtpw6;  // ../RTL/cortexm0ds_logic.v(1606)
  wire Xvxiu6;  // ../RTL/cortexm0ds_logic.v(756)
  wire Xvyhu6;  // ../RTL/cortexm0ds_logic.v(288)
  wire Xvyow6;  // ../RTL/cortexm0ds_logic.v(1313)
  wire Xw3ju6;  // ../RTL/cortexm0ds_logic.v(837)
  wire Xw4iu6;  // ../RTL/cortexm0ds_logic.v(369)
  wire Xw4pw6;  // ../RTL/cortexm0ds_logic.v(1393)
  wire Xwaax6;  // ../RTL/cortexm0ds_logic.v(1633)
  wire Xwbiu6;  // ../RTL/cortexm0ds_logic.v(463)
  wire Xwbpw6;  // ../RTL/cortexm0ds_logic.v(1487)
  wire Xwcow6;  // ../RTL/cortexm0ds_logic.v(1019)
  wire Xwiiu6;  // ../RTL/cortexm0ds_logic.v(556)
  wire Xwjow6;  // ../RTL/cortexm0ds_logic.v(1113)
  wire Xwpiu6;  // ../RTL/cortexm0ds_logic.v(650)
  wire Xwqhu6;  // ../RTL/cortexm0ds_logic.v(182)
  wire Xwqow6;  // ../RTL/cortexm0ds_logic.v(1206)
  wire Xwwiu6;  // ../RTL/cortexm0ds_logic.v(743)
  wire Xwxhu6;  // ../RTL/cortexm0ds_logic.v(275)
  wire Xwxow6;  // ../RTL/cortexm0ds_logic.v(1300)
  wire Xx2ju6;  // ../RTL/cortexm0ds_logic.v(824)
  wire Xx3iu6;  // ../RTL/cortexm0ds_logic.v(356)
  wire Xx3pw6;  // ../RTL/cortexm0ds_logic.v(1380)
  wire Xx6bx6;  // ../RTL/cortexm0ds_logic.v(1691)
  wire Xx9ju6;  // ../RTL/cortexm0ds_logic.v(918)
  wire Xxaiu6;  // ../RTL/cortexm0ds_logic.v(450)
  wire Xxapw6;  // ../RTL/cortexm0ds_logic.v(1474)
  wire Xxbow6;  // ../RTL/cortexm0ds_logic.v(1006)
  wire Xxhiu6;  // ../RTL/cortexm0ds_logic.v(543)
  wire Xxiow6;  // ../RTL/cortexm0ds_logic.v(1100)
  wire Xxlax6;  // ../RTL/cortexm0ds_logic.v(1654)
  wire Xxoiu6;  // ../RTL/cortexm0ds_logic.v(637)
  wire Xxphu6;  // ../RTL/cortexm0ds_logic.v(169)
  wire Xxpow6;  // ../RTL/cortexm0ds_logic.v(1193)
  wire Xxqpw6;  // ../RTL/cortexm0ds_logic.v(1600)
  wire Xxtpw6;  // ../RTL/cortexm0ds_logic.v(1606)
  wire Xxupw6;  // ../RTL/cortexm0ds_logic.v(1608)
  wire Xxviu6;  // ../RTL/cortexm0ds_logic.v(730)
  wire Xxwhu6;  // ../RTL/cortexm0ds_logic.v(262)
  wire Xxwow6;  // ../RTL/cortexm0ds_logic.v(1287)
  wire Xy1ju6;  // ../RTL/cortexm0ds_logic.v(811)
  wire Xy2iu6;  // ../RTL/cortexm0ds_logic.v(343)
  wire Xy2pw6;  // ../RTL/cortexm0ds_logic.v(1367)
  wire Xy8ju6;  // ../RTL/cortexm0ds_logic.v(905)
  wire Xy9iu6;  // ../RTL/cortexm0ds_logic.v(437)
  wire Xy9pw6;  // ../RTL/cortexm0ds_logic.v(1461)
  wire Xyaow6;  // ../RTL/cortexm0ds_logic.v(993)
  wire Xygiu6;  // ../RTL/cortexm0ds_logic.v(530)
  wire Xyhow6;  // ../RTL/cortexm0ds_logic.v(1087)
  wire Xyniu6;  // ../RTL/cortexm0ds_logic.v(624)
  wire Xyohu6;  // ../RTL/cortexm0ds_logic.v(156)
  wire Xyoow6;  // ../RTL/cortexm0ds_logic.v(1180)
  wire Xyuiu6;  // ../RTL/cortexm0ds_logic.v(717)
  wire Xyvhu6;  // ../RTL/cortexm0ds_logic.v(249)
  wire Xyvow6;  // ../RTL/cortexm0ds_logic.v(1274)
  wire Xz0ju6;  // ../RTL/cortexm0ds_logic.v(798)
  wire Xz1iu6;  // ../RTL/cortexm0ds_logic.v(330)
  wire Xz1pw6;  // ../RTL/cortexm0ds_logic.v(1354)
  wire Xz7ju6;  // ../RTL/cortexm0ds_logic.v(892)
  wire Xz8iu6;  // ../RTL/cortexm0ds_logic.v(424)
  wire Xz8pw6;  // ../RTL/cortexm0ds_logic.v(1448)
  wire Xz9ow6;  // ../RTL/cortexm0ds_logic.v(980)
  wire Xzfiu6;  // ../RTL/cortexm0ds_logic.v(517)
  wire Xzgow6;  // ../RTL/cortexm0ds_logic.v(1074)
  wire Xzlax6;  // ../RTL/cortexm0ds_logic.v(1654)
  wire Xzmiu6;  // ../RTL/cortexm0ds_logic.v(611)
  wire Xznow6;  // ../RTL/cortexm0ds_logic.v(1167)
  wire Xztiu6;  // ../RTL/cortexm0ds_logic.v(704)
  wire Xztpw6;  // ../RTL/cortexm0ds_logic.v(1606)
  wire Xzuhu6;  // ../RTL/cortexm0ds_logic.v(236)
  wire Xzuow6;  // ../RTL/cortexm0ds_logic.v(1261)
  wire Y04ju6;  // ../RTL/cortexm0ds_logic.v(839)
  wire Y05iu6;  // ../RTL/cortexm0ds_logic.v(371)
  wire Y05pw6;  // ../RTL/cortexm0ds_logic.v(1395)
  wire Y0ciu6;  // ../RTL/cortexm0ds_logic.v(464)
  wire Y0cpw6;  // ../RTL/cortexm0ds_logic.v(1489)
  wire Y0dow6;  // ../RTL/cortexm0ds_logic.v(1021)
  wire Y0gbx6;  // ../RTL/cortexm0ds_logic.v(1708)
  wire Y0jiu6;  // ../RTL/cortexm0ds_logic.v(558)
  wire Y0kow6;  // ../RTL/cortexm0ds_logic.v(1114)
  wire Y0qiu6;  // ../RTL/cortexm0ds_logic.v(651)
  wire Y0rhu6;  // ../RTL/cortexm0ds_logic.v(183)
  wire Y0row6;  // ../RTL/cortexm0ds_logic.v(1208)
  wire Y0xiu6;  // ../RTL/cortexm0ds_logic.v(745)
  wire Y0yhu6;  // ../RTL/cortexm0ds_logic.v(277)
  wire Y0yow6;  // ../RTL/cortexm0ds_logic.v(1301)
  wire Y13ju6;  // ../RTL/cortexm0ds_logic.v(826)
  wire Y14iu6;  // ../RTL/cortexm0ds_logic.v(358)
  wire Y14pw6;  // ../RTL/cortexm0ds_logic.v(1382)
  wire Y1aju6;  // ../RTL/cortexm0ds_logic.v(919)
  wire Y1biu6;  // ../RTL/cortexm0ds_logic.v(451)
  wire Y1bpw6;  // ../RTL/cortexm0ds_logic.v(1476)
  wire Y1cow6;  // ../RTL/cortexm0ds_logic.v(1008)
  wire Y1iiu6;  // ../RTL/cortexm0ds_logic.v(545)
  wire Y1jow6;  // ../RTL/cortexm0ds_logic.v(1101)
  wire Y1piu6;  // ../RTL/cortexm0ds_logic.v(638)
  wire Y1qhu6;  // ../RTL/cortexm0ds_logic.v(170)
  wire Y1qow6;  // ../RTL/cortexm0ds_logic.v(1195)
  wire Y1wiu6;  // ../RTL/cortexm0ds_logic.v(732)
  wire Y1xhu6;  // ../RTL/cortexm0ds_logic.v(264)
  wire Y1xow6;  // ../RTL/cortexm0ds_logic.v(1288)
  wire Y22ju6;  // ../RTL/cortexm0ds_logic.v(813)
  wire Y23iu6;  // ../RTL/cortexm0ds_logic.v(345)
  wire Y23pw6;  // ../RTL/cortexm0ds_logic.v(1369)
  wire Y29ju6;  // ../RTL/cortexm0ds_logic.v(906)
  wire Y2aiu6;  // ../RTL/cortexm0ds_logic.v(438)
  wire Y2apw6;  // ../RTL/cortexm0ds_logic.v(1463)
  wire Y2bow6;  // ../RTL/cortexm0ds_logic.v(995)
  wire Y2fax6;  // ../RTL/cortexm0ds_logic.v(1641)
  wire Y2hiu6;  // ../RTL/cortexm0ds_logic.v(532)
  wire Y2iow6;  // ../RTL/cortexm0ds_logic.v(1088)
  wire Y2oiu6;  // ../RTL/cortexm0ds_logic.v(625)
  wire Y2phu6;  // ../RTL/cortexm0ds_logic.v(157)
  wire Y2pow6;  // ../RTL/cortexm0ds_logic.v(1182)
  wire Y2viu6;  // ../RTL/cortexm0ds_logic.v(719)
  wire Y2whu6;  // ../RTL/cortexm0ds_logic.v(251)
  wire Y2wow6;  // ../RTL/cortexm0ds_logic.v(1275)
  wire Y31ju6;  // ../RTL/cortexm0ds_logic.v(800)
  wire Y32iu6;  // ../RTL/cortexm0ds_logic.v(332)
  wire Y32pw6;  // ../RTL/cortexm0ds_logic.v(1356)
  wire Y38ju6;  // ../RTL/cortexm0ds_logic.v(893)
  wire Y39iu6;  // ../RTL/cortexm0ds_logic.v(425)
  wire Y39pw6;  // ../RTL/cortexm0ds_logic.v(1450)
  wire Y3aow6;  // ../RTL/cortexm0ds_logic.v(982)
  wire Y3giu6;  // ../RTL/cortexm0ds_logic.v(519)
  wire Y3how6;  // ../RTL/cortexm0ds_logic.v(1075)
  wire Y3niu6;  // ../RTL/cortexm0ds_logic.v(612)
  wire Y3oow6;  // ../RTL/cortexm0ds_logic.v(1169)
  wire Y3uiu6;  // ../RTL/cortexm0ds_logic.v(706)
  wire Y3vhu6;  // ../RTL/cortexm0ds_logic.v(238)
  wire Y3vow6;  // ../RTL/cortexm0ds_logic.v(1262)
  wire Y40ju6;  // ../RTL/cortexm0ds_logic.v(787)
  wire Y41iu6;  // ../RTL/cortexm0ds_logic.v(319)
  wire Y41pw6;  // ../RTL/cortexm0ds_logic.v(1343)
  wire Y47ju6;  // ../RTL/cortexm0ds_logic.v(880)
  wire Y48iu6;  // ../RTL/cortexm0ds_logic.v(412)
  wire Y48pw6;  // ../RTL/cortexm0ds_logic.v(1437)
  wire Y49ow6;  // ../RTL/cortexm0ds_logic.v(969)
  wire Y4fiu6;  // ../RTL/cortexm0ds_logic.v(506)
  wire Y4gow6;  // ../RTL/cortexm0ds_logic.v(1062)
  wire Y4miu6;  // ../RTL/cortexm0ds_logic.v(599)
  wire Y4now6;  // ../RTL/cortexm0ds_logic.v(1156)
  wire Y4tiu6;  // ../RTL/cortexm0ds_logic.v(693)
  wire Y4uhu6;  // ../RTL/cortexm0ds_logic.v(225)
  wire Y4uow6;  // ../RTL/cortexm0ds_logic.v(1249)
  wire Y50iu6;  // ../RTL/cortexm0ds_logic.v(306)
  wire Y50pw6;  // ../RTL/cortexm0ds_logic.v(1330)
  wire Y56ju6;  // ../RTL/cortexm0ds_logic.v(867)
  wire Y57iu6;  // ../RTL/cortexm0ds_logic.v(399)
  wire Y57pw6;  // ../RTL/cortexm0ds_logic.v(1424)
  wire Y58ow6;  // ../RTL/cortexm0ds_logic.v(956)
  wire Y5dax6;  // ../RTL/cortexm0ds_logic.v(1637)
  wire Y5eiu6;  // ../RTL/cortexm0ds_logic.v(493)
  wire Y5fow6;  // ../RTL/cortexm0ds_logic.v(1049)
  wire Y5lhu6;  // ../RTL/cortexm0ds_logic.v(138)
  wire Y5liu6;  // ../RTL/cortexm0ds_logic.v(586)
  wire Y5mow6;  // ../RTL/cortexm0ds_logic.v(1143)
  wire Y5siu6;  // ../RTL/cortexm0ds_logic.v(680)
  wire Y5spw6;  // ../RTL/cortexm0ds_logic.v(1603)
  wire Y5thu6;  // ../RTL/cortexm0ds_logic.v(212)
  wire Y5tow6;  // ../RTL/cortexm0ds_logic.v(1236)
  wire Y5ziu6;  // ../RTL/cortexm0ds_logic.v(774)
  wire Y65ju6;  // ../RTL/cortexm0ds_logic.v(854)
  wire Y66iu6;  // ../RTL/cortexm0ds_logic.v(386)
  wire Y66pw6;  // ../RTL/cortexm0ds_logic.v(1411)
  wire Y67ow6;  // ../RTL/cortexm0ds_logic.v(943)
  wire Y6diu6;  // ../RTL/cortexm0ds_logic.v(480)
  wire Y6dpw6;  // ../RTL/cortexm0ds_logic.v(1504)
  wire Y6eow6;  // ../RTL/cortexm0ds_logic.v(1036)
  wire Y6kiu6;  // ../RTL/cortexm0ds_logic.v(573)
  wire Y6low6;  // ../RTL/cortexm0ds_logic.v(1130)
  wire Y6riu6;  // ../RTL/cortexm0ds_logic.v(667)
  wire Y6shu6;  // ../RTL/cortexm0ds_logic.v(199)
  wire Y6sow6;  // ../RTL/cortexm0ds_logic.v(1223)
  wire Y6yiu6;  // ../RTL/cortexm0ds_logic.v(761)
  wire Y6zhu6;  // ../RTL/cortexm0ds_logic.v(293)
  wire Y6zow6;  // ../RTL/cortexm0ds_logic.v(1317)
  wire Y72bx6;  // ../RTL/cortexm0ds_logic.v(1683)
  wire Y74ju6;  // ../RTL/cortexm0ds_logic.v(841)
  wire Y75iu6;  // ../RTL/cortexm0ds_logic.v(373)
  wire Y75pw6;  // ../RTL/cortexm0ds_logic.v(1398)
  wire Y76ow6;  // ../RTL/cortexm0ds_logic.v(930)
  wire Y7ciu6;  // ../RTL/cortexm0ds_logic.v(467)
  wire Y7cpw6;  // ../RTL/cortexm0ds_logic.v(1491)
  wire Y7dow6;  // ../RTL/cortexm0ds_logic.v(1023)
  wire Y7fhu6;  // ../RTL/cortexm0ds_logic.v(123)
  wire Y7ghu6;  // ../RTL/cortexm0ds_logic.v(126)
  wire Y7jiu6;  // ../RTL/cortexm0ds_logic.v(560)
  wire Y7khu6;  // ../RTL/cortexm0ds_logic.v(136)
  wire Y7kow6;  // ../RTL/cortexm0ds_logic.v(1117)
  wire Y7opw6;  // ../RTL/cortexm0ds_logic.v(1596)
  wire Y7qiu6;  // ../RTL/cortexm0ds_logic.v(654)
  wire Y7rhu6;  // ../RTL/cortexm0ds_logic.v(186)
  wire Y7row6;  // ../RTL/cortexm0ds_logic.v(1210)
  wire Y7upw6;  // ../RTL/cortexm0ds_logic.v(1606)
  wire Y7xiu6;  // ../RTL/cortexm0ds_logic.v(748)
  wire Y7yhu6;  // ../RTL/cortexm0ds_logic.v(280)
  wire Y7yow6;  // ../RTL/cortexm0ds_logic.v(1304)
  wire Y83ju6;  // ../RTL/cortexm0ds_logic.v(828)
  wire Y84iu6;  // ../RTL/cortexm0ds_logic.v(360)
  wire Y84pw6;  // ../RTL/cortexm0ds_logic.v(1385)
  wire Y8aju6;  // ../RTL/cortexm0ds_logic.v(922)
  wire Y8biu6;  // ../RTL/cortexm0ds_logic.v(454)
  wire Y8bpw6;  // ../RTL/cortexm0ds_logic.v(1478)
  wire Y8cow6;  // ../RTL/cortexm0ds_logic.v(1010)
  wire Y8iiu6;  // ../RTL/cortexm0ds_logic.v(547)
  wire Y8jow6;  // ../RTL/cortexm0ds_logic.v(1104)
  wire Y8lpw6;  // ../RTL/cortexm0ds_logic.v(1590)
  wire Y8piu6;  // ../RTL/cortexm0ds_logic.v(641)
  wire Y8qax6;  // ../RTL/cortexm0ds_logic.v(1662)
  wire Y8qhu6;  // ../RTL/cortexm0ds_logic.v(173)
  wire Y8qow6;  // ../RTL/cortexm0ds_logic.v(1197)
  wire Y8wiu6;  // ../RTL/cortexm0ds_logic.v(735)
  wire Y8xhu6;  // ../RTL/cortexm0ds_logic.v(267)
  wire Y8xow6;  // ../RTL/cortexm0ds_logic.v(1291)
  wire Y92ju6;  // ../RTL/cortexm0ds_logic.v(815)
  wire Y93bx6;  // ../RTL/cortexm0ds_logic.v(1685)
  wire Y93iu6;  // ../RTL/cortexm0ds_logic.v(347)
  wire Y93pw6;  // ../RTL/cortexm0ds_logic.v(1372)
  wire Y99ju6;  // ../RTL/cortexm0ds_logic.v(909)
  wire Y9aiu6;  // ../RTL/cortexm0ds_logic.v(441)
  wire Y9apw6;  // ../RTL/cortexm0ds_logic.v(1465)
  wire Y9bow6;  // ../RTL/cortexm0ds_logic.v(997)
  wire Y9hiu6;  // ../RTL/cortexm0ds_logic.v(534)
  wire Y9iow6;  // ../RTL/cortexm0ds_logic.v(1091)
  wire Y9jhu6;  // ../RTL/cortexm0ds_logic.v(133)
  wire Y9oiu6;  // ../RTL/cortexm0ds_logic.v(628)
  wire Y9phu6;  // ../RTL/cortexm0ds_logic.v(160)
  wire Y9pow6;  // ../RTL/cortexm0ds_logic.v(1184)
  wire Y9upw6;  // ../RTL/cortexm0ds_logic.v(1606)
  wire Y9viu6;  // ../RTL/cortexm0ds_logic.v(722)
  wire Y9whu6;  // ../RTL/cortexm0ds_logic.v(254)
  wire Y9wow6;  // ../RTL/cortexm0ds_logic.v(1278)
  wire Ya1ju6;  // ../RTL/cortexm0ds_logic.v(802)
  wire Ya2iu6;  // ../RTL/cortexm0ds_logic.v(334)
  wire Ya2pw6;  // ../RTL/cortexm0ds_logic.v(1359)
  wire Ya8ju6;  // ../RTL/cortexm0ds_logic.v(896)
  wire Ya9iu6;  // ../RTL/cortexm0ds_logic.v(428)
  wire Ya9pw6;  // ../RTL/cortexm0ds_logic.v(1452)
  wire Yaaow6;  // ../RTL/cortexm0ds_logic.v(984)
  wire Yagiu6;  // ../RTL/cortexm0ds_logic.v(521)
  wire Yahow6;  // ../RTL/cortexm0ds_logic.v(1078)
  wire Yaniu6;  // ../RTL/cortexm0ds_logic.v(615)
  wire Yaohu6;  // ../RTL/cortexm0ds_logic.v(147)
  wire Yaoow6;  // ../RTL/cortexm0ds_logic.v(1171)
  wire Yauiu6;  // ../RTL/cortexm0ds_logic.v(709)
  wire Yavhu6;  // ../RTL/cortexm0ds_logic.v(241)
  wire Yavow6;  // ../RTL/cortexm0ds_logic.v(1265)
  wire Yb0ju6;  // ../RTL/cortexm0ds_logic.v(789)
  wire Yb1iu6;  // ../RTL/cortexm0ds_logic.v(321)
  wire Yb1pw6;  // ../RTL/cortexm0ds_logic.v(1346)
  wire Yb7ju6;  // ../RTL/cortexm0ds_logic.v(883)
  wire Yb8iu6;  // ../RTL/cortexm0ds_logic.v(415)
  wire Yb8pw6;  // ../RTL/cortexm0ds_logic.v(1439)
  wire Yb9ow6;  // ../RTL/cortexm0ds_logic.v(971)
  wire Ybfiu6;  // ../RTL/cortexm0ds_logic.v(508)
  wire Ybgow6;  // ../RTL/cortexm0ds_logic.v(1065)
  wire Ybihu6;  // ../RTL/cortexm0ds_logic.v(131)
  wire Ybmiu6;  // ../RTL/cortexm0ds_logic.v(602)
  wire Ybnow6;  // ../RTL/cortexm0ds_logic.v(1158)
  wire Ybtiu6;  // ../RTL/cortexm0ds_logic.v(696)
  wire Ybuhu6;  // ../RTL/cortexm0ds_logic.v(228)
  wire Ybuow6;  // ../RTL/cortexm0ds_logic.v(1252)
  wire Ybupw6;  // ../RTL/cortexm0ds_logic.v(1607)
  wire Yc0iu6;  // ../RTL/cortexm0ds_logic.v(308)
  wire Yc0pw6;  // ../RTL/cortexm0ds_logic.v(1333)
  wire Yc6ju6;  // ../RTL/cortexm0ds_logic.v(870)
  wire Yc7iu6;  // ../RTL/cortexm0ds_logic.v(402)
  wire Yc7pw6;  // ../RTL/cortexm0ds_logic.v(1426)
  wire Yc8ow6;  // ../RTL/cortexm0ds_logic.v(958)
  wire Yceiu6;  // ../RTL/cortexm0ds_logic.v(495)
  wire Ycfow6;  // ../RTL/cortexm0ds_logic.v(1052)
  wire Ycliu6;  // ../RTL/cortexm0ds_logic.v(589)
  wire Ycmow6;  // ../RTL/cortexm0ds_logic.v(1145)
  wire Ycsiu6;  // ../RTL/cortexm0ds_logic.v(683)
  wire Ycthu6;  // ../RTL/cortexm0ds_logic.v(215)
  wire Yctow6;  // ../RTL/cortexm0ds_logic.v(1239)
  wire Ycziu6;  // ../RTL/cortexm0ds_logic.v(776)
  wire Yd5ju6;  // ../RTL/cortexm0ds_logic.v(857)
  wire Yd6iu6;  // ../RTL/cortexm0ds_logic.v(389)
  wire Yd6pw6;  // ../RTL/cortexm0ds_logic.v(1413)
  wire Yd7ow6;  // ../RTL/cortexm0ds_logic.v(945)
  wire Yddiu6;  // ../RTL/cortexm0ds_logic.v(482)
  wire Yddpw6;  // ../RTL/cortexm0ds_logic.v(1507)
  wire Ydeow6;  // ../RTL/cortexm0ds_logic.v(1039)
  wire Ydgax6;  // ../RTL/cortexm0ds_logic.v(1644)
  wire Ydkiu6;  // ../RTL/cortexm0ds_logic.v(576)
  wire Ydlow6;  // ../RTL/cortexm0ds_logic.v(1132)
  wire Ydopw6;  // ../RTL/cortexm0ds_logic.v(1596)
  wire Ydriu6;  // ../RTL/cortexm0ds_logic.v(670)
  wire Ydshu6;  // ../RTL/cortexm0ds_logic.v(202)
  wire Ydsow6;  // ../RTL/cortexm0ds_logic.v(1226)
  wire Ydupw6;  // ../RTL/cortexm0ds_logic.v(1607)
  wire Ydyiu6;  // ../RTL/cortexm0ds_logic.v(763)
  wire Ydzhu6;  // ../RTL/cortexm0ds_logic.v(295)
  wire Ydzow6;  // ../RTL/cortexm0ds_logic.v(1320)
  wire Ye4ju6;  // ../RTL/cortexm0ds_logic.v(844)
  wire Ye5iu6;  // ../RTL/cortexm0ds_logic.v(376)
  wire Ye5pw6;  // ../RTL/cortexm0ds_logic.v(1400)
  wire Ye6ow6;  // ../RTL/cortexm0ds_logic.v(932)
  wire Yeciu6;  // ../RTL/cortexm0ds_logic.v(469)
  wire Yecpw6;  // ../RTL/cortexm0ds_logic.v(1494)
  wire Yedow6;  // ../RTL/cortexm0ds_logic.v(1026)
  wire Yejiu6;  // ../RTL/cortexm0ds_logic.v(563)
  wire Yekow6;  // ../RTL/cortexm0ds_logic.v(1119)
  wire Yenhu6;  // ../RTL/cortexm0ds_logic.v(144)
  wire Yeqiu6;  // ../RTL/cortexm0ds_logic.v(657)
  wire Yerhu6;  // ../RTL/cortexm0ds_logic.v(189)
  wire Yerow6;  // ../RTL/cortexm0ds_logic.v(1213)
  wire Yexiu6;  // ../RTL/cortexm0ds_logic.v(750)
  wire Yeyhu6;  // ../RTL/cortexm0ds_logic.v(282)
  wire Yeyow6;  // ../RTL/cortexm0ds_logic.v(1307)
  wire Yf1qw6;  // ../RTL/cortexm0ds_logic.v(1620)
  wire Yf3ju6;  // ../RTL/cortexm0ds_logic.v(831)
  wire Yf4iu6;  // ../RTL/cortexm0ds_logic.v(363)
  wire Yf4pw6;  // ../RTL/cortexm0ds_logic.v(1387)
  wire Yfaju6;  // ../RTL/cortexm0ds_logic.v(924)
  wire Yfbiu6;  // ../RTL/cortexm0ds_logic.v(456)
  wire Yfbpw6;  // ../RTL/cortexm0ds_logic.v(1481)
  wire Yfcow6;  // ../RTL/cortexm0ds_logic.v(1013)
  wire Yfiiu6;  // ../RTL/cortexm0ds_logic.v(550)
  wire Yfjow6;  // ../RTL/cortexm0ds_logic.v(1106)
  wire Yfpiu6;  // ../RTL/cortexm0ds_logic.v(644)
  wire Yfqhu6;  // ../RTL/cortexm0ds_logic.v(176)
  wire Yfqow6;  // ../RTL/cortexm0ds_logic.v(1200)
  wire Yftpw6;  // ../RTL/cortexm0ds_logic.v(1605)
  wire Yfuax6;  // ../RTL/cortexm0ds_logic.v(1669)
  wire Yfupw6;  // ../RTL/cortexm0ds_logic.v(1607)
  wire Yfwiu6;  // ../RTL/cortexm0ds_logic.v(737)
  wire Yfxhu6;  // ../RTL/cortexm0ds_logic.v(269)
  wire Yfxow6;  // ../RTL/cortexm0ds_logic.v(1294)
  wire Yg2ju6;  // ../RTL/cortexm0ds_logic.v(818)
  wire Yg3iu6;  // ../RTL/cortexm0ds_logic.v(350)
  wire Yg3pw6;  // ../RTL/cortexm0ds_logic.v(1374)
  wire Yg9ju6;  // ../RTL/cortexm0ds_logic.v(911)
  wire Ygaiu6;  // ../RTL/cortexm0ds_logic.v(443)
  wire Ygapw6;  // ../RTL/cortexm0ds_logic.v(1468)
  wire Ygbow6;  // ../RTL/cortexm0ds_logic.v(1000)
  wire Yghiu6;  // ../RTL/cortexm0ds_logic.v(537)
  wire Ygiow6;  // ../RTL/cortexm0ds_logic.v(1093)
  wire Ygoiu6;  // ../RTL/cortexm0ds_logic.v(631)
  wire Ygphu6;  // ../RTL/cortexm0ds_logic.v(163)
  wire Ygpow6;  // ../RTL/cortexm0ds_logic.v(1187)
  wire Ygviu6;  // ../RTL/cortexm0ds_logic.v(724)
  wire Ygwhu6;  // ../RTL/cortexm0ds_logic.v(256)
  wire Ygwow6;  // ../RTL/cortexm0ds_logic.v(1281)
  wire Yh1ju6;  // ../RTL/cortexm0ds_logic.v(805)
  wire Yh2iu6;  // ../RTL/cortexm0ds_logic.v(337)
  wire Yh2pw6;  // ../RTL/cortexm0ds_logic.v(1361)
  wire Yh8ju6;  // ../RTL/cortexm0ds_logic.v(898)
  wire Yh9iu6;  // ../RTL/cortexm0ds_logic.v(430)
  wire Yh9pw6;  // ../RTL/cortexm0ds_logic.v(1455)
  wire Yhaow6;  // ../RTL/cortexm0ds_logic.v(987)
  wire Yhgiu6;  // ../RTL/cortexm0ds_logic.v(524)
  wire Yhhow6;  // ../RTL/cortexm0ds_logic.v(1080)
  wire Yhniu6;  // ../RTL/cortexm0ds_logic.v(618)
  wire Yhohu6;  // ../RTL/cortexm0ds_logic.v(150)
  wire Yhoow6;  // ../RTL/cortexm0ds_logic.v(1174)
  wire Yhuiu6;  // ../RTL/cortexm0ds_logic.v(711)
  wire Yhupw6;  // ../RTL/cortexm0ds_logic.v(1607)
  wire Yhvhu6;  // ../RTL/cortexm0ds_logic.v(243)
  wire Yhvow6;  // ../RTL/cortexm0ds_logic.v(1268)
  wire Yi0ju6;  // ../RTL/cortexm0ds_logic.v(792)
  wire Yi1iu6;  // ../RTL/cortexm0ds_logic.v(324)
  wire Yi1pw6;  // ../RTL/cortexm0ds_logic.v(1348)
  wire Yi7ju6;  // ../RTL/cortexm0ds_logic.v(885)
  wire Yi8iu6;  // ../RTL/cortexm0ds_logic.v(417)
  wire Yi8pw6;  // ../RTL/cortexm0ds_logic.v(1442)
  wire Yi9ow6;  // ../RTL/cortexm0ds_logic.v(974)
  wire Yifiu6;  // ../RTL/cortexm0ds_logic.v(511)
  wire Yigow6;  // ../RTL/cortexm0ds_logic.v(1067)
  wire Yimiu6;  // ../RTL/cortexm0ds_logic.v(605)
  wire Yinow6;  // ../RTL/cortexm0ds_logic.v(1161)
  wire Yitiu6;  // ../RTL/cortexm0ds_logic.v(698)
  wire Yiuhu6;  // ../RTL/cortexm0ds_logic.v(230)
  wire Yiuow6;  // ../RTL/cortexm0ds_logic.v(1255)
  wire Yizpw6;  // ../RTL/cortexm0ds_logic.v(1616)
  wire Yj0iu6;  // ../RTL/cortexm0ds_logic.v(311)
  wire Yj0pw6;  // ../RTL/cortexm0ds_logic.v(1335)
  wire Yj6ju6;  // ../RTL/cortexm0ds_logic.v(872)
  wire Yj7iu6;  // ../RTL/cortexm0ds_logic.v(404)
  wire Yj7pw6;  // ../RTL/cortexm0ds_logic.v(1429)
  wire Yj8ow6;  // ../RTL/cortexm0ds_logic.v(961)
  wire Yjaax6;  // ../RTL/cortexm0ds_logic.v(1632)
  wire Yjeiu6;  // ../RTL/cortexm0ds_logic.v(498)
  wire Yjfow6;  // ../RTL/cortexm0ds_logic.v(1054)
  wire Yjliu6;  // ../RTL/cortexm0ds_logic.v(592)
  wire Yjmow6;  // ../RTL/cortexm0ds_logic.v(1148)
  wire Yjsiu6;  // ../RTL/cortexm0ds_logic.v(685)
  wire Yjthu6;  // ../RTL/cortexm0ds_logic.v(217)
  wire Yjtow6;  // ../RTL/cortexm0ds_logic.v(1242)
  wire Yjupw6;  // ../RTL/cortexm0ds_logic.v(1607)
  wire Yjziu6;  // ../RTL/cortexm0ds_logic.v(779)
  wire Yk5ju6;  // ../RTL/cortexm0ds_logic.v(859)
  wire Yk6iu6;  // ../RTL/cortexm0ds_logic.v(391)
  wire Yk6pw6;  // ../RTL/cortexm0ds_logic.v(1416)
  wire Yk7ow6;  // ../RTL/cortexm0ds_logic.v(948)
  wire Ykdiu6;  // ../RTL/cortexm0ds_logic.v(485)
  wire Ykdpw6;  // ../RTL/cortexm0ds_logic.v(1509)
  wire Ykeow6;  // ../RTL/cortexm0ds_logic.v(1041)
  wire Ykkiu6;  // ../RTL/cortexm0ds_logic.v(579)
  wire Yklow6;  // ../RTL/cortexm0ds_logic.v(1135)
  wire Yklpw6;  // ../RTL/cortexm0ds_logic.v(1591)
  wire Ykriu6;  // ../RTL/cortexm0ds_logic.v(672)
  wire Ykshu6;  // ../RTL/cortexm0ds_logic.v(204)
  wire Yksow6;  // ../RTL/cortexm0ds_logic.v(1229)
  wire Ykyiu6;  // ../RTL/cortexm0ds_logic.v(766)
  wire Ykzhu6;  // ../RTL/cortexm0ds_logic.v(298)
  wire Ykzow6;  // ../RTL/cortexm0ds_logic.v(1322)
  wire Ykzpw6;  // ../RTL/cortexm0ds_logic.v(1616)
  wire Yl4ju6;  // ../RTL/cortexm0ds_logic.v(846)
  wire Yl5iu6;  // ../RTL/cortexm0ds_logic.v(378)
  wire Yl5pw6;  // ../RTL/cortexm0ds_logic.v(1403)
  wire Yl6ow6;  // ../RTL/cortexm0ds_logic.v(935)
  wire Ylciu6;  // ../RTL/cortexm0ds_logic.v(472)
  wire Ylcpw6;  // ../RTL/cortexm0ds_logic.v(1496)
  wire Yldow6;  // ../RTL/cortexm0ds_logic.v(1028)
  wire Yljiu6;  // ../RTL/cortexm0ds_logic.v(566)
  wire Ylkow6;  // ../RTL/cortexm0ds_logic.v(1122)
  wire Ylqiu6;  // ../RTL/cortexm0ds_logic.v(659)
  wire Ylrhu6;  // ../RTL/cortexm0ds_logic.v(191)
  wire Ylrow6;  // ../RTL/cortexm0ds_logic.v(1216)
  wire Ylxiu6;  // ../RTL/cortexm0ds_logic.v(753)
  wire Ylyhu6;  // ../RTL/cortexm0ds_logic.v(285)
  wire Ylyow6;  // ../RTL/cortexm0ds_logic.v(1309)
  wire Ym3ju6;  // ../RTL/cortexm0ds_logic.v(833)
  wire Ym3qw6;  // ../RTL/cortexm0ds_logic.v(1624)
  wire Ym4iu6;  // ../RTL/cortexm0ds_logic.v(365)
  wire Ym4pw6;  // ../RTL/cortexm0ds_logic.v(1390)
  wire Ymaju6;  // ../RTL/cortexm0ds_logic.v(927)
  wire Ymbiu6;  // ../RTL/cortexm0ds_logic.v(459)
  wire Ymbpw6;  // ../RTL/cortexm0ds_logic.v(1483)
  wire Ymcow6;  // ../RTL/cortexm0ds_logic.v(1015)
  wire Ymiiu6;  // ../RTL/cortexm0ds_logic.v(553)
  wire Ymjow6;  // ../RTL/cortexm0ds_logic.v(1109)
  wire Ympiu6;  // ../RTL/cortexm0ds_logic.v(646)
  wire Ymqhu6;  // ../RTL/cortexm0ds_logic.v(178)
  wire Ymqow6;  // ../RTL/cortexm0ds_logic.v(1203)
  wire Ymwiu6;  // ../RTL/cortexm0ds_logic.v(740)
  wire Ymwpw6;  // ../RTL/cortexm0ds_logic.v(1611)
  wire Ymxhu6;  // ../RTL/cortexm0ds_logic.v(272)
  wire Ymxow6;  // ../RTL/cortexm0ds_logic.v(1296)
  wire Ymzpw6;  // ../RTL/cortexm0ds_logic.v(1616)
  wire Yn2ju6;  // ../RTL/cortexm0ds_logic.v(820)
  wire Yn3iu6;  // ../RTL/cortexm0ds_logic.v(352)
  wire Yn3pw6;  // ../RTL/cortexm0ds_logic.v(1377)
  wire Yn9ju6;  // ../RTL/cortexm0ds_logic.v(914)
  wire Ynaiu6;  // ../RTL/cortexm0ds_logic.v(446)
  wire Ynapw6;  // ../RTL/cortexm0ds_logic.v(1470)
  wire Ynbow6;  // ../RTL/cortexm0ds_logic.v(1002)
  wire Ynehu6;  // ../RTL/cortexm0ds_logic.v(122)
  wire Ynhiu6;  // ../RTL/cortexm0ds_logic.v(540)
  wire Yniow6;  // ../RTL/cortexm0ds_logic.v(1096)
  wire Ynoiu6;  // ../RTL/cortexm0ds_logic.v(633)
  wire Ynphu6;  // ../RTL/cortexm0ds_logic.v(165)
  wire Ynpow6;  // ../RTL/cortexm0ds_logic.v(1190)
  wire Ynspw6;  // ../RTL/cortexm0ds_logic.v(1604)
  wire Ynviu6;  // ../RTL/cortexm0ds_logic.v(727)
  wire Ynwhu6;  // ../RTL/cortexm0ds_logic.v(259)
  wire Ynwow6;  // ../RTL/cortexm0ds_logic.v(1283)
  wire Yo1ju6;  // ../RTL/cortexm0ds_logic.v(807)
  wire Yo2iu6;  // ../RTL/cortexm0ds_logic.v(339)
  wire Yo2pw6;  // ../RTL/cortexm0ds_logic.v(1364)
  wire Yo8ju6;  // ../RTL/cortexm0ds_logic.v(901)
  wire Yo9iu6;  // ../RTL/cortexm0ds_logic.v(433)
  wire Yo9pw6;  // ../RTL/cortexm0ds_logic.v(1457)
  wire Yoaow6;  // ../RTL/cortexm0ds_logic.v(989)
  wire Yogax6;  // ../RTL/cortexm0ds_logic.v(1644)
  wire Yogiu6;  // ../RTL/cortexm0ds_logic.v(527)
  wire Yohow6;  // ../RTL/cortexm0ds_logic.v(1083)
  wire Yokhu6;  // ../RTL/cortexm0ds_logic.v(137)
  wire Yoniu6;  // ../RTL/cortexm0ds_logic.v(620)
  wire Yoohu6;  // ../RTL/cortexm0ds_logic.v(152)
  wire Yooow6;  // ../RTL/cortexm0ds_logic.v(1177)
  wire Youiu6;  // ../RTL/cortexm0ds_logic.v(714)
  wire Yovhu6;  // ../RTL/cortexm0ds_logic.v(246)
  wire Yovow6;  // ../RTL/cortexm0ds_logic.v(1270)
  wire Yp0ju6;  // ../RTL/cortexm0ds_logic.v(794)
  wire Yp1iu6;  // ../RTL/cortexm0ds_logic.v(326)
  wire Yp1pw6;  // ../RTL/cortexm0ds_logic.v(1351)
  wire Yp7ju6;  // ../RTL/cortexm0ds_logic.v(888)
  wire Yp8iu6;  // ../RTL/cortexm0ds_logic.v(420)
  wire Yp8pw6;  // ../RTL/cortexm0ds_logic.v(1444)
  wire Yp9ow6;  // ../RTL/cortexm0ds_logic.v(976)
  wire Ypfiu6;  // ../RTL/cortexm0ds_logic.v(514)
  wire Ypgow6;  // ../RTL/cortexm0ds_logic.v(1070)
  wire Ypmhu6;  // ../RTL/cortexm0ds_logic.v(143)
  wire Ypmiu6;  // ../RTL/cortexm0ds_logic.v(607)
  wire Ypnow6;  // ../RTL/cortexm0ds_logic.v(1164)
  wire Ypspw6;  // ../RTL/cortexm0ds_logic.v(1604)
  wire Yptiu6;  // ../RTL/cortexm0ds_logic.v(701)
  wire Ypuhu6;  // ../RTL/cortexm0ds_logic.v(233)
  wire Ypuow6;  // ../RTL/cortexm0ds_logic.v(1257)
  wire Yq0iu6;  // ../RTL/cortexm0ds_logic.v(313)
  wire Yq0pw6;  // ../RTL/cortexm0ds_logic.v(1338)
  wire Yq6ju6;  // ../RTL/cortexm0ds_logic.v(875)
  wire Yq7iu6;  // ../RTL/cortexm0ds_logic.v(407)
  wire Yq7pw6;  // ../RTL/cortexm0ds_logic.v(1431)
  wire Yq8ow6;  // ../RTL/cortexm0ds_logic.v(963)
  wire Yqeiu6;  // ../RTL/cortexm0ds_logic.v(501)
  wire Yqfow6;  // ../RTL/cortexm0ds_logic.v(1057)
  wire Yqjhu6;  // ../RTL/cortexm0ds_logic.v(134)
  wire Yqliu6;  // ../RTL/cortexm0ds_logic.v(594)
  wire Yqmow6;  // ../RTL/cortexm0ds_logic.v(1151)
  wire Yqsiu6;  // ../RTL/cortexm0ds_logic.v(688)
  wire Yqthu6;  // ../RTL/cortexm0ds_logic.v(220)
  wire Yqtow6;  // ../RTL/cortexm0ds_logic.v(1244)
  wire Yqzax6;  // ../RTL/cortexm0ds_logic.v(1679)
  wire Yqziu6;  // ../RTL/cortexm0ds_logic.v(781)
  wire Yr5ju6;  // ../RTL/cortexm0ds_logic.v(862)
  wire Yr6iu6;  // ../RTL/cortexm0ds_logic.v(394)
  wire Yr6pw6;  // ../RTL/cortexm0ds_logic.v(1418)
  wire Yr7ow6;  // ../RTL/cortexm0ds_logic.v(950)
  wire Yrdiu6;  // ../RTL/cortexm0ds_logic.v(488)
  wire Yrdpw6;  // ../RTL/cortexm0ds_logic.v(1512)
  wire Yreow6;  // ../RTL/cortexm0ds_logic.v(1044)
  wire Yrkiu6;  // ../RTL/cortexm0ds_logic.v(581)
  wire Yrlow6;  // ../RTL/cortexm0ds_logic.v(1138)
  wire Yrriu6;  // ../RTL/cortexm0ds_logic.v(675)
  wire Yrshu6;  // ../RTL/cortexm0ds_logic.v(207)
  wire Yrsow6;  // ../RTL/cortexm0ds_logic.v(1231)
  wire Yrspw6;  // ../RTL/cortexm0ds_logic.v(1604)
  wire Yryax6;  // ../RTL/cortexm0ds_logic.v(1677)
  wire Yryiu6;  // ../RTL/cortexm0ds_logic.v(768)
  wire Yrzhu6;  // ../RTL/cortexm0ds_logic.v(300)
  wire Yrzow6;  // ../RTL/cortexm0ds_logic.v(1325)
  wire Ys4ju6;  // ../RTL/cortexm0ds_logic.v(849)
  wire Ys5iu6;  // ../RTL/cortexm0ds_logic.v(381)
  wire Ys5pw6;  // ../RTL/cortexm0ds_logic.v(1405)
  wire Ys6ow6;  // ../RTL/cortexm0ds_logic.v(937)
  wire Ysciu6;  // ../RTL/cortexm0ds_logic.v(475)
  wire Yscpw6;  // ../RTL/cortexm0ds_logic.v(1499)
  wire Ysdow6;  // ../RTL/cortexm0ds_logic.v(1031)
  wire Ysiax6;  // ../RTL/cortexm0ds_logic.v(1648)
  wire Ysihu6;  // ../RTL/cortexm0ds_logic.v(132)
  wire Ysjiu6;  // ../RTL/cortexm0ds_logic.v(568)
  wire Yskow6;  // ../RTL/cortexm0ds_logic.v(1125)
  wire Yslhu6;  // ../RTL/cortexm0ds_logic.v(140)
  wire Ysqiu6;  // ../RTL/cortexm0ds_logic.v(662)
  wire Ysrhu6;  // ../RTL/cortexm0ds_logic.v(194)
  wire Ysrow6;  // ../RTL/cortexm0ds_logic.v(1218)
  wire Ysxiu6;  // ../RTL/cortexm0ds_logic.v(755)
  wire Ysyhu6;  // ../RTL/cortexm0ds_logic.v(287)
  wire Ysyow6;  // ../RTL/cortexm0ds_logic.v(1312)
  wire Yt3ju6;  // ../RTL/cortexm0ds_logic.v(836)
  wire Yt4bx6;  // ../RTL/cortexm0ds_logic.v(1688)
  wire Yt4iu6;  // ../RTL/cortexm0ds_logic.v(368)
  wire Yt4pw6;  // ../RTL/cortexm0ds_logic.v(1392)
  wire Yt8bx6;  // ../RTL/cortexm0ds_logic.v(1695)
  wire Ytbiu6;  // ../RTL/cortexm0ds_logic.v(462)
  wire Ytbpw6;  // ../RTL/cortexm0ds_logic.v(1486)
  wire Ytcow6;  // ../RTL/cortexm0ds_logic.v(1018)
  wire Ytiiu6;  // ../RTL/cortexm0ds_logic.v(555)
  wire Ytjow6;  // ../RTL/cortexm0ds_logic.v(1112)
  wire Ytlax6;  // ../RTL/cortexm0ds_logic.v(1654)
  wire Ytpiu6;  // ../RTL/cortexm0ds_logic.v(649)
  wire Ytqhu6;  // ../RTL/cortexm0ds_logic.v(181)
  wire Ytqow6;  // ../RTL/cortexm0ds_logic.v(1205)
  wire Ytspw6;  // ../RTL/cortexm0ds_logic.v(1604)
  wire Ytwiu6;  // ../RTL/cortexm0ds_logic.v(742)
  wire Ytxhu6;  // ../RTL/cortexm0ds_logic.v(274)
  wire Ytxow6;  // ../RTL/cortexm0ds_logic.v(1299)
  wire Yu2ju6;  // ../RTL/cortexm0ds_logic.v(823)
  wire Yu3iu6;  // ../RTL/cortexm0ds_logic.v(355)
  wire Yu3pw6;  // ../RTL/cortexm0ds_logic.v(1379)
  wire Yu9ju6;  // ../RTL/cortexm0ds_logic.v(917)
  wire Yuaiu6;  // ../RTL/cortexm0ds_logic.v(449)
  wire Yuapw6;  // ../RTL/cortexm0ds_logic.v(1473)
  wire Yubbx6;  // ../RTL/cortexm0ds_logic.v(1700)
  wire Yubow6;  // ../RTL/cortexm0ds_logic.v(1005)
  wire Yuhhu6;  // ../RTL/cortexm0ds_logic.v(129)
  wire Yuhiu6;  // ../RTL/cortexm0ds_logic.v(542)
  wire Yuiow6;  // ../RTL/cortexm0ds_logic.v(1099)
  wire Yuoiu6;  // ../RTL/cortexm0ds_logic.v(636)
  wire Yuphu6;  // ../RTL/cortexm0ds_logic.v(168)
  wire Yupow6;  // ../RTL/cortexm0ds_logic.v(1192)
  wire Yuviu6;  // ../RTL/cortexm0ds_logic.v(729)
  wire Yuwhu6;  // ../RTL/cortexm0ds_logic.v(261)
  wire Yuwow6;  // ../RTL/cortexm0ds_logic.v(1286)
  wire Yv1ju6;  // ../RTL/cortexm0ds_logic.v(810)
  wire Yv2iu6;  // ../RTL/cortexm0ds_logic.v(342)
  wire Yv2pw6;  // ../RTL/cortexm0ds_logic.v(1366)
  wire Yv8ju6;  // ../RTL/cortexm0ds_logic.v(904)
  wire Yv9iu6;  // ../RTL/cortexm0ds_logic.v(436)
  wire Yv9pw6;  // ../RTL/cortexm0ds_logic.v(1460)
  wire Yvabx6;  // ../RTL/cortexm0ds_logic.v(1699)
  wire Yvaow6;  // ../RTL/cortexm0ds_logic.v(992)
  wire Yvgiu6;  // ../RTL/cortexm0ds_logic.v(529)
  wire Yvhow6;  // ../RTL/cortexm0ds_logic.v(1086)
  wire Yvjpw6;  // ../RTL/cortexm0ds_logic.v(1587)
  wire Yvniu6;  // ../RTL/cortexm0ds_logic.v(623)
  wire Yvohu6;  // ../RTL/cortexm0ds_logic.v(155)
  wire Yvoow6;  // ../RTL/cortexm0ds_logic.v(1179)
  wire Yvspw6;  // ../RTL/cortexm0ds_logic.v(1604)
  wire Yvuiu6;  // ../RTL/cortexm0ds_logic.v(716)
  wire Yvvhu6;  // ../RTL/cortexm0ds_logic.v(248)
  wire Yvvow6;  // ../RTL/cortexm0ds_logic.v(1273)
  wire Yw0ju6;  // ../RTL/cortexm0ds_logic.v(797)
  wire Yw1iu6;  // ../RTL/cortexm0ds_logic.v(329)
  wire Yw1pw6;  // ../RTL/cortexm0ds_logic.v(1353)
  wire Yw3bx6;  // ../RTL/cortexm0ds_logic.v(1686)
  wire Yw7ju6;  // ../RTL/cortexm0ds_logic.v(891)
  wire Yw8iu6;  // ../RTL/cortexm0ds_logic.v(423)
  wire Yw8pw6;  // ../RTL/cortexm0ds_logic.v(1447)
  wire Yw9ow6;  // ../RTL/cortexm0ds_logic.v(979)
  wire Ywfiu6;  // ../RTL/cortexm0ds_logic.v(516)
  wire Ywgow6;  // ../RTL/cortexm0ds_logic.v(1073)
  wire Ywmiu6;  // ../RTL/cortexm0ds_logic.v(610)
  wire Ywnow6;  // ../RTL/cortexm0ds_logic.v(1166)
  wire Ywtiu6;  // ../RTL/cortexm0ds_logic.v(703)
  wire Ywuhu6;  // ../RTL/cortexm0ds_logic.v(235)
  wire Ywuow6;  // ../RTL/cortexm0ds_logic.v(1260)
  wire Yx0iu6;  // ../RTL/cortexm0ds_logic.v(316)
  wire Yx0pw6;  // ../RTL/cortexm0ds_logic.v(1340)
  wire Yx6ju6;  // ../RTL/cortexm0ds_logic.v(878)
  wire Yx7iu6;  // ../RTL/cortexm0ds_logic.v(410)
  wire Yx7pw6;  // ../RTL/cortexm0ds_logic.v(1434)
  wire Yx8ow6;  // ../RTL/cortexm0ds_logic.v(966)
  wire Yxdax6;  // ../RTL/cortexm0ds_logic.v(1639)
  wire Yxeiu6;  // ../RTL/cortexm0ds_logic.v(503)
  wire Yxfow6;  // ../RTL/cortexm0ds_logic.v(1060)
  wire Yxliu6;  // ../RTL/cortexm0ds_logic.v(597)
  wire Yxmow6;  // ../RTL/cortexm0ds_logic.v(1153)
  wire Yxrpw6;  // ../RTL/cortexm0ds_logic.v(1602)
  wire Yxsiu6;  // ../RTL/cortexm0ds_logic.v(690)
  wire Yxspw6;  // ../RTL/cortexm0ds_logic.v(1604)
  wire Yxthu6;  // ../RTL/cortexm0ds_logic.v(222)
  wire Yxtow6;  // ../RTL/cortexm0ds_logic.v(1247)
  wire Yxziu6;  // ../RTL/cortexm0ds_logic.v(784)
  wire Yy5ju6;  // ../RTL/cortexm0ds_logic.v(865)
  wire Yy6iu6;  // ../RTL/cortexm0ds_logic.v(397)
  wire Yy6pw6;  // ../RTL/cortexm0ds_logic.v(1421)
  wire Yy7ow6;  // ../RTL/cortexm0ds_logic.v(953)
  wire Yybax6;  // ../RTL/cortexm0ds_logic.v(1635)
  wire Yydiu6;  // ../RTL/cortexm0ds_logic.v(490)
  wire Yydpw6;  // ../RTL/cortexm0ds_logic.v(1515)
  wire Yyeow6;  // ../RTL/cortexm0ds_logic.v(1047)
  wire Yyfhu6;  // ../RTL/cortexm0ds_logic.v(125)
  wire Yyghu6;  // ../RTL/cortexm0ds_logic.v(127)
  wire Yykiu6;  // ../RTL/cortexm0ds_logic.v(584)
  wire Yylow6;  // ../RTL/cortexm0ds_logic.v(1140)
  wire Yyriu6;  // ../RTL/cortexm0ds_logic.v(677)
  wire Yyshu6;  // ../RTL/cortexm0ds_logic.v(209)
  wire Yysow6;  // ../RTL/cortexm0ds_logic.v(1234)
  wire Yyyiu6;  // ../RTL/cortexm0ds_logic.v(771)
  wire Yyzhu6;  // ../RTL/cortexm0ds_logic.v(303)
  wire Yyzow6;  // ../RTL/cortexm0ds_logic.v(1327)
  wire Yz4ju6;  // ../RTL/cortexm0ds_logic.v(852)
  wire Yz5iu6;  // ../RTL/cortexm0ds_logic.v(384)
  wire Yz5pw6;  // ../RTL/cortexm0ds_logic.v(1408)
  wire Yz6ow6;  // ../RTL/cortexm0ds_logic.v(940)
  wire Yzciu6;  // ../RTL/cortexm0ds_logic.v(477)
  wire Yzcpw6;  // ../RTL/cortexm0ds_logic.v(1502)
  wire Yzdow6;  // ../RTL/cortexm0ds_logic.v(1034)
  wire Yzjiu6;  // ../RTL/cortexm0ds_logic.v(571)
  wire Yzkow6;  // ../RTL/cortexm0ds_logic.v(1127)
  wire Yzlpw6;  // ../RTL/cortexm0ds_logic.v(1591)
  wire Yzqiu6;  // ../RTL/cortexm0ds_logic.v(664)
  wire Yzqpw6;  // ../RTL/cortexm0ds_logic.v(1601)
  wire Yzrhu6;  // ../RTL/cortexm0ds_logic.v(196)
  wire Yzrow6;  // ../RTL/cortexm0ds_logic.v(1221)
  wire Yzspw6;  // ../RTL/cortexm0ds_logic.v(1604)
  wire Yzxiu6;  // ../RTL/cortexm0ds_logic.v(758)
  wire Yzyhu6;  // ../RTL/cortexm0ds_logic.v(290)
  wire Yzyow6;  // ../RTL/cortexm0ds_logic.v(1314)
  wire Z01ju6;  // ../RTL/cortexm0ds_logic.v(798)
  wire Z02iu6;  // ../RTL/cortexm0ds_logic.v(330)
  wire Z02pw6;  // ../RTL/cortexm0ds_logic.v(1355)
  wire Z08ju6;  // ../RTL/cortexm0ds_logic.v(892)
  wire Z09iu6;  // ../RTL/cortexm0ds_logic.v(424)
  wire Z09pw6;  // ../RTL/cortexm0ds_logic.v(1448)
  wire Z0aow6;  // ../RTL/cortexm0ds_logic.v(980)
  wire Z0giu6;  // ../RTL/cortexm0ds_logic.v(518)
  wire Z0how6;  // ../RTL/cortexm0ds_logic.v(1074)
  wire Z0niu6;  // ../RTL/cortexm0ds_logic.v(611)
  wire Z0oow6;  // ../RTL/cortexm0ds_logic.v(1168)
  wire Z0uiu6;  // ../RTL/cortexm0ds_logic.v(705)
  wire Z0vhu6;  // ../RTL/cortexm0ds_logic.v(237)
  wire Z0vow6;  // ../RTL/cortexm0ds_logic.v(1261)
  wire Z10ju6;  // ../RTL/cortexm0ds_logic.v(785)
  wire Z11iu6;  // ../RTL/cortexm0ds_logic.v(317)
  wire Z11pw6;  // ../RTL/cortexm0ds_logic.v(1342)
  wire Z17ju6;  // ../RTL/cortexm0ds_logic.v(879)
  wire Z18bx6;  // ../RTL/cortexm0ds_logic.v(1693)
  wire Z18iu6;  // ../RTL/cortexm0ds_logic.v(411)
  wire Z18pw6;  // ../RTL/cortexm0ds_logic.v(1435)
  wire Z19ow6;  // ../RTL/cortexm0ds_logic.v(967)
  wire Z1fiu6;  // ../RTL/cortexm0ds_logic.v(505)
  wire Z1gow6;  // ../RTL/cortexm0ds_logic.v(1061)
  wire Z1miu6;  // ../RTL/cortexm0ds_logic.v(598)
  wire Z1now6;  // ../RTL/cortexm0ds_logic.v(1155)
  wire Z1tiu6;  // ../RTL/cortexm0ds_logic.v(692)
  wire Z1tpw6;  // ../RTL/cortexm0ds_logic.v(1604)
  wire Z1uhu6;  // ../RTL/cortexm0ds_logic.v(224)
  wire Z1uow6;  // ../RTL/cortexm0ds_logic.v(1248)
  wire Z20iu6;  // ../RTL/cortexm0ds_logic.v(304)
  wire Z20pw6;  // ../RTL/cortexm0ds_logic.v(1329)
  wire Z26ju6;  // ../RTL/cortexm0ds_logic.v(866)
  wire Z27iu6;  // ../RTL/cortexm0ds_logic.v(398)
  wire Z27pw6;  // ../RTL/cortexm0ds_logic.v(1422)
  wire Z28ow6;  // ../RTL/cortexm0ds_logic.v(954)
  wire Z2aax6;  // ../RTL/cortexm0ds_logic.v(1631)
  wire Z2eiu6;  // ../RTL/cortexm0ds_logic.v(492)
  wire Z2epw6;  // ../RTL/cortexm0ds_logic.v(1516)
  wire Z2fow6;  // ../RTL/cortexm0ds_logic.v(1048)
  wire Z2liu6;  // ../RTL/cortexm0ds_logic.v(585)
  wire Z2mow6;  // ../RTL/cortexm0ds_logic.v(1142)
  wire Z2siu6;  // ../RTL/cortexm0ds_logic.v(679)
  wire Z2thu6;  // ../RTL/cortexm0ds_logic.v(211)
  wire Z2tow6;  // ../RTL/cortexm0ds_logic.v(1235)
  wire Z2ziu6;  // ../RTL/cortexm0ds_logic.v(772)
  wire Z35ju6;  // ../RTL/cortexm0ds_logic.v(853)
  wire Z36iu6;  // ../RTL/cortexm0ds_logic.v(385)
  wire Z36pw6;  // ../RTL/cortexm0ds_logic.v(1409)
  wire Z37ow6;  // ../RTL/cortexm0ds_logic.v(941)
  wire Z38bx6;  // ../RTL/cortexm0ds_logic.v(1694)
  wire Z3diu6;  // ../RTL/cortexm0ds_logic.v(479)
  wire Z3dpw6;  // ../RTL/cortexm0ds_logic.v(1503)
  wire Z3eow6;  // ../RTL/cortexm0ds_logic.v(1035)
  wire Z3kiu6;  // ../RTL/cortexm0ds_logic.v(572)
  wire Z3low6;  // ../RTL/cortexm0ds_logic.v(1129)
  wire Z3riu6;  // ../RTL/cortexm0ds_logic.v(666)
  wire Z3shu6;  // ../RTL/cortexm0ds_logic.v(198)
  wire Z3sow6;  // ../RTL/cortexm0ds_logic.v(1222)
  wire Z3spw6;  // ../RTL/cortexm0ds_logic.v(1603)
  wire Z3tpw6;  // ../RTL/cortexm0ds_logic.v(1604)
  wire Z3yiu6;  // ../RTL/cortexm0ds_logic.v(759)
  wire Z3zhu6;  // ../RTL/cortexm0ds_logic.v(291)
  wire Z3zow6;  // ../RTL/cortexm0ds_logic.v(1316)
  wire Z44ju6;  // ../RTL/cortexm0ds_logic.v(840)
  wire Z45iu6;  // ../RTL/cortexm0ds_logic.v(372)
  wire Z45pw6;  // ../RTL/cortexm0ds_logic.v(1396)
  wire Z47ax6;  // ../RTL/cortexm0ds_logic.v(1626)
  wire Z4ciu6;  // ../RTL/cortexm0ds_logic.v(466)
  wire Z4cpw6;  // ../RTL/cortexm0ds_logic.v(1490)
  wire Z4dow6;  // ../RTL/cortexm0ds_logic.v(1022)
  wire Z4jiu6;  // ../RTL/cortexm0ds_logic.v(559)
  wire Z4kow6;  // ../RTL/cortexm0ds_logic.v(1116)
  wire Z4qiu6;  // ../RTL/cortexm0ds_logic.v(653)
  wire Z4rhu6;  // ../RTL/cortexm0ds_logic.v(185)
  wire Z4row6;  // ../RTL/cortexm0ds_logic.v(1209)
  wire Z4xiu6;  // ../RTL/cortexm0ds_logic.v(746)
  wire Z4yhu6;  // ../RTL/cortexm0ds_logic.v(278)
  wire Z4yow6;  // ../RTL/cortexm0ds_logic.v(1303)
  wire Z53ju6;  // ../RTL/cortexm0ds_logic.v(827)
  wire Z54iu6;  // ../RTL/cortexm0ds_logic.v(359)
  wire Z54pw6;  // ../RTL/cortexm0ds_logic.v(1383)
  wire Z58bx6;  // ../RTL/cortexm0ds_logic.v(1694)
  wire Z5aju6;  // ../RTL/cortexm0ds_logic.v(921)
  wire Z5biu6;  // ../RTL/cortexm0ds_logic.v(453)
  wire Z5bpw6;  // ../RTL/cortexm0ds_logic.v(1477)
  wire Z5cow6;  // ../RTL/cortexm0ds_logic.v(1009)
  wire Z5iiu6;  // ../RTL/cortexm0ds_logic.v(546)
  wire Z5jow6;  // ../RTL/cortexm0ds_logic.v(1103)
  wire Z5piu6;  // ../RTL/cortexm0ds_logic.v(640)
  wire Z5qhu6;  // ../RTL/cortexm0ds_logic.v(172)
  wire Z5qow6;  // ../RTL/cortexm0ds_logic.v(1196)
  wire Z5tpw6;  // ../RTL/cortexm0ds_logic.v(1604)
  wire Z5wiu6;  // ../RTL/cortexm0ds_logic.v(733)
  wire Z5xhu6;  // ../RTL/cortexm0ds_logic.v(265)
  wire Z5xow6;  // ../RTL/cortexm0ds_logic.v(1290)
  wire Z62ju6;  // ../RTL/cortexm0ds_logic.v(814)
  wire Z63iu6;  // ../RTL/cortexm0ds_logic.v(346)
  wire Z63pw6;  // ../RTL/cortexm0ds_logic.v(1370)
  wire Z67ax6;  // ../RTL/cortexm0ds_logic.v(1626)
  wire Z69ju6;  // ../RTL/cortexm0ds_logic.v(908)
  wire Z6aiu6;  // ../RTL/cortexm0ds_logic.v(440)
  wire Z6apw6;  // ../RTL/cortexm0ds_logic.v(1464)
  wire Z6bow6;  // ../RTL/cortexm0ds_logic.v(996)
  wire Z6hiu6;  // ../RTL/cortexm0ds_logic.v(533)
  wire Z6iow6;  // ../RTL/cortexm0ds_logic.v(1090)
  wire Z6oiu6;  // ../RTL/cortexm0ds_logic.v(627)
  wire Z6phu6;  // ../RTL/cortexm0ds_logic.v(159)
  wire Z6pow6;  // ../RTL/cortexm0ds_logic.v(1183)
  wire Z6qax6;  // ../RTL/cortexm0ds_logic.v(1662)
  wire Z6viu6;  // ../RTL/cortexm0ds_logic.v(720)
  wire Z6whu6;  // ../RTL/cortexm0ds_logic.v(252)
  wire Z6wow6;  // ../RTL/cortexm0ds_logic.v(1277)
  wire Z71bx6;  // ../RTL/cortexm0ds_logic.v(1681)
  wire Z71ju6;  // ../RTL/cortexm0ds_logic.v(801)
  wire Z72iu6;  // ../RTL/cortexm0ds_logic.v(333)
  wire Z72pw6;  // ../RTL/cortexm0ds_logic.v(1357)
  wire Z73qw6;  // ../RTL/cortexm0ds_logic.v(1623)
  wire Z78bx6;  // ../RTL/cortexm0ds_logic.v(1694)
  wire Z78ju6;  // ../RTL/cortexm0ds_logic.v(895)
  wire Z79iu6;  // ../RTL/cortexm0ds_logic.v(427)
  wire Z79pw6;  // ../RTL/cortexm0ds_logic.v(1451)
  wire Z7aow6;  // ../RTL/cortexm0ds_logic.v(983)
  wire Z7giu6;  // ../RTL/cortexm0ds_logic.v(520)
  wire Z7how6;  // ../RTL/cortexm0ds_logic.v(1077)
  wire Z7niu6;  // ../RTL/cortexm0ds_logic.v(614)
  wire Z7oow6;  // ../RTL/cortexm0ds_logic.v(1170)
  wire Z7tpw6;  // ../RTL/cortexm0ds_logic.v(1605)
  wire Z7uiu6;  // ../RTL/cortexm0ds_logic.v(707)
  wire Z7vhu6;  // ../RTL/cortexm0ds_logic.v(239)
  wire Z7vow6;  // ../RTL/cortexm0ds_logic.v(1264)
  wire Z80ju6;  // ../RTL/cortexm0ds_logic.v(788)
  wire Z81iu6;  // ../RTL/cortexm0ds_logic.v(320)
  wire Z81pw6;  // ../RTL/cortexm0ds_logic.v(1344)
  wire Z87ju6;  // ../RTL/cortexm0ds_logic.v(882)
  wire Z88iu6;  // ../RTL/cortexm0ds_logic.v(414)
  wire Z88pw6;  // ../RTL/cortexm0ds_logic.v(1438)
  wire Z89ow6;  // ../RTL/cortexm0ds_logic.v(970)
  wire Z8fiu6;  // ../RTL/cortexm0ds_logic.v(507)
  wire Z8gow6;  // ../RTL/cortexm0ds_logic.v(1064)
  wire Z8jpw6;  // ../RTL/cortexm0ds_logic.v(1586)
  wire Z8miu6;  // ../RTL/cortexm0ds_logic.v(601)
  wire Z8now6;  // ../RTL/cortexm0ds_logic.v(1157)
  wire Z8tiu6;  // ../RTL/cortexm0ds_logic.v(694)
  wire Z8uhu6;  // ../RTL/cortexm0ds_logic.v(226)
  wire Z8uow6;  // ../RTL/cortexm0ds_logic.v(1251)
  wire Z8zpw6;  // ../RTL/cortexm0ds_logic.v(1616)
  wire Z90iu6;  // ../RTL/cortexm0ds_logic.v(307)
  wire Z90pw6;  // ../RTL/cortexm0ds_logic.v(1331)
  wire Z96ju6;  // ../RTL/cortexm0ds_logic.v(869)
  wire Z97iu6;  // ../RTL/cortexm0ds_logic.v(401)
  wire Z97pw6;  // ../RTL/cortexm0ds_logic.v(1425)
  wire Z98bx6;  // ../RTL/cortexm0ds_logic.v(1694)
  wire Z98ow6;  // ../RTL/cortexm0ds_logic.v(957)
  wire Z9abx6;  // ../RTL/cortexm0ds_logic.v(1698)
  wire Z9eiu6;  // ../RTL/cortexm0ds_logic.v(494)
  wire Z9fow6;  // ../RTL/cortexm0ds_logic.v(1051)
  wire Z9liu6;  // ../RTL/cortexm0ds_logic.v(588)
  wire Z9mow6;  // ../RTL/cortexm0ds_logic.v(1144)
  wire Z9opw6;  // ../RTL/cortexm0ds_logic.v(1596)
  wire Z9siu6;  // ../RTL/cortexm0ds_logic.v(681)
  wire Z9thu6;  // ../RTL/cortexm0ds_logic.v(213)
  wire Z9tow6;  // ../RTL/cortexm0ds_logic.v(1238)
  wire Z9tpw6;  // ../RTL/cortexm0ds_logic.v(1605)
  wire Z9ziu6;  // ../RTL/cortexm0ds_logic.v(775)
  wire Za5ju6;  // ../RTL/cortexm0ds_logic.v(856)
  wire Za6iu6;  // ../RTL/cortexm0ds_logic.v(388)
  wire Za6pw6;  // ../RTL/cortexm0ds_logic.v(1412)
  wire Za7ow6;  // ../RTL/cortexm0ds_logic.v(944)
  wire Zadiu6;  // ../RTL/cortexm0ds_logic.v(481)
  wire Zadpw6;  // ../RTL/cortexm0ds_logic.v(1506)
  wire Zaeow6;  // ../RTL/cortexm0ds_logic.v(1038)
  wire Zakiu6;  // ../RTL/cortexm0ds_logic.v(575)
  wire Zalow6;  // ../RTL/cortexm0ds_logic.v(1131)
  wire Zariu6;  // ../RTL/cortexm0ds_logic.v(668)
  wire Zashu6;  // ../RTL/cortexm0ds_logic.v(200)
  wire Zasow6;  // ../RTL/cortexm0ds_logic.v(1225)
  wire Zayiu6;  // ../RTL/cortexm0ds_logic.v(762)
  wire Zazhu6;  // ../RTL/cortexm0ds_logic.v(294)
  wire Zazow6;  // ../RTL/cortexm0ds_logic.v(1318)
  wire Zazpw6;  // ../RTL/cortexm0ds_logic.v(1616)
  wire Zb4ju6;  // ../RTL/cortexm0ds_logic.v(843)
  wire Zb5iu6;  // ../RTL/cortexm0ds_logic.v(375)
  wire Zb5pw6;  // ../RTL/cortexm0ds_logic.v(1399)
  wire Zb6ow6;  // ../RTL/cortexm0ds_logic.v(931)
  wire Zb8bx6;  // ../RTL/cortexm0ds_logic.v(1694)
  wire Zbciu6;  // ../RTL/cortexm0ds_logic.v(468)
  wire Zbcpw6;  // ../RTL/cortexm0ds_logic.v(1493)
  wire Zbdow6;  // ../RTL/cortexm0ds_logic.v(1025)
  wire Zbjiu6;  // ../RTL/cortexm0ds_logic.v(562)
  wire Zbkow6;  // ../RTL/cortexm0ds_logic.v(1118)
  wire Zbmhu6;  // ../RTL/cortexm0ds_logic.v(142)
  wire Zbqiu6;  // ../RTL/cortexm0ds_logic.v(655)
  wire Zbrhu6;  // ../RTL/cortexm0ds_logic.v(187)
  wire Zbrow6;  // ../RTL/cortexm0ds_logic.v(1212)
  wire Zbtpw6;  // ../RTL/cortexm0ds_logic.v(1605)
  wire Zbxiu6;  // ../RTL/cortexm0ds_logic.v(749)
  wire Zbyhu6;  // ../RTL/cortexm0ds_logic.v(281)
  wire Zbyow6;  // ../RTL/cortexm0ds_logic.v(1305)
  wire Zc3ju6;  // ../RTL/cortexm0ds_logic.v(830)
  wire Zc4iu6;  // ../RTL/cortexm0ds_logic.v(362)
  wire Zc4pw6;  // ../RTL/cortexm0ds_logic.v(1386)
  wire Zcaju6;  // ../RTL/cortexm0ds_logic.v(923)
  wire Zcbiu6;  // ../RTL/cortexm0ds_logic.v(455)
  wire Zcbpw6;  // ../RTL/cortexm0ds_logic.v(1480)
  wire Zccow6;  // ../RTL/cortexm0ds_logic.v(1012)
  wire Zciiu6;  // ../RTL/cortexm0ds_logic.v(549)
  wire Zcjow6;  // ../RTL/cortexm0ds_logic.v(1105)
  wire Zcpiu6;  // ../RTL/cortexm0ds_logic.v(642)
  wire Zcqhu6;  // ../RTL/cortexm0ds_logic.v(174)
  wire Zcqow6;  // ../RTL/cortexm0ds_logic.v(1199)
  wire Zcwiu6;  // ../RTL/cortexm0ds_logic.v(736)
  wire Zcxhu6;  // ../RTL/cortexm0ds_logic.v(268)
  wire Zcxow6;  // ../RTL/cortexm0ds_logic.v(1292)
  wire Zczpw6;  // ../RTL/cortexm0ds_logic.v(1616)
  wire Zd2ju6;  // ../RTL/cortexm0ds_logic.v(817)
  wire Zd3iu6;  // ../RTL/cortexm0ds_logic.v(349)
  wire Zd3pw6;  // ../RTL/cortexm0ds_logic.v(1373)
  wire Zd8bx6;  // ../RTL/cortexm0ds_logic.v(1694)
  wire Zd9ju6;  // ../RTL/cortexm0ds_logic.v(910)
  wire Zdaiu6;  // ../RTL/cortexm0ds_logic.v(442)
  wire Zdapw6;  // ../RTL/cortexm0ds_logic.v(1467)
  wire Zdbow6;  // ../RTL/cortexm0ds_logic.v(999)
  wire Zdcbx6;  // ../RTL/cortexm0ds_logic.v(1701)
  wire Zdhax6;  // ../RTL/cortexm0ds_logic.v(1646)
  wire Zdhiu6;  // ../RTL/cortexm0ds_logic.v(536)
  wire Zdiax6;  // ../RTL/cortexm0ds_logic.v(1647)
  wire Zdiow6;  // ../RTL/cortexm0ds_logic.v(1092)
  wire Zdoiu6;  // ../RTL/cortexm0ds_logic.v(629)
  wire Zdphu6;  // ../RTL/cortexm0ds_logic.v(161)
  wire Zdpow6;  // ../RTL/cortexm0ds_logic.v(1186)
  wire Zdtpw6;  // ../RTL/cortexm0ds_logic.v(1605)
  wire Zduax6;  // ../RTL/cortexm0ds_logic.v(1669)
  wire Zdviu6;  // ../RTL/cortexm0ds_logic.v(723)
  wire Zdwhu6;  // ../RTL/cortexm0ds_logic.v(255)
  wire Zdwow6;  // ../RTL/cortexm0ds_logic.v(1279)
  wire Ze1ju6;  // ../RTL/cortexm0ds_logic.v(804)
  wire Ze2iu6;  // ../RTL/cortexm0ds_logic.v(336)
  wire Ze2pw6;  // ../RTL/cortexm0ds_logic.v(1360)
  wire Ze8ju6;  // ../RTL/cortexm0ds_logic.v(897)
  wire Ze9iu6;  // ../RTL/cortexm0ds_logic.v(429)
  wire Ze9pw6;  // ../RTL/cortexm0ds_logic.v(1454)
  wire Zeaow6;  // ../RTL/cortexm0ds_logic.v(986)
  wire Zegiu6;  // ../RTL/cortexm0ds_logic.v(523)
  wire Zehow6;  // ../RTL/cortexm0ds_logic.v(1079)
  wire Zelhu6;  // ../RTL/cortexm0ds_logic.v(139)
  wire Zeniu6;  // ../RTL/cortexm0ds_logic.v(616)
  wire Zeohu6;  // ../RTL/cortexm0ds_logic.v(148)
  wire Zeoow6;  // ../RTL/cortexm0ds_logic.v(1173)
  wire Zeuiu6;  // ../RTL/cortexm0ds_logic.v(710)
  wire Zevhu6;  // ../RTL/cortexm0ds_logic.v(242)
  wire Zevow6;  // ../RTL/cortexm0ds_logic.v(1266)
  wire Zezpw6;  // ../RTL/cortexm0ds_logic.v(1616)
  wire Zf0ju6;  // ../RTL/cortexm0ds_logic.v(791)
  wire Zf1iu6;  // ../RTL/cortexm0ds_logic.v(323)
  wire Zf1pw6;  // ../RTL/cortexm0ds_logic.v(1347)
  wire Zf7ju6;  // ../RTL/cortexm0ds_logic.v(884)
  wire Zf8bx6;  // ../RTL/cortexm0ds_logic.v(1694)
  wire Zf8iu6;  // ../RTL/cortexm0ds_logic.v(416)
  wire Zf8pw6;  // ../RTL/cortexm0ds_logic.v(1441)
  wire Zf9ow6;  // ../RTL/cortexm0ds_logic.v(973)
  wire Zffiu6;  // ../RTL/cortexm0ds_logic.v(510)
  wire Zfgow6;  // ../RTL/cortexm0ds_logic.v(1066)
  wire Zfmiu6;  // ../RTL/cortexm0ds_logic.v(603)
  wire Zfnow6;  // ../RTL/cortexm0ds_logic.v(1160)
  wire Zftiu6;  // ../RTL/cortexm0ds_logic.v(697)
  wire Zfuhu6;  // ../RTL/cortexm0ds_logic.v(229)
  wire Zfuow6;  // ../RTL/cortexm0ds_logic.v(1253)
  wire Zg0iu6;  // ../RTL/cortexm0ds_logic.v(310)
  wire Zg0pw6;  // ../RTL/cortexm0ds_logic.v(1334)
  wire Zg6ju6;  // ../RTL/cortexm0ds_logic.v(871)
  wire Zg7iu6;  // ../RTL/cortexm0ds_logic.v(403)
  wire Zg7pw6;  // ../RTL/cortexm0ds_logic.v(1428)
  wire Zg8ow6;  // ../RTL/cortexm0ds_logic.v(960)
  wire Zgbax6;  // ../RTL/cortexm0ds_logic.v(1634)
  wire Zgeiu6;  // ../RTL/cortexm0ds_logic.v(497)
  wire Zgfax6;  // ../RTL/cortexm0ds_logic.v(1642)
  wire Zgfow6;  // ../RTL/cortexm0ds_logic.v(1053)
  wire Zgliu6;  // ../RTL/cortexm0ds_logic.v(590)
  wire Zgmow6;  // ../RTL/cortexm0ds_logic.v(1147)
  wire Zgsiu6;  // ../RTL/cortexm0ds_logic.v(684)
  wire Zgthu6;  // ../RTL/cortexm0ds_logic.v(216)
  wire Zgtow6;  // ../RTL/cortexm0ds_logic.v(1240)
  wire Zgziu6;  // ../RTL/cortexm0ds_logic.v(778)
  wire Zgzpw6;  // ../RTL/cortexm0ds_logic.v(1616)
  wire Zh5ju6;  // ../RTL/cortexm0ds_logic.v(858)
  wire Zh6iu6;  // ../RTL/cortexm0ds_logic.v(390)
  wire Zh6pw6;  // ../RTL/cortexm0ds_logic.v(1415)
  wire Zh7ow6;  // ../RTL/cortexm0ds_logic.v(947)
  wire Zh8bx6;  // ../RTL/cortexm0ds_logic.v(1694)
  wire Zhdiu6;  // ../RTL/cortexm0ds_logic.v(484)
  wire Zhdpw6;  // ../RTL/cortexm0ds_logic.v(1508)
  wire Zheow6;  // ../RTL/cortexm0ds_logic.v(1040)
  wire Zhkiu6;  // ../RTL/cortexm0ds_logic.v(577)
  wire Zhlow6;  // ../RTL/cortexm0ds_logic.v(1134)
  wire Zhriu6;  // ../RTL/cortexm0ds_logic.v(671)
  wire Zhshu6;  // ../RTL/cortexm0ds_logic.v(203)
  wire Zhsow6;  // ../RTL/cortexm0ds_logic.v(1227)
  wire Zhyiu6;  // ../RTL/cortexm0ds_logic.v(765)
  wire Zhzhu6;  // ../RTL/cortexm0ds_logic.v(297)
  wire Zhzow6;  // ../RTL/cortexm0ds_logic.v(1321)
  wire Zi4ju6;  // ../RTL/cortexm0ds_logic.v(845)
  wire Zi5iu6;  // ../RTL/cortexm0ds_logic.v(377)
  wire Zi5pw6;  // ../RTL/cortexm0ds_logic.v(1402)
  wire Zi6ow6;  // ../RTL/cortexm0ds_logic.v(934)
  wire Ziciu6;  // ../RTL/cortexm0ds_logic.v(471)
  wire Zicpw6;  // ../RTL/cortexm0ds_logic.v(1495)
  wire Zidow6;  // ../RTL/cortexm0ds_logic.v(1027)
  wire Zijiu6;  // ../RTL/cortexm0ds_logic.v(564)
  wire Zikow6;  // ../RTL/cortexm0ds_logic.v(1121)
  wire Ziqiu6;  // ../RTL/cortexm0ds_logic.v(658)
  wire Zirhu6;  // ../RTL/cortexm0ds_logic.v(190)
  wire Zirow6;  // ../RTL/cortexm0ds_logic.v(1214)
  wire Zixiu6;  // ../RTL/cortexm0ds_logic.v(752)
  wire Ziyhu6;  // ../RTL/cortexm0ds_logic.v(284)
  wire Ziyow6;  // ../RTL/cortexm0ds_logic.v(1308)
  wire Zj3ju6;  // ../RTL/cortexm0ds_logic.v(832)
  wire Zj4iu6;  // ../RTL/cortexm0ds_logic.v(364)
  wire Zj4pw6;  // ../RTL/cortexm0ds_logic.v(1389)
  wire Zj8bx6;  // ../RTL/cortexm0ds_logic.v(1694)
  wire Zjaju6;  // ../RTL/cortexm0ds_logic.v(926)
  wire Zjbiu6;  // ../RTL/cortexm0ds_logic.v(458)
  wire Zjbpw6;  // ../RTL/cortexm0ds_logic.v(1482)
  wire Zjcow6;  // ../RTL/cortexm0ds_logic.v(1014)
  wire Zjiiu6;  // ../RTL/cortexm0ds_logic.v(551)
  wire Zjjow6;  // ../RTL/cortexm0ds_logic.v(1108)
  wire Zjpiu6;  // ../RTL/cortexm0ds_logic.v(645)
  wire Zjqhu6;  // ../RTL/cortexm0ds_logic.v(177)
  wire Zjqow6;  // ../RTL/cortexm0ds_logic.v(1201)
  wire Zjwiu6;  // ../RTL/cortexm0ds_logic.v(739)
  wire Zjxhu6;  // ../RTL/cortexm0ds_logic.v(271)
  wire Zjxow6;  // ../RTL/cortexm0ds_logic.v(1295)
  wire Zk2ju6;  // ../RTL/cortexm0ds_logic.v(819)
  wire Zk3iu6;  // ../RTL/cortexm0ds_logic.v(351)
  wire Zk3pw6;  // ../RTL/cortexm0ds_logic.v(1376)
  wire Zk9ju6;  // ../RTL/cortexm0ds_logic.v(913)
  wire Zkaiu6;  // ../RTL/cortexm0ds_logic.v(445)
  wire Zkapw6;  // ../RTL/cortexm0ds_logic.v(1469)
  wire Zkbow6;  // ../RTL/cortexm0ds_logic.v(1001)
  wire Zkhiu6;  // ../RTL/cortexm0ds_logic.v(538)
  wire Zkiow6;  // ../RTL/cortexm0ds_logic.v(1095)
  wire Zkoiu6;  // ../RTL/cortexm0ds_logic.v(632)
  wire Zkphu6;  // ../RTL/cortexm0ds_logic.v(164)
  wire Zkpow6;  // ../RTL/cortexm0ds_logic.v(1188)
  wire Zkviu6;  // ../RTL/cortexm0ds_logic.v(726)
  wire Zkwhu6;  // ../RTL/cortexm0ds_logic.v(258)
  wire Zkwow6;  // ../RTL/cortexm0ds_logic.v(1282)
  wire Zl1ju6;  // ../RTL/cortexm0ds_logic.v(806)
  wire Zl2iu6;  // ../RTL/cortexm0ds_logic.v(338)
  wire Zl2pw6;  // ../RTL/cortexm0ds_logic.v(1363)
  wire Zl8bx6;  // ../RTL/cortexm0ds_logic.v(1694)
  wire Zl8ju6;  // ../RTL/cortexm0ds_logic.v(900)
  wire Zl9bx6;  // ../RTL/cortexm0ds_logic.v(1696)
  wire Zl9pw6;  // ../RTL/cortexm0ds_logic.v(1456)
  wire Zlaow6;  // ../RTL/cortexm0ds_logic.v(988)
  wire Zlghu6;  // ../RTL/cortexm0ds_logic.v(126)
  wire Zlgiu6;  // ../RTL/cortexm0ds_logic.v(525)
  wire Zlhow6;  // ../RTL/cortexm0ds_logic.v(1082)
  wire Zlniu6;  // ../RTL/cortexm0ds_logic.v(619)
  wire Zlohu6;  // ../RTL/cortexm0ds_logic.v(151)
  wire Zloow6;  // ../RTL/cortexm0ds_logic.v(1175)
  wire Zluiu6;  // ../RTL/cortexm0ds_logic.v(713)
  wire Zlvhu6;  // ../RTL/cortexm0ds_logic.v(245)
  wire Zlvow6;  // ../RTL/cortexm0ds_logic.v(1269)
  wire Zm0ju6;  // ../RTL/cortexm0ds_logic.v(793)
  wire Zm1iu6;  // ../RTL/cortexm0ds_logic.v(325)
  wire Zm1pw6;  // ../RTL/cortexm0ds_logic.v(1350)
  wire Zm7ju6;  // ../RTL/cortexm0ds_logic.v(887)
  wire Zm8ax6;  // ../RTL/cortexm0ds_logic.v(1629)
  wire Zm8iu6;  // ../RTL/cortexm0ds_logic.v(419)
  wire Zm8pw6;  // ../RTL/cortexm0ds_logic.v(1443)
  wire Zm9ow6;  // ../RTL/cortexm0ds_logic.v(975)
  wire Zmfiu6;  // ../RTL/cortexm0ds_logic.v(512)
  wire Zmgow6;  // ../RTL/cortexm0ds_logic.v(1069)
  wire Zmmiu6;  // ../RTL/cortexm0ds_logic.v(606)
  wire Zmnow6;  // ../RTL/cortexm0ds_logic.v(1162)
  wire Zmtiu6;  // ../RTL/cortexm0ds_logic.v(700)
  wire Zmuhu6;  // ../RTL/cortexm0ds_logic.v(232)
  wire Zmuow6;  // ../RTL/cortexm0ds_logic.v(1256)
  wire Zn0iu6;  // ../RTL/cortexm0ds_logic.v(312)
  wire Zn0pw6;  // ../RTL/cortexm0ds_logic.v(1337)
  wire Zn6ju6;  // ../RTL/cortexm0ds_logic.v(874)
  wire Zn7iu6;  // ../RTL/cortexm0ds_logic.v(406)
  wire Zn7pw6;  // ../RTL/cortexm0ds_logic.v(1430)
  wire Zn8bx6;  // ../RTL/cortexm0ds_logic.v(1695)
  wire Zn8ow6;  // ../RTL/cortexm0ds_logic.v(962)
  wire Zneiu6;  // ../RTL/cortexm0ds_logic.v(499)
  wire Znfow6;  // ../RTL/cortexm0ds_logic.v(1056)
  wire Znliu6;  // ../RTL/cortexm0ds_logic.v(593)
  wire Znmow6;  // ../RTL/cortexm0ds_logic.v(1149)
  wire Znsiu6;  // ../RTL/cortexm0ds_logic.v(687)
  wire Znthu6;  // ../RTL/cortexm0ds_logic.v(219)
  wire Zntow6;  // ../RTL/cortexm0ds_logic.v(1243)
  wire Znziu6;  // ../RTL/cortexm0ds_logic.v(780)
  wire Zo5ju6;  // ../RTL/cortexm0ds_logic.v(861)
  wire Zo6iu6;  // ../RTL/cortexm0ds_logic.v(393)
  wire Zo6pw6;  // ../RTL/cortexm0ds_logic.v(1417)
  wire Zo7ow6;  // ../RTL/cortexm0ds_logic.v(949)
  wire Zodbx6;  // ../RTL/cortexm0ds_logic.v(1704)
  wire Zodiu6;  // ../RTL/cortexm0ds_logic.v(486)
  wire Zodpw6;  // ../RTL/cortexm0ds_logic.v(1511)
  wire Zoeow6;  // ../RTL/cortexm0ds_logic.v(1043)
  wire Zokiu6;  // ../RTL/cortexm0ds_logic.v(580)
  wire Zolow6;  // ../RTL/cortexm0ds_logic.v(1136)
  wire Zoriu6;  // ../RTL/cortexm0ds_logic.v(674)
  wire Zoshu6;  // ../RTL/cortexm0ds_logic.v(206)
  wire Zosow6;  // ../RTL/cortexm0ds_logic.v(1230)
  wire Zoyiu6;  // ../RTL/cortexm0ds_logic.v(767)
  wire Zozhu6;  // ../RTL/cortexm0ds_logic.v(299)
  wire Zozow6;  // ../RTL/cortexm0ds_logic.v(1324)
  wire Zp4ju6;  // ../RTL/cortexm0ds_logic.v(848)
  wire Zp5iu6;  // ../RTL/cortexm0ds_logic.v(380)
  wire Zp5pw6;  // ../RTL/cortexm0ds_logic.v(1404)
  wire Zp6ow6;  // ../RTL/cortexm0ds_logic.v(936)
  wire Zp8bx6;  // ../RTL/cortexm0ds_logic.v(1695)
  wire Zpciu6;  // ../RTL/cortexm0ds_logic.v(473)
  wire Zpcpw6;  // ../RTL/cortexm0ds_logic.v(1498)
  wire Zpdow6;  // ../RTL/cortexm0ds_logic.v(1030)
  wire Zpjiu6;  // ../RTL/cortexm0ds_logic.v(567)
  wire Zpkow6;  // ../RTL/cortexm0ds_logic.v(1123)
  wire Zpqiu6;  // ../RTL/cortexm0ds_logic.v(661)
  wire Zprhu6;  // ../RTL/cortexm0ds_logic.v(193)
  wire Zprow6;  // ../RTL/cortexm0ds_logic.v(1217)
  wire Zpxiu6;  // ../RTL/cortexm0ds_logic.v(754)
  wire Zpyhu6;  // ../RTL/cortexm0ds_logic.v(286)
  wire Zpyow6;  // ../RTL/cortexm0ds_logic.v(1311)
  wire Zq3ju6;  // ../RTL/cortexm0ds_logic.v(835)
  wire Zq4iu6;  // ../RTL/cortexm0ds_logic.v(367)
  wire Zq4pw6;  // ../RTL/cortexm0ds_logic.v(1391)
  wire Zqaju6;  // ../RTL/cortexm0ds_logic.v(928)
  wire Zqbiu6;  // ../RTL/cortexm0ds_logic.v(460)
  wire Zqbpw6;  // ../RTL/cortexm0ds_logic.v(1485)
  wire Zqcow6;  // ../RTL/cortexm0ds_logic.v(1017)
  wire Zqiax6;  // ../RTL/cortexm0ds_logic.v(1648)
  wire Zqiiu6;  // ../RTL/cortexm0ds_logic.v(554)
  wire Zqjow6;  // ../RTL/cortexm0ds_logic.v(1110)
  wire Zqpiu6;  // ../RTL/cortexm0ds_logic.v(648)
  wire Zqqhu6;  // ../RTL/cortexm0ds_logic.v(180)
  wire Zqqow6;  // ../RTL/cortexm0ds_logic.v(1204)
  wire Zqwiu6;  // ../RTL/cortexm0ds_logic.v(741)
  wire Zqxhu6;  // ../RTL/cortexm0ds_logic.v(273)
  wire Zqxow6;  // ../RTL/cortexm0ds_logic.v(1298)
  wire Zr2ju6;  // ../RTL/cortexm0ds_logic.v(822)
  wire Zr3iu6;  // ../RTL/cortexm0ds_logic.v(354)
  wire Zr3pw6;  // ../RTL/cortexm0ds_logic.v(1378)
  wire Zr7bx6;  // ../RTL/cortexm0ds_logic.v(1693)
  wire Zr8bx6;  // ../RTL/cortexm0ds_logic.v(1695)
  wire Zr9ju6;  // ../RTL/cortexm0ds_logic.v(915)
  wire Zraiu6;  // ../RTL/cortexm0ds_logic.v(447)
  wire Zrapw6;  // ../RTL/cortexm0ds_logic.v(1472)
  wire Zrbow6;  // ../RTL/cortexm0ds_logic.v(1004)
  wire Zrhiu6;  // ../RTL/cortexm0ds_logic.v(541)
  wire Zriow6;  // ../RTL/cortexm0ds_logic.v(1097)
  wire Zrlax6;  // ../RTL/cortexm0ds_logic.v(1654)
  wire Zroiu6;  // ../RTL/cortexm0ds_logic.v(635)
  wire Zrphu6;  // ../RTL/cortexm0ds_logic.v(167)
  wire Zrpow6;  // ../RTL/cortexm0ds_logic.v(1191)
  wire Zrviu6;  // ../RTL/cortexm0ds_logic.v(728)
  wire Zrwhu6;  // ../RTL/cortexm0ds_logic.v(260)
  wire Zrwow6;  // ../RTL/cortexm0ds_logic.v(1285)
  wire Zs1ju6;  // ../RTL/cortexm0ds_logic.v(809)
  wire Zs2iu6;  // ../RTL/cortexm0ds_logic.v(341)
  wire Zs2pw6;  // ../RTL/cortexm0ds_logic.v(1365)
  wire Zs8ju6;  // ../RTL/cortexm0ds_logic.v(902)
  wire Zs9iu6;  // ../RTL/cortexm0ds_logic.v(434)
  wire Zs9pw6;  // ../RTL/cortexm0ds_logic.v(1459)
  wire Zsaow6;  // ../RTL/cortexm0ds_logic.v(991)
  wire Zsgiu6;  // ../RTL/cortexm0ds_logic.v(528)
  wire Zshax6;  // ../RTL/cortexm0ds_logic.v(1646)
  wire Zshow6;  // ../RTL/cortexm0ds_logic.v(1084)
  wire Zslpw6;  // ../RTL/cortexm0ds_logic.v(1591)
  wire Zsniu6;  // ../RTL/cortexm0ds_logic.v(622)
  wire Zsohu6;  // ../RTL/cortexm0ds_logic.v(154)
  wire Zsoow6;  // ../RTL/cortexm0ds_logic.v(1178)
  wire Zsuiu6;  // ../RTL/cortexm0ds_logic.v(715)
  wire Zsvhu6;  // ../RTL/cortexm0ds_logic.v(247)
  wire Zsvow6;  // ../RTL/cortexm0ds_logic.v(1272)
  wire Zszax6;  // ../RTL/cortexm0ds_logic.v(1679)
  wire Zt0ju6;  // ../RTL/cortexm0ds_logic.v(796)
  wire Zt1iu6;  // ../RTL/cortexm0ds_logic.v(328)
  wire Zt1pw6;  // ../RTL/cortexm0ds_logic.v(1352)
  wire Zt7bx6;  // ../RTL/cortexm0ds_logic.v(1693)
  wire Zt7ju6;  // ../RTL/cortexm0ds_logic.v(889)
  wire Zt8iu6;  // ../RTL/cortexm0ds_logic.v(421)
  wire Zt8pw6;  // ../RTL/cortexm0ds_logic.v(1446)
  wire Zt9ow6;  // ../RTL/cortexm0ds_logic.v(978)
  wire Ztfiu6;  // ../RTL/cortexm0ds_logic.v(515)
  wire Ztgbx6;  // ../RTL/cortexm0ds_logic.v(1710)
  wire Ztgow6;  // ../RTL/cortexm0ds_logic.v(1071)
  wire Ztmiu6;  // ../RTL/cortexm0ds_logic.v(609)
  wire Ztnow6;  // ../RTL/cortexm0ds_logic.v(1165)
  wire Zttiu6;  // ../RTL/cortexm0ds_logic.v(702)
  wire Ztuhu6;  // ../RTL/cortexm0ds_logic.v(234)
  wire Ztuow6;  // ../RTL/cortexm0ds_logic.v(1259)
  wire Ztupw6;  // ../RTL/cortexm0ds_logic.v(1607)
  wire Zu0iu6;  // ../RTL/cortexm0ds_logic.v(315)
  wire Zu0pw6;  // ../RTL/cortexm0ds_logic.v(1339)
  wire Zu6ju6;  // ../RTL/cortexm0ds_logic.v(876)
  wire Zu7iu6;  // ../RTL/cortexm0ds_logic.v(408)
  wire Zu7pw6;  // ../RTL/cortexm0ds_logic.v(1433)
  wire Zu8ow6;  // ../RTL/cortexm0ds_logic.v(965)
  wire Zueiu6;  // ../RTL/cortexm0ds_logic.v(502)
  wire Zufow6;  // ../RTL/cortexm0ds_logic.v(1058)
  wire Zuliu6;  // ../RTL/cortexm0ds_logic.v(596)
  wire Zumow6;  // ../RTL/cortexm0ds_logic.v(1152)
  wire Zusiu6;  // ../RTL/cortexm0ds_logic.v(689)
  wire Zuthu6;  // ../RTL/cortexm0ds_logic.v(221)
  wire Zutow6;  // ../RTL/cortexm0ds_logic.v(1246)
  wire Zuziu6;  // ../RTL/cortexm0ds_logic.v(783)
  wire Zv5ju6;  // ../RTL/cortexm0ds_logic.v(863)
  wire Zv6iu6;  // ../RTL/cortexm0ds_logic.v(395)
  wire Zv6pw6;  // ../RTL/cortexm0ds_logic.v(1420)
  wire Zv7bx6;  // ../RTL/cortexm0ds_logic.v(1693)
  wire Zv7ow6;  // ../RTL/cortexm0ds_logic.v(952)
  wire Zvdiu6;  // ../RTL/cortexm0ds_logic.v(489)
  wire Zvdpw6;  // ../RTL/cortexm0ds_logic.v(1513)
  wire Zveow6;  // ../RTL/cortexm0ds_logic.v(1045)
  wire Zvgbx6;  // ../RTL/cortexm0ds_logic.v(1710)
  wire Zvkiu6;  // ../RTL/cortexm0ds_logic.v(583)
  wire Zvlow6;  // ../RTL/cortexm0ds_logic.v(1139)
  wire Zvriu6;  // ../RTL/cortexm0ds_logic.v(676)
  wire Zvrpw6;  // ../RTL/cortexm0ds_logic.v(1602)
  wire Zvshu6;  // ../RTL/cortexm0ds_logic.v(208)
  wire Zvsow6;  // ../RTL/cortexm0ds_logic.v(1233)
  wire Zvyiu6;  // ../RTL/cortexm0ds_logic.v(770)
  wire Zvzhu6;  // ../RTL/cortexm0ds_logic.v(302)
  wire Zvzow6;  // ../RTL/cortexm0ds_logic.v(1326)
  wire Zw4ju6;  // ../RTL/cortexm0ds_logic.v(850)
  wire Zw5iu6;  // ../RTL/cortexm0ds_logic.v(382)
  wire Zw5pw6;  // ../RTL/cortexm0ds_logic.v(1407)
  wire Zw6ow6;  // ../RTL/cortexm0ds_logic.v(939)
  wire Zwciu6;  // ../RTL/cortexm0ds_logic.v(476)
  wire Zwcpw6;  // ../RTL/cortexm0ds_logic.v(1500)
  wire Zwdow6;  // ../RTL/cortexm0ds_logic.v(1032)
  wire Zwjiu6;  // ../RTL/cortexm0ds_logic.v(570)
  wire Zwkow6;  // ../RTL/cortexm0ds_logic.v(1126)
  wire Zwnpw6;  // ../RTL/cortexm0ds_logic.v(1595)
  wire Zwqiu6;  // ../RTL/cortexm0ds_logic.v(663)
  wire Zwrhu6;  // ../RTL/cortexm0ds_logic.v(195)
  wire Zwrow6;  // ../RTL/cortexm0ds_logic.v(1220)
  wire Zwxiu6;  // ../RTL/cortexm0ds_logic.v(757)
  wire Zwyhu6;  // ../RTL/cortexm0ds_logic.v(289)
  wire Zwyow6;  // ../RTL/cortexm0ds_logic.v(1313)
  wire Zx3ju6;  // ../RTL/cortexm0ds_logic.v(837)
  wire Zx4iu6;  // ../RTL/cortexm0ds_logic.v(369)
  wire Zx4pw6;  // ../RTL/cortexm0ds_logic.v(1394)
  wire Zx7bx6;  // ../RTL/cortexm0ds_logic.v(1693)
  wire Zx8ax6;  // ../RTL/cortexm0ds_logic.v(1629)
  wire Zxbiu6;  // ../RTL/cortexm0ds_logic.v(463)
  wire Zxbpw6;  // ../RTL/cortexm0ds_logic.v(1487)
  wire Zxcow6;  // ../RTL/cortexm0ds_logic.v(1019)
  wire Zxiiu6;  // ../RTL/cortexm0ds_logic.v(557)
  wire Zxjow6;  // ../RTL/cortexm0ds_logic.v(1113)
  wire Zxpiu6;  // ../RTL/cortexm0ds_logic.v(650)
  wire Zxqhu6;  // ../RTL/cortexm0ds_logic.v(182)
  wire Zxqow6;  // ../RTL/cortexm0ds_logic.v(1207)
  wire Zxwiu6;  // ../RTL/cortexm0ds_logic.v(744)
  wire Zxxhu6;  // ../RTL/cortexm0ds_logic.v(276)
  wire Zxxow6;  // ../RTL/cortexm0ds_logic.v(1300)
  wire Zy2ju6;  // ../RTL/cortexm0ds_logic.v(824)
  wire Zy3iu6;  // ../RTL/cortexm0ds_logic.v(356)
  wire Zy3pw6;  // ../RTL/cortexm0ds_logic.v(1381)
  wire Zy9ju6;  // ../RTL/cortexm0ds_logic.v(918)
  wire Zyaiu6;  // ../RTL/cortexm0ds_logic.v(450)
  wire Zyapw6;  // ../RTL/cortexm0ds_logic.v(1474)
  wire Zybow6;  // ../RTL/cortexm0ds_logic.v(1006)
  wire Zycbx6;  // ../RTL/cortexm0ds_logic.v(1703)
  wire Zyhiu6;  // ../RTL/cortexm0ds_logic.v(544)
  wire Zyiow6;  // ../RTL/cortexm0ds_logic.v(1100)
  wire Zyoiu6;  // ../RTL/cortexm0ds_logic.v(637)
  wire Zyphu6;  // ../RTL/cortexm0ds_logic.v(169)
  wire Zypow6;  // ../RTL/cortexm0ds_logic.v(1194)
  wire Zyviu6;  // ../RTL/cortexm0ds_logic.v(731)
  wire Zywhu6;  // ../RTL/cortexm0ds_logic.v(263)
  wire Zywow6;  // ../RTL/cortexm0ds_logic.v(1287)
  wire Zz1ju6;  // ../RTL/cortexm0ds_logic.v(811)
  wire Zz2iu6;  // ../RTL/cortexm0ds_logic.v(343)
  wire Zz2pw6;  // ../RTL/cortexm0ds_logic.v(1368)
  wire Zz7bx6;  // ../RTL/cortexm0ds_logic.v(1693)
  wire Zz8ju6;  // ../RTL/cortexm0ds_logic.v(905)
  wire Zz9iu6;  // ../RTL/cortexm0ds_logic.v(437)
  wire Zz9pw6;  // ../RTL/cortexm0ds_logic.v(1461)
  wire Zzaow6;  // ../RTL/cortexm0ds_logic.v(993)
  wire Zzgiu6;  // ../RTL/cortexm0ds_logic.v(531)
  wire Zzhow6;  // ../RTL/cortexm0ds_logic.v(1087)
  wire Zzniu6;  // ../RTL/cortexm0ds_logic.v(624)
  wire Zzohu6;  // ../RTL/cortexm0ds_logic.v(156)
  wire Zzoow6;  // ../RTL/cortexm0ds_logic.v(1181)
  wire Zzuiu6;  // ../RTL/cortexm0ds_logic.v(718)
  wire Zzvhu6;  // ../RTL/cortexm0ds_logic.v(250)
  wire Zzvow6;  // ../RTL/cortexm0ds_logic.v(1274)
  wire n0;
  wire n1;
  wire n10;
  wire n100;
  wire n1000;
  wire n1001;
  wire n1002;
  wire n1003;
  wire n1004;
  wire n1005;
  wire n1006;
  wire n1007;
  wire n1008;
  wire n1009;
  wire n1010;
  wire n1011;
  wire n1012;
  wire n1013;
  wire n1014;
  wire n1015;
  wire n1016;
  wire n1017;
  wire n1018;
  wire n1019;
  wire n102;
  wire n1020;
  wire n1021;
  wire n1022;
  wire n1023;
  wire n1024;
  wire n1025;
  wire n1026;
  wire n1027;
  wire n1028;
  wire n1029;
  wire n103;
  wire n1030;
  wire n1031;
  wire n1032;
  wire n1033;
  wire n1034;
  wire n1035;
  wire n1036;
  wire n1037;
  wire n1038;
  wire n1039;
  wire n104;
  wire n1040;
  wire n1041;
  wire n1042;
  wire n1043;
  wire n1044;
  wire n1045;
  wire n1046;
  wire n1047;
  wire n1048;
  wire n1049;
  wire n105;
  wire n1050;
  wire n1051;
  wire n1052;
  wire n1053;
  wire n1054;
  wire n1055;
  wire n1056;
  wire n1057;
  wire n1058;
  wire n1059;
  wire n106;
  wire n1060;
  wire n1061;
  wire n1062;
  wire n1063;
  wire n1064;
  wire n1065;
  wire n1066;
  wire n1067;
  wire n1068;
  wire n1069;
  wire n107;
  wire n1070;
  wire n1071;
  wire n1072;
  wire n1073;
  wire n1074;
  wire n1075;
  wire n1076;
  wire n1077;
  wire n1078;
  wire n1079;
  wire n108;
  wire n1080;
  wire n1081;
  wire n1082;
  wire n1083;
  wire n1084;
  wire n1085;
  wire n1086;
  wire n1087;
  wire n1088;
  wire n1089;
  wire n109;
  wire n1090;
  wire n1091;
  wire n1092;
  wire n1093;
  wire n1094;
  wire n1095;
  wire n1096;
  wire n1097;
  wire n1098;
  wire n1099;
  wire n11;
  wire n110;
  wire n1100;
  wire n1101;
  wire n1102;
  wire n1103;
  wire n1104;
  wire n1105;
  wire n1106;
  wire n1107;
  wire n1108;
  wire n1109;
  wire n1110;
  wire n1111;
  wire n1112;
  wire n1113;
  wire n1114;
  wire n1115;
  wire n1116;
  wire n1117;
  wire n1118;
  wire n1119;
  wire n1120;
  wire n1121;
  wire n1122;
  wire n1123;
  wire n1124;
  wire n1125;
  wire n1126;
  wire n1127;
  wire n1128;
  wire n1129;
  wire n113;
  wire n1130;
  wire n1131;
  wire n1132;
  wire n1133;
  wire n1134;
  wire n1135;
  wire n1136;
  wire n1137;
  wire n1138;
  wire n1139;
  wire n1140;
  wire n1141;
  wire n1142;
  wire n1143;
  wire n1144;
  wire n1145;
  wire n1146;
  wire n1147;
  wire n1148;
  wire n1149;
  wire n115;
  wire n1150;
  wire n1151;
  wire n1152;
  wire n1153;
  wire n1154;
  wire n1155;
  wire n1156;
  wire n1157;
  wire n1158;
  wire n1159;
  wire n116;
  wire n1160;
  wire n1161;
  wire n1162;
  wire n1163;
  wire n1164;
  wire n1165;
  wire n1166;
  wire n1167;
  wire n1168;
  wire n1169;
  wire n117;
  wire n1170;
  wire n1171;
  wire n1172;
  wire n1173;
  wire n1174;
  wire n1175;
  wire n1176;
  wire n1177;
  wire n1178;
  wire n1179;
  wire n118;
  wire n1180;
  wire n1181;
  wire n1182;
  wire n1183;
  wire n1184;
  wire n1185;
  wire n1186;
  wire n1187;
  wire n1188;
  wire n1189;
  wire n119;
  wire n1190;
  wire n1191;
  wire n1192;
  wire n1193;
  wire n1194;
  wire n1195;
  wire n1196;
  wire n1197;
  wire n1198;
  wire n1199;
  wire n12;
  wire n120;
  wire n1200;
  wire n1201;
  wire n1202;
  wire n1203;
  wire n1204;
  wire n1205;
  wire n1206;
  wire n1207;
  wire n1208;
  wire n1209;
  wire n121;
  wire n1210;
  wire n1211;
  wire n1212;
  wire n1213;
  wire n1214;
  wire n1215;
  wire n1216;
  wire n1217;
  wire n1218;
  wire n1219;
  wire n122;
  wire n1220;
  wire n1221;
  wire n1222;
  wire n1223;
  wire n1224;
  wire n1225;
  wire n1226;
  wire n1227;
  wire n1228;
  wire n1229;
  wire n123;
  wire n1230;
  wire n1231;
  wire n1232;
  wire n1233;
  wire n1234;
  wire n1235;
  wire n1236;
  wire n1237;
  wire n1238;
  wire n1239;
  wire n124;
  wire n1240;
  wire n1241;
  wire n1242;
  wire n1243;
  wire n1244;
  wire n1245;
  wire n1246;
  wire n1247;
  wire n1248;
  wire n1249;
  wire n125;
  wire n1250;
  wire n1251;
  wire n1252;
  wire n1253;
  wire n1254;
  wire n1255;
  wire n1256;
  wire n1257;
  wire n1258;
  wire n1259;
  wire n126;
  wire n1260;
  wire n1261;
  wire n1262;
  wire n1263;
  wire n1264;
  wire n1265;
  wire n1266;
  wire n1267;
  wire n1268;
  wire n1269;
  wire n127;
  wire n1270;
  wire n1271;
  wire n1273;
  wire n1274;
  wire n1275;
  wire n1276;
  wire n1277;
  wire n1278;
  wire n1279;
  wire n128;
  wire n1280;
  wire n1281;
  wire n1282;
  wire n1283;
  wire n1284;
  wire n1285;
  wire n1286;
  wire n1287;
  wire n1288;
  wire n1289;
  wire n129;
  wire n1290;
  wire n1291;
  wire n1292;
  wire n1293;
  wire n1294;
  wire n1295;
  wire n1296;
  wire n1297;
  wire n1298;
  wire n1299;
  wire n13;
  wire n130;
  wire n1300;
  wire n1301;
  wire n1302;
  wire n1303;
  wire n1304;
  wire n1305;
  wire n1306;
  wire n1307;
  wire n1308;
  wire n1309;
  wire n131;
  wire n1310;
  wire n1311;
  wire n1312;
  wire n1313;
  wire n1314;
  wire n1315;
  wire n1316;
  wire n1317;
  wire n1318;
  wire n1319;
  wire n132;
  wire n1320;
  wire n1321;
  wire n1322;
  wire n1323;
  wire n1324;
  wire n1325;
  wire n1326;
  wire n1327;
  wire n1328;
  wire n1329;
  wire n133;
  wire n1330;
  wire n1331;
  wire n1332;
  wire n1333;
  wire n1334;
  wire n1335;
  wire n1336;
  wire n1337;
  wire n1338;
  wire n1339;
  wire n134;
  wire n1340;
  wire n1341;
  wire n1342;
  wire n1343;
  wire n1344;
  wire n1345;
  wire n1346;
  wire n1347;
  wire n1348;
  wire n1349;
  wire n135;
  wire n1350;
  wire n1351;
  wire n1352;
  wire n1353;
  wire n1354;
  wire n1355;
  wire n1356;
  wire n1357;
  wire n1358;
  wire n1359;
  wire n136;
  wire n1360;
  wire n1361;
  wire n1362;
  wire n1363;
  wire n1364;
  wire n1365;
  wire n1366;
  wire n1367;
  wire n1368;
  wire n1369;
  wire n137;
  wire n1370;
  wire n1371;
  wire n1372;
  wire n1373;
  wire n1374;
  wire n1375;
  wire n1376;
  wire n1377;
  wire n1378;
  wire n1379;
  wire n138;
  wire n1380;
  wire n1381;
  wire n1382;
  wire n1383;
  wire n1384;
  wire n1385;
  wire n1386;
  wire n1387;
  wire n1388;
  wire n1389;
  wire n139;
  wire n1390;
  wire n1391;
  wire n1392;
  wire n1393;
  wire n1394;
  wire n1395;
  wire n1396;
  wire n1397;
  wire n1398;
  wire n1399;
  wire n14;
  wire n140;
  wire n1400;
  wire n1401;
  wire n1402;
  wire n1403;
  wire n1404;
  wire n1405;
  wire n1406;
  wire n1407;
  wire n1408;
  wire n1409;
  wire n141;
  wire n1410;
  wire n1411;
  wire n1412;
  wire n1413;
  wire n1414;
  wire n1415;
  wire n1416;
  wire n1417;
  wire n1418;
  wire n1419;
  wire n142;
  wire n1420;
  wire n1421;
  wire n1422;
  wire n1423;
  wire n1424;
  wire n1425;
  wire n1426;
  wire n1427;
  wire n1428;
  wire n1429;
  wire n143;
  wire n1430;
  wire n1431;
  wire n1432;
  wire n1433;
  wire n1434;
  wire n1435;
  wire n1436;
  wire n1437;
  wire n1438;
  wire n1439;
  wire n144;
  wire n1440;
  wire n1441;
  wire n1442;
  wire n1443;
  wire n1444;
  wire n1445;
  wire n1446;
  wire n1447;
  wire n1448;
  wire n1449;
  wire n145;
  wire n1450;
  wire n1451;
  wire n1452;
  wire n1453;
  wire n1454;
  wire n1455;
  wire n1456;
  wire n1457;
  wire n1458;
  wire n1459;
  wire n146;
  wire n1460;
  wire n1461;
  wire n1462;
  wire n1463;
  wire n1464;
  wire n1465;
  wire n1466;
  wire n1467;
  wire n1468;
  wire n1469;
  wire n147;
  wire n1470;
  wire n1471;
  wire n1472;
  wire n1473;
  wire n1474;
  wire n1475;
  wire n1476;
  wire n1477;
  wire n1478;
  wire n1479;
  wire n148;
  wire n1480;
  wire n1481;
  wire n1482;
  wire n1483;
  wire n1484;
  wire n1485;
  wire n1486;
  wire n1487;
  wire n1488;
  wire n1489;
  wire n149;
  wire n1490;
  wire n1491;
  wire n1492;
  wire n1493;
  wire n1494;
  wire n1495;
  wire n1496;
  wire n1497;
  wire n1498;
  wire n1499;
  wire n15;
  wire n150;
  wire n1500;
  wire n1501;
  wire n1502;
  wire n1503;
  wire n1504;
  wire n1505;
  wire n1506;
  wire n1507;
  wire n1508;
  wire n1509;
  wire n151;
  wire n1510;
  wire n1511;
  wire n1512;
  wire n1513;
  wire n1514;
  wire n1515;
  wire n1516;
  wire n1517;
  wire n1518;
  wire n1519;
  wire n152;
  wire n1520;
  wire n1521;
  wire n1522;
  wire n1523;
  wire n1524;
  wire n1525;
  wire n1526;
  wire n1527;
  wire n1528;
  wire n1529;
  wire n153;
  wire n1530;
  wire n1531;
  wire n1532;
  wire n1533;
  wire n1534;
  wire n1535;
  wire n1536;
  wire n1537;
  wire n1538;
  wire n1539;
  wire n154;
  wire n1540;
  wire n1541;
  wire n1542;
  wire n1543;
  wire n1544;
  wire n1545;
  wire n1546;
  wire n1547;
  wire n1548;
  wire n1549;
  wire n155;
  wire n1550;
  wire n1551;
  wire n1552;
  wire n1553;
  wire n1554;
  wire n1555;
  wire n1556;
  wire n1557;
  wire n1558;
  wire n1559;
  wire n156;
  wire n1560;
  wire n1561;
  wire n1562;
  wire n1563;
  wire n1564;
  wire n1565;
  wire n1566;
  wire n1567;
  wire n1568;
  wire n1569;
  wire n157;
  wire n1570;
  wire n1571;
  wire n1572;
  wire n1573;
  wire n1574;
  wire n1575;
  wire n1576;
  wire n1577;
  wire n1578;
  wire n1579;
  wire n158;
  wire n1580;
  wire n1581;
  wire n1582;
  wire n1583;
  wire n1584;
  wire n1585;
  wire n1586;
  wire n1587;
  wire n1588;
  wire n1589;
  wire n159;
  wire n1590;
  wire n1591;
  wire n1592;
  wire n1593;
  wire n1594;
  wire n1595;
  wire n1596;
  wire n1597;
  wire n1598;
  wire n1599;
  wire n16;
  wire n160;
  wire n1600;
  wire n1601;
  wire n1602;
  wire n1603;
  wire n1604;
  wire n1605;
  wire n1606;
  wire n1607;
  wire n1608;
  wire n1609;
  wire n161;
  wire n1610;
  wire n1611;
  wire n1612;
  wire n1613;
  wire n1614;
  wire n1615;
  wire n1616;
  wire n1617;
  wire n1618;
  wire n1619;
  wire n162;
  wire n1620;
  wire n1621;
  wire n1622;
  wire n1623;
  wire n1624;
  wire n1625;
  wire n1626;
  wire n1627;
  wire n1628;
  wire n1629;
  wire n163;
  wire n1630;
  wire n1631;
  wire n1632;
  wire n1633;
  wire n1634;
  wire n1635;
  wire n1636;
  wire n1637;
  wire n1638;
  wire n1639;
  wire n164;
  wire n1640;
  wire n1641;
  wire n1642;
  wire n1643;
  wire n1644;
  wire n1645;
  wire n1646;
  wire n1647;
  wire n1648;
  wire n1649;
  wire n165;
  wire n1650;
  wire n1651;
  wire n1652;
  wire n1653;
  wire n1654;
  wire n1655;
  wire n1656;
  wire n1657;
  wire n1658;
  wire n1659;
  wire n166;
  wire n1660;
  wire n1661;
  wire n1662;
  wire n1663;
  wire n1664;
  wire n1665;
  wire n1666;
  wire n1667;
  wire n1668;
  wire n1669;
  wire n167;
  wire n1670;
  wire n1671;
  wire n1672;
  wire n1673;
  wire n1674;
  wire n1675;
  wire n1676;
  wire n1677;
  wire n1678;
  wire n1679;
  wire n168;
  wire n1680;
  wire n1681;
  wire n1682;
  wire n1683;
  wire n1684;
  wire n1685;
  wire n1686;
  wire n1687;
  wire n1688;
  wire n1689;
  wire n169;
  wire n1690;
  wire n1691;
  wire n1692;
  wire n1693;
  wire n1694;
  wire n1695;
  wire n1696;
  wire n1697;
  wire n1698;
  wire n1699;
  wire n17;
  wire n170;
  wire n1700;
  wire n1701;
  wire n1702;
  wire n1703;
  wire n1704;
  wire n1705;
  wire n1706;
  wire n1707;
  wire n1708;
  wire n1709;
  wire n171;
  wire n1710;
  wire n1711;
  wire n1712;
  wire n1713;
  wire n1714;
  wire n1715;
  wire n1716;
  wire n1717;
  wire n1718;
  wire n1719;
  wire n172;
  wire n1720;
  wire n1721;
  wire n1722;
  wire n1723;
  wire n1724;
  wire n1725;
  wire n1726;
  wire n1727;
  wire n1728;
  wire n1729;
  wire n173;
  wire n1730;
  wire n1731;
  wire n1732;
  wire n1733;
  wire n1734;
  wire n1735;
  wire n1736;
  wire n1737;
  wire n1738;
  wire n1739;
  wire n174;
  wire n1740;
  wire n1741;
  wire n1742;
  wire n1743;
  wire n1744;
  wire n1745;
  wire n1746;
  wire n1747;
  wire n1748;
  wire n1749;
  wire n175;
  wire n1750;
  wire n1751;
  wire n1752;
  wire n1753;
  wire n1754;
  wire n1755;
  wire n1756;
  wire n1757;
  wire n1758;
  wire n1759;
  wire n176;
  wire n1760;
  wire n1761;
  wire n1762;
  wire n1763;
  wire n1764;
  wire n1765;
  wire n1766;
  wire n1767;
  wire n1768;
  wire n1769;
  wire n177;
  wire n1770;
  wire n1771;
  wire n1772;
  wire n1773;
  wire n1774;
  wire n1775;
  wire n1776;
  wire n1777;
  wire n1778;
  wire n1779;
  wire n178;
  wire n1780;
  wire n1781;
  wire n1782;
  wire n1783;
  wire n1784;
  wire n1785;
  wire n1786;
  wire n1787;
  wire n1788;
  wire n1789;
  wire n179;
  wire n1790;
  wire n1791;
  wire n1792;
  wire n1793;
  wire n1794;
  wire n1795;
  wire n1796;
  wire n1797;
  wire n1798;
  wire n1799;
  wire n18;
  wire n180;
  wire n1800;
  wire n1801;
  wire n1802;
  wire n1803;
  wire n1804;
  wire n1805;
  wire n1806;
  wire n1807;
  wire n1808;
  wire n1809;
  wire n181;
  wire n1810;
  wire n1811;
  wire n1812;
  wire n1813;
  wire n1814;
  wire n1815;
  wire n1816;
  wire n1817;
  wire n1818;
  wire n1819;
  wire n182;
  wire n1820;
  wire n1821;
  wire n1822;
  wire n1823;
  wire n1824;
  wire n1825;
  wire n1826;
  wire n1827;
  wire n1828;
  wire n1829;
  wire n183;
  wire n1830;
  wire n1831;
  wire n1832;
  wire n1833;
  wire n1834;
  wire n1835;
  wire n1836;
  wire n1837;
  wire n1838;
  wire n1839;
  wire n184;
  wire n1840;
  wire n1841;
  wire n1842;
  wire n1843;
  wire n1844;
  wire n1845;
  wire n1846;
  wire n1847;
  wire n1848;
  wire n1849;
  wire n185;
  wire n1850;
  wire n1851;
  wire n1852;
  wire n1853;
  wire n1854;
  wire n1855;
  wire n1856;
  wire n1857;
  wire n1858;
  wire n1859;
  wire n186;
  wire n1860;
  wire n1861;
  wire n1862;
  wire n1863;
  wire n1864;
  wire n1865;
  wire n1866;
  wire n1867;
  wire n1868;
  wire n1869;
  wire n187;
  wire n1870;
  wire n1871;
  wire n1872;
  wire n1873;
  wire n1874;
  wire n1875;
  wire n1876;
  wire n1877;
  wire n1878;
  wire n1879;
  wire n188;
  wire n1880;
  wire n1881;
  wire n1882;
  wire n1883;
  wire n1884;
  wire n1885;
  wire n1886;
  wire n1887;
  wire n1888;
  wire n1889;
  wire n189;
  wire n1890;
  wire n1891;
  wire n1892;
  wire n1893;
  wire n1894;
  wire n1895;
  wire n1896;
  wire n1897;
  wire n1898;
  wire n1899;
  wire n19;
  wire n190;
  wire n1900;
  wire n1901;
  wire n1902;
  wire n1903;
  wire n1904;
  wire n1905;
  wire n1906;
  wire n1907;
  wire n1908;
  wire n1909;
  wire n191;
  wire n1910;
  wire n1911;
  wire n1912;
  wire n1913;
  wire n1914;
  wire n1915;
  wire n1916;
  wire n1917;
  wire n1918;
  wire n1919;
  wire n192;
  wire n1920;
  wire n1921;
  wire n1922;
  wire n1923;
  wire n1924;
  wire n1925;
  wire n1926;
  wire n1927;
  wire n1928;
  wire n1929;
  wire n193;
  wire n1930;
  wire n1931;
  wire n1932;
  wire n1933;
  wire n1934;
  wire n1935;
  wire n1936;
  wire n1937;
  wire n1938;
  wire n1939;
  wire n194;
  wire n1940;
  wire n1941;
  wire n1942;
  wire n1943;
  wire n1944;
  wire n1945;
  wire n1946;
  wire n1947;
  wire n1948;
  wire n1949;
  wire n195;
  wire n1950;
  wire n1951;
  wire n1952;
  wire n1953;
  wire n1954;
  wire n1955;
  wire n1956;
  wire n1957;
  wire n1958;
  wire n1959;
  wire n196;
  wire n1960;
  wire n1961;
  wire n1962;
  wire n1963;
  wire n1964;
  wire n1965;
  wire n1966;
  wire n1967;
  wire n1968;
  wire n1969;
  wire n197;
  wire n1970;
  wire n1971;
  wire n1972;
  wire n1973;
  wire n1974;
  wire n1975;
  wire n1976;
  wire n1977;
  wire n1978;
  wire n1979;
  wire n198;
  wire n1980;
  wire n1981;
  wire n1982;
  wire n1983;
  wire n1984;
  wire n1985;
  wire n1986;
  wire n1987;
  wire n1988;
  wire n1989;
  wire n199;
  wire n1990;
  wire n1991;
  wire n1992;
  wire n1993;
  wire n1994;
  wire n1995;
  wire n1996;
  wire n1997;
  wire n1998;
  wire n1999;
  wire n2;
  wire n20;
  wire n200;
  wire n2000;
  wire n2001;
  wire n2002;
  wire n2003;
  wire n2004;
  wire n2005;
  wire n2006;
  wire n2007;
  wire n2008;
  wire n2009;
  wire n201;
  wire n2010;
  wire n2011;
  wire n2012;
  wire n2013;
  wire n2014;
  wire n2015;
  wire n2016;
  wire n2017;
  wire n2018;
  wire n2019;
  wire n202;
  wire n2020;
  wire n2021;
  wire n2022;
  wire n2023;
  wire n2024;
  wire n2025;
  wire n2026;
  wire n2027;
  wire n2028;
  wire n2029;
  wire n203;
  wire n2030;
  wire n2031;
  wire n2032;
  wire n2033;
  wire n2034;
  wire n2035;
  wire n2036;
  wire n2037;
  wire n2038;
  wire n2039;
  wire n204;
  wire n2040;
  wire n2041;
  wire n2042;
  wire n2043;
  wire n2044;
  wire n2045;
  wire n2046;
  wire n2047;
  wire n2048;
  wire n2049;
  wire n205;
  wire n2050;
  wire n2051;
  wire n2052;
  wire n2053;
  wire n2054;
  wire n2055;
  wire n2056;
  wire n2057;
  wire n2058;
  wire n2059;
  wire n206;
  wire n2060;
  wire n2061;
  wire n2062;
  wire n2063;
  wire n2064;
  wire n2065;
  wire n2066;
  wire n2067;
  wire n2068;
  wire n2069;
  wire n207;
  wire n2070;
  wire n2071;
  wire n2072;
  wire n2073;
  wire n2074;
  wire n2075;
  wire n2076;
  wire n2077;
  wire n2078;
  wire n2079;
  wire n208;
  wire n2080;
  wire n2081;
  wire n2082;
  wire n2083;
  wire n2084;
  wire n2085;
  wire n2086;
  wire n2087;
  wire n2088;
  wire n2089;
  wire n209;
  wire n2090;
  wire n2091;
  wire n2092;
  wire n2093;
  wire n2094;
  wire n2095;
  wire n2096;
  wire n2097;
  wire n2098;
  wire n2099;
  wire n21;
  wire n210;
  wire n2100;
  wire n2101;
  wire n2102;
  wire n2103;
  wire n2104;
  wire n2105;
  wire n2106;
  wire n2107;
  wire n2108;
  wire n2109;
  wire n211;
  wire n2110;
  wire n2111;
  wire n2112;
  wire n2113;
  wire n2114;
  wire n2115;
  wire n2116;
  wire n2117;
  wire n2118;
  wire n2119;
  wire n212;
  wire n2120;
  wire n2121;
  wire n2122;
  wire n2123;
  wire n2124;
  wire n2125;
  wire n2126;
  wire n2127;
  wire n2128;
  wire n2129;
  wire n213;
  wire n2130;
  wire n2131;
  wire n2132;
  wire n2133;
  wire n2134;
  wire n2135;
  wire n2136;
  wire n2137;
  wire n2138;
  wire n2139;
  wire n214;
  wire n2140;
  wire n2141;
  wire n2142;
  wire n2143;
  wire n2144;
  wire n2145;
  wire n2146;
  wire n2147;
  wire n2148;
  wire n2149;
  wire n215;
  wire n2150;
  wire n2151;
  wire n2152;
  wire n2153;
  wire n2154;
  wire n2155;
  wire n2156;
  wire n2157;
  wire n2158;
  wire n2159;
  wire n216;
  wire n2160;
  wire n2161;
  wire n2162;
  wire n2163;
  wire n2164;
  wire n2165;
  wire n2166;
  wire n2167;
  wire n2168;
  wire n2169;
  wire n217;
  wire n2170;
  wire n2171;
  wire n2172;
  wire n2173;
  wire n2174;
  wire n2175;
  wire n2176;
  wire n2177;
  wire n2178;
  wire n2179;
  wire n218;
  wire n2180;
  wire n2181;
  wire n2182;
  wire n2183;
  wire n2184;
  wire n2185;
  wire n2186;
  wire n2187;
  wire n2188;
  wire n2189;
  wire n219;
  wire n2190;
  wire n2191;
  wire n2192;
  wire n2193;
  wire n2194;
  wire n2195;
  wire n2196;
  wire n2197;
  wire n2198;
  wire n2199;
  wire n22;
  wire n220;
  wire n2200;
  wire n2201;
  wire n2202;
  wire n2203;
  wire n2204;
  wire n2205;
  wire n2206;
  wire n2207;
  wire n2208;
  wire n2209;
  wire n221;
  wire n2210;
  wire n2211;
  wire n2212;
  wire n2213;
  wire n2214;
  wire n2215;
  wire n2216;
  wire n2217;
  wire n2218;
  wire n2219;
  wire n222;
  wire n2220;
  wire n2221;
  wire n2222;
  wire n2223;
  wire n2224;
  wire n2225;
  wire n2226;
  wire n2227;
  wire n2228;
  wire n2229;
  wire n223;
  wire n2230;
  wire n2231;
  wire n2232;
  wire n2233;
  wire n2234;
  wire n2235;
  wire n2236;
  wire n2237;
  wire n2238;
  wire n2239;
  wire n224;
  wire n2240;
  wire n2241;
  wire n2242;
  wire n2243;
  wire n2244;
  wire n2245;
  wire n2246;
  wire n2247;
  wire n2248;
  wire n2249;
  wire n225;
  wire n2250;
  wire n2251;
  wire n2252;
  wire n2253;
  wire n2254;
  wire n2255;
  wire n2256;
  wire n2257;
  wire n2258;
  wire n2259;
  wire n226;
  wire n2260;
  wire n2261;
  wire n2262;
  wire n2263;
  wire n2264;
  wire n2265;
  wire n2266;
  wire n2267;
  wire n2268;
  wire n2269;
  wire n227;
  wire n2270;
  wire n2271;
  wire n2272;
  wire n2273;
  wire n2274;
  wire n2275;
  wire n2276;
  wire n2277;
  wire n2278;
  wire n2279;
  wire n228;
  wire n2280;
  wire n2281;
  wire n2282;
  wire n2283;
  wire n2284;
  wire n2285;
  wire n2286;
  wire n2287;
  wire n2288;
  wire n2289;
  wire n229;
  wire n2290;
  wire n2291;
  wire n2292;
  wire n2293;
  wire n2294;
  wire n2295;
  wire n2296;
  wire n2297;
  wire n2298;
  wire n2299;
  wire n23;
  wire n230;
  wire n2300;
  wire n2301;
  wire n2302;
  wire n2303;
  wire n2304;
  wire n2305;
  wire n2306;
  wire n2307;
  wire n2308;
  wire n2309;
  wire n231;
  wire n2310;
  wire n2311;
  wire n2312;
  wire n2313;
  wire n2314;
  wire n2315;
  wire n2316;
  wire n2317;
  wire n2318;
  wire n2319;
  wire n232;
  wire n2320;
  wire n2321;
  wire n2322;
  wire n2323;
  wire n2324;
  wire n2325;
  wire n2326;
  wire n2327;
  wire n2328;
  wire n2329;
  wire n233;
  wire n2330;
  wire n2331;
  wire n2332;
  wire n2333;
  wire n2334;
  wire n2335;
  wire n2336;
  wire n2337;
  wire n2338;
  wire n2339;
  wire n234;
  wire n2340;
  wire n2341;
  wire n2342;
  wire n2343;
  wire n2344;
  wire n2345;
  wire n2346;
  wire n2347;
  wire n2348;
  wire n2349;
  wire n235;
  wire n2350;
  wire n2351;
  wire n2352;
  wire n2353;
  wire n2354;
  wire n2355;
  wire n2356;
  wire n2357;
  wire n2358;
  wire n2359;
  wire n236;
  wire n2360;
  wire n2361;
  wire n2362;
  wire n2363;
  wire n2364;
  wire n2365;
  wire n2366;
  wire n2367;
  wire n2368;
  wire n2369;
  wire n237;
  wire n2370;
  wire n2371;
  wire n2372;
  wire n2373;
  wire n2374;
  wire n2375;
  wire n2376;
  wire n2377;
  wire n2378;
  wire n2379;
  wire n238;
  wire n2380;
  wire n2381;
  wire n2382;
  wire n2383;
  wire n2384;
  wire n2385;
  wire n2386;
  wire n2387;
  wire n2388;
  wire n2389;
  wire n239;
  wire n2390;
  wire n2391;
  wire n2392;
  wire n2393;
  wire n2394;
  wire n2395;
  wire n2396;
  wire n2397;
  wire n2398;
  wire n2399;
  wire n24;
  wire n240;
  wire n2400;
  wire n2401;
  wire n2402;
  wire n2403;
  wire n2404;
  wire n2405;
  wire n2406;
  wire n2407;
  wire n2408;
  wire n2409;
  wire n241;
  wire n2410;
  wire n2411;
  wire n2412;
  wire n2413;
  wire n2414;
  wire n2415;
  wire n2416;
  wire n2417;
  wire n2418;
  wire n2419;
  wire n242;
  wire n2420;
  wire n2421;
  wire n2422;
  wire n2423;
  wire n2424;
  wire n2425;
  wire n2426;
  wire n2427;
  wire n2428;
  wire n2429;
  wire n243;
  wire n2430;
  wire n2431;
  wire n2432;
  wire n2433;
  wire n2434;
  wire n2435;
  wire n2436;
  wire n2437;
  wire n2438;
  wire n2439;
  wire n244;
  wire n2440;
  wire n2441;
  wire n2442;
  wire n2443;
  wire n2444;
  wire n2445;
  wire n2446;
  wire n2447;
  wire n2448;
  wire n2449;
  wire n245;
  wire n2450;
  wire n2451;
  wire n2452;
  wire n2453;
  wire n2454;
  wire n2455;
  wire n2456;
  wire n2457;
  wire n2458;
  wire n2459;
  wire n246;
  wire n2460;
  wire n2461;
  wire n2462;
  wire n2463;
  wire n2464;
  wire n2465;
  wire n2466;
  wire n2467;
  wire n2468;
  wire n2469;
  wire n247;
  wire n2470;
  wire n2471;
  wire n2472;
  wire n2473;
  wire n2474;
  wire n2475;
  wire n2476;
  wire n2477;
  wire n2478;
  wire n2479;
  wire n248;
  wire n2480;
  wire n2481;
  wire n2482;
  wire n2483;
  wire n2484;
  wire n2485;
  wire n2486;
  wire n2487;
  wire n2488;
  wire n2489;
  wire n249;
  wire n2490;
  wire n2491;
  wire n2492;
  wire n2493;
  wire n2494;
  wire n2495;
  wire n2496;
  wire n2497;
  wire n2498;
  wire n2499;
  wire n25;
  wire n250;
  wire n2500;
  wire n2501;
  wire n2502;
  wire n2503;
  wire n2504;
  wire n2505;
  wire n2506;
  wire n2507;
  wire n2508;
  wire n2509;
  wire n251;
  wire n2510;
  wire n2511;
  wire n2512;
  wire n2513;
  wire n2514;
  wire n2515;
  wire n2516;
  wire n2517;
  wire n2518;
  wire n2519;
  wire n252;
  wire n2520;
  wire n2521;
  wire n2522;
  wire n2523;
  wire n2524;
  wire n2525;
  wire n2526;
  wire n2527;
  wire n2528;
  wire n2529;
  wire n253;
  wire n2530;
  wire n2531;
  wire n2532;
  wire n2533;
  wire n2534;
  wire n2535;
  wire n2536;
  wire n2537;
  wire n2538;
  wire n2539;
  wire n254;
  wire n2540;
  wire n2541;
  wire n2542;
  wire n2543;
  wire n2544;
  wire n2545;
  wire n2546;
  wire n2547;
  wire n2548;
  wire n2549;
  wire n255;
  wire n2550;
  wire n2551;
  wire n2552;
  wire n2553;
  wire n2554;
  wire n2555;
  wire n2556;
  wire n2557;
  wire n2558;
  wire n2559;
  wire n256;
  wire n2560;
  wire n2561;
  wire n2562;
  wire n2563;
  wire n2564;
  wire n2565;
  wire n2566;
  wire n2567;
  wire n2568;
  wire n2569;
  wire n257;
  wire n2570;
  wire n2571;
  wire n2572;
  wire n2573;
  wire n2574;
  wire n2575;
  wire n2576;
  wire n2577;
  wire n2578;
  wire n2579;
  wire n258;
  wire n2580;
  wire n2581;
  wire n2582;
  wire n2583;
  wire n2584;
  wire n2585;
  wire n2586;
  wire n2587;
  wire n2588;
  wire n2589;
  wire n259;
  wire n2590;
  wire n2591;
  wire n2592;
  wire n2593;
  wire n2594;
  wire n2595;
  wire n2596;
  wire n2597;
  wire n2598;
  wire n2599;
  wire n26;
  wire n260;
  wire n2600;
  wire n2601;
  wire n2602;
  wire n2603;
  wire n2604;
  wire n2605;
  wire n2606;
  wire n2607;
  wire n2608;
  wire n2609;
  wire n261;
  wire n2610;
  wire n2611;
  wire n2612;
  wire n2613;
  wire n2614;
  wire n2615;
  wire n2616;
  wire n2617;
  wire n2618;
  wire n2619;
  wire n262;
  wire n2620;
  wire n2621;
  wire n2622;
  wire n2623;
  wire n2624;
  wire n2625;
  wire n2626;
  wire n2627;
  wire n2628;
  wire n2629;
  wire n263;
  wire n2630;
  wire n2631;
  wire n2632;
  wire n2633;
  wire n2634;
  wire n2635;
  wire n2636;
  wire n2637;
  wire n2638;
  wire n2639;
  wire n264;
  wire n2640;
  wire n2641;
  wire n2642;
  wire n2643;
  wire n2644;
  wire n2645;
  wire n2646;
  wire n2647;
  wire n2648;
  wire n2649;
  wire n265;
  wire n2650;
  wire n2651;
  wire n2652;
  wire n2653;
  wire n2654;
  wire n2655;
  wire n2656;
  wire n2657;
  wire n2658;
  wire n2659;
  wire n266;
  wire n2660;
  wire n2662;
  wire n2663;
  wire n2664;
  wire n2665;
  wire n2666;
  wire n2667;
  wire n2668;
  wire n2669;
  wire n267;
  wire n2670;
  wire n2671;
  wire n2672;
  wire n2673;
  wire n2674;
  wire n2675;
  wire n2676;
  wire n2677;
  wire n2678;
  wire n2679;
  wire n268;
  wire n2680;
  wire n2681;
  wire n2682;
  wire n2683;
  wire n2684;
  wire n2685;
  wire n2686;
  wire n2687;
  wire n2688;
  wire n2689;
  wire n269;
  wire n2690;
  wire n2691;
  wire n2692;
  wire n2693;
  wire n2694;
  wire n2695;
  wire n2696;
  wire n2697;
  wire n2698;
  wire n2699;
  wire n27;
  wire n270;
  wire n2700;
  wire n2701;
  wire n2702;
  wire n2703;
  wire n2704;
  wire n2705;
  wire n2706;
  wire n2707;
  wire n2708;
  wire n2709;
  wire n271;
  wire n2710;
  wire n2711;
  wire n2712;
  wire n2713;
  wire n2714;
  wire n2715;
  wire n2716;
  wire n2717;
  wire n2718;
  wire n2719;
  wire n272;
  wire n2720;
  wire n2721;
  wire n2722;
  wire n2723;
  wire n2724;
  wire n2725;
  wire n2726;
  wire n2727;
  wire n2728;
  wire n2729;
  wire n273;
  wire n2730;
  wire n2731;
  wire n2732;
  wire n2733;
  wire n2734;
  wire n2735;
  wire n2736;
  wire n2737;
  wire n2738;
  wire n2739;
  wire n274;
  wire n2740;
  wire n2741;
  wire n2742;
  wire n2743;
  wire n2744;
  wire n2745;
  wire n2746;
  wire n2747;
  wire n2748;
  wire n2749;
  wire n275;
  wire n2750;
  wire n2751;
  wire n2752;
  wire n2753;
  wire n2754;
  wire n2755;
  wire n2756;
  wire n2757;
  wire n2758;
  wire n2759;
  wire n276;
  wire n2760;
  wire n2761;
  wire n2762;
  wire n2763;
  wire n2764;
  wire n2765;
  wire n2766;
  wire n2767;
  wire n2768;
  wire n2769;
  wire n277;
  wire n2770;
  wire n2771;
  wire n2772;
  wire n2773;
  wire n2774;
  wire n2775;
  wire n2776;
  wire n2777;
  wire n2778;
  wire n2779;
  wire n278;
  wire n2780;
  wire n2781;
  wire n2782;
  wire n2783;
  wire n2784;
  wire n2785;
  wire n2786;
  wire n2787;
  wire n2788;
  wire n2789;
  wire n279;
  wire n2790;
  wire n2791;
  wire n2792;
  wire n2793;
  wire n2794;
  wire n2795;
  wire n2796;
  wire n2797;
  wire n2798;
  wire n2799;
  wire n28;
  wire n280;
  wire n2800;
  wire n2801;
  wire n2802;
  wire n2803;
  wire n2804;
  wire n2805;
  wire n2806;
  wire n2807;
  wire n2808;
  wire n2809;
  wire n281;
  wire n2810;
  wire n2811;
  wire n2812;
  wire n2813;
  wire n2814;
  wire n2815;
  wire n2816;
  wire n2817;
  wire n2818;
  wire n2819;
  wire n282;
  wire n2820;
  wire n2821;
  wire n2822;
  wire n2823;
  wire n2824;
  wire n2825;
  wire n2826;
  wire n2827;
  wire n2828;
  wire n2829;
  wire n283;
  wire n2830;
  wire n2831;
  wire n2832;
  wire n2833;
  wire n2834;
  wire n2835;
  wire n2836;
  wire n2837;
  wire n2838;
  wire n2839;
  wire n284;
  wire n2840;
  wire n2841;
  wire n2842;
  wire n2843;
  wire n2844;
  wire n2845;
  wire n2846;
  wire n2847;
  wire n2848;
  wire n2849;
  wire n285;
  wire n2850;
  wire n2851;
  wire n2852;
  wire n2853;
  wire n2854;
  wire n2855;
  wire n2856;
  wire n2857;
  wire n2858;
  wire n2859;
  wire n286;
  wire n2860;
  wire n2861;
  wire n2862;
  wire n2863;
  wire n2864;
  wire n2865;
  wire n2866;
  wire n2867;
  wire n2868;
  wire n2869;
  wire n287;
  wire n2870;
  wire n2871;
  wire n2872;
  wire n2873;
  wire n2874;
  wire n2875;
  wire n2876;
  wire n2877;
  wire n2878;
  wire n2879;
  wire n288;
  wire n2880;
  wire n2881;
  wire n2882;
  wire n2883;
  wire n2884;
  wire n2885;
  wire n2886;
  wire n2887;
  wire n2888;
  wire n2889;
  wire n289;
  wire n2890;
  wire n2891;
  wire n2892;
  wire n2893;
  wire n2894;
  wire n2895;
  wire n2896;
  wire n2897;
  wire n2898;
  wire n2899;
  wire n29;
  wire n290;
  wire n2900;
  wire n2901;
  wire n2902;
  wire n2903;
  wire n2904;
  wire n2905;
  wire n2906;
  wire n2907;
  wire n2908;
  wire n2909;
  wire n291;
  wire n2910;
  wire n2911;
  wire n2912;
  wire n2913;
  wire n2914;
  wire n2915;
  wire n2916;
  wire n2917;
  wire n2918;
  wire n2919;
  wire n292;
  wire n2920;
  wire n2921;
  wire n2922;
  wire n2923;
  wire n2924;
  wire n2925;
  wire n2926;
  wire n2927;
  wire n2928;
  wire n2929;
  wire n293;
  wire n2930;
  wire n2931;
  wire n2932;
  wire n2933;
  wire n2934;
  wire n2935;
  wire n2936;
  wire n2937;
  wire n2938;
  wire n2939;
  wire n294;
  wire n2940;
  wire n2941;
  wire n2942;
  wire n2943;
  wire n2944;
  wire n2945;
  wire n2946;
  wire n2947;
  wire n2948;
  wire n2949;
  wire n295;
  wire n2950;
  wire n2951;
  wire n2952;
  wire n2953;
  wire n2954;
  wire n2955;
  wire n2956;
  wire n2957;
  wire n2958;
  wire n2959;
  wire n296;
  wire n2960;
  wire n2961;
  wire n2962;
  wire n2963;
  wire n2964;
  wire n2965;
  wire n2966;
  wire n2967;
  wire n2968;
  wire n2969;
  wire n297;
  wire n2970;
  wire n2971;
  wire n2972;
  wire n2973;
  wire n2974;
  wire n2975;
  wire n2976;
  wire n2977;
  wire n2978;
  wire n2979;
  wire n298;
  wire n2980;
  wire n2981;
  wire n2982;
  wire n2983;
  wire n2984;
  wire n2985;
  wire n2986;
  wire n2987;
  wire n2988;
  wire n2989;
  wire n299;
  wire n2990;
  wire n2991;
  wire n2992;
  wire n2993;
  wire n2994;
  wire n2995;
  wire n2996;
  wire n2997;
  wire n2998;
  wire n2999;
  wire n3;
  wire n30;
  wire n300;
  wire n3000;
  wire n3001;
  wire n3002;
  wire n3003;
  wire n3004;
  wire n3005;
  wire n3006;
  wire n3007;
  wire n3008;
  wire n3009;
  wire n301;
  wire n3010;
  wire n3011;
  wire n3012;
  wire n3013;
  wire n3014;
  wire n3015;
  wire n3016;
  wire n3017;
  wire n3018;
  wire n3019;
  wire n302;
  wire n3020;
  wire n3021;
  wire n3022;
  wire n3023;
  wire n3024;
  wire n3025;
  wire n3026;
  wire n3027;
  wire n3028;
  wire n3029;
  wire n303;
  wire n3030;
  wire n3031;
  wire n3032;
  wire n3033;
  wire n3034;
  wire n3035;
  wire n3036;
  wire n3037;
  wire n3038;
  wire n3039;
  wire n304;
  wire n3040;
  wire n3041;
  wire n3042;
  wire n3043;
  wire n3044;
  wire n3045;
  wire n3046;
  wire n3047;
  wire n3048;
  wire n3049;
  wire n305;
  wire n3050;
  wire n3051;
  wire n3052;
  wire n3053;
  wire n3054;
  wire n3055;
  wire n3056;
  wire n3057;
  wire n3058;
  wire n3059;
  wire n306;
  wire n3060;
  wire n3061;
  wire n3062;
  wire n3063;
  wire n3064;
  wire n3065;
  wire n3066;
  wire n3067;
  wire n3068;
  wire n3069;
  wire n307;
  wire n3070;
  wire n3071;
  wire n3072;
  wire n3073;
  wire n3074;
  wire n3075;
  wire n3076;
  wire n3077;
  wire n3078;
  wire n3079;
  wire n308;
  wire n3080;
  wire n3081;
  wire n3082;
  wire n3083;
  wire n3084;
  wire n3085;
  wire n3086;
  wire n3087;
  wire n3088;
  wire n3089;
  wire n309;
  wire n3090;
  wire n3091;
  wire n3092;
  wire n3093;
  wire n3094;
  wire n3095;
  wire n3096;
  wire n3097;
  wire n3098;
  wire n3099;
  wire n31;
  wire n310;
  wire n3100;
  wire n3101;
  wire n3102;
  wire n3103;
  wire n3104;
  wire n3105;
  wire n3106;
  wire n3107;
  wire n3108;
  wire n3109;
  wire n311;
  wire n3110;
  wire n3111;
  wire n3112;
  wire n3113;
  wire n3114;
  wire n3115;
  wire n3116;
  wire n3117;
  wire n3118;
  wire n3119;
  wire n312;
  wire n3120;
  wire n3121;
  wire n3122;
  wire n3123;
  wire n3124;
  wire n3125;
  wire n3126;
  wire n3127;
  wire n3128;
  wire n3129;
  wire n313;
  wire n3130;
  wire n3131;
  wire n3132;
  wire n3133;
  wire n3134;
  wire n3135;
  wire n3136;
  wire n3137;
  wire n3138;
  wire n3139;
  wire n314;
  wire n3140;
  wire n3141;
  wire n3142;
  wire n3143;
  wire n3144;
  wire n3145;
  wire n3146;
  wire n3147;
  wire n3148;
  wire n3149;
  wire n315;
  wire n3150;
  wire n3151;
  wire n3152;
  wire n3153;
  wire n3154;
  wire n3155;
  wire n3156;
  wire n3157;
  wire n3158;
  wire n3159;
  wire n316;
  wire n3160;
  wire n3161;
  wire n3162;
  wire n3163;
  wire n3164;
  wire n3165;
  wire n3166;
  wire n3167;
  wire n3168;
  wire n3169;
  wire n317;
  wire n3170;
  wire n3171;
  wire n3172;
  wire n3173;
  wire n3174;
  wire n3175;
  wire n3176;
  wire n3177;
  wire n3178;
  wire n3179;
  wire n318;
  wire n3180;
  wire n3181;
  wire n3182;
  wire n3183;
  wire n3184;
  wire n3185;
  wire n3186;
  wire n3187;
  wire n3188;
  wire n3189;
  wire n319;
  wire n3190;
  wire n3191;
  wire n3192;
  wire n3193;
  wire n3194;
  wire n3195;
  wire n3196;
  wire n3197;
  wire n3198;
  wire n3199;
  wire n32;
  wire n320;
  wire n3200;
  wire n3201;
  wire n3202;
  wire n3203;
  wire n3204;
  wire n3205;
  wire n3206;
  wire n3207;
  wire n3208;
  wire n3209;
  wire n321;
  wire n3210;
  wire n3211;
  wire n3212;
  wire n3213;
  wire n3214;
  wire n3215;
  wire n3216;
  wire n3217;
  wire n3218;
  wire n3219;
  wire n322;
  wire n3220;
  wire n3221;
  wire n3222;
  wire n3223;
  wire n3224;
  wire n3225;
  wire n3226;
  wire n3227;
  wire n3228;
  wire n3229;
  wire n323;
  wire n3230;
  wire n3231;
  wire n3232;
  wire n3233;
  wire n3234;
  wire n3235;
  wire n3236;
  wire n3237;
  wire n3238;
  wire n3239;
  wire n324;
  wire n3240;
  wire n3241;
  wire n3242;
  wire n3243;
  wire n3244;
  wire n3245;
  wire n3246;
  wire n3247;
  wire n3248;
  wire n3249;
  wire n325;
  wire n3250;
  wire n3251;
  wire n3252;
  wire n3253;
  wire n3254;
  wire n3255;
  wire n3256;
  wire n3257;
  wire n3258;
  wire n3259;
  wire n326;
  wire n3260;
  wire n3261;
  wire n3262;
  wire n3263;
  wire n3264;
  wire n3265;
  wire n3266;
  wire n3267;
  wire n3268;
  wire n3269;
  wire n327;
  wire n3270;
  wire n3271;
  wire n3272;
  wire n3273;
  wire n3274;
  wire n3275;
  wire n3276;
  wire n3277;
  wire n3278;
  wire n3279;
  wire n328;
  wire n3280;
  wire n3281;
  wire n3282;
  wire n3283;
  wire n3284;
  wire n3285;
  wire n3286;
  wire n3287;
  wire n3288;
  wire n3289;
  wire n329;
  wire n3290;
  wire n3291;
  wire n3292;
  wire n3293;
  wire n3294;
  wire n3295;
  wire n3296;
  wire n3297;
  wire n3298;
  wire n3299;
  wire n33;
  wire n330;
  wire n3300;
  wire n3301;
  wire n3302;
  wire n3303;
  wire n3304;
  wire n3305;
  wire n3306;
  wire n3307;
  wire n3308;
  wire n3309;
  wire n331;
  wire n3310;
  wire n3311;
  wire n3312;
  wire n3313;
  wire n3314;
  wire n3315;
  wire n3316;
  wire n3317;
  wire n3318;
  wire n3319;
  wire n332;
  wire n3320;
  wire n3321;
  wire n3322;
  wire n3323;
  wire n3324;
  wire n3325;
  wire n3326;
  wire n3327;
  wire n3328;
  wire n3329;
  wire n333;
  wire n3330;
  wire n3331;
  wire n3332;
  wire n3333;
  wire n3334;
  wire n3335;
  wire n3336;
  wire n3337;
  wire n3338;
  wire n3339;
  wire n334;
  wire n3340;
  wire n3341;
  wire n3342;
  wire n3343;
  wire n3344;
  wire n3345;
  wire n3346;
  wire n3347;
  wire n3348;
  wire n3349;
  wire n335;
  wire n3350;
  wire n3351;
  wire n3352;
  wire n3353;
  wire n3354;
  wire n3355;
  wire n3356;
  wire n3357;
  wire n3358;
  wire n3359;
  wire n336;
  wire n3360;
  wire n3361;
  wire n3362;
  wire n3363;
  wire n3364;
  wire n3365;
  wire n3366;
  wire n3367;
  wire n3368;
  wire n3369;
  wire n337;
  wire n3370;
  wire n3371;
  wire n3372;
  wire n3373;
  wire n3374;
  wire n3375;
  wire n3376;
  wire n3377;
  wire n3378;
  wire n3379;
  wire n338;
  wire n3380;
  wire n3381;
  wire n3382;
  wire n3383;
  wire n3384;
  wire n3385;
  wire n3386;
  wire n3387;
  wire n3388;
  wire n3389;
  wire n339;
  wire n3390;
  wire n3391;
  wire n3392;
  wire n3393;
  wire n3394;
  wire n3395;
  wire n3396;
  wire n3397;
  wire n3398;
  wire n3399;
  wire n34;
  wire n340;
  wire n3400;
  wire n3401;
  wire n3402;
  wire n3403;
  wire n3404;
  wire n3405;
  wire n3406;
  wire n3407;
  wire n3408;
  wire n3409;
  wire n341;
  wire n3410;
  wire n3411;
  wire n3412;
  wire n3413;
  wire n3414;
  wire n3415;
  wire n3416;
  wire n3417;
  wire n3418;
  wire n3419;
  wire n342;
  wire n3420;
  wire n3421;
  wire n3422;
  wire n3423;
  wire n3424;
  wire n3425;
  wire n3426;
  wire n3427;
  wire n3428;
  wire n3429;
  wire n343;
  wire n3430;
  wire n3431;
  wire n3432;
  wire n3433;
  wire n3434;
  wire n3435;
  wire n3436;
  wire n3437;
  wire n3438;
  wire n3439;
  wire n344;
  wire n3440;
  wire n3441;
  wire n3442;
  wire n3443;
  wire n3444;
  wire n3445;
  wire n3446;
  wire n3447;
  wire n3448;
  wire n3449;
  wire n345;
  wire n3450;
  wire n3451;
  wire n3452;
  wire n3453;
  wire n3454;
  wire n3455;
  wire n3456;
  wire n3457;
  wire n3458;
  wire n3459;
  wire n346;
  wire n3460;
  wire n3461;
  wire n3462;
  wire n3463;
  wire n3464;
  wire n3465;
  wire n3466;
  wire n3467;
  wire n3468;
  wire n3469;
  wire n347;
  wire n3470;
  wire n3471;
  wire n3472;
  wire n3473;
  wire n3474;
  wire n3475;
  wire n3476;
  wire n3477;
  wire n3478;
  wire n3479;
  wire n348;
  wire n3480;
  wire n3481;
  wire n3482;
  wire n3483;
  wire n3484;
  wire n3485;
  wire n3486;
  wire n3487;
  wire n3488;
  wire n3489;
  wire n349;
  wire n3490;
  wire n3491;
  wire n3492;
  wire n3493;
  wire n3494;
  wire n3495;
  wire n3496;
  wire n3497;
  wire n3498;
  wire n3499;
  wire n35;
  wire n350;
  wire n3500;
  wire n3501;
  wire n3502;
  wire n3503;
  wire n3504;
  wire n3505;
  wire n3506;
  wire n3507;
  wire n3508;
  wire n3509;
  wire n351;
  wire n3510;
  wire n3511;
  wire n3512;
  wire n3513;
  wire n3514;
  wire n3515;
  wire n3516;
  wire n3517;
  wire n3518;
  wire n3519;
  wire n352;
  wire n3520;
  wire n3521;
  wire n3522;
  wire n3523;
  wire n3524;
  wire n3525;
  wire n3526;
  wire n3527;
  wire n3528;
  wire n3529;
  wire n353;
  wire n3530;
  wire n3531;
  wire n3532;
  wire n3533;
  wire n3534;
  wire n3535;
  wire n3536;
  wire n3537;
  wire n3538;
  wire n3539;
  wire n354;
  wire n3540;
  wire n3541;
  wire n3542;
  wire n3543;
  wire n3544;
  wire n3545;
  wire n3546;
  wire n3547;
  wire n3548;
  wire n3549;
  wire n355;
  wire n3550;
  wire n3551;
  wire n3552;
  wire n3553;
  wire n3554;
  wire n3555;
  wire n3556;
  wire n3557;
  wire n3558;
  wire n3559;
  wire n356;
  wire n3560;
  wire n3561;
  wire n3562;
  wire n3563;
  wire n3564;
  wire n3565;
  wire n3566;
  wire n3567;
  wire n3568;
  wire n3569;
  wire n357;
  wire n3570;
  wire n3571;
  wire n3572;
  wire n3573;
  wire n3574;
  wire n3575;
  wire n3576;
  wire n3577;
  wire n3578;
  wire n3579;
  wire n358;
  wire n3580;
  wire n3581;
  wire n3582;
  wire n3583;
  wire n3584;
  wire n3585;
  wire n3586;
  wire n3587;
  wire n3588;
  wire n3589;
  wire n359;
  wire n3590;
  wire n3591;
  wire n3592;
  wire n3593;
  wire n3594;
  wire n3595;
  wire n3596;
  wire n3597;
  wire n3598;
  wire n3599;
  wire n36;
  wire n360;
  wire n3600;
  wire n3601;
  wire n3602;
  wire n3603;
  wire n3604;
  wire n3605;
  wire n3606;
  wire n3607;
  wire n3608;
  wire n3609;
  wire n361;
  wire n3610;
  wire n3611;
  wire n3612;
  wire n3613;
  wire n3614;
  wire n3615;
  wire n3616;
  wire n3617;
  wire n3618;
  wire n3619;
  wire n362;
  wire n3620;
  wire n3621;
  wire n3622;
  wire n3623;
  wire n3624;
  wire n3625;
  wire n3626;
  wire n3627;
  wire n3628;
  wire n3629;
  wire n363;
  wire n3630;
  wire n3631;
  wire n3632;
  wire n3633;
  wire n3634;
  wire n3635;
  wire n3636;
  wire n3637;
  wire n3638;
  wire n3639;
  wire n364;
  wire n3640;
  wire n3641;
  wire n3642;
  wire n3643;
  wire n3644;
  wire n3645;
  wire n3646;
  wire n3647;
  wire n3648;
  wire n3649;
  wire n365;
  wire n3650;
  wire n3651;
  wire n3652;
  wire n3653;
  wire n3654;
  wire n3655;
  wire n3656;
  wire n3657;
  wire n3658;
  wire n3659;
  wire n366;
  wire n3660;
  wire n3661;
  wire n3662;
  wire n3663;
  wire n3664;
  wire n3665;
  wire n3666;
  wire n3667;
  wire n3668;
  wire n3669;
  wire n367;
  wire n3670;
  wire n3671;
  wire n3672;
  wire n3673;
  wire n3674;
  wire n3675;
  wire n3676;
  wire n3677;
  wire n3678;
  wire n3679;
  wire n368;
  wire n3680;
  wire n3681;
  wire n3682;
  wire n3683;
  wire n3684;
  wire n3685;
  wire n3686;
  wire n3687;
  wire n3688;
  wire n3689;
  wire n369;
  wire n3690;
  wire n3691;
  wire n3692;
  wire n3693;
  wire n3694;
  wire n3695;
  wire n3696;
  wire n3697;
  wire n3698;
  wire n3699;
  wire n37;
  wire n370;
  wire n3700;
  wire n3701;
  wire n3702;
  wire n3703;
  wire n3704;
  wire n3705;
  wire n3706;
  wire n3707;
  wire n3708;
  wire n3709;
  wire n371;
  wire n3710;
  wire n3711;
  wire n3712;
  wire n3713;
  wire n3714;
  wire n3715;
  wire n3716;
  wire n3717;
  wire n3718;
  wire n3719;
  wire n372;
  wire n3720;
  wire n3721;
  wire n3722;
  wire n3723;
  wire n3724;
  wire n3725;
  wire n3726;
  wire n3727;
  wire n3728;
  wire n3729;
  wire n373;
  wire n3730;
  wire n3731;
  wire n3732;
  wire n3733;
  wire n3734;
  wire n3735;
  wire n3736;
  wire n3737;
  wire n3738;
  wire n3739;
  wire n374;
  wire n3740;
  wire n3741;
  wire n3742;
  wire n3743;
  wire n3744;
  wire n3745;
  wire n3746;
  wire n3747;
  wire n3748;
  wire n3749;
  wire n375;
  wire n3750;
  wire n3751;
  wire n3752;
  wire n3753;
  wire n3754;
  wire n3755;
  wire n3756;
  wire n3757;
  wire n3758;
  wire n3759;
  wire n376;
  wire n3760;
  wire n3761;
  wire n3762;
  wire n3763;
  wire n3764;
  wire n3765;
  wire n3766;
  wire n3767;
  wire n3768;
  wire n3769;
  wire n377;
  wire n3770;
  wire n3771;
  wire n3772;
  wire n3773;
  wire n3774;
  wire n3775;
  wire n3776;
  wire n3777;
  wire n3778;
  wire n3779;
  wire n378;
  wire n3780;
  wire n3781;
  wire n3782;
  wire n3783;
  wire n3784;
  wire n3785;
  wire n3786;
  wire n3787;
  wire n3788;
  wire n3789;
  wire n379;
  wire n3790;
  wire n3791;
  wire n3792;
  wire n3793;
  wire n3794;
  wire n3795;
  wire n3796;
  wire n3797;
  wire n3798;
  wire n3799;
  wire n38;
  wire n380;
  wire n3800;
  wire n3801;
  wire n3802;
  wire n3803;
  wire n3804;
  wire n3805;
  wire n3806;
  wire n3807;
  wire n3808;
  wire n3809;
  wire n381;
  wire n3810;
  wire n3811;
  wire n3812;
  wire n3813;
  wire n3814;
  wire n3815;
  wire n3816;
  wire n3817;
  wire n3818;
  wire n3819;
  wire n382;
  wire n3820;
  wire n3821;
  wire n3822;
  wire n3823;
  wire n3824;
  wire n3825;
  wire n3826;
  wire n3827;
  wire n3828;
  wire n3829;
  wire n383;
  wire n3830;
  wire n3831;
  wire n3832;
  wire n3833;
  wire n3834;
  wire n3835;
  wire n3836;
  wire n3837;
  wire n3838;
  wire n3839;
  wire n384;
  wire n3840;
  wire n3841;
  wire n3842;
  wire n3843;
  wire n3844;
  wire n3845;
  wire n3846;
  wire n3847;
  wire n3848;
  wire n3849;
  wire n385;
  wire n3850;
  wire n3851;
  wire n3852;
  wire n3853;
  wire n3854;
  wire n3855;
  wire n3856;
  wire n3857;
  wire n3858;
  wire n3859;
  wire n386;
  wire n3860;
  wire n3861;
  wire n3862;
  wire n3863;
  wire n3864;
  wire n3865;
  wire n3866;
  wire n3867;
  wire n3868;
  wire n3869;
  wire n387;
  wire n3870;
  wire n3871;
  wire n3872;
  wire n3873;
  wire n3874;
  wire n3875;
  wire n3876;
  wire n3877;
  wire n3878;
  wire n3879;
  wire n388;
  wire n3880;
  wire n3881;
  wire n3882;
  wire n3883;
  wire n3884;
  wire n3885;
  wire n3886;
  wire n3887;
  wire n3888;
  wire n3889;
  wire n389;
  wire n3890;
  wire n3891;
  wire n3892;
  wire n3893;
  wire n3894;
  wire n3895;
  wire n3896;
  wire n3897;
  wire n3898;
  wire n3899;
  wire n39;
  wire n390;
  wire n3900;
  wire n3901;
  wire n3902;
  wire n3903;
  wire n3904;
  wire n3905;
  wire n3906;
  wire n3907;
  wire n3908;
  wire n3909;
  wire n391;
  wire n3910;
  wire n3911;
  wire n3912;
  wire n3913;
  wire n3914;
  wire n3915;
  wire n3916;
  wire n3917;
  wire n3918;
  wire n3919;
  wire n392;
  wire n3920;
  wire n3921;
  wire n3922;
  wire n3923;
  wire n3924;
  wire n3925;
  wire n3926;
  wire n3927;
  wire n3928;
  wire n3929;
  wire n393;
  wire n3930;
  wire n3931;
  wire n3932;
  wire n3933;
  wire n3934;
  wire n3935;
  wire n3936;
  wire n3937;
  wire n3938;
  wire n3939;
  wire n394;
  wire n3940;
  wire n3941;
  wire n3942;
  wire n3943;
  wire n3944;
  wire n3945;
  wire n3946;
  wire n3947;
  wire n3948;
  wire n3949;
  wire n395;
  wire n3950;
  wire n3951;
  wire n3952;
  wire n3953;
  wire n3954;
  wire n3955;
  wire n3956;
  wire n3957;
  wire n3958;
  wire n3959;
  wire n396;
  wire n3960;
  wire n3961;
  wire n3962;
  wire n3963;
  wire n3964;
  wire n3965;
  wire n3966;
  wire n3967;
  wire n3968;
  wire n3969;
  wire n397;
  wire n3970;
  wire n3971;
  wire n3972;
  wire n3973;
  wire n3974;
  wire n3975;
  wire n3976;
  wire n3977;
  wire n3978;
  wire n3979;
  wire n398;
  wire n3980;
  wire n3981;
  wire n3982;
  wire n3983;
  wire n3984;
  wire n3985;
  wire n3986;
  wire n3987;
  wire n3988;
  wire n3989;
  wire n399;
  wire n3990;
  wire n3991;
  wire n3992;
  wire n3993;
  wire n3994;
  wire n3995;
  wire n3996;
  wire n3997;
  wire n3998;
  wire n3999;
  wire n4;
  wire n40;
  wire n400;
  wire n4000;
  wire n4001;
  wire n4002;
  wire n4003;
  wire n4004;
  wire n4005;
  wire n4006;
  wire n4007;
  wire n4008;
  wire n4009;
  wire n401;
  wire n4010;
  wire n4011;
  wire n4012;
  wire n4013;
  wire n4014;
  wire n4015;
  wire n4016;
  wire n4017;
  wire n4018;
  wire n4019;
  wire n402;
  wire n4020;
  wire n4021;
  wire n4022;
  wire n4023;
  wire n4024;
  wire n4025;
  wire n4026;
  wire n4027;
  wire n4028;
  wire n4029;
  wire n403;
  wire n4030;
  wire n4031;
  wire n4032;
  wire n4033;
  wire n4034;
  wire n4035;
  wire n4036;
  wire n4037;
  wire n4038;
  wire n4039;
  wire n404;
  wire n4040;
  wire n4041;
  wire n4042;
  wire n4043;
  wire n4044;
  wire n4045;
  wire n4046;
  wire n4047;
  wire n4048;
  wire n4049;
  wire n405;
  wire n4050;
  wire n4051;
  wire n4052;
  wire n4053;
  wire n4054;
  wire n4055;
  wire n4056;
  wire n4057;
  wire n4058;
  wire n4059;
  wire n406;
  wire n4060;
  wire n4061;
  wire n4062;
  wire n4063;
  wire n4064;
  wire n4065;
  wire n4066;
  wire n4067;
  wire n4068;
  wire n4069;
  wire n407;
  wire n4070;
  wire n4071;
  wire n4072;
  wire n4073;
  wire n4074;
  wire n4075;
  wire n4076;
  wire n4077;
  wire n4078;
  wire n4079;
  wire n408;
  wire n4080;
  wire n4081;
  wire n4082;
  wire n4083;
  wire n4084;
  wire n4085;
  wire n4086;
  wire n4087;
  wire n4088;
  wire n4089;
  wire n409;
  wire n4090;
  wire n4091;
  wire n4092;
  wire n4093;
  wire n4094;
  wire n4095;
  wire n4096;
  wire n4097;
  wire n4098;
  wire n4099;
  wire n41;
  wire n410;
  wire n4100;
  wire n4101;
  wire n4102;
  wire n4103;
  wire n4104;
  wire n4105;
  wire n4106;
  wire n4107;
  wire n4108;
  wire n4109;
  wire n411;
  wire n4110;
  wire n4111;
  wire n4112;
  wire n4113;
  wire n4114;
  wire n4115;
  wire n4116;
  wire n4117;
  wire n4118;
  wire n4119;
  wire n412;
  wire n4120;
  wire n4121;
  wire n4122;
  wire n4123;
  wire n4124;
  wire n4125;
  wire n4126;
  wire n4127;
  wire n4128;
  wire n4129;
  wire n413;
  wire n4130;
  wire n4131;
  wire n4132;
  wire n4133;
  wire n4134;
  wire n4135;
  wire n4136;
  wire n4137;
  wire n4138;
  wire n4139;
  wire n414;
  wire n4140;
  wire n4141;
  wire n4142;
  wire n4143;
  wire n4144;
  wire n4145;
  wire n4146;
  wire n4147;
  wire n4148;
  wire n4149;
  wire n415;
  wire n4150;
  wire n4151;
  wire n4152;
  wire n4153;
  wire n4154;
  wire n4155;
  wire n4156;
  wire n4157;
  wire n4158;
  wire n4159;
  wire n416;
  wire n4160;
  wire n4161;
  wire n4162;
  wire n4163;
  wire n4164;
  wire n4165;
  wire n4166;
  wire n4167;
  wire n4168;
  wire n4169;
  wire n417;
  wire n4170;
  wire n4171;
  wire n4172;
  wire n4173;
  wire n4174;
  wire n4175;
  wire n4176;
  wire n4177;
  wire n4178;
  wire n4179;
  wire n418;
  wire n4180;
  wire n4181;
  wire n4182;
  wire n4183;
  wire n4184;
  wire n4185;
  wire n4186;
  wire n4187;
  wire n4188;
  wire n4189;
  wire n419;
  wire n4190;
  wire n4191;
  wire n4192;
  wire n4193;
  wire n4194;
  wire n4195;
  wire n4196;
  wire n4197;
  wire n4198;
  wire n4199;
  wire n42;
  wire n420;
  wire n4200;
  wire n4201;
  wire n4202;
  wire n4203;
  wire n4204;
  wire n4205;
  wire n4206;
  wire n4207;
  wire n4208;
  wire n4209;
  wire n421;
  wire n4210;
  wire n4211;
  wire n4212;
  wire n4213;
  wire n4214;
  wire n4215;
  wire n4216;
  wire n4217;
  wire n4218;
  wire n4219;
  wire n422;
  wire n4220;
  wire n4221;
  wire n4222;
  wire n4223;
  wire n4224;
  wire n4225;
  wire n4226;
  wire n4227;
  wire n4228;
  wire n4229;
  wire n423;
  wire n4230;
  wire n4231;
  wire n4232;
  wire n4233;
  wire n4234;
  wire n4235;
  wire n4236;
  wire n4237;
  wire n4238;
  wire n4239;
  wire n424;
  wire n4240;
  wire n4241;
  wire n4242;
  wire n4243;
  wire n4244;
  wire n4245;
  wire n4246;
  wire n4247;
  wire n4248;
  wire n4249;
  wire n425;
  wire n4250;
  wire n4251;
  wire n4252;
  wire n4253;
  wire n4254;
  wire n4255;
  wire n4256;
  wire n4257;
  wire n4258;
  wire n4259;
  wire n426;
  wire n4260;
  wire n4261;
  wire n4262;
  wire n4263;
  wire n4264;
  wire n4265;
  wire n4266;
  wire n4267;
  wire n4268;
  wire n4269;
  wire n427;
  wire n4270;
  wire n4271;
  wire n4272;
  wire n4273;
  wire n4274;
  wire n4275;
  wire n4276;
  wire n4278;
  wire n4279;
  wire n428;
  wire n4280;
  wire n4281;
  wire n4282;
  wire n4283;
  wire n4284;
  wire n4285;
  wire n4286;
  wire n4287;
  wire n4288;
  wire n4289;
  wire n429;
  wire n4290;
  wire n4291;
  wire n4292;
  wire n4293;
  wire n4294;
  wire n4295;
  wire n4296;
  wire n4297;
  wire n4298;
  wire n4299;
  wire n43;
  wire n430;
  wire n4300;
  wire n4301;
  wire n4302;
  wire n4303;
  wire n4304;
  wire n4305;
  wire n4306;
  wire n4307;
  wire n4308;
  wire n4309;
  wire n431;
  wire n4310;
  wire n4311;
  wire n4312;
  wire n4313;
  wire n4314;
  wire n4315;
  wire n4316;
  wire n4317;
  wire n4318;
  wire n4319;
  wire n432;
  wire n4320;
  wire n4321;
  wire n4322;
  wire n4323;
  wire n4324;
  wire n4325;
  wire n4326;
  wire n4327;
  wire n4328;
  wire n4329;
  wire n433;
  wire n4330;
  wire n4331;
  wire n4332;
  wire n4333;
  wire n4334;
  wire n4335;
  wire n4336;
  wire n4337;
  wire n4338;
  wire n4339;
  wire n434;
  wire n4340;
  wire n4341;
  wire n4342;
  wire n4343;
  wire n4344;
  wire n4345;
  wire n4346;
  wire n4347;
  wire n4348;
  wire n4349;
  wire n435;
  wire n4350;
  wire n4351;
  wire n4352;
  wire n4353;
  wire n4354;
  wire n4355;
  wire n4356;
  wire n4357;
  wire n4358;
  wire n4359;
  wire n436;
  wire n4360;
  wire n4361;
  wire n4362;
  wire n4363;
  wire n4364;
  wire n4365;
  wire n4366;
  wire n4367;
  wire n4368;
  wire n4369;
  wire n437;
  wire n4370;
  wire n4371;
  wire n4372;
  wire n4373;
  wire n4374;
  wire n4375;
  wire n4376;
  wire n4377;
  wire n4378;
  wire n4379;
  wire n438;
  wire n4380;
  wire n4381;
  wire n4382;
  wire n4383;
  wire n4384;
  wire n4385;
  wire n4386;
  wire n4387;
  wire n4388;
  wire n4389;
  wire n439;
  wire n4390;
  wire n4391;
  wire n4392;
  wire n4393;
  wire n4394;
  wire n4395;
  wire n4396;
  wire n4397;
  wire n4398;
  wire n4399;
  wire n44;
  wire n440;
  wire n4400;
  wire n4401;
  wire n4402;
  wire n4403;
  wire n4404;
  wire n4405;
  wire n4406;
  wire n4407;
  wire n4408;
  wire n4409;
  wire n441;
  wire n4410;
  wire n4411;
  wire n4412;
  wire n4413;
  wire n4414;
  wire n4415;
  wire n4416;
  wire n4417;
  wire n4418;
  wire n4419;
  wire n442;
  wire n4420;
  wire n4421;
  wire n4422;
  wire n4423;
  wire n4424;
  wire n4425;
  wire n4426;
  wire n4427;
  wire n4428;
  wire n4429;
  wire n443;
  wire n4430;
  wire n4431;
  wire n4432;
  wire n4433;
  wire n4434;
  wire n4435;
  wire n4436;
  wire n4437;
  wire n4438;
  wire n4439;
  wire n444;
  wire n4440;
  wire n4441;
  wire n4442;
  wire n4443;
  wire n4444;
  wire n4445;
  wire n4446;
  wire n4447;
  wire n4448;
  wire n4449;
  wire n445;
  wire n4450;
  wire n4451;
  wire n4452;
  wire n4453;
  wire n4454;
  wire n4455;
  wire n4456;
  wire n4457;
  wire n4458;
  wire n4459;
  wire n446;
  wire n4460;
  wire n4461;
  wire n4462;
  wire n4463;
  wire n4464;
  wire n4465;
  wire n4466;
  wire n4467;
  wire n4468;
  wire n4469;
  wire n447;
  wire n4470;
  wire n4471;
  wire n4472;
  wire n4473;
  wire n4474;
  wire n4475;
  wire n4476;
  wire n4477;
  wire n4478;
  wire n4479;
  wire n448;
  wire n4480;
  wire n4481;
  wire n4482;
  wire n4483;
  wire n4484;
  wire n4485;
  wire n4486;
  wire n4487;
  wire n4488;
  wire n4489;
  wire n449;
  wire n4490;
  wire n4491;
  wire n4492;
  wire n4493;
  wire n4494;
  wire n4495;
  wire n4496;
  wire n4497;
  wire n4498;
  wire n4499;
  wire n45;
  wire n450;
  wire n4500;
  wire n4501;
  wire n4502;
  wire n4503;
  wire n4504;
  wire n4505;
  wire n4506;
  wire n4507;
  wire n4508;
  wire n4509;
  wire n451;
  wire n4510;
  wire n4511;
  wire n4512;
  wire n4513;
  wire n4514;
  wire n4515;
  wire n4516;
  wire n4517;
  wire n4518;
  wire n4519;
  wire n452;
  wire n4520;
  wire n4521;
  wire n4522;
  wire n4523;
  wire n4524;
  wire n4525;
  wire n4526;
  wire n4527;
  wire n4528;
  wire n4529;
  wire n453;
  wire n4530;
  wire n4531;
  wire n4532;
  wire n4533;
  wire n4534;
  wire n4535;
  wire n4536;
  wire n4537;
  wire n4538;
  wire n4539;
  wire n454;
  wire n4540;
  wire n4541;
  wire n4542;
  wire n4543;
  wire n4544;
  wire n4545;
  wire n4546;
  wire n4547;
  wire n4548;
  wire n4549;
  wire n455;
  wire n4550;
  wire n4551;
  wire n4552;
  wire n4553;
  wire n4554;
  wire n4555;
  wire n4556;
  wire n4557;
  wire n4558;
  wire n4559;
  wire n456;
  wire n4560;
  wire n4561;
  wire n4562;
  wire n4563;
  wire n4564;
  wire n4565;
  wire n4566;
  wire n4567;
  wire n4568;
  wire n4569;
  wire n457;
  wire n4570;
  wire n4571;
  wire n4572;
  wire n4573;
  wire n4574;
  wire n4575;
  wire n4576;
  wire n4577;
  wire n4578;
  wire n4579;
  wire n458;
  wire n4580;
  wire n4581;
  wire n4582;
  wire n4583;
  wire n4584;
  wire n4585;
  wire n4586;
  wire n4587;
  wire n4588;
  wire n4589;
  wire n459;
  wire n4590;
  wire n4591;
  wire n4592;
  wire n4593;
  wire n4594;
  wire n4595;
  wire n4596;
  wire n4597;
  wire n4598;
  wire n4599;
  wire n46;
  wire n460;
  wire n4600;
  wire n4601;
  wire n4602;
  wire n4603;
  wire n4604;
  wire n4605;
  wire n4606;
  wire n4607;
  wire n4608;
  wire n4609;
  wire n461;
  wire n4610;
  wire n4611;
  wire n4612;
  wire n4613;
  wire n4614;
  wire n4615;
  wire n4616;
  wire n4617;
  wire n4618;
  wire n4619;
  wire n462;
  wire n4620;
  wire n4621;
  wire n4622;
  wire n4623;
  wire n4624;
  wire n4625;
  wire n4626;
  wire n4627;
  wire n4628;
  wire n4629;
  wire n463;
  wire n4630;
  wire n4631;
  wire n4632;
  wire n4633;
  wire n4634;
  wire n4635;
  wire n4636;
  wire n4637;
  wire n4638;
  wire n4639;
  wire n464;
  wire n4640;
  wire n4641;
  wire n4642;
  wire n4643;
  wire n4644;
  wire n4645;
  wire n4646;
  wire n4647;
  wire n4648;
  wire n4649;
  wire n465;
  wire n4650;
  wire n4651;
  wire n4652;
  wire n4653;
  wire n4654;
  wire n4655;
  wire n4656;
  wire n4657;
  wire n4658;
  wire n4659;
  wire n466;
  wire n4660;
  wire n4661;
  wire n4662;
  wire n4663;
  wire n4664;
  wire n4665;
  wire n4666;
  wire n4667;
  wire n4668;
  wire n4669;
  wire n467;
  wire n4670;
  wire n4671;
  wire n4672;
  wire n4673;
  wire n4674;
  wire n4675;
  wire n4676;
  wire n4677;
  wire n4678;
  wire n4679;
  wire n468;
  wire n4680;
  wire n4681;
  wire n4682;
  wire n4683;
  wire n4684;
  wire n4685;
  wire n4686;
  wire n4687;
  wire n4688;
  wire n4689;
  wire n469;
  wire n4690;
  wire n4691;
  wire n4692;
  wire n4693;
  wire n4694;
  wire n4695;
  wire n4696;
  wire n4697;
  wire n4698;
  wire n4699;
  wire n47;
  wire n470;
  wire n4700;
  wire n4701;
  wire n4702;
  wire n4703;
  wire n4704;
  wire n4705;
  wire n4706;
  wire n4707;
  wire n4708;
  wire n4709;
  wire n471;
  wire n4710;
  wire n4711;
  wire n4712;
  wire n4713;
  wire n4714;
  wire n4715;
  wire n4716;
  wire n4717;
  wire n4718;
  wire n4719;
  wire n472;
  wire n4720;
  wire n4721;
  wire n4722;
  wire n4723;
  wire n4724;
  wire n4725;
  wire n4726;
  wire n4727;
  wire n4728;
  wire n4729;
  wire n473;
  wire n4730;
  wire n4731;
  wire n4732;
  wire n4733;
  wire n4734;
  wire n4735;
  wire n4736;
  wire n4737;
  wire n4738;
  wire n4739;
  wire n474;
  wire n4740;
  wire n4741;
  wire n4742;
  wire n4743;
  wire n4744;
  wire n4745;
  wire n4746;
  wire n4747;
  wire n4748;
  wire n4749;
  wire n475;
  wire n4750;
  wire n4751;
  wire n4752;
  wire n4753;
  wire n4754;
  wire n4755;
  wire n4756;
  wire n4757;
  wire n4758;
  wire n4759;
  wire n476;
  wire n4760;
  wire n4761;
  wire n4762;
  wire n4763;
  wire n4764;
  wire n4765;
  wire n4766;
  wire n4767;
  wire n4768;
  wire n4769;
  wire n477;
  wire n4770;
  wire n4771;
  wire n4772;
  wire n4773;
  wire n4774;
  wire n4775;
  wire n4776;
  wire n4777;
  wire n4778;
  wire n4779;
  wire n478;
  wire n4780;
  wire n4781;
  wire n4782;
  wire n4783;
  wire n4784;
  wire n4785;
  wire n4786;
  wire n4787;
  wire n4788;
  wire n4789;
  wire n479;
  wire n4790;
  wire n4791;
  wire n4792;
  wire n4793;
  wire n4794;
  wire n4795;
  wire n4796;
  wire n4797;
  wire n4798;
  wire n4799;
  wire n48;
  wire n480;
  wire n4800;
  wire n4801;
  wire n4802;
  wire n4803;
  wire n4804;
  wire n4805;
  wire n4806;
  wire n4807;
  wire n4808;
  wire n4809;
  wire n481;
  wire n4810;
  wire n4811;
  wire n4812;
  wire n4813;
  wire n4814;
  wire n4815;
  wire n4816;
  wire n4817;
  wire n4818;
  wire n4819;
  wire n482;
  wire n4820;
  wire n4821;
  wire n4822;
  wire n4823;
  wire n4824;
  wire n4825;
  wire n4826;
  wire n4827;
  wire n4828;
  wire n4829;
  wire n483;
  wire n4830;
  wire n4831;
  wire n4832;
  wire n4833;
  wire n4834;
  wire n4835;
  wire n4836;
  wire n4837;
  wire n4838;
  wire n4839;
  wire n484;
  wire n4840;
  wire n4841;
  wire n4842;
  wire n4843;
  wire n4844;
  wire n4845;
  wire n4846;
  wire n4847;
  wire n4848;
  wire n4849;
  wire n485;
  wire n4850;
  wire n4851;
  wire n4852;
  wire n4853;
  wire n4854;
  wire n4855;
  wire n4856;
  wire n4857;
  wire n4858;
  wire n4859;
  wire n486;
  wire n4860;
  wire n4861;
  wire n4862;
  wire n4863;
  wire n4864;
  wire n4865;
  wire n4866;
  wire n4867;
  wire n4868;
  wire n4869;
  wire n487;
  wire n4870;
  wire n4871;
  wire n4872;
  wire n4873;
  wire n4874;
  wire n4875;
  wire n4876;
  wire n4877;
  wire n4878;
  wire n4879;
  wire n488;
  wire n4880;
  wire n4881;
  wire n4882;
  wire n4883;
  wire n4884;
  wire n4885;
  wire n4886;
  wire n4887;
  wire n4888;
  wire n4889;
  wire n489;
  wire n4890;
  wire n4891;
  wire n4892;
  wire n4893;
  wire n4894;
  wire n4895;
  wire n4896;
  wire n4897;
  wire n4898;
  wire n4899;
  wire n49;
  wire n490;
  wire n4900;
  wire n4901;
  wire n4902;
  wire n4903;
  wire n4904;
  wire n4905;
  wire n4906;
  wire n4907;
  wire n4908;
  wire n4909;
  wire n491;
  wire n4910;
  wire n4911;
  wire n4912;
  wire n4913;
  wire n4914;
  wire n4915;
  wire n4916;
  wire n4917;
  wire n4918;
  wire n4919;
  wire n492;
  wire n4920;
  wire n4921;
  wire n4922;
  wire n4923;
  wire n4924;
  wire n4925;
  wire n4926;
  wire n4927;
  wire n4928;
  wire n4929;
  wire n493;
  wire n4930;
  wire n4931;
  wire n4932;
  wire n4933;
  wire n4934;
  wire n4935;
  wire n4936;
  wire n4937;
  wire n4938;
  wire n4939;
  wire n494;
  wire n4940;
  wire n4941;
  wire n4942;
  wire n4943;
  wire n4944;
  wire n4945;
  wire n4946;
  wire n4947;
  wire n4948;
  wire n4949;
  wire n495;
  wire n4950;
  wire n4951;
  wire n4952;
  wire n4953;
  wire n4954;
  wire n4955;
  wire n4956;
  wire n4957;
  wire n4958;
  wire n4959;
  wire n496;
  wire n4960;
  wire n4961;
  wire n4962;
  wire n4963;
  wire n4964;
  wire n4965;
  wire n4966;
  wire n4967;
  wire n4968;
  wire n4969;
  wire n497;
  wire n4970;
  wire n4971;
  wire n4972;
  wire n4973;
  wire n4974;
  wire n4975;
  wire n4976;
  wire n4977;
  wire n4978;
  wire n4979;
  wire n498;
  wire n4980;
  wire n4981;
  wire n4982;
  wire n4983;
  wire n4984;
  wire n4985;
  wire n4986;
  wire n4987;
  wire n4988;
  wire n4989;
  wire n499;
  wire n4990;
  wire n4991;
  wire n4992;
  wire n4993;
  wire n4994;
  wire n4995;
  wire n4996;
  wire n4997;
  wire n4998;
  wire n4999;
  wire n5;
  wire n50;
  wire n500;
  wire n5000;
  wire n5001;
  wire n5002;
  wire n5003;
  wire n5004;
  wire n5005;
  wire n5006;
  wire n5007;
  wire n5008;
  wire n5009;
  wire n501;
  wire n5010;
  wire n5011;
  wire n5012;
  wire n5013;
  wire n5014;
  wire n5015;
  wire n5016;
  wire n5017;
  wire n5018;
  wire n5019;
  wire n502;
  wire n5020;
  wire n5021;
  wire n5022;
  wire n5023;
  wire n5024;
  wire n5025;
  wire n5026;
  wire n5027;
  wire n5028;
  wire n5029;
  wire n503;
  wire n5030;
  wire n5031;
  wire n5032;
  wire n5033;
  wire n5034;
  wire n5035;
  wire n5036;
  wire n5037;
  wire n5038;
  wire n5039;
  wire n504;
  wire n5040;
  wire n5041;
  wire n5042;
  wire n5043;
  wire n5044;
  wire n5045;
  wire n5046;
  wire n5047;
  wire n5048;
  wire n5049;
  wire n505;
  wire n5050;
  wire n5051;
  wire n5052;
  wire n5053;
  wire n5054;
  wire n5055;
  wire n5056;
  wire n5057;
  wire n5058;
  wire n5059;
  wire n506;
  wire n5060;
  wire n5061;
  wire n5062;
  wire n5063;
  wire n5064;
  wire n5065;
  wire n5066;
  wire n5067;
  wire n5068;
  wire n5069;
  wire n507;
  wire n5070;
  wire n5071;
  wire n5072;
  wire n5073;
  wire n5074;
  wire n5075;
  wire n5076;
  wire n5077;
  wire n5078;
  wire n5079;
  wire n508;
  wire n5080;
  wire n5081;
  wire n5082;
  wire n5083;
  wire n5084;
  wire n5085;
  wire n5086;
  wire n5087;
  wire n5088;
  wire n5089;
  wire n509;
  wire n5090;
  wire n5091;
  wire n5092;
  wire n5093;
  wire n5094;
  wire n5095;
  wire n5096;
  wire n5097;
  wire n5098;
  wire n5099;
  wire n51;
  wire n510;
  wire n5100;
  wire n5101;
  wire n5102;
  wire n5103;
  wire n5104;
  wire n5105;
  wire n5106;
  wire n5107;
  wire n5108;
  wire n5109;
  wire n511;
  wire n5110;
  wire n5111;
  wire n5112;
  wire n5113;
  wire n5114;
  wire n5115;
  wire n5116;
  wire n5117;
  wire n5118;
  wire n5119;
  wire n512;
  wire n5120;
  wire n5121;
  wire n5122;
  wire n5123;
  wire n5124;
  wire n5125;
  wire n5126;
  wire n5127;
  wire n5128;
  wire n5129;
  wire n513;
  wire n5130;
  wire n5131;
  wire n5132;
  wire n5133;
  wire n5134;
  wire n5135;
  wire n5136;
  wire n5137;
  wire n5138;
  wire n5139;
  wire n514;
  wire n5140;
  wire n5141;
  wire n5142;
  wire n5143;
  wire n5144;
  wire n5145;
  wire n5146;
  wire n5147;
  wire n5148;
  wire n5149;
  wire n515;
  wire n5150;
  wire n5151;
  wire n5152;
  wire n5153;
  wire n5154;
  wire n5155;
  wire n5156;
  wire n5157;
  wire n5158;
  wire n5159;
  wire n516;
  wire n5160;
  wire n5161;
  wire n5162;
  wire n5163;
  wire n5164;
  wire n5165;
  wire n5166;
  wire n5167;
  wire n5168;
  wire n5169;
  wire n517;
  wire n5170;
  wire n5171;
  wire n5172;
  wire n5173;
  wire n5174;
  wire n5175;
  wire n5176;
  wire n5177;
  wire n5178;
  wire n5179;
  wire n518;
  wire n5180;
  wire n5181;
  wire n5182;
  wire n5183;
  wire n5184;
  wire n5185;
  wire n5186;
  wire n5187;
  wire n5188;
  wire n5189;
  wire n519;
  wire n5190;
  wire n5191;
  wire n5192;
  wire n5193;
  wire n5194;
  wire n5195;
  wire n5196;
  wire n5197;
  wire n5198;
  wire n5199;
  wire n52;
  wire n520;
  wire n5201;
  wire n5202;
  wire n5203;
  wire n5204;
  wire n5205;
  wire n5206;
  wire n5207;
  wire n5208;
  wire n5209;
  wire n521;
  wire n5210;
  wire n5211;
  wire n5212;
  wire n5213;
  wire n5214;
  wire n5215;
  wire n5216;
  wire n5217;
  wire n5218;
  wire n5219;
  wire n522;
  wire n5220;
  wire n5221;
  wire n5222;
  wire n5223;
  wire n5224;
  wire n5225;
  wire n5226;
  wire n5227;
  wire n5228;
  wire n5229;
  wire n523;
  wire n5230;
  wire n5231;
  wire n5232;
  wire n5233;
  wire n5234;
  wire n5235;
  wire n5236;
  wire n5237;
  wire n5238;
  wire n5239;
  wire n524;
  wire n5240;
  wire n5241;
  wire n5242;
  wire n5243;
  wire n5244;
  wire n5245;
  wire n5246;
  wire n5247;
  wire n5248;
  wire n5249;
  wire n525;
  wire n5250;
  wire n5251;
  wire n5252;
  wire n5253;
  wire n5254;
  wire n5255;
  wire n5256;
  wire n5257;
  wire n5258;
  wire n5259;
  wire n526;
  wire n5260;
  wire n5261;
  wire n5262;
  wire n5263;
  wire n5264;
  wire n5265;
  wire n5266;
  wire n5267;
  wire n5268;
  wire n5269;
  wire n527;
  wire n5270;
  wire n5271;
  wire n5272;
  wire n5273;
  wire n5274;
  wire n5275;
  wire n5276;
  wire n5277;
  wire n5278;
  wire n5279;
  wire n528;
  wire n5280;
  wire n5281;
  wire n5282;
  wire n5283;
  wire n5284;
  wire n5285;
  wire n5286;
  wire n5287;
  wire n5288;
  wire n5289;
  wire n529;
  wire n5290;
  wire n5291;
  wire n5292;
  wire n5293;
  wire n5294;
  wire n5295;
  wire n5296;
  wire n5297;
  wire n5298;
  wire n5299;
  wire n53;
  wire n530;
  wire n5300;
  wire n5301;
  wire n5302;
  wire n5303;
  wire n5304;
  wire n5305;
  wire n5306;
  wire n5307;
  wire n5308;
  wire n5309;
  wire n531;
  wire n5310;
  wire n5311;
  wire n5312;
  wire n5313;
  wire n5314;
  wire n5315;
  wire n5316;
  wire n5317;
  wire n5318;
  wire n5319;
  wire n532;
  wire n5320;
  wire n5321;
  wire n5322;
  wire n5323;
  wire n5324;
  wire n5325;
  wire n5326;
  wire n5327;
  wire n5328;
  wire n5329;
  wire n533;
  wire n5330;
  wire n5331;
  wire n5332;
  wire n5333;
  wire n5334;
  wire n5335;
  wire n5336;
  wire n5337;
  wire n5338;
  wire n5339;
  wire n534;
  wire n5340;
  wire n5341;
  wire n5342;
  wire n5343;
  wire n5344;
  wire n5345;
  wire n5346;
  wire n5347;
  wire n5348;
  wire n5349;
  wire n535;
  wire n5350;
  wire n5351;
  wire n5352;
  wire n5353;
  wire n5354;
  wire n5355;
  wire n5356;
  wire n5357;
  wire n5358;
  wire n5359;
  wire n536;
  wire n5360;
  wire n5361;
  wire n5362;
  wire n5363;
  wire n5364;
  wire n5365;
  wire n5366;
  wire n5367;
  wire n5368;
  wire n5369;
  wire n537;
  wire n5370;
  wire n5371;
  wire n5372;
  wire n5373;
  wire n5374;
  wire n5375;
  wire n5376;
  wire n5377;
  wire n5378;
  wire n5379;
  wire n538;
  wire n5380;
  wire n5381;
  wire n5382;
  wire n5383;
  wire n5384;
  wire n5385;
  wire n5386;
  wire n5387;
  wire n5388;
  wire n5389;
  wire n539;
  wire n5390;
  wire n5391;
  wire n5392;
  wire n5393;
  wire n5394;
  wire n5395;
  wire n5396;
  wire n5397;
  wire n5398;
  wire n5399;
  wire n54;
  wire n540;
  wire n5400;
  wire n5401;
  wire n5402;
  wire n5403;
  wire n5404;
  wire n5405;
  wire n5406;
  wire n5407;
  wire n5408;
  wire n5409;
  wire n541;
  wire n5410;
  wire n5411;
  wire n5412;
  wire n5413;
  wire n5414;
  wire n5415;
  wire n5416;
  wire n5417;
  wire n5418;
  wire n5419;
  wire n542;
  wire n5420;
  wire n5421;
  wire n5422;
  wire n5423;
  wire n5424;
  wire n5425;
  wire n5426;
  wire n5427;
  wire n5428;
  wire n5429;
  wire n543;
  wire n5430;
  wire n5431;
  wire n5432;
  wire n5433;
  wire n5434;
  wire n5435;
  wire n5436;
  wire n5437;
  wire n5438;
  wire n5439;
  wire n544;
  wire n5440;
  wire n5441;
  wire n5442;
  wire n5443;
  wire n5444;
  wire n5445;
  wire n5446;
  wire n5447;
  wire n5448;
  wire n5449;
  wire n545;
  wire n5450;
  wire n5451;
  wire n5452;
  wire n5453;
  wire n5454;
  wire n5455;
  wire n5456;
  wire n5457;
  wire n5458;
  wire n5459;
  wire n546;
  wire n5460;
  wire n5461;
  wire n5462;
  wire n5463;
  wire n5464;
  wire n5465;
  wire n5466;
  wire n5467;
  wire n5468;
  wire n5469;
  wire n547;
  wire n5470;
  wire n5471;
  wire n5472;
  wire n5473;
  wire n5474;
  wire n5475;
  wire n5476;
  wire n5477;
  wire n5478;
  wire n5479;
  wire n548;
  wire n5480;
  wire n5481;
  wire n5482;
  wire n5483;
  wire n5484;
  wire n5485;
  wire n5486;
  wire n5487;
  wire n5489;
  wire n549;
  wire n5490;
  wire n5491;
  wire n5492;
  wire n5493;
  wire n5494;
  wire n5495;
  wire n5496;
  wire n5497;
  wire n5498;
  wire n5499;
  wire n55;
  wire n550;
  wire n5500;
  wire n5501;
  wire n5502;
  wire n5503;
  wire n5504;
  wire n5505;
  wire n5506;
  wire n5507;
  wire n5508;
  wire n5509;
  wire n551;
  wire n5510;
  wire n5511;
  wire n5512;
  wire n5513;
  wire n5514;
  wire n5515;
  wire n5516;
  wire n5517;
  wire n5518;
  wire n5519;
  wire n552;
  wire n5520;
  wire n5521;
  wire n5522;
  wire n5523;
  wire n5524;
  wire n5525;
  wire n5526;
  wire n5527;
  wire n5528;
  wire n5529;
  wire n553;
  wire n5530;
  wire n5531;
  wire n5532;
  wire n5533;
  wire n5534;
  wire n5535;
  wire n5536;
  wire n5537;
  wire n5538;
  wire n5539;
  wire n554;
  wire n5540;
  wire n5541;
  wire n5542;
  wire n5543;
  wire n5544;
  wire n5545;
  wire n5546;
  wire n5547;
  wire n5548;
  wire n5549;
  wire n555;
  wire n5550;
  wire n5551;
  wire n5552;
  wire n5553;
  wire n5554;
  wire n5555;
  wire n5556;
  wire n5557;
  wire n5558;
  wire n5559;
  wire n556;
  wire n5560;
  wire n5561;
  wire n5562;
  wire n5563;
  wire n5564;
  wire n5565;
  wire n5566;
  wire n5567;
  wire n5568;
  wire n5569;
  wire n557;
  wire n5570;
  wire n5571;
  wire n5572;
  wire n5573;
  wire n5574;
  wire n5575;
  wire n5576;
  wire n5577;
  wire n5578;
  wire n5579;
  wire n558;
  wire n5580;
  wire n5581;
  wire n5582;
  wire n5583;
  wire n5584;
  wire n5585;
  wire n5586;
  wire n5587;
  wire n5588;
  wire n5589;
  wire n559;
  wire n5590;
  wire n5591;
  wire n5592;
  wire n5593;
  wire n5594;
  wire n5595;
  wire n5596;
  wire n5597;
  wire n5598;
  wire n5599;
  wire n56;
  wire n560;
  wire n5600;
  wire n5601;
  wire n5602;
  wire n5603;
  wire n5604;
  wire n5605;
  wire n5606;
  wire n5607;
  wire n5608;
  wire n5609;
  wire n561;
  wire n5610;
  wire n5611;
  wire n5612;
  wire n5613;
  wire n5614;
  wire n5615;
  wire n5616;
  wire n5617;
  wire n5618;
  wire n5619;
  wire n562;
  wire n5620;
  wire n5621;
  wire n5622;
  wire n5623;
  wire n5624;
  wire n5625;
  wire n5626;
  wire n5627;
  wire n5628;
  wire n5629;
  wire n563;
  wire n5630;
  wire n5631;
  wire n5632;
  wire n5633;
  wire n5634;
  wire n5635;
  wire n5636;
  wire n5637;
  wire n5638;
  wire n5639;
  wire n564;
  wire n5640;
  wire n5641;
  wire n5642;
  wire n5643;
  wire n5644;
  wire n5645;
  wire n5646;
  wire n5647;
  wire n5648;
  wire n5649;
  wire n565;
  wire n5650;
  wire n5651;
  wire n5652;
  wire n5653;
  wire n5654;
  wire n5655;
  wire n5656;
  wire n5657;
  wire n5658;
  wire n5659;
  wire n566;
  wire n5660;
  wire n5661;
  wire n5662;
  wire n5663;
  wire n5664;
  wire n5665;
  wire n5666;
  wire n5667;
  wire n5668;
  wire n5669;
  wire n567;
  wire n5670;
  wire n5671;
  wire n5672;
  wire n5673;
  wire n5674;
  wire n5675;
  wire n5676;
  wire n5677;
  wire n5678;
  wire n5679;
  wire n568;
  wire n5680;
  wire n5681;
  wire n5682;
  wire n5683;
  wire n5684;
  wire n5685;
  wire n5686;
  wire n5687;
  wire n5688;
  wire n5689;
  wire n569;
  wire n5690;
  wire n5691;
  wire n5692;
  wire n5693;
  wire n5694;
  wire n5695;
  wire n5696;
  wire n5697;
  wire n5698;
  wire n5699;
  wire n57;
  wire n570;
  wire n5700;
  wire n5701;
  wire n5702;
  wire n5703;
  wire n5704;
  wire n5705;
  wire n5706;
  wire n5707;
  wire n5708;
  wire n5709;
  wire n571;
  wire n5710;
  wire n5711;
  wire n5712;
  wire n5713;
  wire n5714;
  wire n5715;
  wire n5716;
  wire n5717;
  wire n5718;
  wire n5719;
  wire n572;
  wire n5720;
  wire n5721;
  wire n5722;
  wire n5723;
  wire n5724;
  wire n5725;
  wire n5726;
  wire n5727;
  wire n5728;
  wire n5729;
  wire n573;
  wire n5730;
  wire n5731;
  wire n5732;
  wire n5733;
  wire n5734;
  wire n5735;
  wire n5736;
  wire n5737;
  wire n5738;
  wire n5739;
  wire n574;
  wire n5740;
  wire n5741;
  wire n5742;
  wire n5743;
  wire n5744;
  wire n5745;
  wire n5746;
  wire n5747;
  wire n5748;
  wire n5749;
  wire n575;
  wire n5750;
  wire n5751;
  wire n5752;
  wire n5753;
  wire n5754;
  wire n5755;
  wire n5756;
  wire n5757;
  wire n5758;
  wire n5759;
  wire n576;
  wire n5760;
  wire n5761;
  wire n5762;
  wire n5763;
  wire n5764;
  wire n5765;
  wire n5766;
  wire n5767;
  wire n5768;
  wire n5769;
  wire n577;
  wire n5770;
  wire n5771;
  wire n5772;
  wire n5773;
  wire n5774;
  wire n5775;
  wire n5776;
  wire n5777;
  wire n5778;
  wire n5779;
  wire n578;
  wire n5780;
  wire n5781;
  wire n5782;
  wire n5783;
  wire n5784;
  wire n5785;
  wire n5786;
  wire n5787;
  wire n5788;
  wire n5789;
  wire n579;
  wire n5790;
  wire n5791;
  wire n5792;
  wire n5793;
  wire n5794;
  wire n5795;
  wire n5796;
  wire n5797;
  wire n5798;
  wire n5799;
  wire n58;
  wire n580;
  wire n5800;
  wire n5801;
  wire n5802;
  wire n5803;
  wire n5804;
  wire n5805;
  wire n5806;
  wire n5807;
  wire n5808;
  wire n5809;
  wire n581;
  wire n5810;
  wire n5811;
  wire n5812;
  wire n5813;
  wire n5814;
  wire n5815;
  wire n5816;
  wire n5817;
  wire n5818;
  wire n5819;
  wire n582;
  wire n5820;
  wire n5821;
  wire n5822;
  wire n5823;
  wire n5824;
  wire n5825;
  wire n5826;
  wire n5827;
  wire n5828;
  wire n5829;
  wire n583;
  wire n5830;
  wire n5831;
  wire n5832;
  wire n5833;
  wire n5834;
  wire n5835;
  wire n5836;
  wire n5837;
  wire n5838;
  wire n5839;
  wire n584;
  wire n5840;
  wire n5841;
  wire n5842;
  wire n5843;
  wire n5844;
  wire n5845;
  wire n5846;
  wire n5847;
  wire n5848;
  wire n5849;
  wire n585;
  wire n5850;
  wire n5851;
  wire n5852;
  wire n5853;
  wire n5854;
  wire n5855;
  wire n5856;
  wire n5857;
  wire n5858;
  wire n5859;
  wire n586;
  wire n5860;
  wire n5861;
  wire n5862;
  wire n5863;
  wire n5864;
  wire n5865;
  wire n5866;
  wire n5867;
  wire n5868;
  wire n5869;
  wire n587;
  wire n5870;
  wire n5871;
  wire n5872;
  wire n5873;
  wire n5874;
  wire n5875;
  wire n5876;
  wire n5877;
  wire n5878;
  wire n5879;
  wire n588;
  wire n5880;
  wire n5881;
  wire n5882;
  wire n5883;
  wire n5884;
  wire n5885;
  wire n5886;
  wire n5887;
  wire n5888;
  wire n5889;
  wire n589;
  wire n5890;
  wire n5891;
  wire n5892;
  wire n5893;
  wire n5894;
  wire n5895;
  wire n5896;
  wire n5897;
  wire n5898;
  wire n5899;
  wire n59;
  wire n590;
  wire n5900;
  wire n5901;
  wire n5902;
  wire n5903;
  wire n5904;
  wire n5905;
  wire n5906;
  wire n5907;
  wire n5908;
  wire n5909;
  wire n591;
  wire n5910;
  wire n5911;
  wire n5912;
  wire n5913;
  wire n5914;
  wire n5915;
  wire n5916;
  wire n5917;
  wire n5918;
  wire n5919;
  wire n592;
  wire n5920;
  wire n5921;
  wire n5922;
  wire n5923;
  wire n5924;
  wire n5925;
  wire n5926;
  wire n5927;
  wire n5928;
  wire n5929;
  wire n593;
  wire n5930;
  wire n5931;
  wire n5932;
  wire n5933;
  wire n5934;
  wire n5935;
  wire n5936;
  wire n5937;
  wire n5938;
  wire n5939;
  wire n594;
  wire n5940;
  wire n5941;
  wire n5942;
  wire n5943;
  wire n5944;
  wire n5945;
  wire n5946;
  wire n5947;
  wire n5948;
  wire n5949;
  wire n595;
  wire n5950;
  wire n5951;
  wire n5952;
  wire n5953;
  wire n5954;
  wire n5955;
  wire n5956;
  wire n5957;
  wire n5958;
  wire n5959;
  wire n596;
  wire n5960;
  wire n5961;
  wire n5962;
  wire n5963;
  wire n5964;
  wire n5965;
  wire n5966;
  wire n5967;
  wire n5969;
  wire n597;
  wire n5970;
  wire n5971;
  wire n5972;
  wire n5973;
  wire n5974;
  wire n5975;
  wire n5976;
  wire n5977;
  wire n5978;
  wire n5979;
  wire n598;
  wire n5980;
  wire n5981;
  wire n5982;
  wire n5983;
  wire n5984;
  wire n5985;
  wire n5986;
  wire n5987;
  wire n5988;
  wire n5989;
  wire n599;
  wire n5990;
  wire n5991;
  wire n5992;
  wire n5993;
  wire n5994;
  wire n5995;
  wire n5996;
  wire n5997;
  wire n5998;
  wire n5999;
  wire n6;
  wire n60;
  wire n600;
  wire n6000;
  wire n6001;
  wire n6002;
  wire n6003;
  wire n6004;
  wire n6005;
  wire n6006;
  wire n6007;
  wire n6008;
  wire n6009;
  wire n601;
  wire n6010;
  wire n6011;
  wire n6012;
  wire n6013;
  wire n6014;
  wire n6015;
  wire n6016;
  wire n6017;
  wire n6018;
  wire n6019;
  wire n602;
  wire n6020;
  wire n6021;
  wire n6022;
  wire n6023;
  wire n6024;
  wire n6025;
  wire n6026;
  wire n603;
  wire n604;
  wire n605;
  wire n606;
  wire n607;
  wire n608;
  wire n609;
  wire n61;
  wire n610;
  wire n611;
  wire n612;
  wire n613;
  wire n614;
  wire n615;
  wire n616;
  wire n617;
  wire n618;
  wire n619;
  wire n62;
  wire n620;
  wire n621;
  wire n622;
  wire n623;
  wire n624;
  wire n625;
  wire n626;
  wire n627;
  wire n628;
  wire n629;
  wire n63;
  wire n630;
  wire n631;
  wire n632;
  wire n633;
  wire n634;
  wire n635;
  wire n636;
  wire n637;
  wire n638;
  wire n639;
  wire n64;
  wire n640;
  wire n641;
  wire n642;
  wire n643;
  wire n644;
  wire n645;
  wire n646;
  wire n647;
  wire n648;
  wire n649;
  wire n65;
  wire n650;
  wire n651;
  wire n652;
  wire n653;
  wire n654;
  wire n655;
  wire n656;
  wire n657;
  wire n658;
  wire n659;
  wire n66;
  wire n660;
  wire n661;
  wire n662;
  wire n663;
  wire n664;
  wire n665;
  wire n666;
  wire n667;
  wire n668;
  wire n669;
  wire n67;
  wire n670;
  wire n671;
  wire n672;
  wire n673;
  wire n674;
  wire n675;
  wire n676;
  wire n677;
  wire n678;
  wire n679;
  wire n68;
  wire n680;
  wire n681;
  wire n682;
  wire n683;
  wire n684;
  wire n685;
  wire n686;
  wire n687;
  wire n688;
  wire n689;
  wire n69;
  wire n690;
  wire n691;
  wire n692;
  wire n693;
  wire n694;
  wire n695;
  wire n696;
  wire n697;
  wire n698;
  wire n699;
  wire n70;
  wire n700;
  wire n701;
  wire n702;
  wire n703;
  wire n704;
  wire n705;
  wire n706;
  wire n707;
  wire n708;
  wire n709;
  wire n71;
  wire n710;
  wire n711;
  wire n712;
  wire n713;
  wire n714;
  wire n715;
  wire n716;
  wire n717;
  wire n718;
  wire n719;
  wire n72;
  wire n720;
  wire n721;
  wire n722;
  wire n723;
  wire n724;
  wire n725;
  wire n726;
  wire n727;
  wire n728;
  wire n729;
  wire n73;
  wire n730;
  wire n731;
  wire n732;
  wire n733;
  wire n734;
  wire n735;
  wire n736;
  wire n737;
  wire n738;
  wire n739;
  wire n74;
  wire n740;
  wire n741;
  wire n742;
  wire n743;
  wire n744;
  wire n745;
  wire n746;
  wire n747;
  wire n748;
  wire n749;
  wire n75;
  wire n750;
  wire n751;
  wire n752;
  wire n753;
  wire n754;
  wire n755;
  wire n756;
  wire n757;
  wire n758;
  wire n759;
  wire n76;
  wire n760;
  wire n761;
  wire n762;
  wire n763;
  wire n764;
  wire n765;
  wire n766;
  wire n767;
  wire n768;
  wire n769;
  wire n77;
  wire n770;
  wire n771;
  wire n772;
  wire n773;
  wire n774;
  wire n775;
  wire n776;
  wire n777;
  wire n778;
  wire n779;
  wire n78;
  wire n780;
  wire n781;
  wire n782;
  wire n783;
  wire n784;
  wire n785;
  wire n786;
  wire n787;
  wire n788;
  wire n789;
  wire n79;
  wire n790;
  wire n791;
  wire n792;
  wire n793;
  wire n794;
  wire n795;
  wire n796;
  wire n797;
  wire n798;
  wire n799;
  wire n8;
  wire n80;
  wire n800;
  wire n801;
  wire n802;
  wire n803;
  wire n804;
  wire n805;
  wire n806;
  wire n807;
  wire n808;
  wire n809;
  wire n81;
  wire n810;
  wire n811;
  wire n812;
  wire n813;
  wire n814;
  wire n815;
  wire n816;
  wire n817;
  wire n818;
  wire n819;
  wire n82;
  wire n820;
  wire n821;
  wire n822;
  wire n823;
  wire n824;
  wire n825;
  wire n826;
  wire n827;
  wire n828;
  wire n829;
  wire n83;
  wire n830;
  wire n831;
  wire n832;
  wire n833;
  wire n834;
  wire n835;
  wire n836;
  wire n837;
  wire n838;
  wire n839;
  wire n84;
  wire n840;
  wire n841;
  wire n842;
  wire n843;
  wire n844;
  wire n845;
  wire n846;
  wire n847;
  wire n848;
  wire n849;
  wire n85;
  wire n850;
  wire n851;
  wire n852;
  wire n853;
  wire n854;
  wire n855;
  wire n856;
  wire n857;
  wire n858;
  wire n859;
  wire n86;
  wire n860;
  wire n861;
  wire n862;
  wire n863;
  wire n864;
  wire n865;
  wire n866;
  wire n867;
  wire n868;
  wire n869;
  wire n87;
  wire n870;
  wire n871;
  wire n872;
  wire n873;
  wire n874;
  wire n875;
  wire n876;
  wire n877;
  wire n878;
  wire n879;
  wire n88;
  wire n880;
  wire n881;
  wire n882;
  wire n883;
  wire n884;
  wire n885;
  wire n886;
  wire n887;
  wire n888;
  wire n889;
  wire n89;
  wire n890;
  wire n891;
  wire n892;
  wire n893;
  wire n894;
  wire n895;
  wire n896;
  wire n897;
  wire n898;
  wire n899;
  wire n9;
  wire n90;
  wire n900;
  wire n901;
  wire n902;
  wire n903;
  wire n904;
  wire n905;
  wire n906;
  wire n907;
  wire n908;
  wire n909;
  wire n91;
  wire n910;
  wire n911;
  wire n912;
  wire n913;
  wire n914;
  wire n915;
  wire n916;
  wire n917;
  wire n918;
  wire n919;
  wire n92;
  wire n920;
  wire n921;
  wire n922;
  wire n923;
  wire n924;
  wire n925;
  wire n926;
  wire n927;
  wire n928;
  wire n929;
  wire n93;
  wire n930;
  wire n931;
  wire n932;
  wire n933;
  wire n934;
  wire n935;
  wire n936;
  wire n937;
  wire n938;
  wire n939;
  wire n94;
  wire n940;
  wire n941;
  wire n942;
  wire n943;
  wire n944;
  wire n945;
  wire n946;
  wire n947;
  wire n948;
  wire n949;
  wire n95;
  wire n950;
  wire n951;
  wire n952;
  wire n953;
  wire n954;
  wire n955;
  wire n956;
  wire n957;
  wire n958;
  wire n959;
  wire n96;
  wire n960;
  wire n961;
  wire n962;
  wire n963;
  wire n964;
  wire n965;
  wire n966;
  wire n967;
  wire n968;
  wire n969;
  wire n97;
  wire n970;
  wire n971;
  wire n972;
  wire n973;
  wire n974;
  wire n975;
  wire n976;
  wire n977;
  wire n978;
  wire n979;
  wire n98;
  wire n980;
  wire n981;
  wire n982;
  wire n983;
  wire n984;
  wire n985;
  wire n986;
  wire n987;
  wire n988;
  wire n989;
  wire n99;
  wire n990;
  wire n991;
  wire n992;
  wire n993;
  wire n994;
  wire n995;
  wire n996;
  wire n997;
  wire n998;
  wire n999;

  AL_DFF A1qax6_reg (
    .clk(HCLK),
    .d(Mdthu6),
    .reset(1'b0),
    .set(1'b0),
    .q(A1qax6));  // ../RTL/cortexm0ds_logic.v(18823)
  AL_DFF A2spw6_reg (
    .clk(HCLK),
    .d(Cgshu6),
    .reset(1'b0),
    .set(1'b0),
    .q(A2spw6));  // ../RTL/cortexm0ds_logic.v(17639)
  AL_DFF A32qw6_reg (
    .clk(HCLK),
    .d(Fpohu6),
    .reset(1'b0),
    .set(n5973),
    .q(A32qw6));  // ../RTL/cortexm0ds_logic.v(17961)
  AL_DFF A3ipw6_reg (
    .clk(DCLK),
    .d(X3yhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(A3ipw6));  // ../RTL/cortexm0ds_logic.v(17180)
  AL_DFF A3qax6_reg (
    .clk(HCLK),
    .d(Fdthu6),
    .reset(1'b0),
    .set(1'b0),
    .q(A3qax6));  // ../RTL/cortexm0ds_logic.v(18824)
  AL_DFF A5ipw6_reg (
    .clk(SWCLKTCK),
    .d(Nrxhu6),
    .reset(n5972),
    .set(1'b0),
    .q(A5ipw6));  // ../RTL/cortexm0ds_logic.v(17185)
  AL_DFF A5qax6_reg (
    .clk(HCLK),
    .d(Ycthu6),
    .reset(1'b0),
    .set(1'b0),
    .q(A5qax6));  // ../RTL/cortexm0ds_logic.v(18825)
  AL_DFF A6cbx6_reg (
    .clk(SWCLKTCK),
    .d(Qixhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(A6cbx6));  // ../RTL/cortexm0ds_logic.v(19945)
  AL_DFF A7zpw6_reg (
    .clk(HCLK),
    .d(Afshu6),
    .reset(1'b0),
    .set(1'b0),
    .q(A7zpw6));  // ../RTL/cortexm0ds_logic.v(17899)
  AL_DFF Aa2bx6_reg (
    .clk(SCLK),
    .d(C5phu6),
    .reset(n5973),
    .set(1'b0),
    .q(Aa2bx6));  // ../RTL/cortexm0ds_logic.v(19401)
  AL_DFF Ab9ax6_reg (
    .clk(DCLK),
    .d(Wnvhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Ab9ax6));  // ../RTL/cortexm0ds_logic.v(18163)
  AL_DFF Acebx6_reg (
    .clk(DCLK),
    .d(Hpwhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Acebx6));  // ../RTL/cortexm0ds_logic.v(19991)
  AL_DFF Acuax6_reg (
    .clk(HCLK),
    .d(Drshu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Acuax6));  // ../RTL/cortexm0ds_logic.v(18901)
  AL_DFF Ad7ax6_reg (
    .clk(DCLK),
    .d(Gdxhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Ad7ax6));  // ../RTL/cortexm0ds_logic.v(18091)
  AL_DFF Ahdax6_reg (
    .clk(DCLK),
    .d(Zrwhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Ahdax6));  // ../RTL/cortexm0ds_logic.v(18289)
  AL_DFF Ahdbx6_reg (
    .clk(SWCLKTCK),
    .d(Gkxhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Ahdbx6));  // ../RTL/cortexm0ds_logic.v(19975)
  AL_DFF Ahlpw6_reg (
    .clk(SWCLKTCK),
    .d(Zehpw6[6]),
    .reset(1'b0),
    .set(n5972),
    .q(Ahlpw6));  // ../RTL/cortexm0ds_logic.v(17362)
  AL_DFF Amupw6_reg (
    .clk(SCLK),
    .d(Iauhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Amupw6));  // ../RTL/cortexm0ds_logic.v(17710)
  AL_DFF Aniax6_reg (
    .clk(HCLK),
    .d(G1vhu6),
    .reset(n5973),
    .set(1'b0),
    .q(Aniax6));  // ../RTL/cortexm0ds_logic.v(18613)
  AL_DFF Aoeax6_reg (
    .clk(DCLK),
    .d(Wfwhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Aoeax6));  // ../RTL/cortexm0ds_logic.v(18317)
  AL_DFF Apcax6_reg (
    .clk(DCLK),
    .d(Lywhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Apcax6));  // ../RTL/cortexm0ds_logic.v(18269)
  AL_DFF Aqlax6_reg (
    .clk(HCLK),
    .d(Tlshu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Aqlax6));  // ../RTL/cortexm0ds_logic.v(18745)
  AL_DFF Ar1bx6_reg (
    .clk(SCLK),
    .d(Vruhu6),
    .reset(n5973),
    .set(1'b0),
    .q(Ar1bx6));  // ../RTL/cortexm0ds_logic.v(19347)
  AL_DFF Arnpw6_reg (
    .clk(HCLK),
    .d(Kgphu6),
    .reset(1'b0),
    .set(n5973),
    .q(Arnpw6));  // ../RTL/cortexm0ds_logic.v(17475)
  AL_DFF Asupw6_reg (
    .clk(HCLK),
    .d(Hfshu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Asupw6));  // ../RTL/cortexm0ds_logic.v(17718)
  AL_DFF At2bx6_reg (
    .clk(SCLK),
    .d(Ipthu6),
    .reset(n5973),
    .set(1'b0),
    .q(At2bx6));  // ../RTL/cortexm0ds_logic.v(19455)
  AL_DFF Aujpw6_reg (
    .clk(HCLK),
    .d(Axohu6),
    .reset(n5973),
    .set(1'b0),
    .q(Aujpw6));  // ../RTL/cortexm0ds_logic.v(17271)
  AL_DFF Aurpw6_reg (
    .clk(HCLK),
    .d(Kdshu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Aurpw6));  // ../RTL/cortexm0ds_logic.v(17630)
  AL_DFF Auyax6_reg (
    .clk(HCLK),
    .d(Euthu6),
    .reset(n5973),
    .set(1'b0),
    .q(Auyax6));  // ../RTL/cortexm0ds_logic.v(19041)
  AL_DFF Avzax6_reg (
    .clk(HCLK),
    .d(Qluhu6),
    .reset(n5973),
    .set(1'b0),
    .q(Avzax6));  // ../RTL/cortexm0ds_logic.v(19149)
  AL_DFF Aw4bx6_reg (
    .clk(HCLK),
    .d(V6uhu6),
    .reset(n5973),
    .set(1'b0),
    .q(Aw4bx6));  // ../RTL/cortexm0ds_logic.v(19671)
  AL_DFF Awupw6_reg (
    .clk(HCLK),
    .d(Xrohu6),
    .reset(1'b0),
    .set(n5973),
    .q(Awupw6));  // ../RTL/cortexm0ds_logic.v(17729)
  AL_DFF Az3bx6_reg (
    .clk(HCLK),
    .d(M5uhu6),
    .reset(n5973),
    .set(1'b0),
    .q(Az3bx6));  // ../RTL/cortexm0ds_logic.v(19575)
  AL_DFF Azpax6_reg (
    .clk(HCLK),
    .d(Tdthu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Azpax6));  // ../RTL/cortexm0ds_logic.v(18822)
  AL_DFF B0spw6_reg (
    .clk(HCLK),
    .d(Vfshu6),
    .reset(1'b0),
    .set(1'b0),
    .q(B0spw6));  // ../RTL/cortexm0ds_logic.v(17638)
  AL_DFF B3gbx6_reg (
    .clk(HCLK),
    .d(Bvuhu6),
    .reset(n5973),
    .set(1'b0),
    .q(B3gbx6));  // ../RTL/cortexm0ds_logic.v(20037)
  AL_DFF B4uax6_reg (
    .clk(HCLK),
    .d(Nathu6),
    .reset(1'b0),
    .set(1'b0),
    .q(B4uax6));  // ../RTL/cortexm0ds_logic.v(18897)
  AL_DFF B5zpw6_reg (
    .clk(HCLK),
    .d(Pjshu6),
    .reset(1'b0),
    .set(1'b0),
    .q(B5zpw6));  // ../RTL/cortexm0ds_logic.v(17898)
  AL_DFF B6uax6_reg (
    .clk(HCLK),
    .d(Gathu6),
    .reset(1'b0),
    .set(1'b0),
    .q(B6uax6));  // ../RTL/cortexm0ds_logic.v(18898)
  AL_DFF B79bx6_reg (
    .clk(DCLK),
    .d(Iexhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(B79bx6));  // ../RTL/cortexm0ds_logic.v(19810)
  AL_DFF B7lpw6_reg (
    .clk(SWCLKTCK),
    .d(Fwohu6),
    .reset(n5972),
    .set(1'b0),
    .q(B7lpw6));  // ../RTL/cortexm0ds_logic.v(17331)
  AL_DFF B8uax6_reg (
    .clk(HCLK),
    .d(Z9thu6),
    .reset(1'b0),
    .set(1'b0),
    .q(B8uax6));  // ../RTL/cortexm0ds_logic.v(18899)
  AL_DFF B9eax6_reg (
    .clk(DCLK),
    .d(Lkwhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(B9eax6));  // ../RTL/cortexm0ds_logic.v(18304)
  AL_DFF B9jbx6_reg (
    .clk(DCLK),
    .d(Zdwhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(B9jbx6));  // ../RTL/cortexm0ds_logic.v(20186)
  AL_DFF Bauax6_reg (
    .clk(HCLK),
    .d(S9thu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Bauax6));  // ../RTL/cortexm0ds_logic.v(18900)
  AL_DFF Bbjpw6_reg (
    .clk(HCLK),
    .d(Z5qhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Bbjpw6));  // ../RTL/cortexm0ds_logic.v(17232)
  AL_DFF Bc3bx6_reg (
    .clk(SCLK),
    .d(Qyohu6),
    .reset(n5973),
    .set(1'b0),
    .q(Bc3bx6));  // ../RTL/cortexm0ds_logic.v(19509)
  AL_DFF Bcabx6_reg (
    .clk(HCLK),
    .d(Nvthu6),
    .reset(n5973),
    .set(1'b0),
    .q(Bcabx6));  // ../RTL/cortexm0ds_logic.v(19885)
  AL_DFF Bccax6_reg (
    .clk(DCLK),
    .d(J5whu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Bccax6));  // ../RTL/cortexm0ds_logic.v(18257)
  AL_DFF Bcdbx6_reg (
    .clk(SWCLKTCK),
    .d(Pzxhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Bcdbx6));  // ../RTL/cortexm0ds_logic.v(19972)
  AL_DFF Bcgax6_reg (
    .clk(DCLK),
    .d(Uzwhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Bcgax6));  // ../RTL/cortexm0ds_logic.v(18404)
  AL_DFF Bciax6_reg (
    .clk(SCLK),
    .d(P2vhu6),
    .reset(n5973),
    .set(1'b0),
    .q(Bciax6));  // ../RTL/cortexm0ds_logic.v(18577)
  AL_DFF Bclpw6_reg (
    .clk(SWCLKTCK),
    .d(Zehpw6[0]),
    .reset(n5972),
    .set(1'b0),
    .q(Bclpw6));  // ../RTL/cortexm0ds_logic.v(17344)
  AL_DFF Bdjpw6_reg (
    .clk(HCLK),
    .d(D8qhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Bdjpw6));  // ../RTL/cortexm0ds_logic.v(17233)
  AL_DFF Bf3qw6_reg (
    .clk(DCLK),
    .d(P7xhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Bf3qw6));  // ../RTL/cortexm0ds_logic.v(18033)
  AL_DFF Bfjpw6_reg (
    .clk(HCLK),
    .d(Ksrhu6),
    .reset(1'b0),
    .set(n5973),
    .q(Bfjpw6));  // ../RTL/cortexm0ds_logic.v(17238)
  AL_DFF Biaax6_reg (
    .clk(DCLK),
    .d(Twvhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Biaax6));  // ../RTL/cortexm0ds_logic.v(18186)
  AL_DFF Bk7ax6_reg (
    .clk(SWCLKTCK),
    .d(Cpxhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Bk7ax6));  // ../RTL/cortexm0ds_logic.v(18100)
  AL_DFF Bngax6_reg (
    .clk(DCLK),
    .d(Erwhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Bngax6));  // ../RTL/cortexm0ds_logic.v(18410)
  AL_DFF Bolax6_reg (
    .clk(HCLK),
    .d(Pqshu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Bolax6));  // ../RTL/cortexm0ds_logic.v(18744)
  AL_DFF Bp2qw6_reg (
    .clk(SWCLKTCK),
    .d(Xixhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Bp2qw6));  // ../RTL/cortexm0ds_logic.v(17999)
  AL_DFF Bq9ax6_reg (
    .clk(DCLK),
    .d(Qkvhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Bq9ax6));  // ../RTL/cortexm0ds_logic.v(18171)
  AL_DFF Bsrpw6_reg (
    .clk(HCLK),
    .d(Wcshu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Bsrpw6));  // ../RTL/cortexm0ds_logic.v(17629)
  AL_DFF Bt2qw6_reg (
    .clk(DCLK),
    .d(I0xhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Bt2qw6));  // ../RTL/cortexm0ds_logic.v(18006)
  AL_DFF Btbbx6_reg (
    .clk(DCLK),
    .d(Hwwhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Btbbx6));  // ../RTL/cortexm0ds_logic.v(19938)
  AL_DFF Bu6bx6_reg (
    .clk(DCLK),
    .d(Vbphu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Bu6bx6));  // ../RTL/cortexm0ds_logic.v(19762)
  AL_DFF Buabx6_reg (
    .clk(DCLK),
    .d(Mvwhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Buabx6));  // ../RTL/cortexm0ds_logic.v(19895)
  AL_DFF Bvaax6_reg (
    .clk(DCLK),
    .d(Buvhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Bvaax6));  // ../RTL/cortexm0ds_logic.v(18193)
  AL_DFF Bvfbx6_reg (
    .clk(DCLK),
    .d(Jbxhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Bvfbx6));  // ../RTL/cortexm0ds_logic.v(20019)
  AL_DFF Bwdax6_reg (
    .clk(DCLK),
    .d(Dnwhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Bwdax6));  // ../RTL/cortexm0ds_logic.v(18297)
  AL_DFF Bx2qw6_reg (
    .clk(SWCLKTCK),
    .d(Bsxhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Bx2qw6));  // ../RTL/cortexm0ds_logic.v(18008)
  AL_DFF Bxbax6_reg (
    .clk(DCLK),
    .d(P8whu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Bxbax6));  // ../RTL/cortexm0ds_logic.v(18249)
  AL_DFF Bxpax6_reg (
    .clk(HCLK),
    .d(Aethu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Bxpax6));  // ../RTL/cortexm0ds_logic.v(18821)
  AL_DFF C07bx6_reg (
    .clk(HCLK),
    .d(V3qhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(C07bx6));  // ../RTL/cortexm0ds_logic.v(19765)
  AL_DFF C10bx6_reg (
    .clk(HCLK),
    .d(Pouhu6),
    .reset(n5973),
    .set(1'b0),
    .q(C10bx6));  // ../RTL/cortexm0ds_logic.v(19167)
  AL_DFF C14bx6_reg (
    .clk(HCLK),
    .d(Y4uhu6),
    .reset(n5973),
    .set(1'b0),
    .q(C14bx6));  // ../RTL/cortexm0ds_logic.v(19581)
  AL_DFF C1fax6_reg (
    .clk(DCLK),
    .d(Xcwhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(C1fax6));  // ../RTL/cortexm0ds_logic.v(18324)
  AL_DFF C1wpw6_reg (
    .clk(HCLK),
    .d(Hyuhu6),
    .reset(n5973),
    .set(1'b0),
    .q(C1wpw6));  // ../RTL/cortexm0ds_logic.v(17800)
  AL_DFF C27bx6_reg (
    .clk(HCLK),
    .d(Nzphu6),
    .reset(1'b0),
    .set(1'b0),
    .q(C27bx6));  // ../RTL/cortexm0ds_logic.v(19766)
  AL_DFF C2uax6_reg (
    .clk(HCLK),
    .d(Uathu6),
    .reset(1'b0),
    .set(1'b0),
    .q(C2uax6));  // ../RTL/cortexm0ds_logic.v(18896)
  AL_DFF C2ypw6_reg (
    .clk(SWCLKTCK),
    .d(Ymxhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(C2ypw6));  // ../RTL/cortexm0ds_logic.v(17858)
  AL_DFF C30bx6_reg (
    .clk(HCLK),
    .d(Wouhu6),
    .reset(n5973),
    .set(1'b0),
    .q(C30bx6));  // ../RTL/cortexm0ds_logic.v(19173)
  AL_DFF C37ax6_reg (
    .clk(HCLK),
    .d(Roohu6),
    .reset(1'b0),
    .set(n5973),
    .q(C37ax6));  // ../RTL/cortexm0ds_logic.v(18085)
  AL_DFF C3wpw6_reg (
    .clk(HCLK),
    .d(Tbvhu6),
    .reset(n5973),
    .set(1'b0),
    .q(C3wpw6));  // ../RTL/cortexm0ds_logic.v(17806)
  AL_DFF C3zpw6_reg (
    .clk(HCLK),
    .d(Eoshu6),
    .reset(1'b0),
    .set(1'b0),
    .q(C3zpw6));  // ../RTL/cortexm0ds_logic.v(17897)
  AL_DFF C47bx6_reg (
    .clk(HCLK),
    .d(Uzphu6),
    .reset(1'b0),
    .set(1'b0),
    .q(C47bx6));  // ../RTL/cortexm0ds_logic.v(19767)
  AL_DFF C4dax6_reg (
    .clk(DCLK),
    .d(Kuwhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(C4dax6));  // ../RTL/cortexm0ds_logic.v(18277)
  AL_DFF C50bx6_reg (
    .clk(HCLK),
    .d(Kpuhu6),
    .reset(n5973),
    .set(1'b0),
    .q(C50bx6));  // ../RTL/cortexm0ds_logic.v(19179)
  AL_DFF C5gbx6_reg (
    .clk(HCLK),
    .d(Nuuhu6),
    .reset(n5973),
    .set(1'b0),
    .q(C5gbx6));  // ../RTL/cortexm0ds_logic.v(20043)
  AL_DFF C5wpw6_reg (
    .clk(HCLK),
    .d(Kmqhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(C5wpw6));  // ../RTL/cortexm0ds_logic.v(17808)
  AL_DFF C67bx6_reg (
    .clk(HCLK),
    .d(B0qhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(C67bx6));  // ../RTL/cortexm0ds_logic.v(19768)
  AL_DFF C72qw6_reg (
    .clk(SWCLKTCK),
    .d(T1yhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(C72qw6));  // ../RTL/cortexm0ds_logic.v(17964)
  AL_DFF C7wpw6_reg (
    .clk(HCLK),
    .d(Rmqhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(C7wpw6));  // ../RTL/cortexm0ds_logic.v(17809)
  AL_DFF C87bx6_reg (
    .clk(HCLK),
    .d(I0qhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(C87bx6));  // ../RTL/cortexm0ds_logic.v(19769)
  AL_DFF C9wpw6_reg (
    .clk(HCLK),
    .d(Tnqhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(C9wpw6));  // ../RTL/cortexm0ds_logic.v(17810)
  AL_DFF Ca1bx6_reg (
    .clk(SCLK),
    .d(Snthu6),
    .reset(n5973),
    .set(1'b0),
    .q(Ca1bx6));  // ../RTL/cortexm0ds_logic.v(19299)
  AL_DFF Ca7bx6_reg (
    .clk(HCLK),
    .d(P0qhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Ca7bx6));  // ../RTL/cortexm0ds_logic.v(19770)
  AL_DFF Cbwpw6_reg (
    .clk(HCLK),
    .d(Hoqhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Cbwpw6));  // ../RTL/cortexm0ds_logic.v(17811)
  AL_DFF Cc2bx6_reg (
    .clk(SCLK),
    .d(Ltuhu6),
    .reset(n5973),
    .set(1'b0),
    .q(Cc2bx6));  // ../RTL/cortexm0ds_logic.v(19407)
  AL_DFF Cc7bx6_reg (
    .clk(HCLK),
    .d(W0qhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Cc7bx6));  // ../RTL/cortexm0ds_logic.v(19771)
  AL_DFF Cccbx6_reg (
    .clk(DCLK),
    .d(N0whu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Cccbx6));  // ../RTL/cortexm0ds_logic.v(19948)
  AL_DFF Cchax6_reg (
    .clk(HCLK),
    .d(Umohu6),
    .reset(1'b0),
    .set(n5973),
    .q(Cchax6));  // ../RTL/cortexm0ds_logic.v(18483)
  AL_DFF Cdwpw6_reg (
    .clk(HCLK),
    .d(Voqhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Cdwpw6));  // ../RTL/cortexm0ds_logic.v(17812)
  AL_DFF Ce7bx6_reg (
    .clk(HCLK),
    .d(D1qhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Ce7bx6));  // ../RTL/cortexm0ds_logic.v(19772)
  AL_DFF Ceabx6_reg (
    .clk(DCLK),
    .d(Ldphu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Ceabx6));  // ../RTL/cortexm0ds_logic.v(19887)
  AL_DFF Cfvpw6_reg (
    .clk(SWCLKTCK),
    .d(Nkxhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Cfvpw6));  // ../RTL/cortexm0ds_logic.v(17775)
  AL_DFF Cfwpw6_reg (
    .clk(HCLK),
    .d(Lqqhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Cfwpw6));  // ../RTL/cortexm0ds_logic.v(17813)
  AL_DFF Cg7bx6_reg (
    .clk(HCLK),
    .d(K1qhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Cg7bx6));  // ../RTL/cortexm0ds_logic.v(19773)
  AL_DFF Cglax6_reg (
    .clk(HCLK),
    .d(Nwshu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Cglax6));  // ../RTL/cortexm0ds_logic.v(18740)
  AL_DFF Chwpw6_reg (
    .clk(HCLK),
    .d(Sqqhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Chwpw6));  // ../RTL/cortexm0ds_logic.v(17814)
  AL_DFF Ci7bx6_reg (
    .clk(HCLK),
    .d(R1qhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Ci7bx6));  // ../RTL/cortexm0ds_logic.v(19774)
  AL_DFF Cilax6_reg (
    .clk(HCLK),
    .d(Gwshu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Cilax6));  // ../RTL/cortexm0ds_logic.v(18741)
  AL_DFF Cjqpw6_reg (
    .clk(SWCLKTCK),
    .d(Yfxhu6),
    .reset(n5972),
    .set(1'b0),
    .q(Cjqpw6));  // ../RTL/cortexm0ds_logic.v(17566)
  AL_DFF Cjwpw6_reg (
    .clk(DCLK),
    .d(Maphu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Cjwpw6));  // ../RTL/cortexm0ds_logic.v(17815)
  AL_DFF Ck7bx6_reg (
    .clk(HCLK),
    .d(Y1qhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Ck7bx6));  // ../RTL/cortexm0ds_logic.v(19775)
  AL_DFF Cklax6_reg (
    .clk(HCLK),
    .d(Zvshu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Cklax6));  // ../RTL/cortexm0ds_logic.v(18742)
  AL_DFF Cm7bx6_reg (
    .clk(HCLK),
    .d(F2qhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Cm7bx6));  // ../RTL/cortexm0ds_logic.v(19776)
  AL_DFF Cmlax6_reg (
    .clk(HCLK),
    .d(Svshu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Cmlax6));  // ../RTL/cortexm0ds_logic.v(18743)
  AL_DFF Cncbx6_reg (
    .clk(DCLK),
    .d(U7phu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Cncbx6));  // ../RTL/cortexm0ds_logic.v(19954)
  AL_DFF Cndbx6_reg (
    .clk(DCLK),
    .d(Xyvhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Cndbx6));  // ../RTL/cortexm0ds_logic.v(19978)
  AL_DFF Co7bx6_reg (
    .clk(HCLK),
    .d(M2qhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Co7bx6));  // ../RTL/cortexm0ds_logic.v(19777)
  AL_DFF Cokbx6_reg (
    .clk(SCLK),
    .d(Raohu6),
    .reset(n5973),
    .set(1'b0),
    .q(Cokbx6));  // ../RTL/cortexm0ds_logic.v(20266)
  AL_DFF Coupw6_reg (
    .clk(SCLK),
    .d(S8uhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Coupw6));  // ../RTL/cortexm0ds_logic.v(17711)
  AL_DFF Cq3qw6_reg (
    .clk(DCLK),
    .d(M9xhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Cq3qw6));  // ../RTL/cortexm0ds_logic.v(18045)
  AL_DFF Cq7bx6_reg (
    .clk(HCLK),
    .d(Vcohu6),
    .reset(1'b0),
    .set(n5973),
    .q(Cq7bx6));  // ../RTL/cortexm0ds_logic.v(19782)
  AL_DFF Cqrpw6_reg (
    .clk(HCLK),
    .d(Icshu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Cqrpw6));  // ../RTL/cortexm0ds_logic.v(17628)
  AL_DFF Cs6bx6_reg (
    .clk(HCLK),
    .d(Imphu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Cs6bx6));  // ../RTL/cortexm0ds_logic.v(19761)
  AL_DFF Cvpax6_reg (
    .clk(HCLK),
    .d(Hethu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Cvpax6));  // ../RTL/cortexm0ds_logic.v(18820)
  AL_DFF Cwyax6_reg (
    .clk(HCLK),
    .d(Xtthu6),
    .reset(n5973),
    .set(1'b0),
    .q(Cwyax6));  // ../RTL/cortexm0ds_logic.v(19047)
  AL_DFF Cxcbx6_reg (
    .clk(DCLK),
    .d(Tawhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Cxcbx6));  // ../RTL/cortexm0ds_logic.v(19964)
  AL_DFF Cxzax6_reg (
    .clk(HCLK),
    .d(Lmuhu6),
    .reset(n5973),
    .set(1'b0),
    .q(Cxzax6));  // ../RTL/cortexm0ds_logic.v(19155)
  AL_DFF Cy4bx6_reg (
    .clk(HCLK),
    .d(O6uhu6),
    .reset(n5973),
    .set(1'b0),
    .q(Cy4bx6));  // ../RTL/cortexm0ds_logic.v(19677)
  AL_DFF Cydbx6_reg (
    .clk(DCLK),
    .d(K9phu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Cydbx6));  // ../RTL/cortexm0ds_logic.v(19984)
  AL_DFF Czzax6_reg (
    .clk(HCLK),
    .d(Nnuhu6),
    .reset(n5973),
    .set(1'b0),
    .q(Czzax6));  // ../RTL/cortexm0ds_logic.v(19161)
  AL_DFF D0uax6_reg (
    .clk(HCLK),
    .d(Bbthu6),
    .reset(1'b0),
    .set(1'b0),
    .q(D0uax6));  // ../RTL/cortexm0ds_logic.v(18895)
  AL_DFF D12qw6_reg (
    .clk(HCLK),
    .d(Mpohu6),
    .reset(1'b0),
    .set(n5973),
    .q(D12qw6));  // ../RTL/cortexm0ds_logic.v(17955)
  AL_DFF D1aax6_reg (
    .clk(DCLK),
    .d(D2whu6),
    .reset(1'b0),
    .set(1'b0),
    .q(D1aax6));  // ../RTL/cortexm0ds_logic.v(18177)
  AL_DFF D1zpw6_reg (
    .clk(HCLK),
    .d(Atshu6),
    .reset(1'b0),
    .set(1'b0),
    .q(D1zpw6));  // ../RTL/cortexm0ds_logic.v(17896)
  AL_DFF D2opw6_reg (
    .clk(SWCLKTCK),
    .d(Wsxhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(D2opw6));  // ../RTL/cortexm0ds_logic.v(17492)
  AL_DFF D2rpw6_reg (
    .clk(SWCLKTCK),
    .d(Cixhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(D2rpw6));  // ../RTL/cortexm0ds_logic.v(17596)
  AL_DFF D43qw6_reg (
    .clk(DCLK),
    .d(T2xhu6),
    .reset(n5974),
    .set(1'b0),
    .q(D43qw6));  // ../RTL/cortexm0ds_logic.v(18021)
  AL_DFF D46bx6_reg (
    .clk(HCLK),
    .d(Carhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(D46bx6));  // ../RTL/cortexm0ds_logic.v(19749)
  AL_DFF D66bx6_reg (
    .clk(HCLK),
    .d(N5rhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(D66bx6));  // ../RTL/cortexm0ds_logic.v(19750)
  AL_DFF D70bx6_reg (
    .clk(HCLK),
    .d(Rpuhu6),
    .reset(n5973),
    .set(1'b0),
    .q(D70bx6));  // ../RTL/cortexm0ds_logic.v(19185)
  AL_DFF D7gbx6_reg (
    .clk(HCLK),
    .d(Vkuhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(D7gbx6));  // ../RTL/cortexm0ds_logic.v(20045)
  AL_DFF D86bx6_reg (
    .clk(HCLK),
    .d(Y0rhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(D86bx6));  // ../RTL/cortexm0ds_logic.v(19751)
  AL_DFF D99ax6_reg (
    .clk(DCLK),
    .d(Fpvhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(D99ax6));  // ../RTL/cortexm0ds_logic.v(18162)
  AL_DFF Da6bx6_reg (
    .clk(HCLK),
    .d(Jwqhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Da6bx6));  // ../RTL/cortexm0ds_logic.v(19752)
  AL_DFF Daebx6_reg (
    .clk(DCLK),
    .d(Fhwhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Daebx6));  // ../RTL/cortexm0ds_logic.v(19990)
  AL_DFF Daiax6_reg (
    .clk(HCLK),
    .d(Ajohu6),
    .reset(n5973),
    .set(1'b0),
    .q(Daiax6));  // ../RTL/cortexm0ds_logic.v(18571)
  AL_DFF Dc6bx6_reg (
    .clk(HCLK),
    .d(Urqhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Dc6bx6));  // ../RTL/cortexm0ds_logic.v(19753)
  AL_DFF De6bx6_reg (
    .clk(HCLK),
    .d(Fnqhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(De6bx6));  // ../RTL/cortexm0ds_logic.v(19754)
  AL_DFF Delax6_reg (
    .clk(HCLK),
    .d(Uwshu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Delax6));  // ../RTL/cortexm0ds_logic.v(18739)
  AL_DFF Dfbax6_reg (
    .clk(DCLK),
    .d(R2whu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Dfbax6));  // ../RTL/cortexm0ds_logic.v(18224)
  AL_DFF Dg2qw6_reg (
    .clk(DCLK),
    .d(G6xhu6),
    .reset(n5974),
    .set(1'b0),
    .q(Dg2qw6));  // ../RTL/cortexm0ds_logic.v(17983)
  AL_DFF Dg6bx6_reg (
    .clk(HCLK),
    .d(Beqhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Dg6bx6));  // ../RTL/cortexm0ds_logic.v(19755)
  AL_DFF Di3qw6_reg (
    .clk(DCLK),
    .d(A3xhu6),
    .reset(n5974),
    .set(1'b0),
    .q(Di3qw6));  // ../RTL/cortexm0ds_logic.v(18039)
  AL_DFF Di6bx6_reg (
    .clk(HCLK),
    .d(M9qhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Di6bx6));  // ../RTL/cortexm0ds_logic.v(19756)
  AL_DFF Dk6bx6_reg (
    .clk(HCLK),
    .d(X4qhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Dk6bx6));  // ../RTL/cortexm0ds_logic.v(19757)
  AL_DFF Dk9bx6_reg (
    .clk(DCLK),
    .d(Glwhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Dk9bx6));  // ../RTL/cortexm0ds_logic.v(19817)
  AL_DFF Dm6bx6_reg (
    .clk(HCLK),
    .d(K8qhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Dm6bx6));  // ../RTL/cortexm0ds_logic.v(19758)
  AL_DFF Dmeax6_reg (
    .clk(DCLK),
    .d(Kgwhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Dmeax6));  // ../RTL/cortexm0ds_logic.v(18316)
  AL_DFF Dncax6_reg (
    .clk(DCLK),
    .d(Nzwhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Dncax6));  // ../RTL/cortexm0ds_logic.v(18268)
  AL_DFF Do6bx6_reg (
    .clk(HCLK),
    .d(Tvphu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Do6bx6));  // ../RTL/cortexm0ds_logic.v(19759)
  AL_DFF Dorpw6_reg (
    .clk(HCLK),
    .d(Nbshu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Dorpw6));  // ../RTL/cortexm0ds_logic.v(17627)
  AL_DFF Dpwpw6_reg (
    .clk(DCLK),
    .d(Zcxhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Dpwpw6));  // ../RTL/cortexm0ds_logic.v(17818)
  AL_DFF Dq6bx6_reg (
    .clk(HCLK),
    .d(Xqphu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Dq6bx6));  // ../RTL/cortexm0ds_logic.v(19760)
  AL_DFF Dqkbx6_reg (
    .clk(SWCLKTCK),
    .d(I5nhu6),
    .reset(n5972),
    .set(1'b0),
    .q(Dqkbx6));  // ../RTL/cortexm0ds_logic.v(20272)
  AL_DFF Drcbx6_reg (
    .clk(SWCLKTCK),
    .d(Jixhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Drcbx6));  // ../RTL/cortexm0ds_logic.v(19961)
  AL_DFF Drhax6_reg (
    .clk(HCLK),
    .d(Qkohu6),
    .reset(1'b0),
    .set(n5973),
    .q(Drhax6));  // ../RTL/cortexm0ds_logic.v(18531)
  AL_DFF Dt1bx6_reg (
    .clk(SCLK),
    .d(I1phu6),
    .reset(n5973),
    .set(1'b0),
    .q(Dt1bx6));  // ../RTL/cortexm0ds_logic.v(19353)
  AL_DFF Dtpax6_reg (
    .clk(HCLK),
    .d(Fophu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Dtpax6));  // ../RTL/cortexm0ds_logic.v(18819)
  AL_DFF Dugax6_reg (
    .clk(DCLK),
    .d(Wexhu6),
    .reset(n5974),
    .set(1'b0),
    .q(Dugax6));  // ../RTL/cortexm0ds_logic.v(18423)
  AL_DFF Dv2bx6_reg (
    .clk(SCLK),
    .d(Nwdpw6),
    .reset(n5973),
    .set(1'b0),
    .q(Dv2bx6));  // ../RTL/cortexm0ds_logic.v(19461)
  AL_DFF Dxvpw6_reg (
    .clk(HCLK),
    .d(Gfvhu6),
    .reset(1'b0),
    .set(n5973),
    .q(Dxvpw6));  // ../RTL/cortexm0ds_logic.v(17793)
  AL_DFF Dzvpw6_reg (
    .clk(HCLK),
    .d(Aqohu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Dzvpw6));  // ../RTL/cortexm0ds_logic.v(17795)
  AL_DFF E05bx6_reg (
    .clk(HCLK),
    .d(Ozthu6),
    .reset(n5973),
    .set(1'b0),
    .q(E05bx6));  // ../RTL/cortexm0ds_logic.v(19683)
  AL_DFF E1npw6_reg (
    .clk(HCLK),
    .d(Gxrhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(E1npw6));  // ../RTL/cortexm0ds_logic.v(17448)
  AL_DFF E34bx6_reg (
    .clk(HCLK),
    .d(R4uhu6),
    .reset(n5973),
    .set(1'b0),
    .q(E34bx6));  // ../RTL/cortexm0ds_logic.v(19587)
  AL_DFF E3npw6_reg (
    .clk(HCLK),
    .d(Ysrhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(E3npw6));  // ../RTL/cortexm0ds_logic.v(17449)
  AL_DFF E5npw6_reg (
    .clk(HCLK),
    .d(H9rhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(E5npw6));  // ../RTL/cortexm0ds_logic.v(17450)
  AL_DFF E5pax6_reg (
    .clk(HCLK),
    .d(Klrhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(E5pax6));  // ../RTL/cortexm0ds_logic.v(18807)
  AL_DFF E6iax6_reg (
    .clk(SCLK),
    .d(H5vhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(E6iax6));  // ../RTL/cortexm0ds_logic.v(18565)
  AL_DFF E7npw6_reg (
    .clk(HCLK),
    .d(S4rhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(E7npw6));  // ../RTL/cortexm0ds_logic.v(17451)
  AL_DFF E7pax6_reg (
    .clk(HCLK),
    .d(Zbrhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(E7pax6));  // ../RTL/cortexm0ds_logic.v(18808)
  AL_DFF E8iax6_reg (
    .clk(SCLK),
    .d(D3vhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(E8iax6));  // ../RTL/cortexm0ds_logic.v(18566)
  AL_DFF E90bx6_reg (
    .clk(HCLK),
    .d(Ypuhu6),
    .reset(n5973),
    .set(1'b0),
    .q(E90bx6));  // ../RTL/cortexm0ds_logic.v(19191)
  AL_DFF E97ax6_reg (
    .clk(SWCLKTCK),
    .d(Sxxhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(E97ax6));  // ../RTL/cortexm0ds_logic.v(18089)
  AL_DFF E9npw6_reg (
    .clk(HCLK),
    .d(R8qhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(E9npw6));  // ../RTL/cortexm0ds_logic.v(17452)
  AL_DFF E9pax6_reg (
    .clk(HCLK),
    .d(K7rhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(E9pax6));  // ../RTL/cortexm0ds_logic.v(18809)
  AL_DFF Eafax6_reg (
    .clk(DCLK),
    .d(K1xhu6),
    .reset(n5974),
    .set(1'b0),
    .q(Eafax6));  // ../RTL/cortexm0ds_logic.v(18343)
  AL_DFF Eagax6_reg (
    .clk(DCLK),
    .d(Srwhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Eagax6));  // ../RTL/cortexm0ds_logic.v(18403)
  AL_DFF Ebnpw6_reg (
    .clk(HCLK),
    .d(C4qhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Ebnpw6));  // ../RTL/cortexm0ds_logic.v(17453)
  AL_DFF Ebpax6_reg (
    .clk(HCLK),
    .d(V2rhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Ebpax6));  // ../RTL/cortexm0ds_logic.v(18810)
  AL_DFF Eclax6_reg (
    .clk(HCLK),
    .d(Bxshu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Eclax6));  // ../RTL/cortexm0ds_logic.v(18738)
  AL_DFF Ectax6_reg (
    .clk(HCLK),
    .d(Ylrhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Ectax6));  // ../RTL/cortexm0ds_logic.v(18883)
  AL_DFF Ednpw6_reg (
    .clk(HCLK),
    .d(Rgphu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Ednpw6));  // ../RTL/cortexm0ds_logic.v(17454)
  AL_DFF Edpax6_reg (
    .clk(HCLK),
    .d(Gyqhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Edpax6));  // ../RTL/cortexm0ds_logic.v(18811)
  AL_DFF Ee3bx6_reg (
    .clk(SCLK),
    .d(Q6vhu6),
    .reset(n5973),
    .set(1'b0),
    .q(Ee3bx6));  // ../RTL/cortexm0ds_logic.v(19515)
  AL_DFF Eetax6_reg (
    .clk(HCLK),
    .d(Ncrhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Eetax6));  // ../RTL/cortexm0ds_logic.v(18884)
  AL_DFF Efdax6_reg (
    .clk(DCLK),
    .d(Gswhu6),
    .reset(n5974),
    .set(1'b0),
    .q(Efdax6));  // ../RTL/cortexm0ds_logic.v(18287)
  AL_DFF Efnpw6_reg (
    .clk(HCLK),
    .d(Pxshu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Efnpw6));  // ../RTL/cortexm0ds_logic.v(17455)
  AL_DFF Efpax6_reg (
    .clk(HCLK),
    .d(Rtqhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Efpax6));  // ../RTL/cortexm0ds_logic.v(18812)
  AL_DFF Egaax6_reg (
    .clk(DCLK),
    .d(Axvhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Egaax6));  // ../RTL/cortexm0ds_logic.v(18185)
  AL_DFF Eghbx6_reg (
    .clk(SCLK),
    .d(Asthu6),
    .reset(n5973),
    .set(1'b0),
    .q(Eghbx6));  // ../RTL/cortexm0ds_logic.v(20112)
  AL_DFF Egtax6_reg (
    .clk(HCLK),
    .d(Y7rhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Egtax6));  // ../RTL/cortexm0ds_logic.v(18885)
  AL_DFF Ehnpw6_reg (
    .clk(HCLK),
    .d(Cdvhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Ehnpw6));  // ../RTL/cortexm0ds_logic.v(17456)
  AL_DFF Ehpax6_reg (
    .clk(HCLK),
    .d(Cpqhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Ehpax6));  // ../RTL/cortexm0ds_logic.v(18813)
  AL_DFF Ehqpw6_reg (
    .clk(SWCLKTCK),
    .d(Fgxhu6),
    .reset(n5972),
    .set(1'b0),
    .q(Ehqpw6));  // ../RTL/cortexm0ds_logic.v(17560)
  AL_DFF Eitax6_reg (
    .clk(HCLK),
    .d(J3rhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Eitax6));  // ../RTL/cortexm0ds_logic.v(18886)
  AL_DFF Ejnpw6_reg (
    .clk(HCLK),
    .d(Jdvhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Ejnpw6));  // ../RTL/cortexm0ds_logic.v(17457)
  AL_DFF Ejpax6_reg (
    .clk(HCLK),
    .d(Yfqhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Ejpax6));  // ../RTL/cortexm0ds_logic.v(18814)
  AL_DFF Ektax6_reg (
    .clk(HCLK),
    .d(Uyqhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Ektax6));  // ../RTL/cortexm0ds_logic.v(18887)
  AL_DFF Elgax6_reg (
    .clk(DCLK),
    .d(Cjwhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Elgax6));  // ../RTL/cortexm0ds_logic.v(18409)
  AL_DFF Eliax6_reg (
    .clk(HCLK),
    .d(W2vhu6),
    .reset(1'b0),
    .set(n5973),
    .q(Eliax6));  // ../RTL/cortexm0ds_logic.v(18607)
  AL_DFF Elnpw6_reg (
    .clk(HCLK),
    .d(Yjthu6),
    .reset(n5973),
    .set(1'b0),
    .q(Elnpw6));  // ../RTL/cortexm0ds_logic.v(17462)
  AL_DFF Elpax6_reg (
    .clk(HCLK),
    .d(Jbqhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Elpax6));  // ../RTL/cortexm0ds_logic.v(18815)
  AL_DFF Emrpw6_reg (
    .clk(HCLK),
    .d(Gbshu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Emrpw6));  // ../RTL/cortexm0ds_logic.v(17626)
  AL_DFF Emtax6_reg (
    .clk(HCLK),
    .d(Fuqhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Emtax6));  // ../RTL/cortexm0ds_logic.v(18888)
  AL_DFF Enpax6_reg (
    .clk(HCLK),
    .d(U6qhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Enpax6));  // ../RTL/cortexm0ds_logic.v(18816)
  AL_DFF Eotax6_reg (
    .clk(HCLK),
    .d(Qpqhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Eotax6));  // ../RTL/cortexm0ds_logic.v(18889)
  AL_DFF Eppax6_reg (
    .clk(HCLK),
    .d(Qxphu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Eppax6));  // ../RTL/cortexm0ds_logic.v(18817)
  AL_DFF Eqtax6_reg (
    .clk(HCLK),
    .d(Mgqhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Eqtax6));  // ../RTL/cortexm0ds_logic.v(18890)
  AL_DFF Equpw6_reg (
    .clk(HCLK),
    .d(Esohu6),
    .reset(1'b0),
    .set(n5973),
    .q(Equpw6));  // ../RTL/cortexm0ds_logic.v(17716)
  AL_DFF Erbbx6_reg (
    .clk(DCLK),
    .d(Fowhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Erbbx6));  // ../RTL/cortexm0ds_logic.v(19937)
  AL_DFF Erpax6_reg (
    .clk(HCLK),
    .d(Usphu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Erpax6));  // ../RTL/cortexm0ds_logic.v(18818)
  AL_DFF Esabx6_reg (
    .clk(DCLK),
    .d(Knwhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Esabx6));  // ../RTL/cortexm0ds_logic.v(19894)
  AL_DFF Estax6_reg (
    .clk(HCLK),
    .d(Xbqhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Estax6));  // ../RTL/cortexm0ds_logic.v(18891)
  AL_DFF Etfbx6_reg (
    .clk(DCLK),
    .d(Qxwhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Etfbx6));  // ../RTL/cortexm0ds_logic.v(20018)
  AL_DFF Eudax6_reg (
    .clk(DCLK),
    .d(Rnwhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Eudax6));  // ../RTL/cortexm0ds_logic.v(18296)
  AL_DFF Eutax6_reg (
    .clk(HCLK),
    .d(I7qhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Eutax6));  // ../RTL/cortexm0ds_logic.v(18892)
  AL_DFF Evbax6_reg (
    .clk(DCLK),
    .d(Y9whu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Evbax6));  // ../RTL/cortexm0ds_logic.v(18248)
  AL_DFF Evhpw6_reg (
    .clk(SWCLKTCK),
    .d(1'b1),
    .reset(n5971),
    .set(1'b0),
    .q(Evhpw6));  // ../RTL/cortexm0ds_logic.v(17154)
  AL_DFF Evypw6_reg (
    .clk(HCLK),
    .d(I4thu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Evypw6));  // ../RTL/cortexm0ds_logic.v(17893)
  AL_DFF Ewtax6_reg (
    .clk(HCLK),
    .d(Eyphu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Ewtax6));  // ../RTL/cortexm0ds_logic.v(18893)
  AL_DFF Exypw6_reg (
    .clk(HCLK),
    .d(B4thu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Exypw6));  // ../RTL/cortexm0ds_logic.v(17894)
  AL_DFF Eytax6_reg (
    .clk(HCLK),
    .d(Tophu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Eytax6));  // ../RTL/cortexm0ds_logic.v(18894)
  AL_DFF Eyyax6_reg (
    .clk(HCLK),
    .d(Qtthu6),
    .reset(n5973),
    .set(1'b0),
    .q(Eyyax6));  // ../RTL/cortexm0ds_logic.v(19053)
  AL_DFF Ez1qw6_reg (
    .clk(HCLK),
    .d(Btphu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Ez1qw6));  // ../RTL/cortexm0ds_logic.v(17950)
  AL_DFF Ezypw6_reg (
    .clk(HCLK),
    .d(N3thu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Ezypw6));  // ../RTL/cortexm0ds_logic.v(17895)
  AL_DFF F17ax6_reg (
    .clk(HCLK),
    .d(Rjthu6),
    .reset(n5973),
    .set(1'b0),
    .q(F17ax6));  // ../RTL/cortexm0ds_logic.v(18079)
  AL_DFF F1pax6_reg (
    .clk(HCLK),
    .d(Jvrhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(F1pax6));  // ../RTL/cortexm0ds_logic.v(18805)
  AL_DFF F26bx6_reg (
    .clk(HCLK),
    .d(Ruphu6),
    .reset(1'b0),
    .set(n5973),
    .q(F26bx6));  // ../RTL/cortexm0ds_logic.v(19747)
  AL_DFF F2dax6_reg (
    .clk(DCLK),
    .d(Yuwhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(F2dax6));  // ../RTL/cortexm0ds_logic.v(18276)
  AL_DFF F2tax6_reg (
    .clk(HCLK),
    .d(J9shu6),
    .reset(1'b0),
    .set(1'b0),
    .q(F2tax6));  // ../RTL/cortexm0ds_logic.v(18878)
  AL_DFF F3pax6_reg (
    .clk(HCLK),
    .d(Zprhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(F3pax6));  // ../RTL/cortexm0ds_logic.v(18806)
  AL_DFF F4iax6_reg (
    .clk(SCLK),
    .d(I2vhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(F4iax6));  // ../RTL/cortexm0ds_logic.v(18564)
  AL_DFF F4ibx6_reg (
    .clk(DCLK),
    .d(Uephu6),
    .reset(n5974),
    .set(1'b0),
    .q(F4ibx6));  // ../RTL/cortexm0ds_logic.v(20159)
  AL_DFF F4tax6_reg (
    .clk(HCLK),
    .d(U4shu6),
    .reset(1'b0),
    .set(1'b0),
    .q(F4tax6));  // ../RTL/cortexm0ds_logic.v(18879)
  AL_DFF F59bx6_reg (
    .clk(DCLK),
    .d(Ruwhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(F59bx6));  // ../RTL/cortexm0ds_logic.v(19809)
  AL_DFF F6dbx6_reg (
    .clk(HCLK),
    .d(Dsrhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(F6dbx6));  // ../RTL/cortexm0ds_logic.v(19969)
  AL_DFF F6tax6_reg (
    .clk(HCLK),
    .d(F0shu6),
    .reset(1'b0),
    .set(1'b0),
    .q(F6tax6));  // ../RTL/cortexm0ds_logic.v(18880)
  AL_DFF F7eax6_reg (
    .clk(DCLK),
    .d(Skwhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(F7eax6));  // ../RTL/cortexm0ds_logic.v(18303)
  AL_DFF F7jbx6_reg (
    .clk(DCLK),
    .d(X5whu6),
    .reset(1'b0),
    .set(1'b0),
    .q(F7jbx6));  // ../RTL/cortexm0ds_logic.v(20185)
  AL_DFF F8cbx6_reg (
    .clk(HCLK),
    .d(W5shu6),
    .reset(1'b0),
    .set(1'b0),
    .q(F8cbx6));  // ../RTL/cortexm0ds_logic.v(19946)
  AL_DFF F8dbx6_reg (
    .clk(DCLK),
    .d(P8phu6),
    .reset(1'b0),
    .set(1'b0),
    .q(F8dbx6));  // ../RTL/cortexm0ds_logic.v(19970)
  AL_DFF F8tax6_reg (
    .clk(HCLK),
    .d(Xvrhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(F8tax6));  // ../RTL/cortexm0ds_logic.v(18881)
  AL_DFF F9gbx6_reg (
    .clk(SCLK),
    .d(Z8uhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(F9gbx6));  // ../RTL/cortexm0ds_logic.v(20046)
  AL_DFF F9vpw6_reg (
    .clk(HCLK),
    .d(Hqohu6),
    .reset(n5973),
    .set(1'b0),
    .q(F9vpw6));  // ../RTL/cortexm0ds_logic.v(17771)
  AL_DFF Facax6_reg (
    .clk(DCLK),
    .d(Q5whu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Facax6));  // ../RTL/cortexm0ds_logic.v(18256)
  AL_DFF Facbx6_reg (
    .clk(DCLK),
    .d(Tpvhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Facbx6));  // ../RTL/cortexm0ds_logic.v(19947)
  AL_DFF Fahax6_reg (
    .clk(HCLK),
    .d(Bnohu6),
    .reset(1'b0),
    .set(n5973),
    .q(Fahax6));  // ../RTL/cortexm0ds_logic.v(18477)
  AL_DFF Fatax6_reg (
    .clk(HCLK),
    .d(Nqrhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Fatax6));  // ../RTL/cortexm0ds_logic.v(18882)
  AL_DFF Fb0bx6_reg (
    .clk(HCLK),
    .d(Fquhu6),
    .reset(n5973),
    .set(1'b0),
    .q(Fb0bx6));  // ../RTL/cortexm0ds_logic.v(19197)
  AL_DFF Fc1bx6_reg (
    .clk(SCLK),
    .d(F3phu6),
    .reset(n5973),
    .set(1'b0),
    .q(Fc1bx6));  // ../RTL/cortexm0ds_logic.v(19305)
  AL_DFF Fe2bx6_reg (
    .clk(SCLK),
    .d(N0phu6),
    .reset(n5973),
    .set(1'b0),
    .q(Fe2bx6));  // ../RTL/cortexm0ds_logic.v(19413)
  AL_DFF Fj8ax6_reg (
    .clk(SWCLKTCK),
    .d(Dmxhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Fj8ax6));  // ../RTL/cortexm0ds_logic.v(18123)
  AL_DFF Fjdbx6_reg (
    .clk(HCLK),
    .d(A9rhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Fjdbx6));  // ../RTL/cortexm0ds_logic.v(19976)
  AL_DFF Fkrpw6_reg (
    .clk(HCLK),
    .d(Ssohu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Fkrpw6));  // ../RTL/cortexm0ds_logic.v(17625)
  AL_DFF Fl2qw6_reg (
    .clk(DCLK),
    .d(B8phu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Fl2qw6));  // ../RTL/cortexm0ds_logic.v(17997)
  AL_DFF Fldbx6_reg (
    .clk(DCLK),
    .d(Dovhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Fldbx6));  // ../RTL/cortexm0ds_logic.v(19977)
  AL_DFF Fm7ax6_reg (
    .clk(DCLK),
    .d(P0xhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Fm7ax6));  // ../RTL/cortexm0ds_logic.v(18101)
  AL_DFF Fnnpw6_reg (
    .clk(SCLK),
    .d(Puohu6),
    .reset(1'b0),
    .set(n5973),
    .q(Fnnpw6));  // ../RTL/cortexm0ds_logic.v(17468)
  AL_DFF Fo9ax6_reg (
    .clk(DCLK),
    .d(Xkvhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Fo9ax6));  // ../RTL/cortexm0ds_logic.v(18170)
  AL_DFF Fpnpw6_reg (
    .clk(HCLK),
    .d(Iuohu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Fpnpw6));  // ../RTL/cortexm0ds_logic.v(17470)
  AL_DFF Ftaax6_reg (
    .clk(DCLK),
    .d(Iuvhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Ftaax6));  // ../RTL/cortexm0ds_logic.v(18192)
  AL_DFF Ftypw6_reg (
    .clk(HCLK),
    .d(P4thu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Ftypw6));  // ../RTL/cortexm0ds_logic.v(17892)
  AL_DFF Fvcbx6_reg (
    .clk(DCLK),
    .d(U0whu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Fvcbx6));  // ../RTL/cortexm0ds_logic.v(19963)
  AL_DFF Fvoax6_reg (
    .clk(HCLK),
    .d(V8shu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Fvoax6));  // ../RTL/cortexm0ds_logic.v(18802)
  AL_DFF Fx1qw6_reg (
    .clk(HCLK),
    .d(Nsphu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Fx1qw6));  // ../RTL/cortexm0ds_logic.v(17949)
  AL_DFF Fxoax6_reg (
    .clk(HCLK),
    .d(G4shu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Fxoax6));  // ../RTL/cortexm0ds_logic.v(18803)
  AL_DFF Fzmpw6_reg (
    .clk(HCLK),
    .d(Kkshu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Fzmpw6));  // ../RTL/cortexm0ds_logic.v(17447)
  AL_DFF Fzoax6_reg (
    .clk(HCLK),
    .d(Rzrhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Fzoax6));  // ../RTL/cortexm0ds_logic.v(18804)
  AL_DFF G0tax6_reg (
    .clk(HCLK),
    .d(Feshu6),
    .reset(1'b0),
    .set(1'b0),
    .q(G0tax6));  // ../RTL/cortexm0ds_logic.v(18877)
  AL_DFF G0zax6_reg (
    .clk(HCLK),
    .d(Vlthu6),
    .reset(n5973),
    .set(1'b0),
    .q(G0zax6));  // ../RTL/cortexm0ds_logic.v(19059)
  AL_DFF G25bx6_reg (
    .clk(HCLK),
    .d(Hzthu6),
    .reset(n5973),
    .set(1'b0),
    .q(G25bx6));  // ../RTL/cortexm0ds_logic.v(19689)
  AL_DFF G2iax6_reg (
    .clk(SCLK),
    .d(B2vhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(G2iax6));  // ../RTL/cortexm0ds_logic.v(18563)
  AL_DFF G54bx6_reg (
    .clk(HCLK),
    .d(K4uhu6),
    .reset(n5973),
    .set(1'b0),
    .q(G54bx6));  // ../RTL/cortexm0ds_logic.v(19593)
  AL_DFF G79ax6_reg (
    .clk(DCLK),
    .d(Mpvhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(G79ax6));  // ../RTL/cortexm0ds_logic.v(18161)
  AL_DFF G8ebx6_reg (
    .clk(DCLK),
    .d(D9whu6),
    .reset(1'b0),
    .set(1'b0),
    .q(G8ebx6));  // ../RTL/cortexm0ds_logic.v(19989)
  AL_DFF Gbvpw6_reg (
    .clk(DCLK),
    .d(R9phu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Gbvpw6));  // ../RTL/cortexm0ds_logic.v(17773)
  AL_DFF Gc1qw6_reg (
    .clk(SWCLKTCK),
    .d(Mnxhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Gc1qw6));  // ../RTL/cortexm0ds_logic.v(17938)
  AL_DFF Gd0bx6_reg (
    .clk(HCLK),
    .d(Tquhu6),
    .reset(n5973),
    .set(1'b0),
    .q(Gd0bx6));  // ../RTL/cortexm0ds_logic.v(19203)
  AL_DFF Ggabx6_reg (
    .clk(DCLK),
    .d(Hbphu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Ggabx6));  // ../RTL/cortexm0ds_logic.v(19888)
  AL_DFF Gihbx6_reg (
    .clk(SCLK),
    .d(H4phu6),
    .reset(n5973),
    .set(1'b0),
    .q(Gihbx6));  // ../RTL/cortexm0ds_logic.v(20118)
  AL_DFF Gkeax6_reg (
    .clk(DCLK),
    .d(Rgwhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Gkeax6));  // ../RTL/cortexm0ds_logic.v(18315)
  AL_DFF Gl1qw6_reg (
    .clk(SWCLKTCK),
    .d(Fnxhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Gl1qw6));  // ../RTL/cortexm0ds_logic.v(17943)
  AL_DFF Gnqpw6_reg (
    .clk(SWCLKTCK),
    .d(Ahxhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Gnqpw6));  // ../RTL/cortexm0ds_logic.v(17574)
  AL_DFF Golpw6_reg (
    .clk(SWCLKTCK),
    .d(Yvohu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Golpw6));  // ../RTL/cortexm0ds_logic.v(17382)
  AL_DFF Gp6ax6_reg (
    .clk(HCLK),
    .d(L2thu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Gp6ax6));  // ../RTL/cortexm0ds_logic.v(18064)
  AL_DFF Gpqpw6_reg (
    .clk(SWCLKTCK),
    .d(Qpxhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Gpqpw6));  // ../RTL/cortexm0ds_logic.v(17575)
  AL_DFF Gr2qw6_reg (
    .clk(DCLK),
    .d(W0xhu6),
    .reset(n5974),
    .set(1'b0),
    .q(Gr2qw6));  // ../RTL/cortexm0ds_logic.v(18004)
  AL_DFF Gr6ax6_reg (
    .clk(HCLK),
    .d(U3thu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Gr6ax6));  // ../RTL/cortexm0ds_logic.v(18065)
  AL_DFF Gt6ax6_reg (
    .clk(HCLK),
    .d(X8thu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Gt6ax6));  // ../RTL/cortexm0ds_logic.v(18066)
  AL_DFF Gtoax6_reg (
    .clk(HCLK),
    .d(Rdshu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Gtoax6));  // ../RTL/cortexm0ds_logic.v(18801)
  AL_DFF Gv1bx6_reg (
    .clk(SCLK),
    .d(Zgthu6),
    .reset(n5973),
    .set(1'b0),
    .q(Gv1bx6));  // ../RTL/cortexm0ds_logic.v(19359)
  AL_DFF Gv1qw6_reg (
    .clk(HCLK),
    .d(Zrphu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Gv1qw6));  // ../RTL/cortexm0ds_logic.v(17948)
  AL_DFF Gv6ax6_reg (
    .clk(HCLK),
    .d(W9vhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Gv6ax6));  // ../RTL/cortexm0ds_logic.v(18067)
  AL_DFF Gvmpw6_reg (
    .clk(HCLK),
    .d(Ocvhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Gvmpw6));  // ../RTL/cortexm0ds_logic.v(17445)
  AL_DFF Gw6bx6_reg (
    .clk(SWCLKTCK),
    .d(Qwxhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Gw6bx6));  // ../RTL/cortexm0ds_logic.v(19763)
  AL_DFF Gwwpw6_reg (
    .clk(SWCLKTCK),
    .d(Ukxhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Gwwpw6));  // ../RTL/cortexm0ds_logic.v(17827)
  AL_DFF Gwxpw6_reg (
    .clk(HCLK),
    .d(Gzphu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Gwxpw6));  // ../RTL/cortexm0ds_logic.v(17855)
  AL_DFF Gx2bx6_reg (
    .clk(SCLK),
    .d(Wpthu6),
    .reset(n5973),
    .set(1'b0),
    .q(Gx2bx6));  // ../RTL/cortexm0ds_logic.v(19467)
  AL_DFF Gx6ax6_reg (
    .clk(HCLK),
    .d(Davhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Gx6ax6));  // ../RTL/cortexm0ds_logic.v(18068)
  AL_DFF Gxmpw6_reg (
    .clk(HCLK),
    .d(Gpshu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Gxmpw6));  // ../RTL/cortexm0ds_logic.v(17446)
  AL_DFF Gylpw6_reg (
    .clk(SWCLKTCK),
    .d(Ktxhu6),
    .reset(n5972),
    .set(1'b0),
    .q(Gylpw6));  // ../RTL/cortexm0ds_logic.v(17402)
  AL_DFF Gyxpw6_reg (
    .clk(DCLK),
    .d(Ccphu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Gyxpw6));  // ../RTL/cortexm0ds_logic.v(17856)
  AL_DFF Gz6ax6_reg (
    .clk(HCLK),
    .d(Mkthu6),
    .reset(n5973),
    .set(1'b0),
    .q(Gz6ax6));  // ../RTL/cortexm0ds_logic.v(18073)
  AL_DFF Gzeax6_reg (
    .clk(DCLK),
    .d(Ldwhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Gzeax6));  // ../RTL/cortexm0ds_logic.v(18323)
  AL_DFF H0ebx6_reg (
    .clk(SWCLKTCK),
    .d(Zjxhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(H0ebx6));  // ../RTL/cortexm0ds_logic.v(19985)
  AL_DFF H3lpw6_reg (
    .clk(DCLK),
    .d(L6phu6),
    .reset(1'b0),
    .set(1'b0),
    .q(H3lpw6));  // ../RTL/cortexm0ds_logic.v(17325)
  AL_DFF H4bax6_reg (
    .clk(DCLK),
    .d(T3whu6),
    .reset(n5974),
    .set(1'b0),
    .q(H4bax6));  // ../RTL/cortexm0ds_logic.v(18217)
  AL_DFF H4ypw6_reg (
    .clk(DCLK),
    .d(Pexhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(H4ypw6));  // ../RTL/cortexm0ds_logic.v(17859)
  AL_DFF H4zax6_reg (
    .clk(HCLK),
    .d(S1uhu6),
    .reset(n5973),
    .set(1'b0),
    .q(H4zax6));  // ../RTL/cortexm0ds_logic.v(19071)
  AL_DFF H7hbx6_reg (
    .clk(DCLK),
    .d(Cbxhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(H7hbx6));  // ../RTL/cortexm0ds_logic.v(20103)
  AL_DFF H8gax6_reg (
    .clk(DCLK),
    .d(Qjwhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(H8gax6));  // ../RTL/cortexm0ds_logic.v(18402)
  AL_DFF Halax6_reg (
    .clk(HCLK),
    .d(Z7vhu6),
    .reset(n5973),
    .set(1'b0),
    .q(Halax6));  // ../RTL/cortexm0ds_logic.v(18736)
  AL_DFF Hbgbx6_reg (
    .clk(HCLK),
    .d(J7uhu6),
    .reset(n5973),
    .set(1'b0),
    .q(Hbgbx6));  // ../RTL/cortexm0ds_logic.v(20051)
  AL_DFF Hdbax6_reg (
    .clk(DCLK),
    .d(K2whu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Hdbax6));  // ../RTL/cortexm0ds_logic.v(18223)
  AL_DFF Hdfax6_reg (
    .clk(DCLK),
    .d(D1xhu6),
    .reset(n5974),
    .set(1'b0),
    .q(Hdfax6));  // ../RTL/cortexm0ds_logic.v(18355)
  AL_DFF Heaax6_reg (
    .clk(DCLK),
    .d(Oxvhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Heaax6));  // ../RTL/cortexm0ds_logic.v(18184)
  AL_DFF Hf0bx6_reg (
    .clk(HCLK),
    .d(Hruhu6),
    .reset(n5973),
    .set(1'b0),
    .q(Hf0bx6));  // ../RTL/cortexm0ds_logic.v(19209)
  AL_DFF Hg3bx6_reg (
    .clk(SCLK),
    .d(Cyohu6),
    .reset(n5973),
    .set(1'b0),
    .q(Hg3bx6));  // ../RTL/cortexm0ds_logic.v(19521)
  AL_DFF Hg7ax6_reg (
    .clk(DCLK),
    .d(Gephu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Hg7ax6));  // ../RTL/cortexm0ds_logic.v(18098)
  AL_DFF Hgrpw6_reg (
    .clk(HCLK),
    .d(X4xhu6),
    .reset(1'b0),
    .set(n5973),
    .q(Hgrpw6));  // ../RTL/cortexm0ds_logic.v(17617)
  AL_DFF Hhvpw6_reg (
    .clk(HCLK),
    .d(Akuhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Hhvpw6));  // ../RTL/cortexm0ds_logic.v(17776)
  AL_DFF Hi9bx6_reg (
    .clk(DCLK),
    .d(Edwhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Hi9bx6));  // ../RTL/cortexm0ds_logic.v(19816)
  AL_DFF Hirpw6_reg (
    .clk(HCLK),
    .d(Zsohu6),
    .reset(n5973),
    .set(1'b0),
    .q(Hirpw6));  // ../RTL/cortexm0ds_logic.v(17623)
  AL_DFF Hjgax6_reg (
    .clk(DCLK),
    .d(Abwhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Hjgax6));  // ../RTL/cortexm0ds_logic.v(18408)
  AL_DFF Hkxpw6_reg (
    .clk(HCLK),
    .d(Yuphu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Hkxpw6));  // ../RTL/cortexm0ds_logic.v(17849)
  AL_DFF Hlcax6_reg (
    .clk(DCLK),
    .d(B0xhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Hlcax6));  // ../RTL/cortexm0ds_logic.v(18267)
  AL_DFF Hlwpw6_reg (
    .clk(SWCLKTCK),
    .d(Zxxhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Hlwpw6));  // ../RTL/cortexm0ds_logic.v(17816)
  AL_DFF Hmbax6_reg (
    .clk(DCLK),
    .d(Oyuhu6),
    .reset(n5974),
    .set(1'b0),
    .q(Hmbax6));  // ../RTL/cortexm0ds_logic.v(18237)
  AL_DFF Hmxpw6_reg (
    .clk(HCLK),
    .d(Fvphu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Hmxpw6));  // ../RTL/cortexm0ds_logic.v(17850)
  AL_DFF Hoxpw6_reg (
    .clk(HCLK),
    .d(Hwphu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Hoxpw6));  // ../RTL/cortexm0ds_logic.v(17851)
  AL_DFF Hpbbx6_reg (
    .clk(DCLK),
    .d(Dgwhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Hpbbx6));  // ../RTL/cortexm0ds_logic.v(19936)
  AL_DFF Hpcbx6_reg (
    .clk(SWCLKTCK),
    .d(Mgxhu6),
    .reset(n5972),
    .set(1'b0),
    .q(Hpcbx6));  // ../RTL/cortexm0ds_logic.v(19959)
  AL_DFF Hphax6_reg (
    .clk(HCLK),
    .d(Xkohu6),
    .reset(1'b0),
    .set(n5973),
    .q(Hphax6));  // ../RTL/cortexm0ds_logic.v(18525)
  AL_DFF Hqabx6_reg (
    .clk(DCLK),
    .d(Ifwhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Hqabx6));  // ../RTL/cortexm0ds_logic.v(19893)
  AL_DFF Hqxpw6_reg (
    .clk(HCLK),
    .d(Vwphu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Hqxpw6));  // ../RTL/cortexm0ds_logic.v(17852)
  AL_DFF Hrfbx6_reg (
    .clk(DCLK),
    .d(Opwhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Hrfbx6));  // ../RTL/cortexm0ds_logic.v(20017)
  AL_DFF Hroax6_reg (
    .clk(HCLK),
    .d(Gishu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Hroax6));  // ../RTL/cortexm0ds_logic.v(18800)
  AL_DFF Hsdax6_reg (
    .clk(DCLK),
    .d(Ynwhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Hsdax6));  // ../RTL/cortexm0ds_logic.v(18295)
  AL_DFF Hsxpw6_reg (
    .clk(HCLK),
    .d(Jxphu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Hsxpw6));  // ../RTL/cortexm0ds_logic.v(17853)
  AL_DFF Ht1qw6_reg (
    .clk(HCLK),
    .d(Lrphu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Ht1qw6));  // ../RTL/cortexm0ds_logic.v(17947)
  AL_DFF Htbax6_reg (
    .clk(DCLK),
    .d(Fawhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Htbax6));  // ../RTL/cortexm0ds_logic.v(18247)
  AL_DFF Htmpw6_reg (
    .clk(HCLK),
    .d(Wuohu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Htmpw6));  // ../RTL/cortexm0ds_logic.v(17444)
  AL_DFF Huxpw6_reg (
    .clk(HCLK),
    .d(Zyphu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Huxpw6));  // ../RTL/cortexm0ds_logic.v(17854)
  AL_DFF Hw8ax6_reg (
    .clk(DCLK),
    .d(Y1xhu6),
    .reset(n5974),
    .set(1'b0),
    .q(Hw8ax6));  // ../RTL/cortexm0ds_logic.v(18139)
  AL_DFF Hwhpw6_reg (
    .clk(SWCLKTCK),
    .d(Qmdhu6),
    .reset(n5971),
    .set(1'b0),
    .q(Hwhpw6));  // ../RTL/cortexm0ds_logic.v(17160)
  AL_DFF Hysax6_reg (
    .clk(HCLK),
    .d(Uishu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Hysax6));  // ../RTL/cortexm0ds_logic.v(18876)
  AL_DFF Hz9ax6_reg (
    .clk(DCLK),
    .d(Ajvhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Hz9ax6));  // ../RTL/cortexm0ds_logic.v(18176)
  AL_DFF I0dax6_reg (
    .clk(DCLK),
    .d(Fvwhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(I0dax6));  // ../RTL/cortexm0ds_logic.v(18275)
  AL_DFF I0opw6_reg (
    .clk(SWCLKTCK),
    .d(Q3yhu6),
    .reset(n5972),
    .set(1'b0),
    .q(I0opw6));  // ../RTL/cortexm0ds_logic.v(17490)
  AL_DFF I1lpw6_reg (
    .clk(HCLK),
    .d(Qdvhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(I1lpw6));  // ../RTL/cortexm0ds_logic.v(17324)
  AL_DFF I1qpw6_reg (
    .clk(HCLK),
    .d(O9rhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(I1qpw6));  // ../RTL/cortexm0ds_logic.v(17548)
  AL_DFF I2zax6_reg (
    .clk(HCLK),
    .d(Olthu6),
    .reset(n5973),
    .set(1'b0),
    .q(I2zax6));  // ../RTL/cortexm0ds_logic.v(19065)
  AL_DFF I3qpw6_reg (
    .clk(HCLK),
    .d(Z4rhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(I3qpw6));  // ../RTL/cortexm0ds_logic.v(17549)
  AL_DFF I45bx6_reg (
    .clk(HCLK),
    .d(Azthu6),
    .reset(n5973),
    .set(1'b0),
    .q(I45bx6));  // ../RTL/cortexm0ds_logic.v(19695)
  AL_DFF I4rpw6_reg (
    .clk(SWCLKTCK),
    .d(Hhxhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(I4rpw6));  // ../RTL/cortexm0ds_logic.v(17597)
  AL_DFF I5qpw6_reg (
    .clk(HCLK),
    .d(Y8qhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(I5qpw6));  // ../RTL/cortexm0ds_logic.v(17550)
  AL_DFF I5xax6_reg (
    .clk(HCLK),
    .d(Hcvhu6),
    .reset(n5973),
    .set(1'b0),
    .q(I5xax6));  // ../RTL/cortexm0ds_logic.v(18956)
  AL_DFF I74bx6_reg (
    .clk(HCLK),
    .d(Kxthu6),
    .reset(n5973),
    .set(1'b0),
    .q(I74bx6));  // ../RTL/cortexm0ds_logic.v(19599)
  AL_DFF I7qpw6_reg (
    .clk(HCLK),
    .d(J4qhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(I7qpw6));  // ../RTL/cortexm0ds_logic.v(17551)
  AL_DFF I8hax6_reg (
    .clk(HCLK),
    .d(Inohu6),
    .reset(1'b0),
    .set(n5973),
    .q(I8hax6));  // ../RTL/cortexm0ds_logic.v(18471)
  AL_DFF I8lax6_reg (
    .clk(HCLK),
    .d(Qdohu6),
    .reset(n5973),
    .set(1'b0),
    .q(I8lax6));  // ../RTL/cortexm0ds_logic.v(18730)
  AL_DFF I9qpw6_reg (
    .clk(HCLK),
    .d(Ygphu6),
    .reset(1'b0),
    .set(1'b0),
    .q(I9qpw6));  // ../RTL/cortexm0ds_logic.v(17552)
  AL_DFF Ibqpw6_reg (
    .clk(HCLK),
    .d(Zkphu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Ibqpw6));  // ../RTL/cortexm0ds_logic.v(17553)
  AL_DFF Iddax6_reg (
    .clk(DCLK),
    .d(Nswhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Iddax6));  // ../RTL/cortexm0ds_logic.v(18282)
  AL_DFF Idqpw6_reg (
    .clk(DCLK),
    .d(G7phu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Idqpw6));  // ../RTL/cortexm0ds_logic.v(17554)
  AL_DFF Ie1bx6_reg (
    .clk(SCLK),
    .d(Znthu6),
    .reset(n5973),
    .set(1'b0),
    .q(Ie1bx6));  // ../RTL/cortexm0ds_logic.v(19311)
  AL_DFF Iekax6_reg (
    .clk(HCLK),
    .d(Xfthu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Iekax6));  // ../RTL/cortexm0ds_logic.v(18701)
  AL_DFF Ig2bx6_reg (
    .clk(SCLK),
    .d(Ztuhu6),
    .reset(n5973),
    .set(1'b0),
    .q(Ig2bx6));  // ../RTL/cortexm0ds_logic.v(19419)
  AL_DFF Ih0bx6_reg (
    .clk(HCLK),
    .d(Oruhu6),
    .reset(n5973),
    .set(1'b0),
    .q(Ih0bx6));  // ../RTL/cortexm0ds_logic.v(19215)
  AL_DFF Iixpw6_reg (
    .clk(HCLK),
    .d(Q4xhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Iixpw6));  // ../RTL/cortexm0ds_logic.v(17848)
  AL_DFF Ijiax6_reg (
    .clk(HCLK),
    .d(Ctthu6),
    .reset(n5973),
    .set(1'b0),
    .q(Ijiax6));  // ../RTL/cortexm0ds_logic.v(18601)
  AL_DFF Ikhbx6_reg (
    .clk(HCLK),
    .d(Gnuhu6),
    .reset(n5973),
    .set(1'b0),
    .q(Ikhbx6));  // ../RTL/cortexm0ds_logic.v(20124)
  AL_DFF Im9ax6_reg (
    .clk(DCLK),
    .d(Llvhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Im9ax6));  // ../RTL/cortexm0ds_logic.v(18169)
  AL_DFF Imhbx6_reg (
    .clk(HCLK),
    .d(Zfuhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Imhbx6));  // ../RTL/cortexm0ds_logic.v(20126)
  AL_DFF Ipoax6_reg (
    .clk(HCLK),
    .d(Vmshu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Ipoax6));  // ../RTL/cortexm0ds_logic.v(18799)
  AL_DFF Ir1qw6_reg (
    .clk(HCLK),
    .d(Jqphu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Ir1qw6));  // ../RTL/cortexm0ds_logic.v(17946)
  AL_DFF Irmpw6_reg (
    .clk(HCLK),
    .d(Uhthu6),
    .reset(1'b0),
    .set(n5973),
    .q(Irmpw6));  // ../RTL/cortexm0ds_logic.v(17442)
  AL_DFF Isjpw6_reg (
    .clk(DCLK),
    .d(E5xhu6),
    .reset(n5974),
    .set(1'b0),
    .q(Isjpw6));  // ../RTL/cortexm0ds_logic.v(17265)
  AL_DFF Itcbx6_reg (
    .clk(DCLK),
    .d(Aqvhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Itcbx6));  // ../RTL/cortexm0ds_logic.v(19962)
  AL_DFF Iwsax6_reg (
    .clk(HCLK),
    .d(Jnshu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Iwsax6));  // ../RTL/cortexm0ds_logic.v(18875)
  AL_DFF Ixppw6_reg (
    .clk(HCLK),
    .d(Nxrhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Ixppw6));  // ../RTL/cortexm0ds_logic.v(17546)
  AL_DFF Izppw6_reg (
    .clk(HCLK),
    .d(Ftrhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Izppw6));  // ../RTL/cortexm0ds_logic.v(17547)
  AL_DFF J06bx6_reg (
    .clk(HCLK),
    .d(Cdohu6),
    .reset(1'b0),
    .set(n5973),
    .q(J06bx6));  // ../RTL/cortexm0ds_logic.v(19741)
  AL_DFF J0gax6_reg (
    .clk(SWCLKTCK),
    .d(Tuxhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(J0gax6));  // ../RTL/cortexm0ds_logic.v(18398)
  AL_DFF J0iax6_reg (
    .clk(HCLK),
    .d(Hjohu6),
    .reset(1'b0),
    .set(n5973),
    .q(J0iax6));  // ../RTL/cortexm0ds_logic.v(18561)
  AL_DFF J39bx6_reg (
    .clk(DCLK),
    .d(Pmwhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(J39bx6));  // ../RTL/cortexm0ds_logic.v(19808)
  AL_DFF J3xax6_reg (
    .clk(HCLK),
    .d(Kcthu6),
    .reset(1'b0),
    .set(1'b0),
    .q(J3xax6));  // ../RTL/cortexm0ds_logic.v(18951)
  AL_DFF J4cbx6_reg (
    .clk(SWCLKTCK),
    .d(R0yhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(J4cbx6));  // ../RTL/cortexm0ds_logic.v(19944)
  AL_DFF J59ax6_reg (
    .clk(DCLK),
    .d(Vqvhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(J59ax6));  // ../RTL/cortexm0ds_logic.v(18160)
  AL_DFF J5eax6_reg (
    .clk(DCLK),
    .d(Zkwhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(J5eax6));  // ../RTL/cortexm0ds_logic.v(18302)
  AL_DFF J5jbx6_reg (
    .clk(DCLK),
    .d(Yvvhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(J5jbx6));  // ../RTL/cortexm0ds_logic.v(20184)
  AL_DFF J6ebx6_reg (
    .clk(DCLK),
    .d(Ezvhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(J6ebx6));  // ../RTL/cortexm0ds_logic.v(19988)
  AL_DFF J6zax6_reg (
    .clk(HCLK),
    .d(L1uhu6),
    .reset(n5973),
    .set(1'b0),
    .q(J6zax6));  // ../RTL/cortexm0ds_logic.v(19077)
  AL_DFF J7xax6_reg (
    .clk(HCLK),
    .d(Cluhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(J7xax6));  // ../RTL/cortexm0ds_logic.v(18958)
  AL_DFF J8cax6_reg (
    .clk(DCLK),
    .d(E6whu6),
    .reset(1'b0),
    .set(1'b0),
    .q(J8cax6));  // ../RTL/cortexm0ds_logic.v(18255)
  AL_DFF Jckax6_reg (
    .clk(HCLK),
    .d(Pithu6),
    .reset(1'b0),
    .set(n5973),
    .q(Jckax6));  // ../RTL/cortexm0ds_logic.v(18699)
  AL_DFF Jdgbx6_reg (
    .clk(HCLK),
    .d(F5uhu6),
    .reset(n5973),
    .set(1'b0),
    .q(Jdgbx6));  // ../RTL/cortexm0ds_logic.v(20057)
  AL_DFF Jfdbx6_reg (
    .clk(SWCLKTCK),
    .d(Bzxhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Jfdbx6));  // ../RTL/cortexm0ds_logic.v(19974)
  AL_DFF Jflpw6_reg (
    .clk(SWCLKTCK),
    .d(Zehpw6[3]),
    .reset(n5972),
    .set(1'b0),
    .q(Jflpw6));  // ../RTL/cortexm0ds_logic.v(17356)
  AL_DFF Jgxpw6_reg (
    .clk(HCLK),
    .d(Iithu6),
    .reset(1'b0),
    .set(n5973),
    .q(Jgxpw6));  // ../RTL/cortexm0ds_logic.v(17846)
  AL_DFF Jhebx6_reg (
    .clk(DCLK),
    .d(D9phu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Jhebx6));  // ../RTL/cortexm0ds_logic.v(19994)
  AL_DFF Jieax6_reg (
    .clk(DCLK),
    .d(Aiwhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Jieax6));  // ../RTL/cortexm0ds_logic.v(18314)
  AL_DFF Jj0bx6_reg (
    .clk(HCLK),
    .d(Csuhu6),
    .reset(n5973),
    .set(1'b0),
    .q(Jj0bx6));  // ../RTL/cortexm0ds_logic.v(19221)
  AL_DFF Jjvpw6_reg (
    .clk(HCLK),
    .d(D0rhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Jjvpw6));  // ../RTL/cortexm0ds_logic.v(17777)
  AL_DFF Jl3qw6_reg (
    .clk(DCLK),
    .d(Lcxhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Jl3qw6));  // ../RTL/cortexm0ds_logic.v(18042)
  AL_DFF Jlvpw6_reg (
    .clk(HCLK),
    .d(K0rhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Jlvpw6));  // ../RTL/cortexm0ds_logic.v(17778)
  AL_DFF Jnoax6_reg (
    .clk(HCLK),
    .d(Rrshu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Jnoax6));  // ../RTL/cortexm0ds_logic.v(18798)
  AL_DFF Jnvpw6_reg (
    .clk(HCLK),
    .d(M1rhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Jnvpw6));  // ../RTL/cortexm0ds_logic.v(17779)
  AL_DFF Johbx6_reg (
    .clk(SCLK),
    .d(Vduhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Johbx6));  // ../RTL/cortexm0ds_logic.v(20127)
  AL_DFF Jp1qw6_reg (
    .clk(HCLK),
    .d(Cqphu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Jp1qw6));  // ../RTL/cortexm0ds_logic.v(17945)
  AL_DFF Jp9bx6_reg (
    .clk(SCLK),
    .d(Osthu6),
    .reset(n5973),
    .set(1'b0),
    .q(Jp9bx6));  // ../RTL/cortexm0ds_logic.v(19824)
  AL_DFF Jpmpw6_reg (
    .clk(SCLK),
    .d(N1vhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Jpmpw6));  // ../RTL/cortexm0ds_logic.v(17437)
  AL_DFF Jpvpw6_reg (
    .clk(HCLK),
    .d(A2rhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Jpvpw6));  // ../RTL/cortexm0ds_logic.v(17780)
  AL_DFF Jraax6_reg (
    .clk(DCLK),
    .d(Puvhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Jraax6));  // ../RTL/cortexm0ds_logic.v(18191)
  AL_DFF Jrvpw6_reg (
    .clk(HCLK),
    .d(O2rhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Jrvpw6));  // ../RTL/cortexm0ds_logic.v(17781)
  AL_DFF Jrypw6_reg (
    .clk(HCLK),
    .d(P9vhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Jrypw6));  // ../RTL/cortexm0ds_logic.v(17891)
  AL_DFF Jtvpw6_reg (
    .clk(HCLK),
    .d(E4rhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Jtvpw6));  // ../RTL/cortexm0ds_logic.v(17782)
  AL_DFF Jusax6_reg (
    .clk(HCLK),
    .d(Fsshu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Jusax6));  // ../RTL/cortexm0ds_logic.v(18874)
  AL_DFF Jvkpw6_reg (
    .clk(SWCLKTCK),
    .d(Ejxhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Jvkpw6));  // ../RTL/cortexm0ds_logic.v(17311)
  AL_DFF Jvppw6_reg (
    .clk(HCLK),
    .d(Rkshu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Jvppw6));  // ../RTL/cortexm0ds_logic.v(17545)
  AL_DFF Jvvpw6_reg (
    .clk(DCLK),
    .d(Dhvhu6),
    .reset(n5974),
    .set(1'b0),
    .q(Jvvpw6));  // ../RTL/cortexm0ds_logic.v(17787)
  AL_DFF Jx1bx6_reg (
    .clk(SCLK),
    .d(P1phu6),
    .reset(n5973),
    .set(1'b0),
    .q(Jx1bx6));  // ../RTL/cortexm0ds_logic.v(19365)
  AL_DFF Jxgax6_reg (
    .clk(DCLK),
    .d(V3xhu6),
    .reset(1'b0),
    .set(n5974),
    .q(Jxgax6));  // ../RTL/cortexm0ds_logic.v(18435)
  AL_DFF Jy5bx6_reg (
    .clk(HCLK),
    .d(Njrhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Jy5bx6));  // ../RTL/cortexm0ds_logic.v(19736)
  AL_DFF Jz2bx6_reg (
    .clk(SCLK),
    .d(Lzohu6),
    .reset(n5973),
    .set(1'b0),
    .q(Jz2bx6));  // ../RTL/cortexm0ds_logic.v(19473)
  AL_DFF K1xax6_reg (
    .clk(HCLK),
    .d(Rcthu6),
    .reset(1'b0),
    .set(1'b0),
    .q(K1xax6));  // ../RTL/cortexm0ds_logic.v(18950)
  AL_DFF K5hbx6_reg (
    .clk(DCLK),
    .d(Xxwhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(K5hbx6));  // ../RTL/cortexm0ds_logic.v(20102)
  AL_DFF K65bx6_reg (
    .clk(HCLK),
    .d(Mythu6),
    .reset(n5973),
    .set(1'b0),
    .q(K65bx6));  // ../RTL/cortexm0ds_logic.v(19701)
  AL_DFF K6gax6_reg (
    .clk(DCLK),
    .d(Obwhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(K6gax6));  // ../RTL/cortexm0ds_logic.v(18401)
  AL_DFF K7vpw6_reg (
    .clk(DCLK),
    .d(Vyuhu6),
    .reset(1'b0),
    .set(n5974),
    .q(K7vpw6));  // ../RTL/cortexm0ds_logic.v(17765)
  AL_DFF K94bx6_reg (
    .clk(HCLK),
    .d(Dxthu6),
    .reset(n5973),
    .set(1'b0),
    .q(K94bx6));  // ../RTL/cortexm0ds_logic.v(19605)
  AL_DFF Kadbx6_reg (
    .clk(SWCLKTCK),
    .d(Wzxhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Kadbx6));  // ../RTL/cortexm0ds_logic.v(19971)
  AL_DFF Kakax6_reg (
    .clk(HCLK),
    .d(Seohu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Kakax6));  // ../RTL/cortexm0ds_logic.v(18694)
  AL_DFF Kalpw6_reg (
    .clk(SWCLKTCK),
    .d(Zehpw6[2]),
    .reset(1'b0),
    .set(n5972),
    .q(Kalpw6));  // ../RTL/cortexm0ds_logic.v(17338)
  AL_DFF Kcaax6_reg (
    .clk(DCLK),
    .d(Vxvhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Kcaax6));  // ../RTL/cortexm0ds_logic.v(18183)
  AL_DFF Ke1qw6_reg (
    .clk(DCLK),
    .d(U6xhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Ke1qw6));  // ../RTL/cortexm0ds_logic.v(17939)
  AL_DFF Kfoax6_reg (
    .clk(HCLK),
    .d(H7thu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Kfoax6));  // ../RTL/cortexm0ds_logic.v(18794)
  AL_DFF Khgax6_reg (
    .clk(DCLK),
    .d(B1whu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Khgax6));  // ../RTL/cortexm0ds_logic.v(18407)
  AL_DFF Khoax6_reg (
    .clk(HCLK),
    .d(A7thu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Khoax6));  // ../RTL/cortexm0ds_logic.v(18795)
  AL_DFF Ki3bx6_reg (
    .clk(SCLK),
    .d(Hsthu6),
    .reset(n5973),
    .set(1'b0),
    .q(Ki3bx6));  // ../RTL/cortexm0ds_logic.v(19527)
  AL_DFF Kjoax6_reg (
    .clk(HCLK),
    .d(T6thu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Kjoax6));  // ../RTL/cortexm0ds_logic.v(18796)
  AL_DFF Kkjpw6_reg (
    .clk(HCLK),
    .d(Ourhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Kkjpw6));  // ../RTL/cortexm0ds_logic.v(17247)
  AL_DFF Kl0bx6_reg (
    .clk(HCLK),
    .d(Qsuhu6),
    .reset(n5973),
    .set(1'b0),
    .q(Kl0bx6));  // ../RTL/cortexm0ds_logic.v(19227)
  AL_DFF Kl8ax6_reg (
    .clk(DCLK),
    .d(Udxhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Kl8ax6));  // ../RTL/cortexm0ds_logic.v(18124)
  AL_DFF Kloax6_reg (
    .clk(HCLK),
    .d(M6thu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Kloax6));  // ../RTL/cortexm0ds_logic.v(18797)
  AL_DFF Kmjpw6_reg (
    .clk(HCLK),
    .d(Zwrhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Kmjpw6));  // ../RTL/cortexm0ds_logic.v(17248)
  AL_DFF Kmsax6_reg (
    .clk(HCLK),
    .d(Tzshu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Kmsax6));  // ../RTL/cortexm0ds_logic.v(18870)
  AL_DFF Kn1qw6_reg (
    .clk(HCLK),
    .d(Kuphu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Kn1qw6));  // ../RTL/cortexm0ds_logic.v(17944)
  AL_DFF Kn2qw6_reg (
    .clk(SWCLKTCK),
    .d(K0yhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Kn2qw6));  // ../RTL/cortexm0ds_logic.v(17998)
  AL_DFF Knbbx6_reg (
    .clk(DCLK),
    .d(B8whu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Knbbx6));  // ../RTL/cortexm0ds_logic.v(19935)
  AL_DFF Knhax6_reg (
    .clk(HCLK),
    .d(Elohu6),
    .reset(1'b0),
    .set(n5973),
    .q(Knhax6));  // ../RTL/cortexm0ds_logic.v(18519)
  AL_DFF Koabx6_reg (
    .clk(DCLK),
    .d(G7whu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Koabx6));  // ../RTL/cortexm0ds_logic.v(19892)
  AL_DFF Kojpw6_reg (
    .clk(HCLK),
    .d(Mxuhu6),
    .reset(n5973),
    .set(1'b0),
    .q(Kojpw6));  // ../RTL/cortexm0ds_logic.v(17253)
  AL_DFF Kosax6_reg (
    .clk(HCLK),
    .d(Mzshu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Kosax6));  // ../RTL/cortexm0ds_logic.v(18871)
  AL_DFF Kpfbx6_reg (
    .clk(DCLK),
    .d(Mhwhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Kpfbx6));  // ../RTL/cortexm0ds_logic.v(20016)
  AL_DFF Kqdax6_reg (
    .clk(DCLK),
    .d(Mowhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Kqdax6));  // ../RTL/cortexm0ds_logic.v(18294)
  AL_DFF Kqhbx6_reg (
    .clk(HCLK),
    .d(Jtthu6),
    .reset(n5973),
    .set(1'b0),
    .q(Kqhbx6));  // ../RTL/cortexm0ds_logic.v(20132)
  AL_DFF Kqsax6_reg (
    .clk(HCLK),
    .d(Fzshu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Kqsax6));  // ../RTL/cortexm0ds_logic.v(18872)
  AL_DFF Krbax6_reg (
    .clk(DCLK),
    .d(Hbwhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Krbax6));  // ../RTL/cortexm0ds_logic.v(18246)
  AL_DFF Krlpw6_reg (
    .clk(SWCLKTCK),
    .d(Kvohu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Krlpw6));  // ../RTL/cortexm0ds_logic.v(17384)
  AL_DFF Ksgax6_reg (
    .clk(DCLK),
    .d(Kfxhu6),
    .reset(n5974),
    .set(1'b0),
    .q(Ksgax6));  // ../RTL/cortexm0ds_logic.v(18417)
  AL_DFF Kshbx6_reg (
    .clk(SCLK),
    .d(Trthu6),
    .reset(n5973),
    .set(1'b0),
    .q(Kshbx6));  // ../RTL/cortexm0ds_logic.v(20138)
  AL_DFF Kssax6_reg (
    .clk(HCLK),
    .d(Yyshu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Kssax6));  // ../RTL/cortexm0ds_logic.v(18873)
  AL_DFF Kswpw6_reg (
    .clk(DCLK),
    .d(Y9phu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Kswpw6));  // ../RTL/cortexm0ds_logic.v(17825)
  AL_DFF Ktppw6_reg (
    .clk(HCLK),
    .d(Npshu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Ktppw6));  // ../RTL/cortexm0ds_logic.v(17544)
  AL_DFF Kwlpw6_reg (
    .clk(SWCLKTCK),
    .d(Tgxhu6),
    .reset(n5972),
    .set(1'b0),
    .q(Kwlpw6));  // ../RTL/cortexm0ds_logic.v(17396)
  AL_DFF Kxeax6_reg (
    .clk(DCLK),
    .d(Sdwhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Kxeax6));  // ../RTL/cortexm0ds_logic.v(18322)
  AL_DFF Kxhpw6_reg (
    .clk(SWCLKTCK),
    .d(Pndhu6),
    .reset(n5971),
    .set(1'b0),
    .q(Kxhpw6));  // ../RTL/cortexm0ds_logic.v(17166)
  AL_DFF Kzabx6_reg (
    .clk(SCLK),
    .d(Jeuhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Kzabx6));  // ../RTL/cortexm0ds_logic.v(19903)
  AL_DFF L03qw6_reg (
    .clk(SWCLKTCK),
    .d(Voxhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(L03qw6));  // ../RTL/cortexm0ds_logic.v(18015)
  AL_DFF L0ypw6_reg (
    .clk(SWCLKTCK),
    .d(Jwxhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(L0ypw6));  // ../RTL/cortexm0ds_logic.v(17857)
  AL_DFF L1bbx6_reg (
    .clk(HCLK),
    .d(Smuhu6),
    .reset(n5973),
    .set(1'b0),
    .q(L1bbx6));  // ../RTL/cortexm0ds_logic.v(19908)
  AL_DFF L2bax6_reg (
    .clk(DCLK),
    .d(Zsvhu6),
    .reset(n5974),
    .set(1'b0),
    .q(L2bax6));  // ../RTL/cortexm0ds_logic.v(18211)
  AL_DFF L3bbx6_reg (
    .clk(SCLK),
    .d(Jmthu6),
    .reset(n5973),
    .set(1'b0),
    .q(L3bbx6));  // ../RTL/cortexm0ds_logic.v(19914)
  AL_DFF L4lax6_reg (
    .clk(SCLK),
    .d(Wfphu6),
    .reset(1'b0),
    .set(n5973),
    .q(L4lax6));  // ../RTL/cortexm0ds_logic.v(18718)
  AL_DFF L5lpw6_reg (
    .clk(SWCLKTCK),
    .d(Zqxhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(L5lpw6));  // ../RTL/cortexm0ds_logic.v(17326)
  AL_DFF L6hax6_reg (
    .clk(HCLK),
    .d(Pnohu6),
    .reset(1'b0),
    .set(n5973),
    .q(L6hax6));  // ../RTL/cortexm0ds_logic.v(18465)
  AL_DFF L6lax6_reg (
    .clk(HCLK),
    .d(Xdohu6),
    .reset(1'b0),
    .set(n5973),
    .q(L6lax6));  // ../RTL/cortexm0ds_logic.v(18724)
  AL_DFF L8kax6_reg (
    .clk(HCLK),
    .d(Zeohu6),
    .reset(1'b0),
    .set(1'b0),
    .q(L8kax6));  // ../RTL/cortexm0ds_logic.v(18693)
  AL_DFF L8zax6_reg (
    .clk(HCLK),
    .d(E1uhu6),
    .reset(n5973),
    .set(1'b0),
    .q(L8zax6));  // ../RTL/cortexm0ds_logic.v(19083)
  AL_DFF L9bbx6_reg (
    .clk(DCLK),
    .d(Nephu6),
    .reset(1'b0),
    .set(1'b0),
    .q(L9bbx6));  // ../RTL/cortexm0ds_logic.v(19928)
  AL_DFF L9xax6_reg (
    .clk(HCLK),
    .d(Yiuhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(L9xax6));  // ../RTL/cortexm0ds_logic.v(18959)
  AL_DFF Lbbax6_reg (
    .clk(DCLK),
    .d(Lsvhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Lbbax6));  // ../RTL/cortexm0ds_logic.v(18222)
  AL_DFF Ldoax6_reg (
    .clk(HCLK),
    .d(O7thu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Ldoax6));  // ../RTL/cortexm0ds_logic.v(18793)
  AL_DFF Ldvpw6_reg (
    .clk(SWCLKTCK),
    .d(Uyxhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Ldvpw6));  // ../RTL/cortexm0ds_logic.v(17774)
  AL_DFF Ldwax6_reg (
    .clk(HCLK),
    .d(Rlrhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Ldwax6));  // ../RTL/cortexm0ds_logic.v(18938)
  AL_DFF Le2qw6_reg (
    .clk(DCLK),
    .d(F2xhu6),
    .reset(n5974),
    .set(1'b0),
    .q(Le2qw6));  // ../RTL/cortexm0ds_logic.v(17977)
  AL_DFF Lerpw6_reg (
    .clk(HCLK),
    .d(Gtohu6),
    .reset(1'b0),
    .set(n5973),
    .q(Lerpw6));  // ../RTL/cortexm0ds_logic.v(17611)
  AL_DFF Lfgbx6_reg (
    .clk(HCLK),
    .d(B3uhu6),
    .reset(n5973),
    .set(1'b0),
    .q(Lfgbx6));  // ../RTL/cortexm0ds_logic.v(20063)
  AL_DFF Lfppw6_reg (
    .clk(HCLK),
    .d(Kzrhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Lfppw6));  // ../RTL/cortexm0ds_logic.v(17537)
  AL_DFF Lfwax6_reg (
    .clk(HCLK),
    .d(Gcrhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Lfwax6));  // ../RTL/cortexm0ds_logic.v(18939)
  AL_DFF Lg1bx6_reg (
    .clk(SCLK),
    .d(Y2phu6),
    .reset(n5973),
    .set(1'b0),
    .q(Lg1bx6));  // ../RTL/cortexm0ds_logic.v(19317)
  AL_DFF Lg9bx6_reg (
    .clk(DCLK),
    .d(C5whu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Lg9bx6));  // ../RTL/cortexm0ds_logic.v(19815)
  AL_DFF Lgkax6_reg (
    .clk(HCLK),
    .d(Qfthu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Lgkax6));  // ../RTL/cortexm0ds_logic.v(18702)
  AL_DFF Lhbbx6_reg (
    .clk(SWCLKTCK),
    .d(Blxhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Lhbbx6));  // ../RTL/cortexm0ds_logic.v(19932)
  AL_DFF Lhppw6_reg (
    .clk(HCLK),
    .d(Cvrhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Lhppw6));  // ../RTL/cortexm0ds_logic.v(17538)
  AL_DFF Lhwax6_reg (
    .clk(HCLK),
    .d(R7rhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Lhwax6));  // ../RTL/cortexm0ds_logic.v(18940)
  AL_DFF Li2bx6_reg (
    .clk(SCLK),
    .d(G0phu6),
    .reset(n5973),
    .set(1'b0),
    .q(Li2bx6));  // ../RTL/cortexm0ds_logic.v(19425)
  AL_DFF Li7ax6_reg (
    .clk(SWCLKTCK),
    .d(Urxhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Li7ax6));  // ../RTL/cortexm0ds_logic.v(18099)
  AL_DFF Liabx6_reg (
    .clk(SWCLKTCK),
    .d(Wlxhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Liabx6));  // ../RTL/cortexm0ds_logic.v(19889)
  AL_DFF Ljcax6_reg (
    .clk(DCLK),
    .d(A4whu6),
    .reset(n5974),
    .set(1'b0),
    .q(Ljcax6));  // ../RTL/cortexm0ds_logic.v(18265)
  AL_DFF Ljppw6_reg (
    .clk(HCLK),
    .d(Sbrhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Ljppw6));  // ../RTL/cortexm0ds_logic.v(17539)
  AL_DFF Ljwax6_reg (
    .clk(HCLK),
    .d(C3rhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Ljwax6));  // ../RTL/cortexm0ds_logic.v(18941)
  AL_DFF Lk9ax6_reg (
    .clk(DCLK),
    .d(Zlvhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Lk9ax6));  // ../RTL/cortexm0ds_logic.v(18168)
  AL_DFF Lksax6_reg (
    .clk(HCLK),
    .d(A0thu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Lksax6));  // ../RTL/cortexm0ds_logic.v(18869)
  AL_DFF Llppw6_reg (
    .clk(HCLK),
    .d(D7rhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Llppw6));  // ../RTL/cortexm0ds_logic.v(17540)
  AL_DFF Llwax6_reg (
    .clk(HCLK),
    .d(Nyqhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Llwax6));  // ../RTL/cortexm0ds_logic.v(18942)
  AL_DFF Lmkbx6_reg (
    .clk(DCLK),
    .d(Pfphu6),
    .reset(n5974),
    .set(1'b0),
    .q(Lmkbx6));  // ../RTL/cortexm0ds_logic.v(20260)
  AL_DFF Ln0bx6_reg (
    .clk(HCLK),
    .d(Etuhu6),
    .reset(n5973),
    .set(1'b0),
    .q(Ln0bx6));  // ../RTL/cortexm0ds_logic.v(19233)
  AL_DFF Lnppw6_reg (
    .clk(HCLK),
    .d(Cbqhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Lnppw6));  // ../RTL/cortexm0ds_logic.v(17541)
  AL_DFF Lnwax6_reg (
    .clk(HCLK),
    .d(Ytqhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Lnwax6));  // ../RTL/cortexm0ds_logic.v(18943)
  AL_DFF Lp7ax6_reg (
    .clk(HCLK),
    .d(Xluhu6),
    .reset(n5973),
    .set(1'b0),
    .q(Lp7ax6));  // ../RTL/cortexm0ds_logic.v(18107)
  AL_DFF Lpppw6_reg (
    .clk(HCLK),
    .d(N6qhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Lpppw6));  // ../RTL/cortexm0ds_logic.v(17542)
  AL_DFF Lpwax6_reg (
    .clk(HCLK),
    .d(Jpqhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Lpwax6));  // ../RTL/cortexm0ds_logic.v(18944)
  AL_DFF Lqjpw6_reg (
    .clk(HCLK),
    .d(Hxohu6),
    .reset(1'b0),
    .set(n5973),
    .q(Lqjpw6));  // ../RTL/cortexm0ds_logic.v(17259)
  AL_DFF Lr9bx6_reg (
    .clk(SCLK),
    .d(T3phu6),
    .reset(n5973),
    .set(1'b0),
    .q(Lr9bx6));  // ../RTL/cortexm0ds_logic.v(19830)
  AL_DFF Lrppw6_reg (
    .clk(HCLK),
    .d(Zevhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Lrppw6));  // ../RTL/cortexm0ds_logic.v(17543)
  AL_DFF Lrwax6_reg (
    .clk(HCLK),
    .d(Fgqhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Lrwax6));  // ../RTL/cortexm0ds_logic.v(18945)
  AL_DFF Ltwax6_reg (
    .clk(HCLK),
    .d(Qbqhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Ltwax6));  // ../RTL/cortexm0ds_logic.v(18946)
  AL_DFF Lvwax6_reg (
    .clk(HCLK),
    .d(B7qhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Lvwax6));  // ../RTL/cortexm0ds_logic.v(18947)
  AL_DFF Lx9ax6_reg (
    .clk(DCLK),
    .d(Hjvhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Lx9ax6));  // ../RTL/cortexm0ds_logic.v(18175)
  AL_DFF Lxwax6_reg (
    .clk(HCLK),
    .d(Xxphu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Lxwax6));  // ../RTL/cortexm0ds_logic.v(18948)
  AL_DFF Lycax6_reg (
    .clk(DCLK),
    .d(Tvwhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Lycax6));  // ../RTL/cortexm0ds_logic.v(18274)
  AL_DFF Lywpw6_reg (
    .clk(HCLK),
    .d(Tjuhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Lywpw6));  // ../RTL/cortexm0ds_logic.v(17828)
  AL_DFF Lzwax6_reg (
    .clk(HCLK),
    .d(Mophu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Lzwax6));  // ../RTL/cortexm0ds_logic.v(18949)
  AL_DFF M13bx6_reg (
    .clk(SCLK),
    .d(Dqthu6),
    .reset(n5973),
    .set(1'b0),
    .q(M13bx6));  // ../RTL/cortexm0ds_logic.v(19479)
  AL_DFF M2ebx6_reg (
    .clk(HCLK),
    .d(Pdrhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(M2ebx6));  // ../RTL/cortexm0ds_logic.v(19986)
  AL_DFF M2lax6_reg (
    .clk(HCLK),
    .d(Sevhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(M2lax6));  // ../RTL/cortexm0ds_logic.v(18713)
  AL_DFF M3wax6_reg (
    .clk(HCLK),
    .d(C9shu6),
    .reset(1'b0),
    .set(1'b0),
    .q(M3wax6));  // ../RTL/cortexm0ds_logic.v(18933)
  AL_DFF M4ebx6_reg (
    .clk(DCLK),
    .d(Kovhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(M4ebx6));  // ../RTL/cortexm0ds_logic.v(19987)
  AL_DFF M5wax6_reg (
    .clk(HCLK),
    .d(N4shu6),
    .reset(1'b0),
    .set(1'b0),
    .q(M5wax6));  // ../RTL/cortexm0ds_logic.v(18934)
  AL_DFF M6cax6_reg (
    .clk(DCLK),
    .d(S6whu6),
    .reset(1'b0),
    .set(1'b0),
    .q(M6cax6));  // ../RTL/cortexm0ds_logic.v(18254)
  AL_DFF M6kax6_reg (
    .clk(HCLK),
    .d(Gfohu6),
    .reset(1'b0),
    .set(1'b0),
    .q(M6kax6));  // ../RTL/cortexm0ds_logic.v(18692)
  AL_DFF M6rpw6_reg (
    .clk(HCLK),
    .d(Jluhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(M6rpw6));  // ../RTL/cortexm0ds_logic.v(17598)
  AL_DFF M7wax6_reg (
    .clk(HCLK),
    .d(Yzrhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(M7wax6));  // ../RTL/cortexm0ds_logic.v(18935)
  AL_DFF M81qw6_reg (
    .clk(DCLK),
    .d(Qcphu6),
    .reset(1'b0),
    .set(1'b0),
    .q(M81qw6));  // ../RTL/cortexm0ds_logic.v(17936)
  AL_DFF M85bx6_reg (
    .clk(HCLK),
    .d(Fythu6),
    .reset(n5973),
    .set(1'b0),
    .q(M85bx6));  // ../RTL/cortexm0ds_logic.v(19707)
  AL_DFF M8fax6_reg (
    .clk(DCLK),
    .d(Czuhu6),
    .reset(n5974),
    .set(1'b0),
    .q(M8fax6));  // ../RTL/cortexm0ds_logic.v(18337)
  AL_DFF M8ipw6_reg (
    .clk(SWCLKTCK),
    .d(Jpxhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(M8ipw6));  // ../RTL/cortexm0ds_logic.v(17188)
  AL_DFF M9wax6_reg (
    .clk(HCLK),
    .d(Qvrhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(M9wax6));  // ../RTL/cortexm0ds_logic.v(18936)
  AL_DFF Mb4bx6_reg (
    .clk(HCLK),
    .d(Wwthu6),
    .reset(n5973),
    .set(1'b0),
    .q(Mb4bx6));  // ../RTL/cortexm0ds_logic.v(19611)
  AL_DFF Mbdax6_reg (
    .clk(DCLK),
    .d(Uswhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Mbdax6));  // ../RTL/cortexm0ds_logic.v(18281)
  AL_DFF Mboax6_reg (
    .clk(HCLK),
    .d(V7thu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Mboax6));  // ../RTL/cortexm0ds_logic.v(18792)
  AL_DFF Mbwax6_reg (
    .clk(HCLK),
    .d(Gqrhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Mbwax6));  // ../RTL/cortexm0ds_logic.v(18937)
  AL_DFF Mdppw6_reg (
    .clk(HCLK),
    .d(Omshu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Mdppw6));  // ../RTL/cortexm0ds_logic.v(17536)
  AL_DFF Mfyax6_reg (
    .clk(HCLK),
    .d(W3uhu6),
    .reset(n5973),
    .set(1'b0),
    .q(Mfyax6));  // ../RTL/cortexm0ds_logic.v(18999)
  AL_DFF Mgeax6_reg (
    .clk(DCLK),
    .d(Hiwhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Mgeax6));  // ../RTL/cortexm0ds_logic.v(18313)
  AL_DFF Mh1qw6_reg (
    .clk(DCLK),
    .d(Jcphu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Mh1qw6));  // ../RTL/cortexm0ds_logic.v(17941)
  AL_DFF Misax6_reg (
    .clk(HCLK),
    .d(H0thu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Misax6));  // ../RTL/cortexm0ds_logic.v(18868)
  AL_DFF Mjmpw6_reg (
    .clk(HCLK),
    .d(Wyrhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Mjmpw6));  // ../RTL/cortexm0ds_logic.v(17429)
  AL_DFF Mk3bx6_reg (
    .clk(SCLK),
    .d(A4phu6),
    .reset(n5973),
    .set(1'b0),
    .q(Mk3bx6));  // ../RTL/cortexm0ds_logic.v(19533)
  AL_DFF Mlmpw6_reg (
    .clk(HCLK),
    .d(O1shu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Mlmpw6));  // ../RTL/cortexm0ds_logic.v(17430)
  AL_DFF Mnmpw6_reg (
    .clk(HCLK),
    .d(Xmthu6),
    .reset(n5973),
    .set(1'b0),
    .q(Mnmpw6));  // ../RTL/cortexm0ds_logic.v(17435)
  AL_DFF Mp0bx6_reg (
    .clk(HCLK),
    .d(Stuhu6),
    .reset(n5973),
    .set(1'b0),
    .q(Mp0bx6));  // ../RTL/cortexm0ds_logic.v(19239)
  AL_DFF Ms5bx6_reg (
    .clk(HCLK),
    .d(Lirhu6),
    .reset(n5973),
    .set(1'b0),
    .q(Ms5bx6));  // ../RTL/cortexm0ds_logic.v(19727)
  AL_DFF Muhbx6_reg (
    .clk(SCLK),
    .d(O4phu6),
    .reset(n5973),
    .set(1'b0),
    .q(Muhbx6));  // ../RTL/cortexm0ds_logic.v(20144)
  AL_DFF Mw5bx6_reg (
    .clk(HCLK),
    .d(Jdohu6),
    .reset(1'b0),
    .set(n5973),
    .q(Mw5bx6));  // ../RTL/cortexm0ds_logic.v(19734)
  AL_DFF Mz1bx6_reg (
    .clk(SCLK),
    .d(Jsuhu6),
    .reset(n5973),
    .set(1'b0),
    .q(Mz1bx6));  // ../RTL/cortexm0ds_logic.v(19371)
  AL_DFF N0cbx6_reg (
    .clk(DCLK),
    .d(N7phu6),
    .reset(1'b0),
    .set(1'b0),
    .q(N0cbx6));  // ../RTL/cortexm0ds_logic.v(19942)
  AL_DFF N0lax6_reg (
    .clk(HCLK),
    .d(Eevhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(N0lax6));  // ../RTL/cortexm0ds_logic.v(18712)
  AL_DFF N0xpw6_reg (
    .clk(SCLK),
    .d(Bauhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(N0xpw6));  // ../RTL/cortexm0ds_logic.v(17829)
  AL_DFF N19bx6_reg (
    .clk(DCLK),
    .d(Newhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(N19bx6));  // ../RTL/cortexm0ds_logic.v(19807)
  AL_DFF N1oax6_reg (
    .clk(HCLK),
    .d(Tgqhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(N1oax6));  // ../RTL/cortexm0ds_logic.v(18787)
  AL_DFF N1wax6_reg (
    .clk(HCLK),
    .d(Ydshu6),
    .reset(1'b0),
    .set(1'b0),
    .q(N1wax6));  // ../RTL/cortexm0ds_logic.v(18932)
  AL_DFF N39ax6_reg (
    .clk(DCLK),
    .d(Jrvhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(N39ax6));  // ../RTL/cortexm0ds_logic.v(18159)
  AL_DFF N3eax6_reg (
    .clk(DCLK),
    .d(Nlwhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(N3eax6));  // ../RTL/cortexm0ds_logic.v(18301)
  AL_DFF N3hbx6_reg (
    .clk(DCLK),
    .d(Vpwhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(N3hbx6));  // ../RTL/cortexm0ds_logic.v(20101)
  AL_DFF N3jbx6_reg (
    .clk(DCLK),
    .d(Elvhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(N3jbx6));  // ../RTL/cortexm0ds_logic.v(20183)
  AL_DFF N3oax6_reg (
    .clk(HCLK),
    .d(Ecqhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(N3oax6));  // ../RTL/cortexm0ds_logic.v(18788)
  AL_DFF N4gax6_reg (
    .clk(DCLK),
    .d(W1whu6),
    .reset(1'b0),
    .set(1'b0),
    .q(N4gax6));  // ../RTL/cortexm0ds_logic.v(18400)
  AL_DFF N4kax6_reg (
    .clk(HCLK),
    .d(Djthu6),
    .reset(1'b0),
    .set(n5973),
    .q(N4kax6));  // ../RTL/cortexm0ds_logic.v(18690)
  AL_DFF N5bbx6_reg (
    .clk(SCLK),
    .d(V4phu6),
    .reset(n5973),
    .set(1'b0),
    .q(N5bbx6));  // ../RTL/cortexm0ds_logic.v(19920)
  AL_DFF N5oax6_reg (
    .clk(HCLK),
    .d(P7qhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(N5oax6));  // ../RTL/cortexm0ds_logic.v(18789)
  AL_DFF N61qw6_reg (
    .clk(HCLK),
    .d(Vpphu6),
    .reset(1'b0),
    .set(1'b0),
    .q(N61qw6));  // ../RTL/cortexm0ds_logic.v(17935)
  AL_DFF N7oax6_reg (
    .clk(HCLK),
    .d(Lyphu6),
    .reset(1'b0),
    .set(1'b0),
    .q(N7oax6));  // ../RTL/cortexm0ds_logic.v(18790)
  AL_DFF N7ppw6_reg (
    .clk(HCLK),
    .d(Q8thu6),
    .reset(1'b0),
    .set(1'b0),
    .q(N7ppw6));  // ../RTL/cortexm0ds_logic.v(17533)
  AL_DFF N8rpw6_reg (
    .clk(SCLK),
    .d(Xeuhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(N8rpw6));  // ../RTL/cortexm0ds_logic.v(17599)
  AL_DFF N9oax6_reg (
    .clk(HCLK),
    .d(Apphu6),
    .reset(1'b0),
    .set(1'b0),
    .q(N9oax6));  // ../RTL/cortexm0ds_logic.v(18791)
  AL_DFF N9ppw6_reg (
    .clk(HCLK),
    .d(J8thu6),
    .reset(1'b0),
    .set(1'b0),
    .q(N9ppw6));  // ../RTL/cortexm0ds_logic.v(17534)
  AL_DFF Naaax6_reg (
    .clk(DCLK),
    .d(Jyvhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Naaax6));  // ../RTL/cortexm0ds_logic.v(18182)
  AL_DFF Nazax6_reg (
    .clk(HCLK),
    .d(Q0uhu6),
    .reset(n5973),
    .set(1'b0),
    .q(Nazax6));  // ../RTL/cortexm0ds_logic.v(19089)
  AL_DFF Nbppw6_reg (
    .clk(HCLK),
    .d(Krshu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Nbppw6));  // ../RTL/cortexm0ds_logic.v(17535)
  AL_DFF Nbxax6_reg (
    .clk(SCLK),
    .d(Wauhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Nbxax6));  // ../RTL/cortexm0ds_logic.v(18960)
  AL_DFF Nckbx6_reg (
    .clk(DCLK),
    .d(Xcphu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Nckbx6));  // ../RTL/cortexm0ds_logic.v(20246)
  AL_DFF Nd3qw6_reg (
    .clk(DCLK),
    .d(B7xhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Nd3qw6));  // ../RTL/cortexm0ds_logic.v(18032)
  AL_DFF Nfgax6_reg (
    .clk(DCLK),
    .d(Hqvhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Nfgax6));  // ../RTL/cortexm0ds_logic.v(18406)
  AL_DFF Nfnax6_reg (
    .clk(HCLK),
    .d(Q9shu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Nfnax6));  // ../RTL/cortexm0ds_logic.v(18776)
  AL_DFF Nfqpw6_reg (
    .clk(SWCLKTCK),
    .d(F1yhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Nfqpw6));  // ../RTL/cortexm0ds_logic.v(17555)
  AL_DFF Ngsax6_reg (
    .clk(HCLK),
    .d(Pmphu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Ngsax6));  // ../RTL/cortexm0ds_logic.v(18867)
  AL_DFF Nhgbx6_reg (
    .clk(HCLK),
    .d(X0uhu6),
    .reset(n5973),
    .set(1'b0),
    .q(Nhgbx6));  // ../RTL/cortexm0ds_logic.v(20069)
  AL_DFF Nhnax6_reg (
    .clk(HCLK),
    .d(B5shu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Nhnax6));  // ../RTL/cortexm0ds_logic.v(18777)
  AL_DFF Ni5bx6_reg (
    .clk(HCLK),
    .d(F7shu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Ni5bx6));  // ../RTL/cortexm0ds_logic.v(19718)
  AL_DFF Nj2qw6_reg (
    .clk(DCLK),
    .d(E7vhu6),
    .reset(1'b0),
    .set(n5974),
    .q(Nj2qw6));  // ../RTL/cortexm0ds_logic.v(17995)
  AL_DFF Njnax6_reg (
    .clk(HCLK),
    .d(M0shu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Njnax6));  // ../RTL/cortexm0ds_logic.v(18778)
  AL_DFF Nk5bx6_reg (
    .clk(HCLK),
    .d(Q2shu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Nk5bx6));  // ../RTL/cortexm0ds_logic.v(19719)
  AL_DFF Nlbbx6_reg (
    .clk(DCLK),
    .d(Cyvhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Nlbbx6));  // ../RTL/cortexm0ds_logic.v(19934)
  AL_DFF Nlcbx6_reg (
    .clk(DCLK),
    .d(Haxhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Nlcbx6));  // ../RTL/cortexm0ds_logic.v(19953)
  AL_DFF Nlhax6_reg (
    .clk(HCLK),
    .d(Llohu6),
    .reset(1'b0),
    .set(n5973),
    .q(Nlhax6));  // ../RTL/cortexm0ds_logic.v(18513)
  AL_DFF Nlnax6_reg (
    .clk(HCLK),
    .d(Ewrhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Nlnax6));  // ../RTL/cortexm0ds_logic.v(18779)
  AL_DFF Nm5bx6_reg (
    .clk(HCLK),
    .d(Byrhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Nm5bx6));  // ../RTL/cortexm0ds_logic.v(19720)
  AL_DFF Nmabx6_reg (
    .clk(DCLK),
    .d(Hxvhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Nmabx6));  // ../RTL/cortexm0ds_logic.v(19891)
  AL_DFF Nmfax6_reg (
    .clk(SWCLKTCK),
    .d(Xpxhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Nmfax6));  // ../RTL/cortexm0ds_logic.v(18361)
  AL_DFF Nnfbx6_reg (
    .clk(DCLK),
    .d(K9whu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Nnfbx6));  // ../RTL/cortexm0ds_logic.v(20015)
  AL_DFF Nnnax6_reg (
    .clk(HCLK),
    .d(Fmrhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Nnnax6));  // ../RTL/cortexm0ds_logic.v(18780)
  AL_DFF No3qw6_reg (
    .clk(DCLK),
    .d(Vaxhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(No3qw6));  // ../RTL/cortexm0ds_logic.v(18044)
  AL_DFF No5bx6_reg (
    .clk(HCLK),
    .d(Ttrhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(No5bx6));  // ../RTL/cortexm0ds_logic.v(19721)
  AL_DFF Nodax6_reg (
    .clk(DCLK),
    .d(Towhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Nodax6));  // ../RTL/cortexm0ds_logic.v(18293)
  AL_DFF Npaax6_reg (
    .clk(DCLK),
    .d(Wuvhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Npaax6));  // ../RTL/cortexm0ds_logic.v(18190)
  AL_DFF Npnax6_reg (
    .clk(HCLK),
    .d(Ucrhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Npnax6));  // ../RTL/cortexm0ds_logic.v(18781)
  AL_DFF Npypw6_reg (
    .clk(HCLK),
    .d(Brrhu6),
    .reset(n5973),
    .set(1'b0),
    .q(Npypw6));  // ../RTL/cortexm0ds_logic.v(17889)
  AL_DFF Nq5bx6_reg (
    .clk(HCLK),
    .d(Corhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Nq5bx6));  // ../RTL/cortexm0ds_logic.v(19722)
  AL_DFF Nr0bx6_reg (
    .clk(HCLK),
    .d(Guuhu6),
    .reset(n5973),
    .set(1'b0),
    .q(Nr0bx6));  // ../RTL/cortexm0ds_logic.v(19245)
  AL_DFF Nr7ax6_reg (
    .clk(SCLK),
    .d(U9uhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Nr7ax6));  // ../RTL/cortexm0ds_logic.v(18109)
  AL_DFF Nrkpw6_reg (
    .clk(DCLK),
    .d(I8phu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Nrkpw6));  // ../RTL/cortexm0ds_logic.v(17309)
  AL_DFF Nrnax6_reg (
    .clk(HCLK),
    .d(F8rhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Nrnax6));  // ../RTL/cortexm0ds_logic.v(18782)
  AL_DFF Nrqpw6_reg (
    .clk(SWCLKTCK),
    .d(Eqxhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Nrqpw6));  // ../RTL/cortexm0ds_logic.v(17576)
  AL_DFF Ns8ax6_reg (
    .clk(SWCLKTCK),
    .d(Kmxhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Ns8ax6));  // ../RTL/cortexm0ds_logic.v(18133)
  AL_DFF Nt9bx6_reg (
    .clk(HCLK),
    .d(Bouhu6),
    .reset(n5973),
    .set(1'b0),
    .q(Nt9bx6));  // ../RTL/cortexm0ds_logic.v(19836)
  AL_DFF Ntnax6_reg (
    .clk(HCLK),
    .d(Q3rhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Ntnax6));  // ../RTL/cortexm0ds_logic.v(18783)
  AL_DFF Nu5bx6_reg (
    .clk(HCLK),
    .d(Irrhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Nu5bx6));  // ../RTL/cortexm0ds_logic.v(19729)
  AL_DFF Nv3qw6_reg (
    .clk(SWCLKTCK),
    .d(Vhxhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Nv3qw6));  // ../RTL/cortexm0ds_logic.v(18048)
  AL_DFF Nv9bx6_reg (
    .clk(HCLK),
    .d(Unuhu6),
    .reset(n5973),
    .set(1'b0),
    .q(Nv9bx6));  // ../RTL/cortexm0ds_logic.v(19842)
  AL_DFF Nvnax6_reg (
    .clk(HCLK),
    .d(Bzqhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Nvnax6));  // ../RTL/cortexm0ds_logic.v(18784)
  AL_DFF Nwbbx6_reg (
    .clk(HCLK),
    .d(Anrhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Nwbbx6));  // ../RTL/cortexm0ds_logic.v(19940)
  AL_DFF Nwdbx6_reg (
    .clk(DCLK),
    .d(Xbxhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Nwdbx6));  // ../RTL/cortexm0ds_logic.v(19983)
  AL_DFF Nxabx6_reg (
    .clk(HCLK),
    .d(Ocohu6),
    .reset(1'b0),
    .set(n5973),
    .q(Nxabx6));  // ../RTL/cortexm0ds_logic.v(19901)
  AL_DFF Nxnax6_reg (
    .clk(HCLK),
    .d(Muqhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Nxnax6));  // ../RTL/cortexm0ds_logic.v(18785)
  AL_DFF Nybbx6_reg (
    .clk(HCLK),
    .d(H1shu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Nybbx6));  // ../RTL/cortexm0ds_logic.v(19941)
  AL_DFF Nyhax6_reg (
    .clk(HCLK),
    .d(Ojohu6),
    .reset(1'b0),
    .set(n5973),
    .q(Nyhax6));  // ../RTL/cortexm0ds_logic.v(18555)
  AL_DFF Nyhpw6_reg (
    .clk(SWCLKTCK),
    .d(CDBGPWRUPACK),
    .reset(n5972),
    .set(1'b0),
    .q(Nyhpw6));  // ../RTL/cortexm0ds_logic.v(17172)
  AL_DFF Nznax6_reg (
    .clk(HCLK),
    .d(Xpqhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Nznax6));  // ../RTL/cortexm0ds_logic.v(18786)
  AL_DFF O0sax6_reg (
    .clk(HCLK),
    .d(Qwqhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(O0sax6));  // ../RTL/cortexm0ds_logic.v(18859)
  AL_DFF O1jbx6_reg (
    .clk(HCLK),
    .d(Duphu6),
    .reset(1'b0),
    .set(1'b0),
    .q(O1jbx6));  // ../RTL/cortexm0ds_logic.v(20182)
  AL_DFF O1mpw6_reg (
    .clk(SWCLKTCK),
    .d(Tnxhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(O1mpw6));  // ../RTL/cortexm0ds_logic.v(17405)
  AL_DFF O1ppw6_reg (
    .clk(HCLK),
    .d(Aaqhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(O1ppw6));  // ../RTL/cortexm0ds_logic.v(17530)
  AL_DFF O2kax6_reg (
    .clk(HCLK),
    .d(Nfohu6),
    .reset(1'b0),
    .set(1'b0),
    .q(O2kax6));  // ../RTL/cortexm0ds_logic.v(18685)
  AL_DFF O2sax6_reg (
    .clk(HCLK),
    .d(Bsqhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(O2sax6));  // ../RTL/cortexm0ds_logic.v(18860)
  AL_DFF O3ppw6_reg (
    .clk(HCLK),
    .d(L5qhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(O3ppw6));  // ../RTL/cortexm0ds_logic.v(17531)
  AL_DFF O41qw6_reg (
    .clk(HCLK),
    .d(Opphu6),
    .reset(1'b0),
    .set(1'b0),
    .q(O41qw6));  // ../RTL/cortexm0ds_logic.v(17934)
  AL_DFF O4hax6_reg (
    .clk(HCLK),
    .d(Wnohu6),
    .reset(1'b0),
    .set(n5973),
    .q(O4hax6));  // ../RTL/cortexm0ds_logic.v(18459)
  AL_DFF O4sax6_reg (
    .clk(HCLK),
    .d(Mnqhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(O4sax6));  // ../RTL/cortexm0ds_logic.v(18861)
  AL_DFF O5ppw6_reg (
    .clk(HCLK),
    .d(E9thu6),
    .reset(1'b0),
    .set(1'b0),
    .q(O5ppw6));  // ../RTL/cortexm0ds_logic.v(17532)
  AL_DFF O6sax6_reg (
    .clk(HCLK),
    .d(Ieqhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(O6sax6));  // ../RTL/cortexm0ds_logic.v(18862)
  AL_DFF O8sax6_reg (
    .clk(HCLK),
    .d(T9qhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(O8sax6));  // ../RTL/cortexm0ds_logic.v(18863)
  AL_DFF Oa5bx6_reg (
    .clk(HCLK),
    .d(Yxthu6),
    .reset(n5973),
    .set(1'b0),
    .q(Oa5bx6));  // ../RTL/cortexm0ds_logic.v(19713)
  AL_DFF Oarpw6_reg (
    .clk(SCLK),
    .d(Qeuhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Oarpw6));  // ../RTL/cortexm0ds_logic.v(17600)
  AL_DFF Oasax6_reg (
    .clk(HCLK),
    .d(E5qhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Oasax6));  // ../RTL/cortexm0ds_logic.v(18864)
  AL_DFF Ocsax6_reg (
    .clk(HCLK),
    .d(Awphu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Ocsax6));  // ../RTL/cortexm0ds_logic.v(18865)
  AL_DFF Od4bx6_reg (
    .clk(HCLK),
    .d(Iwthu6),
    .reset(n5973),
    .set(1'b0),
    .q(Od4bx6));  // ../RTL/cortexm0ds_logic.v(19617)
  AL_DFF Odnax6_reg (
    .clk(HCLK),
    .d(Meshu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Odnax6));  // ../RTL/cortexm0ds_logic.v(18775)
  AL_DFF Oesax6_reg (
    .clk(HCLK),
    .d(Erphu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Oesax6));  // ../RTL/cortexm0ds_logic.v(18866)
  AL_DFF Ofmpw6_reg (
    .clk(HCLK),
    .d(Whuhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Ofmpw6));  // ../RTL/cortexm0ds_logic.v(17422)
  AL_DFF Og5bx6_reg (
    .clk(HCLK),
    .d(Bcshu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Og5bx6));  // ../RTL/cortexm0ds_logic.v(19717)
  AL_DFF Oh8ax6_reg (
    .clk(SWCLKTCK),
    .d(Exxhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Oh8ax6));  // ../RTL/cortexm0ds_logic.v(18122)
  AL_DFF Ohyax6_reg (
    .clk(HCLK),
    .d(P3uhu6),
    .reset(n5973),
    .set(1'b0),
    .q(Ohyax6));  // ../RTL/cortexm0ds_logic.v(19005)
  AL_DFF Oi1bx6_reg (
    .clk(SCLK),
    .d(Nothu6),
    .reset(n5973),
    .set(1'b0),
    .q(Oi1bx6));  // ../RTL/cortexm0ds_logic.v(19323)
  AL_DFF Oi9ax6_reg (
    .clk(DCLK),
    .d(Gmvhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Oi9ax6));  // ../RTL/cortexm0ds_logic.v(18167)
  AL_DFF Oikax6_reg (
    .clk(HCLK),
    .d(Jfthu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Oikax6));  // ../RTL/cortexm0ds_logic.v(18703)
  AL_DFF Ojebx6_reg (
    .clk(SWCLKTCK),
    .d(Sjxhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Ojebx6));  // ../RTL/cortexm0ds_logic.v(19995)
  AL_DFF Ok2bx6_reg (
    .clk(SCLK),
    .d(Ppthu6),
    .reset(n5973),
    .set(1'b0),
    .q(Ok2bx6));  // ../RTL/cortexm0ds_logic.v(19431)
  AL_DFF Okfax6_reg (
    .clk(SWCLKTCK),
    .d(Isxhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Okfax6));  // ../RTL/cortexm0ds_logic.v(18360)
  AL_DFF Om3bx6_reg (
    .clk(SCLK),
    .d(Vsthu6),
    .reset(n5973),
    .set(1'b0),
    .q(Om3bx6));  // ../RTL/cortexm0ds_logic.v(19539)
  AL_DFF Onypw6_reg (
    .clk(HCLK),
    .d(Uqrhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Onypw6));  // ../RTL/cortexm0ds_logic.v(17884)
  AL_DFF Opbax6_reg (
    .clk(DCLK),
    .d(Vbwhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Opbax6));  // ../RTL/cortexm0ds_logic.v(18245)
  AL_DFF Osrax6_reg (
    .clk(HCLK),
    .d(Ujrhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Osrax6));  // ../RTL/cortexm0ds_logic.v(18855)
  AL_DFF Ot0bx6_reg (
    .clk(HCLK),
    .d(Wvuhu6),
    .reset(n5973),
    .set(1'b0),
    .q(Ot0bx6));  // ../RTL/cortexm0ds_logic.v(19251)
  AL_DFF Otopw6_reg (
    .clk(HCLK),
    .d(Iyrhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Otopw6));  // ../RTL/cortexm0ds_logic.v(17526)
  AL_DFF Oulpw6_reg (
    .clk(SWCLKTCK),
    .d(Sqxhu6),
    .reset(n5972),
    .set(1'b0),
    .q(Oulpw6));  // ../RTL/cortexm0ds_logic.v(17390)
  AL_DFF Ourax6_reg (
    .clk(HCLK),
    .d(Jarhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Ourax6));  // ../RTL/cortexm0ds_logic.v(18856)
  AL_DFF Oveax6_reg (
    .clk(DCLK),
    .d(Gewhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Oveax6));  // ../RTL/cortexm0ds_logic.v(18321)
  AL_DFF Ovopw6_reg (
    .clk(HCLK),
    .d(Aurhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Ovopw6));  // ../RTL/cortexm0ds_logic.v(17527)
  AL_DFF Owcax6_reg (
    .clk(DCLK),
    .d(Awwhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Owcax6));  // ../RTL/cortexm0ds_logic.v(18273)
  AL_DFF Owhbx6_reg (
    .clk(HCLK),
    .d(Zmuhu6),
    .reset(n5973),
    .set(1'b0),
    .q(Owhbx6));  // ../RTL/cortexm0ds_logic.v(20150)
  AL_DFF Owrax6_reg (
    .clk(HCLK),
    .d(U5rhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Owrax6));  // ../RTL/cortexm0ds_logic.v(18857)
  AL_DFF Ox9bx6_reg (
    .clk(HCLK),
    .d(Nguhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Ox9bx6));  // ../RTL/cortexm0ds_logic.v(19844)
  AL_DFF Oxkpw6_reg (
    .clk(HCLK),
    .d(Dwuhu6),
    .reset(n5973),
    .set(1'b0),
    .q(Oxkpw6));  // ../RTL/cortexm0ds_logic.v(17316)
  AL_DFF Oxopw6_reg (
    .clk(HCLK),
    .d(Qarhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Oxopw6));  // ../RTL/cortexm0ds_logic.v(17528)
  AL_DFF Oyhbx6_reg (
    .clk(HCLK),
    .d(Sfuhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Oyhbx6));  // ../RTL/cortexm0ds_logic.v(20152)
  AL_DFF Oykax6_reg (
    .clk(HCLK),
    .d(C8thu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Oykax6));  // ../RTL/cortexm0ds_logic.v(18711)
  AL_DFF Oyrax6_reg (
    .clk(HCLK),
    .d(F1rhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Oyrax6));  // ../RTL/cortexm0ds_logic.v(18858)
  AL_DFF Ozopw6_reg (
    .clk(HCLK),
    .d(B6rhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Ozopw6));  // ../RTL/cortexm0ds_logic.v(17529)
  AL_DFF Ozvax6_reg (
    .clk(HCLK),
    .d(Nishu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Ozvax6));  // ../RTL/cortexm0ds_logic.v(18931)
  AL_DFF P0bax6_reg (
    .clk(DCLK),
    .d(Gtvhu6),
    .reset(n5974),
    .set(1'b0),
    .q(P0bax6));  // ../RTL/cortexm0ds_logic.v(18205)
  AL_DFF P0ibx6_reg (
    .clk(SCLK),
    .d(Ceuhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(P0ibx6));  // ../RTL/cortexm0ds_logic.v(20153)
  AL_DFF P0kax6_reg (
    .clk(HCLK),
    .d(V5vhu6),
    .reset(1'b0),
    .set(n5973),
    .q(P0kax6));  // ../RTL/cortexm0ds_logic.v(18683)
  AL_DFF P12bx6_reg (
    .clk(SCLK),
    .d(B1phu6),
    .reset(n5973),
    .set(1'b0),
    .q(P12bx6));  // ../RTL/cortexm0ds_logic.v(19377)
  AL_DFF P14qw6_reg (
    .clk(HCLK),
    .d(Wgvhu6),
    .reset(1'b0),
    .set(n5973),
    .q(P14qw6));  // ../RTL/cortexm0ds_logic.v(18060)
  AL_DFF P21qw6_reg (
    .clk(HCLK),
    .d(Ynphu6),
    .reset(1'b0),
    .set(1'b0),
    .q(P21qw6));  // ../RTL/cortexm0ds_logic.v(17933)
  AL_DFF P23qw6_reg (
    .clk(DCLK),
    .d(D8xhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(P23qw6));  // ../RTL/cortexm0ds_logic.v(18016)
  AL_DFF P2xpw6_reg (
    .clk(HCLK),
    .d(Ovqhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(P2xpw6));  // ../RTL/cortexm0ds_logic.v(17830)
  AL_DFF P33bx6_reg (
    .clk(SCLK),
    .d(Ezohu6),
    .reset(n5973),
    .set(1'b0),
    .q(P33bx6));  // ../RTL/cortexm0ds_logic.v(19485)
  AL_DFF P34qw6_reg (
    .clk(HCLK),
    .d(Xushu6),
    .reset(1'b0),
    .set(1'b0),
    .q(P34qw6));  // ../RTL/cortexm0ds_logic.v(18062)
  AL_DFF P4cax6_reg (
    .clk(DCLK),
    .d(Z6whu6),
    .reset(1'b0),
    .set(1'b0),
    .q(P4cax6));  // ../RTL/cortexm0ds_logic.v(18253)
  AL_DFF P4xpw6_reg (
    .clk(HCLK),
    .d(Vvqhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(P4xpw6));  // ../RTL/cortexm0ds_logic.v(17831)
  AL_DFF P54qw6_reg (
    .clk(HCLK),
    .d(Dyshu6),
    .reset(1'b0),
    .set(1'b0),
    .q(P54qw6));  // ../RTL/cortexm0ds_logic.v(18063)
  AL_DFF P5vpw6_reg (
    .clk(HCLK),
    .d(Oqohu6),
    .reset(1'b0),
    .set(n5973),
    .q(P5vpw6));  // ../RTL/cortexm0ds_logic.v(17759)
  AL_DFF P6xpw6_reg (
    .clk(HCLK),
    .d(Xwqhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(P6xpw6));  // ../RTL/cortexm0ds_logic.v(17832)
  AL_DFF P7bbx6_reg (
    .clk(HCLK),
    .d(Hcohu6),
    .reset(1'b0),
    .set(n5973),
    .q(P7bbx6));  // ../RTL/cortexm0ds_logic.v(19926)
  AL_DFF P8xpw6_reg (
    .clk(HCLK),
    .d(Lxqhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(P8xpw6));  // ../RTL/cortexm0ds_logic.v(17833)
  AL_DFF P93qw6_reg (
    .clk(SWCLKTCK),
    .d(Ooxhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(P93qw6));  // ../RTL/cortexm0ds_logic.v(18025)
  AL_DFF P9bax6_reg (
    .clk(DCLK),
    .d(Esvhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(P9bax6));  // ../RTL/cortexm0ds_logic.v(18221)
  AL_DFF Paxpw6_reg (
    .clk(HCLK),
    .d(Zxqhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Paxpw6));  // ../RTL/cortexm0ds_logic.v(17834)
  AL_DFF Pbbbx6_reg (
    .clk(HCLK),
    .d(Hvqhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Pbbbx6));  // ../RTL/cortexm0ds_logic.v(19929)
  AL_DFF Pbnax6_reg (
    .clk(HCLK),
    .d(Bjshu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Pbnax6));  // ../RTL/cortexm0ds_logic.v(18774)
  AL_DFF Pcrpw6_reg (
    .clk(HCLK),
    .d(S0vhu6),
    .reset(1'b0),
    .set(n5973),
    .q(Pcrpw6));  // ../RTL/cortexm0ds_logic.v(17605)
  AL_DFF Pcxpw6_reg (
    .clk(HCLK),
    .d(Pzqhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Pcxpw6));  // ../RTL/cortexm0ds_logic.v(17835)
  AL_DFF Pczax6_reg (
    .clk(HCLK),
    .d(J0uhu6),
    .reset(n5973),
    .set(1'b0),
    .q(Pczax6));  // ../RTL/cortexm0ds_logic.v(19095)
  AL_DFF Pdbbx6_reg (
    .clk(DCLK),
    .d(Faphu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Pdbbx6));  // ../RTL/cortexm0ds_logic.v(19930)
  AL_DFF Pdmpw6_reg (
    .clk(HCLK),
    .d(Otshu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Pdmpw6));  // ../RTL/cortexm0ds_logic.v(17421)
  AL_DFF Pdxax6_reg (
    .clk(HCLK),
    .d(Riuhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Pdxax6));  // ../RTL/cortexm0ds_logic.v(18961)
  AL_DFF Pdyax6_reg (
    .clk(SCLK),
    .d(Npghu6),
    .reset(n5973),
    .set(1'b0),
    .q(Pdyax6));  // ../RTL/cortexm0ds_logic.v(18993)
  AL_DFF Pe5bx6_reg (
    .clk(HCLK),
    .d(Qgshu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Pe5bx6));  // ../RTL/cortexm0ds_logic.v(19716)
  AL_DFF Pe7ax6_reg (
    .clk(DCLK),
    .d(M2xhu6),
    .reset(n5974),
    .set(1'b0),
    .q(Pe7ax6));  // ../RTL/cortexm0ds_logic.v(18096)
  AL_DFF Pe9bx6_reg (
    .clk(DCLK),
    .d(Dvvhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Pe9bx6));  // ../RTL/cortexm0ds_logic.v(19814)
  AL_DFF Peeax6_reg (
    .clk(DCLK),
    .d(Jjwhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Peeax6));  // ../RTL/cortexm0ds_logic.v(18312)
  AL_DFF Pejbx6_reg (
    .clk(HCLK),
    .d(Lkphu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Pejbx6));  // ../RTL/cortexm0ds_logic.v(20189)
  AL_DFF Pexpw6_reg (
    .clk(DCLK),
    .d(Khvhu6),
    .reset(n5974),
    .set(1'b0),
    .q(Pexpw6));  // ../RTL/cortexm0ds_logic.v(17840)
  AL_DFF Pg3qw6_reg (
    .clk(DCLK),
    .d(W7xhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Pg3qw6));  // ../RTL/cortexm0ds_logic.v(18034)
  AL_DFF Pgjbx6_reg (
    .clk(SCLK),
    .d(Lnthu6),
    .reset(n5973),
    .set(1'b0),
    .q(Pgjbx6));  // ../RTL/cortexm0ds_logic.v(20194)
  AL_DFF Phcax6_reg (
    .clk(DCLK),
    .d(H4whu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Phcax6));  // ../RTL/cortexm0ds_logic.v(18260)
  AL_DFF Pifax6_reg (
    .clk(SWCLKTCK),
    .d(Avxhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Pifax6));  // ../RTL/cortexm0ds_logic.v(18359)
  AL_DFF Pjgbx6_reg (
    .clk(HCLK),
    .d(Tythu6),
    .reset(n5973),
    .set(1'b0),
    .q(Pjgbx6));  // ../RTL/cortexm0ds_logic.v(20075)
  AL_DFF Pkkbx6_reg (
    .clk(DCLK),
    .d(Ssvhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Pkkbx6));  // ../RTL/cortexm0ds_logic.v(20255)
  AL_DFF Plypw6_reg (
    .clk(HCLK),
    .d(Sprhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Plypw6));  // ../RTL/cortexm0ds_logic.v(17883)
  AL_DFF Pmlpw6_reg (
    .clk(SWCLKTCK),
    .d(Zehpw6[5]),
    .reset(n5972),
    .set(1'b0),
    .q(Pmlpw6));  // ../RTL/cortexm0ds_logic.v(17380)
  AL_DFF Pqrax6_reg (
    .clk(HCLK),
    .d(Jorhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Pqrax6));  // ../RTL/cortexm0ds_logic.v(18854)
  AL_DFF Propw6_reg (
    .clk(HCLK),
    .d(Mlshu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Propw6));  // ../RTL/cortexm0ds_logic.v(17525)
  AL_DFF Pt7ax6_reg (
    .clk(SCLK),
    .d(Ybuhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Pt7ax6));  // ../RTL/cortexm0ds_logic.v(18110)
  AL_DFF Puwpw6_reg (
    .clk(SWCLKTCK),
    .d(Nyxhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Puwpw6));  // ../RTL/cortexm0ds_logic.v(17826)
  AL_DFF Pv0bx6_reg (
    .clk(HCLK),
    .d(Kwuhu6),
    .reset(n5973),
    .set(1'b0),
    .q(Pv0bx6));  // ../RTL/cortexm0ds_logic.v(19257)
  AL_DFF Pv9ax6_reg (
    .clk(DCLK),
    .d(Ojvhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Pv9ax6));  // ../RTL/cortexm0ds_logic.v(18174)
  AL_DFF Pwkax6_reg (
    .clk(HCLK),
    .d(Ixshu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Pwkax6));  // ../RTL/cortexm0ds_logic.v(18710)
  AL_DFF Pxvax6_reg (
    .clk(HCLK),
    .d(Cnshu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Pxvax6));  // ../RTL/cortexm0ds_logic.v(18930)
  AL_DFF Pz9bx6_reg (
    .clk(HCLK),
    .d(L8uhu6),
    .reset(n5973),
    .set(1'b0),
    .q(Pz9bx6));  // ../RTL/cortexm0ds_logic.v(19849)
  AL_DFF Pzibx6_reg (
    .clk(HCLK),
    .d(Wtphu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Pzibx6));  // ../RTL/cortexm0ds_logic.v(20181)
  AL_DFF Pzkpw6_reg (
    .clk(HCLK),
    .d(Nfvhu6),
    .reset(1'b0),
    .set(n5973),
    .q(Pzkpw6));  // ../RTL/cortexm0ds_logic.v(17322)
  AL_DFF Q01qw6_reg (
    .clk(HCLK),
    .d(Knphu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Q01qw6));  // ../RTL/cortexm0ds_logic.v(17932)
  AL_DFF Q1hbx6_reg (
    .clk(DCLK),
    .d(Thwhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Q1hbx6));  // ../RTL/cortexm0ds_logic.v(20100)
  AL_DFF Q2gax6_reg (
    .clk(DCLK),
    .d(Crvhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Q2gax6));  // ../RTL/cortexm0ds_logic.v(18399)
  AL_DFF Q2ibx6_reg (
    .clk(DCLK),
    .d(Oaxhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Q2ibx6));  // ../RTL/cortexm0ds_logic.v(20154)
  AL_DFF Q4dbx6_reg (
    .clk(DCLK),
    .d(Aaxhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Q4dbx6));  // ../RTL/cortexm0ds_logic.v(19968)
  AL_DFF Q6fax6_reg (
    .clk(DCLK),
    .d(Ccwhu6),
    .reset(n5974),
    .set(1'b0),
    .q(Q6fax6));  // ../RTL/cortexm0ds_logic.v(18331)
  AL_DFF Q89bx6_reg (
    .clk(SWCLKTCK),
    .d(Aoxhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Q89bx6));  // ../RTL/cortexm0ds_logic.v(19811)
  AL_DFF Q8aax6_reg (
    .clk(DCLK),
    .d(Qyvhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Q8aax6));  // ../RTL/cortexm0ds_logic.v(18181)
  AL_DFF Q9dax6_reg (
    .clk(DCLK),
    .d(Btwhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Q9dax6));  // ../RTL/cortexm0ds_logic.v(18280)
  AL_DFF Q9nax6_reg (
    .clk(HCLK),
    .d(Qnshu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Q9nax6));  // ../RTL/cortexm0ds_logic.v(18773)
  AL_DFF Qa1qw6_reg (
    .clk(SWCLKTCK),
    .d(Vvxhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Qa1qw6));  // ../RTL/cortexm0ds_logic.v(17937)
  AL_DFF Qaipw6_reg (
    .clk(SCLK),
    .d(Sgthu6),
    .reset(n5973),
    .set(1'b0),
    .q(Qaipw6));  // ../RTL/cortexm0ds_logic.v(17193)
  AL_DFF Qakbx6_reg (
    .clk(HCLK),
    .d(Rqthu6),
    .reset(n5973),
    .set(1'b0),
    .q(Qakbx6));  // ../RTL/cortexm0ds_logic.v(20244)
  AL_DFF Qbmpw6_reg (
    .clk(HCLK),
    .d(Wqshu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Qbmpw6));  // ../RTL/cortexm0ds_logic.v(17420)
  AL_DFF Qc5bx6_reg (
    .clk(HCLK),
    .d(Loshu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Qc5bx6));  // ../RTL/cortexm0ds_logic.v(19715)
  AL_DFF Qehbx6_reg (
    .clk(DCLK),
    .d(Y8xhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Qehbx6));  // ../RTL/cortexm0ds_logic.v(20107)
  AL_DFF Qf4bx6_reg (
    .clk(HCLK),
    .d(Bwthu6),
    .reset(n5973),
    .set(1'b0),
    .q(Qf4bx6));  // ../RTL/cortexm0ds_logic.v(19623)
  AL_DFF Qhmpw6_reg (
    .clk(HCLK),
    .d(Mrthu6),
    .reset(n5973),
    .set(1'b0),
    .q(Qhmpw6));  // ../RTL/cortexm0ds_logic.v(17427)
  AL_DFF Qijpw6_reg (
    .clk(HCLK),
    .d(Bgvhu6),
    .reset(n5973),
    .set(1'b0),
    .q(Qijpw6));  // ../RTL/cortexm0ds_logic.v(17245)
  AL_DFF Qirax6_reg (
    .clk(HCLK),
    .d(Zashu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Qirax6));  // ../RTL/cortexm0ds_logic.v(18850)
  AL_DFF Qj1qw6_reg (
    .clk(SWCLKTCK),
    .d(Cwxhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Qj1qw6));  // ../RTL/cortexm0ds_logic.v(17942)
  AL_DFF Qjbbx6_reg (
    .clk(DCLK),
    .d(Invhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Qjbbx6));  // ../RTL/cortexm0ds_logic.v(19933)
  AL_DFF Qjcbx6_reg (
    .clk(DCLK),
    .d(Sywhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Qjcbx6));  // ../RTL/cortexm0ds_logic.v(19952)
  AL_DFF Qjhax6_reg (
    .clk(HCLK),
    .d(Slohu6),
    .reset(1'b0),
    .set(n5973),
    .q(Qjhax6));  // ../RTL/cortexm0ds_logic.v(18507)
  AL_DFF Qjyax6_reg (
    .clk(HCLK),
    .d(I3uhu6),
    .reset(n5973),
    .set(1'b0),
    .q(Qjyax6));  // ../RTL/cortexm0ds_logic.v(19011)
  AL_DFF Qjypw6_reg (
    .clk(HCLK),
    .d(Eprhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Qjypw6));  // ../RTL/cortexm0ds_logic.v(17882)
  AL_DFF Qkabx6_reg (
    .clk(DCLK),
    .d(Nmvhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Qkabx6));  // ../RTL/cortexm0ds_logic.v(19890)
  AL_DFF Qkrax6_reg (
    .clk(HCLK),
    .d(Rsrhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Qkrax6));  // ../RTL/cortexm0ds_logic.v(18851)
  AL_DFF Qlfbx6_reg (
    .clk(DCLK),
    .d(Lzvhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Qlfbx6));  // ../RTL/cortexm0ds_logic.v(20014)
  AL_DFF Qlopw6_reg (
    .clk(HCLK),
    .d(Qushu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Qlopw6));  // ../RTL/cortexm0ds_logic.v(17522)
  AL_DFF Qmdax6_reg (
    .clk(DCLK),
    .d(Cqwhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Qmdax6));  // ../RTL/cortexm0ds_logic.v(18292)
  AL_DFF Qmrax6_reg (
    .clk(HCLK),
    .d(Wrrhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Qmrax6));  // ../RTL/cortexm0ds_logic.v(18852)
  AL_DFF Qnopw6_reg (
    .clk(HCLK),
    .d(Jushu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Qnopw6));  // ../RTL/cortexm0ds_logic.v(17523)
  AL_DFF Qo3bx6_reg (
    .clk(SCLK),
    .d(M3phu6),
    .reset(n5973),
    .set(1'b0),
    .q(Qo3bx6));  // ../RTL/cortexm0ds_logic.v(19545)
  AL_DFF Qorax6_reg (
    .clk(HCLK),
    .d(Prrhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Qorax6));  // ../RTL/cortexm0ds_logic.v(18853)
  AL_DFF Qpopw6_reg (
    .clk(HCLK),
    .d(Iqshu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Qpopw6));  // ../RTL/cortexm0ds_logic.v(17524)
  AL_DFF Qsfax6_reg (
    .clk(DCLK),
    .d(Muxhu6),
    .reset(n5974),
    .set(1'b0),
    .q(Qsfax6));  // ../RTL/cortexm0ds_logic.v(18378)
  AL_DFF Qudbx6_reg (
    .clk(DCLK),
    .d(Cxwhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Qudbx6));  // ../RTL/cortexm0ds_logic.v(19982)
  AL_DFF Qufax6_reg (
    .clk(SWCLKTCK),
    .d(Dtnhu6),
    .reset(n5972),
    .set(1'b0),
    .q(Qufax6));  // ../RTL/cortexm0ds_logic.v(18384)
  AL_DFF Qukax6_reg (
    .clk(HCLK),
    .d(Cushu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Qukax6));  // ../RTL/cortexm0ds_logic.v(18709)
  AL_DFF Qvvax6_reg (
    .clk(HCLK),
    .d(Yrshu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Qvvax6));  // ../RTL/cortexm0ds_logic.v(18929)
  AL_DFF Qwfax6_reg (
    .clk(SWCLKTCK),
    .d(S3ohu6),
    .reset(n5972),
    .set(1'b0),
    .q(Qwfax6));  // ../RTL/cortexm0ds_logic.v(18390)
  AL_DFF Qwfbx6_reg (
    .clk(DCLK),
    .d(W8phu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Qwfbx6));  // ../RTL/cortexm0ds_logic.v(20020)
  AL_DFF Qx0bx6_reg (
    .clk(HCLK),
    .d(Ywuhu6),
    .reset(n5973),
    .set(1'b0),
    .q(Qx0bx6));  // ../RTL/cortexm0ds_logic.v(19263)
  AL_DFF Qxibx6_reg (
    .clk(HCLK),
    .d(Ptphu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Qxibx6));  // ../RTL/cortexm0ds_logic.v(20180)
  AL_DFF Qyjax6_reg (
    .clk(HCLK),
    .d(Ufohu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Qyjax6));  // ../RTL/cortexm0ds_logic.v(18678)
  AL_DFF Qynpw6_reg (
    .clk(SWCLKTCK),
    .d(Hvxhu6),
    .reset(n5972),
    .set(1'b0),
    .q(P13iu6));  // ../RTL/cortexm0ds_logic.v(17484)
  AL_DFF R19ax6_reg (
    .clk(DCLK),
    .d(L5xhu6),
    .reset(n5974),
    .set(1'b0),
    .q(R19ax6));  // ../RTL/cortexm0ds_logic.v(18157)
  AL_DFF R1abx6_reg (
    .clk(HCLK),
    .d(H6uhu6),
    .reset(n5973),
    .set(1'b0),
    .q(R1abx6));  // ../RTL/cortexm0ds_logic.v(19855)
  AL_DFF R1eax6_reg (
    .clk(DCLK),
    .d(Ulwhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(R1eax6));  // ../RTL/cortexm0ds_logic.v(18300)
  AL_DFF R2hax6_reg (
    .clk(HCLK),
    .d(Doohu6),
    .reset(1'b0),
    .set(n5973),
    .q(R2hax6));  // ../RTL/cortexm0ds_logic.v(18453)
  AL_DFF R3vpw6_reg (
    .clk(HCLK),
    .d(Vqohu6),
    .reset(n5973),
    .set(1'b0),
    .q(R3vpw6));  // ../RTL/cortexm0ds_logic.v(17753)
  AL_DFF R7ibx6_reg (
    .clk(HCLK),
    .d(Fhphu6),
    .reset(1'b0),
    .set(1'b0),
    .q(R7ibx6));  // ../RTL/cortexm0ds_logic.v(20167)
  AL_DFF R7kpw6_reg (
    .clk(HCLK),
    .d(Kiuhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(R7kpw6));  // ../RTL/cortexm0ds_logic.v(17289)
  AL_DFF R7nax6_reg (
    .clk(HCLK),
    .d(Msshu6),
    .reset(1'b0),
    .set(1'b0),
    .q(R7nax6));  // ../RTL/cortexm0ds_logic.v(18772)
  AL_DFF R9ibx6_reg (
    .clk(HCLK),
    .d(Mhphu6),
    .reset(1'b0),
    .set(1'b0),
    .q(R9ibx6));  // ../RTL/cortexm0ds_logic.v(20168)
  AL_DFF R9mpw6_reg (
    .clk(HCLK),
    .d(L7vhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(R9mpw6));  // ../RTL/cortexm0ds_logic.v(17419)
  AL_DFF R9yax6_reg (
    .clk(HCLK),
    .d(Mbvhu6),
    .reset(n5973),
    .set(1'b0),
    .q(R9yax6));  // ../RTL/cortexm0ds_logic.v(18981)
  AL_DFF Ra2qw6_reg (
    .clk(SWCLKTCK),
    .d(Ohxhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Ra2qw6));  // ../RTL/cortexm0ds_logic.v(17971)
  AL_DFF Rbibx6_reg (
    .clk(HCLK),
    .d(Thphu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Rbibx6));  // ../RTL/cortexm0ds_logic.v(20169)
  AL_DFF Rdibx6_reg (
    .clk(HCLK),
    .d(Aiphu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Rdibx6));  // ../RTL/cortexm0ds_logic.v(20170)
  AL_DFF Rdkpw6_reg (
    .clk(HCLK),
    .d(Ebrhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Rdkpw6));  // ../RTL/cortexm0ds_logic.v(17297)
  AL_DFF Rekbx6_reg (
    .clk(HCLK),
    .d(Yaohu6),
    .reset(n5973),
    .set(1'b0),
    .q(Rekbx6));  // ../RTL/cortexm0ds_logic.v(20251)
  AL_DFF Rezax6_reg (
    .clk(HCLK),
    .d(C0uhu6),
    .reset(n5973),
    .set(1'b0),
    .q(Rezax6));  // ../RTL/cortexm0ds_logic.v(19101)
  AL_DFF Rfibx6_reg (
    .clk(HCLK),
    .d(Hiphu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Rfibx6));  // ../RTL/cortexm0ds_logic.v(20171)
  AL_DFF Rfkpw6_reg (
    .clk(HCLK),
    .d(Idrhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Rfkpw6));  // ../RTL/cortexm0ds_logic.v(17298)
  AL_DFF Rfxax6_reg (
    .clk(SCLK),
    .d(Dbuhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Rfxax6));  // ../RTL/cortexm0ds_logic.v(18962)
  AL_DFF Rg9ax6_reg (
    .clk(DCLK),
    .d(Umvhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Rg9ax6));  // ../RTL/cortexm0ds_logic.v(18166)
  AL_DFF Rgrax6_reg (
    .clk(HCLK),
    .d(Zoshu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Rgrax6));  // ../RTL/cortexm0ds_logic.v(18849)
  AL_DFF Rhibx6_reg (
    .clk(HCLK),
    .d(Viphu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Rhibx6));  // ../RTL/cortexm0ds_logic.v(20172)
  AL_DFF Rhkpw6_reg (
    .clk(HCLK),
    .d(Okuhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Rhkpw6));  // ../RTL/cortexm0ds_logic.v(17299)
  AL_DFF Rhypw6_reg (
    .clk(HCLK),
    .d(Qorhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Rhypw6));  // ../RTL/cortexm0ds_logic.v(17881)
  AL_DFF Rijbx6_reg (
    .clk(SCLK),
    .d(Uwdpw6),
    .reset(n5973),
    .set(1'b0),
    .q(Rijbx6));  // ../RTL/cortexm0ds_logic.v(20200)
  AL_DFF Rilpw6_reg (
    .clk(SWCLKTCK),
    .d(Ovxhu6),
    .reset(1'b0),
    .set(n5972),
    .q(Rilpw6));  // ../RTL/cortexm0ds_logic.v(17368)
  AL_DFF Rjibx6_reg (
    .clk(HCLK),
    .d(Cjphu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Rjibx6));  // ../RTL/cortexm0ds_logic.v(20173)
  AL_DFF Rjopw6_reg (
    .clk(HCLK),
    .d(Evshu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Rjopw6));  // ../RTL/cortexm0ds_logic.v(17521)
  AL_DFF Rk1bx6_reg (
    .clk(SCLK),
    .d(K2phu6),
    .reset(n5973),
    .set(1'b0),
    .q(Rk1bx6));  // ../RTL/cortexm0ds_logic.v(19329)
  AL_DFF Rkbax6_reg (
    .clk(DCLK),
    .d(Ifphu6),
    .reset(n5974),
    .set(1'b0),
    .q(Rkbax6));  // ../RTL/cortexm0ds_logic.v(18231)
  AL_DFF Rkkax6_reg (
    .clk(HCLK),
    .d(Cfthu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Rkkax6));  // ../RTL/cortexm0ds_logic.v(18704)
  AL_DFF Rlgbx6_reg (
    .clk(HCLK),
    .d(Pwthu6),
    .reset(n5973),
    .set(1'b0),
    .q(Rlgbx6));  // ../RTL/cortexm0ds_logic.v(20081)
  AL_DFF Rlibx6_reg (
    .clk(HCLK),
    .d(Jjphu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Rlibx6));  // ../RTL/cortexm0ds_logic.v(20174)
  AL_DFF Rm2bx6_reg (
    .clk(SCLK),
    .d(Gwdpw6),
    .reset(n5973),
    .set(1'b0),
    .q(Rm2bx6));  // ../RTL/cortexm0ds_logic.v(19437)
  AL_DFF Rnaax6_reg (
    .clk(DCLK),
    .d(Kvvhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Rnaax6));  // ../RTL/cortexm0ds_logic.v(18189)
  AL_DFF Rnibx6_reg (
    .clk(HCLK),
    .d(Qjphu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Rnibx6));  // ../RTL/cortexm0ds_logic.v(20175)
  AL_DFF Rnvax6_reg (
    .clk(HCLK),
    .d(R5thu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Rnvax6));  // ../RTL/cortexm0ds_logic.v(18925)
  AL_DFF Ro8ax6_reg (
    .clk(DCLK),
    .d(Obphu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Ro8ax6));  // ../RTL/cortexm0ds_logic.v(18131)
  AL_DFF Rpibx6_reg (
    .clk(HCLK),
    .d(Xjphu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Rpibx6));  // ../RTL/cortexm0ds_logic.v(20176)
  AL_DFF Rpvax6_reg (
    .clk(HCLK),
    .d(K5thu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Rpvax6));  // ../RTL/cortexm0ds_logic.v(18926)
  AL_DFF Rq0qw6_reg (
    .clk(HCLK),
    .d(Bhuhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Rq0qw6));  // ../RTL/cortexm0ds_logic.v(17927)
  AL_DFF Rr3qw6_reg (
    .clk(DCLK),
    .d(Z6phu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Rr3qw6));  // ../RTL/cortexm0ds_logic.v(18046)
  AL_DFF Rribx6_reg (
    .clk(HCLK),
    .d(Ekphu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Rribx6));  // ../RTL/cortexm0ds_logic.v(20177)
  AL_DFF Rrvax6_reg (
    .clk(HCLK),
    .d(D5thu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Rrvax6));  // ../RTL/cortexm0ds_logic.v(18927)
  AL_DFF Rskax6_reg (
    .clk(HCLK),
    .d(Oethu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Rskax6));  // ../RTL/cortexm0ds_logic.v(18708)
  AL_DFF Rteax6_reg (
    .clk(DCLK),
    .d(Uewhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Rteax6));  // ../RTL/cortexm0ds_logic.v(18320)
  AL_DFF Rtibx6_reg (
    .clk(HCLK),
    .d(Skphu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Rtibx6));  // ../RTL/cortexm0ds_logic.v(20178)
  AL_DFF Rtvax6_reg (
    .clk(HCLK),
    .d(W4thu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Rtvax6));  // ../RTL/cortexm0ds_logic.v(18928)
  AL_DFF Rucax6_reg (
    .clk(DCLK),
    .d(Owwhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Rucax6));  // ../RTL/cortexm0ds_logic.v(18272)
  AL_DFF Rv7ax6_reg (
    .clk(SCLK),
    .d(Hduhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Rv7ax6));  // ../RTL/cortexm0ds_logic.v(18111)
  AL_DFF Rvibx6_reg (
    .clk(HCLK),
    .d(Itphu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Rvibx6));  // ../RTL/cortexm0ds_logic.v(20179)
  AL_DFF Rwhax6_reg (
    .clk(HCLK),
    .d(Vjohu6),
    .reset(1'b0),
    .set(n5973),
    .q(Rwhax6));  // ../RTL/cortexm0ds_logic.v(18549)
  AL_DFF Rwjax6_reg (
    .clk(HCLK),
    .d(Jzuhu6),
    .reset(1'b0),
    .set(n5973),
    .q(Rwjax6));  // ../RTL/cortexm0ds_logic.v(18676)
  AL_DFF Ry0qw6_reg (
    .clk(HCLK),
    .d(Wmphu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Ry0qw6));  // ../RTL/cortexm0ds_logic.v(17931)
  AL_DFF Ry2qw6_reg (
    .clk(SWCLKTCK),
    .d(J3yhu6),
    .reset(n5972),
    .set(1'b0),
    .q(Ry2qw6));  // ../RTL/cortexm0ds_logic.v(18013)
  AL_DFF Ryfax6_reg (
    .clk(SWCLKTCK),
    .d(Rtxhu6),
    .reset(n5972),
    .set(1'b0),
    .q(Ryfax6));  // ../RTL/cortexm0ds_logic.v(18396)
  AL_DFF Rz0bx6_reg (
    .clk(HCLK),
    .d(Ayuhu6),
    .reset(n5973),
    .set(1'b0),
    .q(Rz0bx6));  // ../RTL/cortexm0ds_logic.v(19269)
  AL_DFF Rz8bx6_reg (
    .clk(DCLK),
    .d(L6whu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Rz8bx6));  // ../RTL/cortexm0ds_logic.v(19806)
  AL_DFF S0kbx6_reg (
    .clk(HCLK),
    .d(Acvhu6),
    .reset(n5973),
    .set(1'b0),
    .q(S0kbx6));  // ../RTL/cortexm0ds_logic.v(20219)
  AL_DFF S11bx6_reg (
    .clk(SCLK),
    .d(Mivhu6),
    .reset(n5973),
    .set(1'b0),
    .q(S11bx6));  // ../RTL/cortexm0ds_logic.v(19275)
  AL_DFF S18ax6_reg (
    .clk(HCLK),
    .d(Peqhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(S18ax6));  // ../RTL/cortexm0ds_logic.v(18114)
  AL_DFF S1nax6_reg (
    .clk(HCLK),
    .d(C1thu6),
    .reset(1'b0),
    .set(1'b0),
    .q(S1nax6));  // ../RTL/cortexm0ds_logic.v(18769)
  AL_DFF S2cax6_reg (
    .clk(DCLK),
    .d(N7whu6),
    .reset(1'b0),
    .set(1'b0),
    .q(S2cax6));  // ../RTL/cortexm0ds_logic.v(18252)
  AL_DFF S2cbx6_reg (
    .clk(SWCLKTCK),
    .d(Y0yhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(S2cbx6));  // ../RTL/cortexm0ds_logic.v(19943)
  AL_DFF S32bx6_reg (
    .clk(SCLK),
    .d(Xsuhu6),
    .reset(n5973),
    .set(1'b0),
    .q(S32bx6));  // ../RTL/cortexm0ds_logic.v(19383)
  AL_DFF S38ax6_reg (
    .clk(HCLK),
    .d(Dfqhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(S38ax6));  // ../RTL/cortexm0ds_logic.v(18115)
  AL_DFF S3mpw6_reg (
    .clk(HCLK),
    .d(Gvthu6),
    .reset(n5973),
    .set(1'b0),
    .q(S3mpw6));  // ../RTL/cortexm0ds_logic.v(17410)
  AL_DFF S3nax6_reg (
    .clk(HCLK),
    .d(V0thu6),
    .reset(1'b0),
    .set(1'b0),
    .q(S3nax6));  // ../RTL/cortexm0ds_logic.v(18770)
  AL_DFF S4kbx6_reg (
    .clk(HCLK),
    .d(Levhu6),
    .reset(n5973),
    .set(1'b0),
    .q(S4kbx6));  // ../RTL/cortexm0ds_logic.v(20231)
  AL_DFF S53bx6_reg (
    .clk(SCLK),
    .d(Kqthu6),
    .reset(n5973),
    .set(1'b0),
    .q(S53bx6));  // ../RTL/cortexm0ds_logic.v(19491)
  AL_DFF S58ax6_reg (
    .clk(HCLK),
    .d(Rfqhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(S58ax6));  // ../RTL/cortexm0ds_logic.v(18116)
  AL_DFF S5kpw6_reg (
    .clk(HCLK),
    .d(Soshu6),
    .reset(1'b0),
    .set(1'b0),
    .q(S5kpw6));  // ../RTL/cortexm0ds_logic.v(17288)
  AL_DFF S5nax6_reg (
    .clk(HCLK),
    .d(O0thu6),
    .reset(1'b0),
    .set(1'b0),
    .q(S5nax6));  // ../RTL/cortexm0ds_logic.v(18771)
  AL_DFF S78ax6_reg (
    .clk(HCLK),
    .d(Ahqhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(S78ax6));  // ../RTL/cortexm0ds_logic.v(18117)
  AL_DFF S7mpw6_reg (
    .clk(HCLK),
    .d(Nhthu6),
    .reset(1'b0),
    .set(n5973),
    .q(S7mpw6));  // ../RTL/cortexm0ds_logic.v(17417)
  AL_DFF S7yax6_reg (
    .clk(HCLK),
    .d(Flshu6),
    .reset(1'b0),
    .set(1'b0),
    .q(S7yax6));  // ../RTL/cortexm0ds_logic.v(18976)
  AL_DFF S98ax6_reg (
    .clk(HCLK),
    .d(Hhqhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(S98ax6));  // ../RTL/cortexm0ds_logic.v(18118)
  AL_DFF Sb8ax6_reg (
    .clk(HCLK),
    .d(Ohqhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Sb8ax6));  // ../RTL/cortexm0ds_logic.v(18119)
  AL_DFF Sbfax6_reg (
    .clk(DCLK),
    .d(R1xhu6),
    .reset(n5974),
    .set(1'b0),
    .q(Sbfax6));  // ../RTL/cortexm0ds_logic.v(18349)
  AL_DFF Sbyax6_reg (
    .clk(SCLK),
    .d(Yqthu6),
    .reset(n5973),
    .set(1'b0),
    .q(Sbyax6));  // ../RTL/cortexm0ds_logic.v(18987)
  AL_DFF Sd8ax6_reg (
    .clk(DCLK),
    .d(Abphu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Sd8ax6));  // ../RTL/cortexm0ds_logic.v(18120)
  AL_DFF Sddbx6_reg (
    .clk(SWCLKTCK),
    .d(Izxhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Sddbx6));  // ../RTL/cortexm0ds_logic.v(19973)
  AL_DFF Sdlpw6_reg (
    .clk(SWCLKTCK),
    .d(Zehpw6[1]),
    .reset(1'b0),
    .set(n5972),
    .q(Sdlpw6));  // ../RTL/cortexm0ds_logic.v(17350)
  AL_DFF Sejax6_reg (
    .clk(HCLK),
    .d(Khohu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Sejax6));  // ../RTL/cortexm0ds_logic.v(18648)
  AL_DFF Serax6_reg (
    .clk(HCLK),
    .d(Vtshu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Serax6));  // ../RTL/cortexm0ds_logic.v(18848)
  AL_DFF Sfypw6_reg (
    .clk(HCLK),
    .d(Onrhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Sfypw6));  // ../RTL/cortexm0ds_logic.v(17880)
  AL_DFF Sgjax6_reg (
    .clk(HCLK),
    .d(Dhohu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Sgjax6));  // ../RTL/cortexm0ds_logic.v(18649)
  AL_DFF Sh4bx6_reg (
    .clk(HCLK),
    .d(Uvthu6),
    .reset(n5973),
    .set(1'b0),
    .q(Sh4bx6));  // ../RTL/cortexm0ds_logic.v(19629)
  AL_DFF Shopw6_reg (
    .clk(HCLK),
    .d(Ntohu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Shopw6));  // ../RTL/cortexm0ds_logic.v(17520)
  AL_DFF Sijax6_reg (
    .clk(HCLK),
    .d(Wgohu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Sijax6));  // ../RTL/cortexm0ds_logic.v(18650)
  AL_DFF Skjax6_reg (
    .clk(HCLK),
    .d(E0vhu6),
    .reset(1'b0),
    .set(n5973),
    .q(Skjax6));  // ../RTL/cortexm0ds_logic.v(18655)
  AL_DFF Slvax6_reg (
    .clk(HCLK),
    .d(Y5thu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Slvax6));  // ../RTL/cortexm0ds_logic.v(18924)
  AL_DFF Slyax6_reg (
    .clk(HCLK),
    .d(U2uhu6),
    .reset(n5973),
    .set(1'b0),
    .q(Slyax6));  // ../RTL/cortexm0ds_logic.v(19017)
  AL_DFF Smjax6_reg (
    .clk(HCLK),
    .d(Pgohu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Smjax6));  // ../RTL/cortexm0ds_logic.v(18657)
  AL_DFF Sn4bx6_reg (
    .clk(HCLK),
    .d(E8uhu6),
    .reset(n5973),
    .set(1'b0),
    .q(Sn4bx6));  // ../RTL/cortexm0ds_logic.v(19647)
  AL_DFF So0qw6_reg (
    .clk(HCLK),
    .d(Hpphu6),
    .reset(1'b0),
    .set(1'b0),
    .q(So0qw6));  // ../RTL/cortexm0ds_logic.v(17926)
  AL_DFF Sojax6_reg (
    .clk(HCLK),
    .d(Xzuhu6),
    .reset(1'b0),
    .set(n5973),
    .q(Sojax6));  // ../RTL/cortexm0ds_logic.v(18662)
  AL_DFF Sq3bx6_reg (
    .clk(SCLK),
    .d(Enthu6),
    .reset(n5973),
    .set(1'b0),
    .q(Sq3bx6));  // ../RTL/cortexm0ds_logic.v(19551)
  AL_DFF Sqfax6_reg (
    .clk(DCLK),
    .d(Pkhpw6[0]),
    .reset(n5974),
    .set(1'b0),
    .q(Sqfax6));  // ../RTL/cortexm0ds_logic.v(18372)
  AL_DFF Sqjax6_reg (
    .clk(HCLK),
    .d(Igohu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Sqjax6));  // ../RTL/cortexm0ds_logic.v(18664)
  AL_DFF Sqkax6_reg (
    .clk(HCLK),
    .d(Pgvhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Sqkax6));  // ../RTL/cortexm0ds_logic.v(18707)
  AL_DFF Sqwpw6_reg (
    .clk(DCLK),
    .d(O3xhu6),
    .reset(n5974),
    .set(1'b0),
    .q(Sqwpw6));  // ../RTL/cortexm0ds_logic.v(17823)
  AL_DFF Ss0qw6_reg (
    .clk(SCLK),
    .d(Tcuhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Ss0qw6));  // ../RTL/cortexm0ds_logic.v(17928)
  AL_DFF Ssjax6_reg (
    .clk(HCLK),
    .d(Qzuhu6),
    .reset(1'b0),
    .set(n5973),
    .q(Ssjax6));  // ../RTL/cortexm0ds_logic.v(18669)
  AL_DFF Stkpw6_reg (
    .clk(SWCLKTCK),
    .d(D0yhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Stkpw6));  // ../RTL/cortexm0ds_logic.v(17310)
  AL_DFF Su8ax6_reg (
    .clk(DCLK),
    .d(Bexhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Su8ax6));  // ../RTL/cortexm0ds_logic.v(18134)
  AL_DFF Sujax6_reg (
    .clk(HCLK),
    .d(Bgohu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Sujax6));  // ../RTL/cortexm0ds_logic.v(18671)
  AL_DFF Sw0qw6_reg (
    .clk(HCLK),
    .d(Ulphu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Sw0qw6));  // ../RTL/cortexm0ds_logic.v(17930)
  AL_DFF Swjbx6_reg (
    .clk(HCLK),
    .d(Fbohu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Swjbx6));  // ../RTL/cortexm0ds_logic.v(20213)
  AL_DFF Sx3qw6_reg (
    .clk(HCLK),
    .d(Ufvhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Sx3qw6));  // ../RTL/cortexm0ds_logic.v(18049)
  AL_DFF Sx7ax6_reg (
    .clk(HCLK),
    .d(Gdqhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Sx7ax6));  // ../RTL/cortexm0ds_logic.v(18112)
  AL_DFF Syjbx6_reg (
    .clk(HCLK),
    .d(Wzqhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Syjbx6));  // ../RTL/cortexm0ds_logic.v(20214)
  AL_DFF Sz3qw6_reg (
    .clk(HCLK),
    .d(Yoohu6),
    .reset(1'b0),
    .set(n5973),
    .q(Sz3qw6));  // ../RTL/cortexm0ds_logic.v(18054)
  AL_DFF Sz7ax6_reg (
    .clk(HCLK),
    .d(Ndqhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Sz7ax6));  // ../RTL/cortexm0ds_logic.v(18113)
  AL_DFF Szmax6_reg (
    .clk(HCLK),
    .d(J1thu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Szmax6));  // ../RTL/cortexm0ds_logic.v(18768)
  AL_DFF T00qw6_reg (
    .clk(HCLK),
    .d(T0shu6),
    .reset(1'b0),
    .set(1'b0),
    .q(T00qw6));  // ../RTL/cortexm0ds_logic.v(17914)
  AL_DFF T0ipw6_reg (
    .clk(SWCLKTCK),
    .d(O5ohu6),
    .reset(n5972),
    .set(1'b0),
    .q(T0ipw6));  // ../RTL/cortexm0ds_logic.v(17178)
  AL_DFF T1fbx6_reg (
    .clk(HCLK),
    .d(Tfrhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(T1fbx6));  // ../RTL/cortexm0ds_logic.v(20004)
  AL_DFF T1vpw6_reg (
    .clk(HCLK),
    .d(Crohu6),
    .reset(n5973),
    .set(1'b0),
    .q(T1vpw6));  // ../RTL/cortexm0ds_logic.v(17747)
  AL_DFF T20qw6_reg (
    .clk(HCLK),
    .d(Lwrhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(T20qw6));  // ../RTL/cortexm0ds_logic.v(17915)
  AL_DFF T2dbx6_reg (
    .clk(DCLK),
    .d(Zywhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(T2dbx6));  // ../RTL/cortexm0ds_logic.v(19967)
  AL_DFF T2kbx6_reg (
    .clk(SCLK),
    .d(Kjthu6),
    .reset(n5973),
    .set(1'b0),
    .q(T2kbx6));  // ../RTL/cortexm0ds_logic.v(20225)
  AL_DFF T3abx6_reg (
    .clk(HCLK),
    .d(D4uhu6),
    .reset(n5973),
    .set(1'b0),
    .q(T3abx6));  // ../RTL/cortexm0ds_logic.v(19861)
  AL_DFF T3fbx6_reg (
    .clk(HCLK),
    .d(Agrhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(T3fbx6));  // ../RTL/cortexm0ds_logic.v(20005)
  AL_DFF T3kpw6_reg (
    .clk(HCLK),
    .d(Amshu6),
    .reset(1'b0),
    .set(1'b0),
    .q(T3kpw6));  // ../RTL/cortexm0ds_logic.v(17287)
  AL_DFF T3opw6_reg (
    .clk(SWCLKTCK),
    .d(Hoxhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(T3opw6));  // ../RTL/cortexm0ds_logic.v(17493)
  AL_DFF T40qw6_reg (
    .clk(HCLK),
    .d(Mmrhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(T40qw6));  // ../RTL/cortexm0ds_logic.v(17916)
  AL_DFF T5fbx6_reg (
    .clk(HCLK),
    .d(Hgrhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(T5fbx6));  // ../RTL/cortexm0ds_logic.v(20006)
  AL_DFF T5mpw6_reg (
    .clk(SCLK),
    .d(Z0vhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(T5mpw6));  // ../RTL/cortexm0ds_logic.v(17412)
  AL_DFF T5yax6_reg (
    .clk(HCLK),
    .d(Htshu6),
    .reset(1'b0),
    .set(1'b0),
    .q(T5yax6));  // ../RTL/cortexm0ds_logic.v(18975)
  AL_DFF T60qw6_reg (
    .clk(HCLK),
    .d(Bdrhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(T60qw6));  // ../RTL/cortexm0ds_logic.v(17917)
  AL_DFF T6aax6_reg (
    .clk(DCLK),
    .d(Zzvhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(T6aax6));  // ../RTL/cortexm0ds_logic.v(18180)
  AL_DFF T6kbx6_reg (
    .clk(HCLK),
    .d(L4rhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(T6kbx6));  // ../RTL/cortexm0ds_logic.v(20233)
  AL_DFF T7bax6_reg (
    .clk(DCLK),
    .d(Xrvhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(T7bax6));  // ../RTL/cortexm0ds_logic.v(18220)
  AL_DFF T7fbx6_reg (
    .clk(HCLK),
    .d(Ogrhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(T7fbx6));  // ../RTL/cortexm0ds_logic.v(20007)
  AL_DFF T80qw6_reg (
    .clk(HCLK),
    .d(M8rhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(T80qw6));  // ../RTL/cortexm0ds_logic.v(17918)
  AL_DFF T82qw6_reg (
    .clk(SWCLKTCK),
    .d(Lqxhu6),
    .reset(n5972),
    .set(1'b0),
    .q(T82qw6));  // ../RTL/cortexm0ds_logic.v(17969)
  AL_DFF T8kbx6_reg (
    .clk(HCLK),
    .d(G8vhu6),
    .reset(n5973),
    .set(1'b0),
    .q(T8kbx6));  // ../RTL/cortexm0ds_logic.v(20238)
  AL_DFF T9fbx6_reg (
    .clk(HCLK),
    .d(Vgrhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(T9fbx6));  // ../RTL/cortexm0ds_logic.v(20008)
  AL_DFF T9kpw6_reg (
    .clk(SCLK),
    .d(Kbuhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(T9kpw6));  // ../RTL/cortexm0ds_logic.v(17290)
  AL_DFF Ta0qw6_reg (
    .clk(HCLK),
    .d(X3rhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Ta0qw6));  // ../RTL/cortexm0ds_logic.v(17919)
  AL_DFF Tajax6_reg (
    .clk(HCLK),
    .d(Yhohu6),
    .reset(1'b0),
    .set(n5973),
    .q(Tajax6));  // ../RTL/cortexm0ds_logic.v(18645)
  AL_DFF Tb3qw6_reg (
    .clk(DCLK),
    .d(Dfxhu6),
    .reset(n5974),
    .set(1'b0),
    .q(Tb3qw6));  // ../RTL/cortexm0ds_logic.v(18030)
  AL_DFF Tbfbx6_reg (
    .clk(HCLK),
    .d(Chrhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Tbfbx6));  // ../RTL/cortexm0ds_logic.v(20009)
  AL_DFF Tc0qw6_reg (
    .clk(HCLK),
    .d(Izqhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Tc0qw6));  // ../RTL/cortexm0ds_logic.v(17920)
  AL_DFF Tc9bx6_reg (
    .clk(DCLK),
    .d(Jkvhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Tc9bx6));  // ../RTL/cortexm0ds_logic.v(19813)
  AL_DFF Tceax6_reg (
    .clk(DCLK),
    .d(Xjwhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Tceax6));  // ../RTL/cortexm0ds_logic.v(18311)
  AL_DFF Tchbx6_reg (
    .clk(DCLK),
    .d(I1whu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Tchbx6));  // ../RTL/cortexm0ds_logic.v(20106)
  AL_DFF Tcipw6_reg (
    .clk(SCLK),
    .d(Jyohu6),
    .reset(n5973),
    .set(1'b0),
    .q(Tcipw6));  // ../RTL/cortexm0ds_logic.v(17199)
  AL_DFF Tcjax6_reg (
    .clk(HCLK),
    .d(Rhohu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Tcjax6));  // ../RTL/cortexm0ds_logic.v(18647)
  AL_DFF Tcjbx6_reg (
    .clk(DCLK),
    .d(Duwhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Tcjbx6));  // ../RTL/cortexm0ds_logic.v(20188)
  AL_DFF Tcrax6_reg (
    .clk(HCLK),
    .d(Bmphu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Tcrax6));  // ../RTL/cortexm0ds_logic.v(18847)
  AL_DFF Tdfbx6_reg (
    .clk(HCLK),
    .d(Jhrhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Tdfbx6));  // ../RTL/cortexm0ds_logic.v(20010)
  AL_DFF Tdypw6_reg (
    .clk(HCLK),
    .d(Hnrhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Tdypw6));  // ../RTL/cortexm0ds_logic.v(17879)
  AL_DFF Te0qw6_reg (
    .clk(HCLK),
    .d(Tuqhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Te0qw6));  // ../RTL/cortexm0ds_logic.v(17921)
  AL_DFF Tfcax6_reg (
    .clk(DCLK),
    .d(O4whu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Tfcax6));  // ../RTL/cortexm0ds_logic.v(18259)
  AL_DFF Tffbx6_reg (
    .clk(HCLK),
    .d(Qhrhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Tffbx6));  // ../RTL/cortexm0ds_logic.v(20011)
  AL_DFF Tg0qw6_reg (
    .clk(HCLK),
    .d(Eqqhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Tg0qw6));  // ../RTL/cortexm0ds_logic.v(17922)
  AL_DFF Tgkbx6_reg (
    .clk(HCLK),
    .d(Lashu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Tgkbx6));  // ../RTL/cortexm0ds_logic.v(20253)
  AL_DFF Tgzax6_reg (
    .clk(HCLK),
    .d(Ravhu6),
    .reset(n5973),
    .set(1'b0),
    .q(Tgzax6));  // ../RTL/cortexm0ds_logic.v(19107)
  AL_DFF Thcbx6_reg (
    .clk(DCLK),
    .d(Qqwhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Thcbx6));  // ../RTL/cortexm0ds_logic.v(19951)
  AL_DFF Thfbx6_reg (
    .clk(HCLK),
    .d(Xhrhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Thfbx6));  // ../RTL/cortexm0ds_logic.v(20012)
  AL_DFF Thhax6_reg (
    .clk(HCLK),
    .d(Zlohu6),
    .reset(1'b0),
    .set(n5973),
    .q(Thhax6));  // ../RTL/cortexm0ds_logic.v(18501)
  AL_DFF Thiax6_reg (
    .clk(DCLK),
    .d(Frthu6),
    .reset(n5974),
    .set(1'b0),
    .q(Thiax6));  // ../RTL/cortexm0ds_logic.v(18595)
  AL_DFF Thxax6_reg (
    .clk(HCLK),
    .d(Uguhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Thxax6));  // ../RTL/cortexm0ds_logic.v(18963)
  AL_DFF Ti0qw6_reg (
    .clk(HCLK),
    .d(Lcqhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Ti0qw6));  // ../RTL/cortexm0ds_logic.v(17923)
  AL_DFF Tikbx6_reg (
    .clk(DCLK),
    .d(M3whu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Tikbx6));  // ../RTL/cortexm0ds_logic.v(20254)
  AL_DFF Tjfbx6_reg (
    .clk(DCLK),
    .d(Rovhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Tjfbx6));  // ../RTL/cortexm0ds_logic.v(20013)
  AL_DFF Tjkpw6_reg (
    .clk(SCLK),
    .d(G9uhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Tjkpw6));  // ../RTL/cortexm0ds_logic.v(17300)
  AL_DFF Tjvax6_reg (
    .clk(HCLK),
    .d(F6thu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Tjvax6));  // ../RTL/cortexm0ds_logic.v(18923)
  AL_DFF Tk0qw6_reg (
    .clk(HCLK),
    .d(W7qhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Tk0qw6));  // ../RTL/cortexm0ds_logic.v(17924)
  AL_DFF Tkdax6_reg (
    .clk(DCLK),
    .d(Jqwhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Tkdax6));  // ../RTL/cortexm0ds_logic.v(18291)
  AL_DFF Tkjbx6_reg (
    .clk(HCLK),
    .d(Dpuhu6),
    .reset(n5973),
    .set(1'b0),
    .q(Tkjbx6));  // ../RTL/cortexm0ds_logic.v(20206)
  AL_DFF Tl4bx6_reg (
    .clk(HCLK),
    .d(Hlthu6),
    .reset(n5973),
    .set(1'b0),
    .q(Tl4bx6));  // ../RTL/cortexm0ds_logic.v(19641)
  AL_DFF Tlebx6_reg (
    .clk(HCLK),
    .d(Eirhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Tlebx6));  // ../RTL/cortexm0ds_logic.v(19996)
  AL_DFF Tm0qw6_reg (
    .clk(HCLK),
    .d(Syphu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Tm0qw6));  // ../RTL/cortexm0ds_logic.v(17925)
  AL_DFF Tmjbx6_reg (
    .clk(HCLK),
    .d(Ihuhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Tmjbx6));  // ../RTL/cortexm0ds_logic.v(20208)
  AL_DFF Tnebx6_reg (
    .clk(HCLK),
    .d(Wdrhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Tnebx6));  // ../RTL/cortexm0ds_logic.v(19997)
  AL_DFF Tngbx6_reg (
    .clk(HCLK),
    .d(Luthu6),
    .reset(n5973),
    .set(1'b0),
    .q(Tngbx6));  // ../RTL/cortexm0ds_logic.v(20087)
  AL_DFF Tokax6_reg (
    .clk(HCLK),
    .d(Eeohu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Tokax6));  // ../RTL/cortexm0ds_logic.v(18706)
  AL_DFF Tpebx6_reg (
    .clk(HCLK),
    .d(Derhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Tpebx6));  // ../RTL/cortexm0ds_logic.v(19998)
  AL_DFF Tptpw6_reg (
    .clk(HCLK),
    .d(Phuhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Tptpw6));  // ../RTL/cortexm0ds_logic.v(17689)
  AL_DFF Trebx6_reg (
    .clk(HCLK),
    .d(Kerhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Trebx6));  // ../RTL/cortexm0ds_logic.v(19999)
  AL_DFF Tsdbx6_reg (
    .clk(DCLK),
    .d(Apwhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Tsdbx6));  // ../RTL/cortexm0ds_logic.v(19981)
  AL_DFF Tt9ax6_reg (
    .clk(DCLK),
    .d(Vjvhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Tt9ax6));  // ../RTL/cortexm0ds_logic.v(18173)
  AL_DFF Ttebx6_reg (
    .clk(HCLK),
    .d(Rerhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Ttebx6));  // ../RTL/cortexm0ds_logic.v(20000)
  AL_DFF Tu0qw6_reg (
    .clk(HCLK),
    .d(Nlphu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Tu0qw6));  // ../RTL/cortexm0ds_logic.v(17929)
  AL_DFF Tujbx6_reg (
    .clk(HCLK),
    .d(Mbohu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Tujbx6));  // ../RTL/cortexm0ds_logic.v(20212)
  AL_DFF Tvebx6_reg (
    .clk(HCLK),
    .d(Yerhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Tvebx6));  // ../RTL/cortexm0ds_logic.v(20001)
  AL_DFF Twzpw6_reg (
    .clk(HCLK),
    .d(X9shu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Twzpw6));  // ../RTL/cortexm0ds_logic.v(17912)
  AL_DFF Txebx6_reg (
    .clk(HCLK),
    .d(Ffrhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Txebx6));  // ../RTL/cortexm0ds_logic.v(20002)
  AL_DFF Txmax6_reg (
    .clk(HCLK),
    .d(Q1thu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Txmax6));  // ../RTL/cortexm0ds_logic.v(18767)
  AL_DFF Tyaax6_reg (
    .clk(DCLK),
    .d(Ntvhu6),
    .reset(n5974),
    .set(1'b0),
    .q(Tyaax6));  // ../RTL/cortexm0ds_logic.v(18199)
  AL_DFF Tyipw6_reg (
    .clk(HCLK),
    .d(Diuhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Tyipw6));  // ../RTL/cortexm0ds_logic.v(17226)
  AL_DFF Tyzpw6_reg (
    .clk(HCLK),
    .d(I5shu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Tyzpw6));  // ../RTL/cortexm0ds_logic.v(17913)
  AL_DFF Tzebx6_reg (
    .clk(HCLK),
    .d(Mfrhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Tzebx6));  // ../RTL/cortexm0ds_logic.v(20003)
  AL_DFF Tzgbx6_reg (
    .clk(DCLK),
    .d(R9whu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Tzgbx6));  // ../RTL/cortexm0ds_logic.v(20099)
  AL_DFF U0hax6_reg (
    .clk(HCLK),
    .d(Koohu6),
    .reset(1'b0),
    .set(n5973),
    .q(U0hax6));  // ../RTL/cortexm0ds_logic.v(18447)
  AL_DFF U0rax6_reg (
    .clk(HCLK),
    .d(Ymqhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(U0rax6));  // ../RTL/cortexm0ds_logic.v(18841)
  AL_DFF U1kpw6_reg (
    .clk(HCLK),
    .d(Vethu6),
    .reset(1'b0),
    .set(1'b0),
    .q(U1kpw6));  // ../RTL/cortexm0ds_logic.v(17286)
  AL_DFF U2rax6_reg (
    .clk(HCLK),
    .d(Udqhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(U2rax6));  // ../RTL/cortexm0ds_logic.v(18842)
  AL_DFF U31bx6_reg (
    .clk(SCLK),
    .d(J5phu6),
    .reset(n5973),
    .set(1'b0),
    .q(U31bx6));  // ../RTL/cortexm0ds_logic.v(19281)
  AL_DFF U3yax6_reg (
    .clk(HCLK),
    .d(Bqshu6),
    .reset(1'b0),
    .set(1'b0),
    .q(U3yax6));  // ../RTL/cortexm0ds_logic.v(18974)
  AL_DFF U4fax6_reg (
    .clk(DCLK),
    .d(Jcwhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(U4fax6));  // ../RTL/cortexm0ds_logic.v(18326)
  AL_DFF U4rax6_reg (
    .clk(HCLK),
    .d(F9qhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(U4rax6));  // ../RTL/cortexm0ds_logic.v(18843)
  AL_DFF U6rax6_reg (
    .clk(HCLK),
    .d(Q4qhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(U6rax6));  // ../RTL/cortexm0ds_logic.v(18844)
  AL_DFF U7dax6_reg (
    .clk(DCLK),
    .d(Ptwhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(U7dax6));  // ../RTL/cortexm0ds_logic.v(18279)
  AL_DFF U8jax6_reg (
    .clk(HCLK),
    .d(Fiohu6),
    .reset(n5973),
    .set(1'b0),
    .q(U8jax6));  // ../RTL/cortexm0ds_logic.v(18639)
  AL_DFF U8rax6_reg (
    .clk(HCLK),
    .d(Mvphu6),
    .reset(1'b0),
    .set(1'b0),
    .q(U8rax6));  // ../RTL/cortexm0ds_logic.v(18845)
  AL_DFF U9ypw6_reg (
    .clk(HCLK),
    .d(Rhvhu6),
    .reset(1'b0),
    .set(n5973),
    .q(U9ypw6));  // ../RTL/cortexm0ds_logic.v(17876)
  AL_DFF Ua9bx6_reg (
    .clk(HCLK),
    .d(Wjshu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Ua9bx6));  // ../RTL/cortexm0ds_logic.v(19812)
  AL_DFF Uarax6_reg (
    .clk(HCLK),
    .d(Qqphu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Uarax6));  // ../RTL/cortexm0ds_logic.v(18846)
  AL_DFF Ubypw6_reg (
    .clk(HCLK),
    .d(Tpohu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Ubypw6));  // ../RTL/cortexm0ds_logic.v(17878)
  AL_DFF Ue9ax6_reg (
    .clk(DCLK),
    .d(Bnvhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Ue9ax6));  // ../RTL/cortexm0ds_logic.v(18165)
  AL_DFF Ufbbx6_reg (
    .clk(SWCLKTCK),
    .d(Gyxhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Ufbbx6));  // ../RTL/cortexm0ds_logic.v(19931)
  AL_DFF Ufebx6_reg (
    .clk(DCLK),
    .d(Qbxhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Ufebx6));  // ../RTL/cortexm0ds_logic.v(19993)
  AL_DFF Ufopw6_reg (
    .clk(HCLK),
    .d(Utohu6),
    .reset(n5973),
    .set(1'b0),
    .q(Ufopw6));  // ../RTL/cortexm0ds_logic.v(17518)
  AL_DFF Uh2qw6_reg (
    .clk(DCLK),
    .d(Ghthu6),
    .reset(n5974),
    .set(1'b0),
    .q(Uh2qw6));  // ../RTL/cortexm0ds_logic.v(17989)
  AL_DFF Uhvax6_reg (
    .clk(HCLK),
    .d(Rnphu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Uhvax6));  // ../RTL/cortexm0ds_logic.v(18922)
  AL_DFF Uizax6_reg (
    .clk(HCLK),
    .d(Txuhu6),
    .reset(n5973),
    .set(1'b0),
    .q(Uizax6));  // ../RTL/cortexm0ds_logic.v(19113)
  AL_DFF Uj4bx6_reg (
    .clk(HCLK),
    .d(Althu6),
    .reset(n5973),
    .set(1'b0),
    .q(Uj4bx6));  // ../RTL/cortexm0ds_logic.v(19635)
  AL_DFF Ujspw6_reg (
    .clk(HCLK),
    .d(Fjuhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Ujspw6));  // ../RTL/cortexm0ds_logic.v(17658)
  AL_DFF Ujxax6_reg (
    .clk(SCLK),
    .d(Aduhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Ujxax6));  // ../RTL/cortexm0ds_logic.v(18964)
  AL_DFF Um1bx6_reg (
    .clk(SCLK),
    .d(Uothu6),
    .reset(n5973),
    .set(1'b0),
    .q(Um1bx6));  // ../RTL/cortexm0ds_logic.v(19335)
  AL_DFF Umkax6_reg (
    .clk(HCLK),
    .d(Leohu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Umkax6));  // ../RTL/cortexm0ds_logic.v(18705)
  AL_DFF Untpw6_reg (
    .clk(HCLK),
    .d(I9vhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Untpw6));  // ../RTL/cortexm0ds_logic.v(17688)
  AL_DFF Unyax6_reg (
    .clk(HCLK),
    .d(N2uhu6),
    .reset(n5973),
    .set(1'b0),
    .q(Unyax6));  // ../RTL/cortexm0ds_logic.v(19023)
  AL_DFF Uo2bx6_reg (
    .clk(SCLK),
    .d(Pvuhu6),
    .reset(n5973),
    .set(1'b0),
    .q(Uo2bx6));  // ../RTL/cortexm0ds_logic.v(19443)
  AL_DFF Uofax6_reg (
    .clk(DCLK),
    .d(Pkhpw6[1]),
    .reset(n5974),
    .set(1'b0),
    .q(Uofax6));  // ../RTL/cortexm0ds_logic.v(18366)
  AL_DFF Uoipw6_reg (
    .clk(HCLK),
    .d(Wxshu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Uoipw6));  // ../RTL/cortexm0ds_logic.v(17216)
  AL_DFF Uojbx6_reg (
    .clk(SCLK),
    .d(Mcuhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Uojbx6));  // ../RTL/cortexm0ds_logic.v(20209)
  AL_DFF Uoqax6_reg (
    .clk(HCLK),
    .d(Gjrhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Uoqax6));  // ../RTL/cortexm0ds_logic.v(18835)
  AL_DFF Up4bx6_reg (
    .clk(HCLK),
    .d(X7uhu6),
    .reset(n5973),
    .set(1'b0),
    .q(Up4bx6));  // ../RTL/cortexm0ds_logic.v(19653)
  AL_DFF Uqipw6_reg (
    .clk(HCLK),
    .d(Oiphu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Uqipw6));  // ../RTL/cortexm0ds_logic.v(17217)
  AL_DFF Uqqax6_reg (
    .clk(HCLK),
    .d(V9rhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Uqqax6));  // ../RTL/cortexm0ds_logic.v(18836)
  AL_DFF Ureax6_reg (
    .clk(DCLK),
    .d(Bfwhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Ureax6));  // ../RTL/cortexm0ds_logic.v(18319)
  AL_DFF Urgbx6_reg (
    .clk(SWCLKTCK),
    .d(Ljxhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Urgbx6));  // ../RTL/cortexm0ds_logic.v(20095)
  AL_DFF Us3bx6_reg (
    .clk(SCLK),
    .d(Bxdpw6),
    .reset(n5973),
    .set(1'b0),
    .q(Us3bx6));  // ../RTL/cortexm0ds_logic.v(19557)
  AL_DFF Uscax6_reg (
    .clk(DCLK),
    .d(Vwwhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Uscax6));  // ../RTL/cortexm0ds_logic.v(18271)
  AL_DFF Usipw6_reg (
    .clk(HCLK),
    .d(Fxuhu6),
    .reset(n5973),
    .set(1'b0),
    .q(Usipw6));  // ../RTL/cortexm0ds_logic.v(17222)
  AL_DFF Usjbx6_reg (
    .clk(HCLK),
    .d(Tbohu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Usjbx6));  // ../RTL/cortexm0ds_logic.v(20211)
  AL_DFF Usnpw6_reg (
    .clk(HCLK),
    .d(Dgphu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Usnpw6));  // ../RTL/cortexm0ds_logic.v(17477)
  AL_DFF Usqax6_reg (
    .clk(HCLK),
    .d(G5rhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Usqax6));  // ../RTL/cortexm0ds_logic.v(18837)
  AL_DFF Utqpw6_reg (
    .clk(SWCLKTCK),
    .d(Fuxhu6),
    .reset(n5972),
    .set(1'b0),
    .q(Utqpw6));  // ../RTL/cortexm0ds_logic.v(17581)
  AL_DFF Uunpw6_reg (
    .clk(DCLK),
    .d(H2yhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Uunpw6));  // ../RTL/cortexm0ds_logic.v(17478)
  AL_DFF Uuqax6_reg (
    .clk(HCLK),
    .d(R0rhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Uuqax6));  // ../RTL/cortexm0ds_logic.v(18838)
  AL_DFF Uuzpw6_reg (
    .clk(HCLK),
    .d(Teshu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Uuzpw6));  // ../RTL/cortexm0ds_logic.v(17911)
  AL_DFF Uvmax6_reg (
    .clk(HCLK),
    .d(X1thu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Uvmax6));  // ../RTL/cortexm0ds_logic.v(18766)
  AL_DFF Uwipw6_reg (
    .clk(HCLK),
    .d(Igvhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Uwipw6));  // ../RTL/cortexm0ds_logic.v(17225)
  AL_DFF Uwqax6_reg (
    .clk(HCLK),
    .d(Cwqhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Uwqax6));  // ../RTL/cortexm0ds_logic.v(18839)
  AL_DFF Ux8bx6_reg (
    .clk(DCLK),
    .d(Mwvhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Ux8bx6));  // ../RTL/cortexm0ds_logic.v(19805)
  AL_DFF Uyqax6_reg (
    .clk(HCLK),
    .d(Nrqhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Uyqax6));  // ../RTL/cortexm0ds_logic.v(18840)
  AL_DFF V0cax6_reg (
    .clk(DCLK),
    .d(U7whu6),
    .reset(1'b0),
    .set(1'b0),
    .q(V0cax6));  // ../RTL/cortexm0ds_logic.v(18251)
  AL_DFF V0jpw6_reg (
    .clk(SCLK),
    .d(Rbuhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(V0jpw6));  // ../RTL/cortexm0ds_logic.v(17227)
  AL_DFF V1vax6_reg (
    .clk(HCLK),
    .d(Sxqhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(V1vax6));  // ../RTL/cortexm0ds_logic.v(18914)
  AL_DFF V1yax6_reg (
    .clk(HCLK),
    .d(Ibthu6),
    .reset(1'b0),
    .set(1'b0),
    .q(V1yax6));  // ../RTL/cortexm0ds_logic.v(18973)
  AL_DFF V3vax6_reg (
    .clk(HCLK),
    .d(Dtqhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(V3vax6));  // ../RTL/cortexm0ds_logic.v(18915)
  AL_DFF V52bx6_reg (
    .clk(SCLK),
    .d(U0phu6),
    .reset(n5973),
    .set(1'b0),
    .q(V52bx6));  // ../RTL/cortexm0ds_logic.v(19389)
  AL_DFF V53qw6_reg (
    .clk(DCLK),
    .d(Sdphu6),
    .reset(1'b0),
    .set(1'b0),
    .q(V53qw6));  // ../RTL/cortexm0ds_logic.v(18023)
  AL_DFF V5abx6_reg (
    .clk(HCLK),
    .d(Z1uhu6),
    .reset(n5973),
    .set(1'b0),
    .q(V5abx6));  // ../RTL/cortexm0ds_logic.v(19867)
  AL_DFF V5vax6_reg (
    .clk(HCLK),
    .d(Ooqhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(V5vax6));  // ../RTL/cortexm0ds_logic.v(18916)
  AL_DFF V6jax6_reg (
    .clk(HCLK),
    .d(Miohu6),
    .reset(1'b0),
    .set(1'b0),
    .q(V6jax6));  // ../RTL/cortexm0ds_logic.v(18634)
  AL_DFF V73bx6_reg (
    .clk(SCLK),
    .d(Xyohu6),
    .reset(n5973),
    .set(1'b0),
    .q(V73bx6));  // ../RTL/cortexm0ds_logic.v(19497)
  AL_DFF V7vax6_reg (
    .clk(HCLK),
    .d(Kfqhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(V7vax6));  // ../RTL/cortexm0ds_logic.v(18917)
  AL_DFF V9vax6_reg (
    .clk(HCLK),
    .d(Vaqhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(V9vax6));  // ../RTL/cortexm0ds_logic.v(18918)
  AL_DFF Va7ax6_reg (
    .clk(SWCLKTCK),
    .d(Plxhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Va7ax6));  // ../RTL/cortexm0ds_logic.v(18090)
  AL_DFF Vbkpw6_reg (
    .clk(HCLK),
    .d(C6vhu6),
    .reset(n5973),
    .set(1'b0),
    .q(Vbkpw6));  // ../RTL/cortexm0ds_logic.v(17295)
  AL_DFF Vbspw6_reg (
    .clk(HCLK),
    .d(Zuthu6),
    .reset(n5973),
    .set(1'b0),
    .q(Vbspw6));  // ../RTL/cortexm0ds_logic.v(17648)
  AL_DFF Vbvax6_reg (
    .clk(HCLK),
    .d(G6qhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Vbvax6));  // ../RTL/cortexm0ds_logic.v(18919)
  AL_DFF Vdvax6_reg (
    .clk(HCLK),
    .d(Cxphu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Vdvax6));  // ../RTL/cortexm0ds_logic.v(18920)
  AL_DFF Vefax6_reg (
    .clk(DCLK),
    .d(Edphu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Vefax6));  // ../RTL/cortexm0ds_logic.v(18357)
  AL_DFF Veqax6_reg (
    .clk(HCLK),
    .d(Y6shu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Veqax6));  // ../RTL/cortexm0ds_logic.v(18830)
  AL_DFF Vfvax6_reg (
    .clk(HCLK),
    .d(Gsphu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Vfvax6));  // ../RTL/cortexm0ds_logic.v(18921)
  AL_DFF Vgjpw6_reg (
    .clk(HCLK),
    .d(Oxohu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Vgjpw6));  // ../RTL/cortexm0ds_logic.v(17240)
  AL_DFF Vgqax6_reg (
    .clk(HCLK),
    .d(J2shu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Vgqax6));  // ../RTL/cortexm0ds_logic.v(18831)
  AL_DFF Vhspw6_reg (
    .clk(HCLK),
    .d(Lsohu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Vhspw6));  // ../RTL/cortexm0ds_logic.v(17657)
  AL_DFF Vibax6_reg (
    .clk(DCLK),
    .d(F3whu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Vibax6));  // ../RTL/cortexm0ds_logic.v(18226)
  AL_DFF Viqax6_reg (
    .clk(HCLK),
    .d(Uxrhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Viqax6));  // ../RTL/cortexm0ds_logic.v(18832)
  AL_DFF Vj3qw6_reg (
    .clk(DCLK),
    .d(R8xhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Vj3qw6));  // ../RTL/cortexm0ds_logic.v(18041)
  AL_DFF Vkqax6_reg (
    .clk(HCLK),
    .d(Mtrhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Vkqax6));  // ../RTL/cortexm0ds_logic.v(18833)
  AL_DFF Vkzax6_reg (
    .clk(HCLK),
    .d(Ivuhu6),
    .reset(n5973),
    .set(1'b0),
    .q(Vkzax6));  // ../RTL/cortexm0ds_logic.v(19119)
  AL_DFF Vlaax6_reg (
    .clk(DCLK),
    .d(Rvvhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Vlaax6));  // ../RTL/cortexm0ds_logic.v(18188)
  AL_DFF Vlkpw6_reg (
    .clk(HCLK),
    .d(Oaqhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Vlkpw6));  // ../RTL/cortexm0ds_logic.v(17301)
  AL_DFF Vltpw6_reg (
    .clk(HCLK),
    .d(B9vhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Vltpw6));  // ../RTL/cortexm0ds_logic.v(17687)
  AL_DFF Vlxax6_reg (
    .clk(HCLK),
    .d(Lfuhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Vlxax6));  // ../RTL/cortexm0ds_logic.v(18965)
  AL_DFF Vmipw6_reg (
    .clk(HCLK),
    .d(Vxohu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Vmipw6));  // ../RTL/cortexm0ds_logic.v(17215)
  AL_DFF Vmqax6_reg (
    .clk(HCLK),
    .d(Vnrhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Vmqax6));  // ../RTL/cortexm0ds_logic.v(18834)
  AL_DFF Vn9bx6_reg (
    .clk(DCLK),
    .d(I7xhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Vn9bx6));  // ../RTL/cortexm0ds_logic.v(19819)
  AL_DFF Vnkpw6_reg (
    .clk(HCLK),
    .d(Scqhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Vnkpw6));  // ../RTL/cortexm0ds_logic.v(17302)
  AL_DFF Vpgbx6_reg (
    .clk(HCLK),
    .d(Tkthu6),
    .reset(n5973),
    .set(1'b0),
    .q(Vpgbx6));  // ../RTL/cortexm0ds_logic.v(20093)
  AL_DFF Vpkpw6_reg (
    .clk(DCLK),
    .d(Bfphu6),
    .reset(n5974),
    .set(1'b0),
    .q(Vpkpw6));  // ../RTL/cortexm0ds_logic.v(17307)
  AL_DFF Vplpw6_reg (
    .clk(SWCLKTCK),
    .d(Rvohu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Vplpw6));  // ../RTL/cortexm0ds_logic.v(17383)
  AL_DFF Vqgax6_reg (
    .clk(DCLK),
    .d(T9xhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Vqgax6));  // ../RTL/cortexm0ds_logic.v(18412)
  AL_DFF Vqjbx6_reg (
    .clk(HCLK),
    .d(Acohu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Vqjbx6));  // ../RTL/cortexm0ds_logic.v(20210)
  AL_DFF Vrtpw6_reg (
    .clk(SCLK),
    .d(Fcuhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Vrtpw6));  // ../RTL/cortexm0ds_logic.v(17690)
  AL_DFF Vszpw6_reg (
    .clk(HCLK),
    .d(Ijshu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Vszpw6));  // ../RTL/cortexm0ds_logic.v(17910)
  AL_DFF Vtmax6_reg (
    .clk(HCLK),
    .d(Dnphu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Vtmax6));  // ../RTL/cortexm0ds_logic.v(18765)
  AL_DFF Vtuax6_reg (
    .clk(HCLK),
    .d(Wkrhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Vtuax6));  // ../RTL/cortexm0ds_logic.v(18910)
  AL_DFF Vuhax6_reg (
    .clk(HCLK),
    .d(Ckohu6),
    .reset(1'b0),
    .set(n5973),
    .q(Vuhax6));  // ../RTL/cortexm0ds_logic.v(18543)
  AL_DFF Vuipw6_reg (
    .clk(HCLK),
    .d(Kyshu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Vuipw6));  // ../RTL/cortexm0ds_logic.v(17224)
  AL_DFF Vvuax6_reg (
    .clk(HCLK),
    .d(Lbrhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Vvuax6));  // ../RTL/cortexm0ds_logic.v(18911)
  AL_DFF Vvxax6_reg (
    .clk(HCLK),
    .d(Dcthu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Vvxax6));  // ../RTL/cortexm0ds_logic.v(18970)
  AL_DFF Vxuax6_reg (
    .clk(HCLK),
    .d(W6rhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Vxuax6));  // ../RTL/cortexm0ds_logic.v(18912)
  AL_DFF Vxxax6_reg (
    .clk(HCLK),
    .d(Wbthu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Vxxax6));  // ../RTL/cortexm0ds_logic.v(18971)
  AL_DFF Vyfbx6_reg (
    .clk(SCLK),
    .d(Uuuhu6),
    .reset(n5973),
    .set(1'b0),
    .q(Vyfbx6));  // ../RTL/cortexm0ds_logic.v(20025)
  AL_DFF Vygax6_reg (
    .clk(HCLK),
    .d(U8vhu6),
    .reset(n5973),
    .set(1'b0),
    .q(Vygax6));  // ../RTL/cortexm0ds_logic.v(18441)
  AL_DFF Vz8ax6_reg (
    .clk(DCLK),
    .d(S5xhu6),
    .reset(n5974),
    .set(1'b0),
    .q(Vz8ax6));  // ../RTL/cortexm0ds_logic.v(18151)
  AL_DFF Vzdax6_reg (
    .clk(DCLK),
    .d(Imwhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Vzdax6));  // ../RTL/cortexm0ds_logic.v(18299)
  AL_DFF Vzjpw6_reg (
    .clk(SCLK),
    .d(Fivhu6),
    .reset(n5973),
    .set(1'b0),
    .q(Vzjpw6));  // ../RTL/cortexm0ds_logic.v(17284)
  AL_DFF Vzuax6_reg (
    .clk(HCLK),
    .d(H2rhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Vzuax6));  // ../RTL/cortexm0ds_logic.v(18913)
  AL_DFF Vzupw6_reg (
    .clk(HCLK),
    .d(Jrohu6),
    .reset(n5973),
    .set(1'b0),
    .q(Vzupw6));  // ../RTL/cortexm0ds_logic.v(17741)
  AL_DFF Vzxax6_reg (
    .clk(HCLK),
    .d(Pbthu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Vzxax6));  // ../RTL/cortexm0ds_logic.v(18972)
  AL_DFF W0dbx6_reg (
    .clk(DCLK),
    .d(Xqwhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(W0dbx6));  // ../RTL/cortexm0ds_logic.v(19966)
  AL_DFF W0jax6_reg (
    .clk(SCLK),
    .d(T4vhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(W0jax6));  // ../RTL/cortexm0ds_logic.v(18626)
  AL_DFF W2jax6_reg (
    .clk(SCLK),
    .d(A5vhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(W2jax6));  // ../RTL/cortexm0ds_logic.v(18627)
  AL_DFF W4aax6_reg (
    .clk(DCLK),
    .d(G0whu6),
    .reset(1'b0),
    .set(1'b0),
    .q(W4aax6));  // ../RTL/cortexm0ds_logic.v(18179)
  AL_DFF W4jax6_reg (
    .clk(HCLK),
    .d(Withu6),
    .reset(1'b0),
    .set(n5973),
    .q(W4jax6));  // ../RTL/cortexm0ds_logic.v(18632)
  AL_DFF W51bx6_reg (
    .clk(SCLK),
    .d(Gothu6),
    .reset(n5973),
    .set(1'b0),
    .q(W51bx6));  // ../RTL/cortexm0ds_logic.v(19287)
  AL_DFF W5max6_reg (
    .clk(HCLK),
    .d(Ikrhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(W5max6));  // ../RTL/cortexm0ds_logic.v(18753)
  AL_DFF W5ypw6_reg (
    .clk(HCLK),
    .d(Yavhu6),
    .reset(n5973),
    .set(1'b0),
    .q(W5ypw6));  // ../RTL/cortexm0ds_logic.v(17864)
  AL_DFF W6ipw6_reg (
    .clk(SWCLKTCK),
    .d(Grxhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(W6ipw6));  // ../RTL/cortexm0ds_logic.v(17187)
  AL_DFF W7max6_reg (
    .clk(HCLK),
    .d(Xarhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(W7max6));  // ../RTL/cortexm0ds_logic.v(18754)
  AL_DFF W8hbx6_reg (
    .clk(SCLK),
    .d(Yhvhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(W8hbx6));  // ../RTL/cortexm0ds_logic.v(20104)
  AL_DFF W9max6_reg (
    .clk(HCLK),
    .d(I6rhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(W9max6));  // ../RTL/cortexm0ds_logic.v(18755)
  AL_DFF W9spw6_reg (
    .clk(HCLK),
    .d(Dkshu6),
    .reset(1'b0),
    .set(1'b0),
    .q(W9spw6));  // ../RTL/cortexm0ds_logic.v(17643)
  AL_DFF Wahbx6_reg (
    .clk(DCLK),
    .d(Oqvhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Wahbx6));  // ../RTL/cortexm0ds_logic.v(20105)
  AL_DFF Wbmax6_reg (
    .clk(HCLK),
    .d(T1rhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Wbmax6));  // ../RTL/cortexm0ds_logic.v(18756)
  AL_DFF Wc2qw6_reg (
    .clk(DCLK),
    .d(F9xhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Wc2qw6));  // ../RTL/cortexm0ds_logic.v(17972)
  AL_DFF Wcqax6_reg (
    .clk(HCLK),
    .d(Ubshu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Wcqax6));  // ../RTL/cortexm0ds_logic.v(18829)
  AL_DFF Wdmax6_reg (
    .clk(HCLK),
    .d(Exqhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Wdmax6));  // ../RTL/cortexm0ds_logic.v(18757)
  AL_DFF Weipw6_reg (
    .clk(HCLK),
    .d(Vcvhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Weipw6));  // ../RTL/cortexm0ds_logic.v(17201)
  AL_DFF Wfcbx6_reg (
    .clk(DCLK),
    .d(Oiwhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Wfcbx6));  // ../RTL/cortexm0ds_logic.v(19950)
  AL_DFF Wfhax6_reg (
    .clk(HCLK),
    .d(Gmohu6),
    .reset(1'b0),
    .set(n5973),
    .q(Wfhax6));  // ../RTL/cortexm0ds_logic.v(18495)
  AL_DFF Wfmax6_reg (
    .clk(HCLK),
    .d(Psqhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Wfmax6));  // ../RTL/cortexm0ds_logic.v(18758)
  AL_DFF Wfspw6_reg (
    .clk(HCLK),
    .d(S7vhu6),
    .reset(1'b0),
    .set(n5973),
    .q(Wfspw6));  // ../RTL/cortexm0ds_logic.v(17655)
  AL_DFF Wgipw6_reg (
    .clk(HCLK),
    .d(Fkthu6),
    .reset(n5973),
    .set(1'b0),
    .q(Wgipw6));  // ../RTL/cortexm0ds_logic.v(17206)
  AL_DFF Whmax6_reg (
    .clk(HCLK),
    .d(Aoqhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Whmax6));  // ../RTL/cortexm0ds_logic.v(18759)
  AL_DFF Widax6_reg (
    .clk(DCLK),
    .d(Lrwhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Widax6));  // ../RTL/cortexm0ds_logic.v(18290)
  AL_DFF Wjmax6_reg (
    .clk(HCLK),
    .d(Weqhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Wjmax6));  // ../RTL/cortexm0ds_logic.v(18760)
  AL_DFF Wjtpw6_reg (
    .clk(HCLK),
    .d(L9thu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Wjtpw6));  // ../RTL/cortexm0ds_logic.v(17686)
  AL_DFF Wjuax6_reg (
    .clk(HCLK),
    .d(H8shu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Wjuax6));  // ../RTL/cortexm0ds_logic.v(18905)
  AL_DFF Wkipw6_reg (
    .clk(HCLK),
    .d(Bithu6),
    .reset(1'b0),
    .set(n5973),
    .q(Wkipw6));  // ../RTL/cortexm0ds_logic.v(17213)
  AL_DFF Wlmax6_reg (
    .clk(HCLK),
    .d(Haqhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Wlmax6));  // ../RTL/cortexm0ds_logic.v(18761)
  AL_DFF Wlspw6_reg (
    .clk(SCLK),
    .d(Pauhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Wlspw6));  // ../RTL/cortexm0ds_logic.v(17659)
  AL_DFF Wluax6_reg (
    .clk(HCLK),
    .d(S3shu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Wluax6));  // ../RTL/cortexm0ds_logic.v(18906)
  AL_DFF Wmzax6_reg (
    .clk(HCLK),
    .d(Aruhu6),
    .reset(n5973),
    .set(1'b0),
    .q(Wmzax6));  // ../RTL/cortexm0ds_logic.v(19125)
  AL_DFF Wnmax6_reg (
    .clk(HCLK),
    .d(S5qhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Wnmax6));  // ../RTL/cortexm0ds_logic.v(18762)
  AL_DFF Wnuax6_reg (
    .clk(HCLK),
    .d(Dzrhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Wnuax6));  // ../RTL/cortexm0ds_logic.v(18907)
  AL_DFF Wnxax6_reg (
    .clk(HCLK),
    .d(Efuhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Wnxax6));  // ../RTL/cortexm0ds_logic.v(18966)
  AL_DFF Woiax6_reg (
    .clk(SCLK),
    .d(Bpthu6),
    .reset(n5973),
    .set(1'b0),
    .q(Woiax6));  // ../RTL/cortexm0ds_logic.v(18619)
  AL_DFF Wpmax6_reg (
    .clk(HCLK),
    .d(Owphu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Wpmax6));  // ../RTL/cortexm0ds_logic.v(18763)
  AL_DFF Wpuax6_reg (
    .clk(HCLK),
    .d(Vurhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Wpuax6));  // ../RTL/cortexm0ds_logic.v(18908)
  AL_DFF Wpyax6_reg (
    .clk(HCLK),
    .d(G2uhu6),
    .reset(n5973),
    .set(1'b0),
    .q(Wpyax6));  // ../RTL/cortexm0ds_logic.v(19029)
  AL_DFF Wq8ax6_reg (
    .clk(SWCLKTCK),
    .d(Xwxhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Wq8ax6));  // ../RTL/cortexm0ds_logic.v(18132)
  AL_DFF Wqdbx6_reg (
    .clk(DCLK),
    .d(Ygwhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Wqdbx6));  // ../RTL/cortexm0ds_logic.v(19980)
  AL_DFF Wqzpw6_reg (
    .clk(HCLK),
    .d(Xnshu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Wqzpw6));  // ../RTL/cortexm0ds_logic.v(17909)
  AL_DFF Wr4bx6_reg (
    .clk(HCLK),
    .d(Q7uhu6),
    .reset(n5973),
    .set(1'b0),
    .q(Wr4bx6));  // ../RTL/cortexm0ds_logic.v(19659)
  AL_DFF Wrmax6_reg (
    .clk(HCLK),
    .d(Srphu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Wrmax6));  // ../RTL/cortexm0ds_logic.v(18764)
  AL_DFF Wruax6_reg (
    .clk(HCLK),
    .d(Lprhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Wruax6));  // ../RTL/cortexm0ds_logic.v(18909)
  AL_DFF Wt3qw6_reg (
    .clk(SWCLKTCK),
    .d(M1yhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Wt3qw6));  // ../RTL/cortexm0ds_logic.v(18047)
  AL_DFF Wtxax6_reg (
    .clk(HCLK),
    .d(Lgthu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Wtxax6));  // ../RTL/cortexm0ds_logic.v(18969)
  AL_DFF Wu3bx6_reg (
    .clk(HCLK),
    .d(A6uhu6),
    .reset(n5973),
    .set(1'b0),
    .q(Wu3bx6));  // ../RTL/cortexm0ds_logic.v(19563)
  AL_DFF Wvgax6_reg (
    .clk(DCLK),
    .d(C4xhu6),
    .reset(n5974),
    .set(1'b0),
    .q(Wvgax6));  // ../RTL/cortexm0ds_logic.v(18429)
  AL_DFF Wwiax6_reg (
    .clk(SCLK),
    .d(F4vhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Wwiax6));  // ../RTL/cortexm0ds_logic.v(18624)
  AL_DFF Wxgbx6_reg (
    .clk(DCLK),
    .d(Szvhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Wxgbx6));  // ../RTL/cortexm0ds_logic.v(20098)
  AL_DFF Wxjpw6_reg (
    .clk(HCLK),
    .d(Mwohu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Wxjpw6));  // ../RTL/cortexm0ds_logic.v(17279)
  AL_DFF Wyiax6_reg (
    .clk(SCLK),
    .d(M4vhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Wyiax6));  // ../RTL/cortexm0ds_logic.v(18625)
  AL_DFF X1max6_reg (
    .clk(HCLK),
    .d(Hurhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(X1max6));  // ../RTL/cortexm0ds_logic.v(18751)
  AL_DFF X1upw6_reg (
    .clk(HCLK),
    .d(Z3shu6),
    .reset(1'b0),
    .set(1'b0),
    .q(X1upw6));  // ../RTL/cortexm0ds_logic.v(17695)
  AL_DFF X2jpw6_reg (
    .clk(HCLK),
    .d(P6rhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(X2jpw6));  // ../RTL/cortexm0ds_logic.v(17228)
  AL_DFF X3max6_reg (
    .clk(HCLK),
    .d(Xorhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(X3max6));  // ../RTL/cortexm0ds_logic.v(18752)
  AL_DFF X3upw6_reg (
    .clk(HCLK),
    .d(D6shu6),
    .reset(1'b0),
    .set(1'b0),
    .q(X3upw6));  // ../RTL/cortexm0ds_logic.v(17696)
  AL_DFF X42qw6_reg (
    .clk(DCLK),
    .d(S6phu6),
    .reset(1'b0),
    .set(1'b0),
    .q(X42qw6));  // ../RTL/cortexm0ds_logic.v(17963)
  AL_DFF X4jpw6_reg (
    .clk(HCLK),
    .d(T8rhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(X4jpw6));  // ../RTL/cortexm0ds_logic.v(17229)
  AL_DFF X5bax6_reg (
    .clk(DCLK),
    .d(Qrvhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(X5bax6));  // ../RTL/cortexm0ds_logic.v(18219)
  AL_DFF X5ibx6_reg (
    .clk(HCLK),
    .d(Glphu6),
    .reset(n5973),
    .set(1'b0),
    .q(X5ibx6));  // ../RTL/cortexm0ds_logic.v(20165)
  AL_DFF X5opw6_reg (
    .clk(HCLK),
    .d(Gguhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(X5opw6));  // ../RTL/cortexm0ds_logic.v(17494)
  AL_DFF X5upw6_reg (
    .clk(HCLK),
    .d(Rwuhu6),
    .reset(n5973),
    .set(1'b0),
    .q(X5upw6));  // ../RTL/cortexm0ds_logic.v(17701)
  AL_DFF X6jpw6_reg (
    .clk(HCLK),
    .d(Hkuhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(X6jpw6));  // ../RTL/cortexm0ds_logic.v(17230)
  AL_DFF X7abx6_reg (
    .clk(HCLK),
    .d(Vzthu6),
    .reset(n5973),
    .set(1'b0),
    .q(X7abx6));  // ../RTL/cortexm0ds_logic.v(19873)
  AL_DFF X7spw6_reg (
    .clk(HCLK),
    .d(Zhshu6),
    .reset(1'b0),
    .set(1'b0),
    .q(X7spw6));  // ../RTL/cortexm0ds_logic.v(17642)
  AL_DFF X7ypw6_reg (
    .clk(HCLK),
    .d(L0vhu6),
    .reset(n5973),
    .set(1'b0),
    .q(X7ypw6));  // ../RTL/cortexm0ds_logic.v(17870)
  AL_DFF Xaeax6_reg (
    .clk(DCLK),
    .d(Ekwhu6),
    .reset(n5974),
    .set(1'b0),
    .q(Xaeax6));  // ../RTL/cortexm0ds_logic.v(18309)
  AL_DFF Xajbx6_reg (
    .clk(DCLK),
    .d(Bmwhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Xajbx6));  // ../RTL/cortexm0ds_logic.v(20187)
  AL_DFF Xaqax6_reg (
    .clk(HCLK),
    .d(Jgshu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Xaqax6));  // ../RTL/cortexm0ds_logic.v(18828)
  AL_DFF Xbopw6_reg (
    .clk(SCLK),
    .d(N8vhu6),
    .reset(1'b0),
    .set(n5973),
    .q(Xbopw6));  // ../RTL/cortexm0ds_logic.v(17506)
  AL_DFF Xc9ax6_reg (
    .clk(DCLK),
    .d(Pnvhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Xc9ax6));  // ../RTL/cortexm0ds_logic.v(18164)
  AL_DFF Xdcax6_reg (
    .clk(DCLK),
    .d(V4whu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Xdcax6));  // ../RTL/cortexm0ds_logic.v(18258)
  AL_DFF Xdebx6_reg (
    .clk(DCLK),
    .d(Jxwhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Xdebx6));  // ../RTL/cortexm0ds_logic.v(19992)
  AL_DFF Xdspw6_reg (
    .clk(SCLK),
    .d(O5vhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Xdspw6));  // ../RTL/cortexm0ds_logic.v(17650)
  AL_DFF Xf8ax6_reg (
    .clk(SWCLKTCK),
    .d(Lxxhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Xf8ax6));  // ../RTL/cortexm0ds_logic.v(18121)
  AL_DFF Xfiax6_reg (
    .clk(HCLK),
    .d(Xdvhu6),
    .reset(n5973),
    .set(1'b0),
    .q(Xfiax6));  // ../RTL/cortexm0ds_logic.v(18589)
  AL_DFF Xhtpw6_reg (
    .clk(HCLK),
    .d(Ryshu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Xhtpw6));  // ../RTL/cortexm0ds_logic.v(17685)
  AL_DFF Xhuax6_reg (
    .clk(HCLK),
    .d(Ddshu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Xhuax6));  // ../RTL/cortexm0ds_logic.v(18904)
  AL_DFF Xiipw6_reg (
    .clk(SCLK),
    .d(U1vhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Xiipw6));  // ../RTL/cortexm0ds_logic.v(17208)
  AL_DFF Xkqpw6_reg (
    .clk(SWCLKTCK),
    .d(Ytxhu6),
    .reset(n5972),
    .set(1'b0),
    .q(Xkqpw6));  // ../RTL/cortexm0ds_logic.v(17572)
  AL_DFF Xn7ax6_reg (
    .clk(DCLK),
    .d(K8xhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Xn7ax6));  // ../RTL/cortexm0ds_logic.v(18102)
  AL_DFF Xnbax6_reg (
    .clk(DCLK),
    .d(X6vhu6),
    .reset(n5974),
    .set(1'b0),
    .q(Xnbax6));  // ../RTL/cortexm0ds_logic.v(18243)
  AL_DFF Xo1bx6_reg (
    .clk(SCLK),
    .d(D2phu6),
    .reset(n5973),
    .set(1'b0),
    .q(Xo1bx6));  // ../RTL/cortexm0ds_logic.v(19341)
  AL_DFF Xozax6_reg (
    .clk(HCLK),
    .d(Mquhu6),
    .reset(n5973),
    .set(1'b0),
    .q(Xozax6));  // ../RTL/cortexm0ds_logic.v(19131)
  AL_DFF Xozpw6_reg (
    .clk(HCLK),
    .d(Tsshu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Xozpw6));  // ../RTL/cortexm0ds_logic.v(17908)
  AL_DFF Xpeax6_reg (
    .clk(DCLK),
    .d(Pfwhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Xpeax6));  // ../RTL/cortexm0ds_logic.v(18318)
  AL_DFF Xpxax6_reg (
    .clk(HCLK),
    .d(Zcqhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Xpxax6));  // ../RTL/cortexm0ds_logic.v(18967)
  AL_DFF Xq2bx6_reg (
    .clk(SCLK),
    .d(Szohu6),
    .reset(n5973),
    .set(1'b0),
    .q(Xq2bx6));  // ../RTL/cortexm0ds_logic.v(19449)
  AL_DFF Xqcax6_reg (
    .clk(DCLK),
    .d(Eywhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Xqcax6));  // ../RTL/cortexm0ds_logic.v(18270)
  AL_DFF Xr9ax6_reg (
    .clk(DCLK),
    .d(Ckvhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Xr9ax6));  // ../RTL/cortexm0ds_logic.v(18172)
  AL_DFF Xrxax6_reg (
    .clk(HCLK),
    .d(Egthu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Xrxax6));  // ../RTL/cortexm0ds_logic.v(18968)
  AL_DFF Xttpw6_reg (
    .clk(HCLK),
    .d(V1shu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Xttpw6));  // ../RTL/cortexm0ds_logic.v(17691)
  AL_DFF Xu2qw6_reg (
    .clk(DCLK),
    .d(Zdphu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Xu2qw6));  // ../RTL/cortexm0ds_logic.v(18007)
  AL_DFF Xuiax6_reg (
    .clk(SCLK),
    .d(Y3vhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Xuiax6));  // ../RTL/cortexm0ds_logic.v(18623)
  AL_DFF Xv8bx6_reg (
    .clk(DCLK),
    .d(Slvhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Xv8bx6));  // ../RTL/cortexm0ds_logic.v(19804)
  AL_DFF Xvlax6_reg (
    .clk(HCLK),
    .d(T7shu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Xvlax6));  // ../RTL/cortexm0ds_logic.v(18748)
  AL_DFF Xvqpw6_reg (
    .clk(DCLK),
    .d(G2ohu6),
    .reset(n5974),
    .set(1'b0),
    .q(Xvqpw6));  // ../RTL/cortexm0ds_logic.v(17587)
  AL_DFF Xvtpw6_reg (
    .clk(HCLK),
    .d(C2shu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Xvtpw6));  // ../RTL/cortexm0ds_logic.v(17692)
  AL_DFF Xwaax6_reg (
    .clk(DCLK),
    .d(Utvhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Xwaax6));  // ../RTL/cortexm0ds_logic.v(18194)
  AL_DFF Xx6bx6_reg (
    .clk(SWCLKTCK),
    .d(Rmxhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Xx6bx6));  // ../RTL/cortexm0ds_logic.v(19764)
  AL_DFF Xxlax6_reg (
    .clk(HCLK),
    .d(E3shu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Xxlax6));  // ../RTL/cortexm0ds_logic.v(18749)
  AL_DFF Xxqpw6_reg (
    .clk(DCLK),
    .d(Q7ohu6),
    .reset(n5974),
    .set(1'b0),
    .q(Xxqpw6));  // ../RTL/cortexm0ds_logic.v(17593)
  AL_DFF Xxtpw6_reg (
    .clk(HCLK),
    .d(X2shu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Xxtpw6));  // ../RTL/cortexm0ds_logic.v(17693)
  AL_DFF Xxupw6_reg (
    .clk(HCLK),
    .d(Qrohu6),
    .reset(n5973),
    .set(1'b0),
    .q(Xxupw6));  // ../RTL/cortexm0ds_logic.v(17735)
  AL_DFF Xzlax6_reg (
    .clk(HCLK),
    .d(Pyrhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Xzlax6));  // ../RTL/cortexm0ds_logic.v(18750)
  AL_DFF Xztpw6_reg (
    .clk(HCLK),
    .d(L3shu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Xztpw6));  // ../RTL/cortexm0ds_logic.v(17694)
  AL_DFF Y0gbx6_reg (
    .clk(SCLK),
    .d(Zzohu6),
    .reset(n5973),
    .set(1'b0),
    .q(Y0gbx6));  // ../RTL/cortexm0ds_logic.v(20031)
  AL_DFF Y2fax6_reg (
    .clk(DCLK),
    .d(Qcwhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Y2fax6));  // ../RTL/cortexm0ds_logic.v(18325)
  AL_DFF Y5dax6_reg (
    .clk(DCLK),
    .d(Wtwhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Y5dax6));  // ../RTL/cortexm0ds_logic.v(18278)
  AL_DFF Y5spw6_reg (
    .clk(HCLK),
    .d(Lhshu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Y5spw6));  // ../RTL/cortexm0ds_logic.v(17641)
  AL_DFF Y72bx6_reg (
    .clk(SCLK),
    .d(Cmthu6),
    .reset(n5973),
    .set(1'b0),
    .q(Y72bx6));  // ../RTL/cortexm0ds_logic.v(19395)
  AL_DFF Y7opw6_reg (
    .clk(SCLK),
    .d(Oduhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Y7opw6));  // ../RTL/cortexm0ds_logic.v(17495)
  AL_DFF Y7upw6_reg (
    .clk(HCLK),
    .d(Zqqhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Y7upw6));  // ../RTL/cortexm0ds_logic.v(17703)
  AL_DFF Y8lpw6_reg (
    .clk(SWCLKTCK),
    .d(Rfxhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Y8lpw6));  // ../RTL/cortexm0ds_logic.v(17333)
  AL_DFF Y8qax6_reg (
    .clk(HCLK),
    .d(Ykshu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Y8qax6));  // ../RTL/cortexm0ds_logic.v(18827)
  AL_DFF Y93bx6_reg (
    .clk(SCLK),
    .d(J6vhu6),
    .reset(n5973),
    .set(1'b0),
    .q(Y93bx6));  // ../RTL/cortexm0ds_logic.v(19503)
  AL_DFF Y9upw6_reg (
    .clk(HCLK),
    .d(Grqhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Y9upw6));  // ../RTL/cortexm0ds_logic.v(17704)
  AL_DFF Ybupw6_reg (
    .clk(HCLK),
    .d(Isqhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Ybupw6));  // ../RTL/cortexm0ds_logic.v(17705)
  AL_DFF Ydgax6_reg (
    .clk(DCLK),
    .d(O2yhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Ydgax6));  // ../RTL/cortexm0ds_logic.v(18405)
  AL_DFF Ydopw6_reg (
    .clk(HCLK),
    .d(Buohu6),
    .reset(n5973),
    .set(1'b0),
    .q(Ydopw6));  // ../RTL/cortexm0ds_logic.v(17512)
  AL_DFF Ydupw6_reg (
    .clk(HCLK),
    .d(Wsqhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Ydupw6));  // ../RTL/cortexm0ds_logic.v(17706)
  AL_DFF Yf1qw6_reg (
    .clk(DCLK),
    .d(N6xhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Yf1qw6));  // ../RTL/cortexm0ds_logic.v(17940)
  AL_DFF Yftpw6_reg (
    .clk(HCLK),
    .d(Lvshu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Yftpw6));  // ../RTL/cortexm0ds_logic.v(17684)
  AL_DFF Yfuax6_reg (
    .clk(HCLK),
    .d(Shshu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Yfuax6));  // ../RTL/cortexm0ds_logic.v(18903)
  AL_DFF Yfupw6_reg (
    .clk(HCLK),
    .d(Ktqhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Yfupw6));  // ../RTL/cortexm0ds_logic.v(17707)
  AL_DFF Yhupw6_reg (
    .clk(HCLK),
    .d(Avqhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Yhupw6));  // ../RTL/cortexm0ds_logic.v(17708)
  AL_DFF Yizpw6_reg (
    .clk(HCLK),
    .d(Z2thu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Yizpw6));  // ../RTL/cortexm0ds_logic.v(17905)
  AL_DFF Yjaax6_reg (
    .clk(DCLK),
    .d(Fwvhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Yjaax6));  // ../RTL/cortexm0ds_logic.v(18187)
  AL_DFF Yjupw6_reg (
    .clk(HCLK),
    .d(Mjuhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Yjupw6));  // ../RTL/cortexm0ds_logic.v(17709)
  AL_DFF Yklpw6_reg (
    .clk(SWCLKTCK),
    .d(Zehpw6[4]),
    .reset(n5972),
    .set(1'b0),
    .q(Yklpw6));  // ../RTL/cortexm0ds_logic.v(17374)
  AL_DFF Ykzpw6_reg (
    .clk(HCLK),
    .d(S2thu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Ykzpw6));  // ../RTL/cortexm0ds_logic.v(17906)
  AL_DFF Ym3qw6_reg (
    .clk(DCLK),
    .d(Ecxhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Ym3qw6));  // ../RTL/cortexm0ds_logic.v(18043)
  AL_DFF Ymwpw6_reg (
    .clk(SWCLKTCK),
    .d(Ilxhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Ymwpw6));  // ../RTL/cortexm0ds_logic.v(17817)
  AL_DFF Ymzpw6_reg (
    .clk(HCLK),
    .d(E2thu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Ymzpw6));  // ../RTL/cortexm0ds_logic.v(17907)
  AL_DFF Ynspw6_reg (
    .clk(HCLK),
    .d(K6shu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Ynspw6));  // ../RTL/cortexm0ds_logic.v(17660)
  AL_DFF Yogax6_reg (
    .clk(DCLK),
    .d(Gzwhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Yogax6));  // ../RTL/cortexm0ds_logic.v(18411)
  AL_DFF Ypspw6_reg (
    .clk(HCLK),
    .d(R6shu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Ypspw6));  // ../RTL/cortexm0ds_logic.v(17661)
  AL_DFF Yqzax6_reg (
    .clk(HCLK),
    .d(Iouhu6),
    .reset(n5973),
    .set(1'b0),
    .q(Yqzax6));  // ../RTL/cortexm0ds_logic.v(19137)
  AL_DFF Yrspw6_reg (
    .clk(HCLK),
    .d(M7shu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Yrspw6));  // ../RTL/cortexm0ds_logic.v(17662)
  AL_DFF Yryax6_reg (
    .clk(HCLK),
    .d(Suthu6),
    .reset(n5973),
    .set(1'b0),
    .q(Yryax6));  // ../RTL/cortexm0ds_logic.v(19035)
  AL_DFF Ysiax6_reg (
    .clk(SCLK),
    .d(R3vhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Ysiax6));  // ../RTL/cortexm0ds_logic.v(18622)
  AL_DFF Yt4bx6_reg (
    .clk(HCLK),
    .d(C7uhu6),
    .reset(n5973),
    .set(1'b0),
    .q(Yt4bx6));  // ../RTL/cortexm0ds_logic.v(19665)
  AL_DFF Yt8bx6_reg (
    .clk(HCLK),
    .d(O3qhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Yt8bx6));  // ../RTL/cortexm0ds_logic.v(19803)
  AL_DFF Ytlax6_reg (
    .clk(HCLK),
    .d(Pcshu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Ytlax6));  // ../RTL/cortexm0ds_logic.v(18747)
  AL_DFF Ytspw6_reg (
    .clk(HCLK),
    .d(A8shu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Ytspw6));  // ../RTL/cortexm0ds_logic.v(17663)
  AL_DFF Yubbx6_reg (
    .clk(DCLK),
    .d(Scxhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Yubbx6));  // ../RTL/cortexm0ds_logic.v(19939)
  AL_DFF Yvabx6_reg (
    .clk(DCLK),
    .d(Ndxhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Yvabx6));  // ../RTL/cortexm0ds_logic.v(19896)
  AL_DFF Yvjpw6_reg (
    .clk(HCLK),
    .d(Twohu6),
    .reset(n5973),
    .set(1'b0),
    .q(Yvjpw6));  // ../RTL/cortexm0ds_logic.v(17277)
  AL_DFF Yvspw6_reg (
    .clk(HCLK),
    .d(O8shu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Yvspw6));  // ../RTL/cortexm0ds_logic.v(17664)
  AL_DFF Yw3bx6_reg (
    .clk(HCLK),
    .d(T5uhu6),
    .reset(n5973),
    .set(1'b0),
    .q(Yw3bx6));  // ../RTL/cortexm0ds_logic.v(19569)
  AL_DFF Yxdax6_reg (
    .clk(DCLK),
    .d(Wmwhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Yxdax6));  // ../RTL/cortexm0ds_logic.v(18298)
  AL_DFF Yxrpw6_reg (
    .clk(SCLK),
    .d(W1phu6),
    .reset(n5973),
    .set(1'b0),
    .q(Yxrpw6));  // ../RTL/cortexm0ds_logic.v(17636)
  AL_DFF Yxspw6_reg (
    .clk(HCLK),
    .d(Sashu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Yxspw6));  // ../RTL/cortexm0ds_logic.v(17665)
  AL_DFF Yybax6_reg (
    .clk(DCLK),
    .d(I8whu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Yybax6));  // ../RTL/cortexm0ds_logic.v(18250)
  AL_DFF Yzlpw6_reg (
    .clk(SWCLKTCK),
    .d(C3yhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Yzlpw6));  // ../RTL/cortexm0ds_logic.v(17404)
  AL_DFF Yzqpw6_reg (
    .clk(SWCLKTCK),
    .d(V2yhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Yzqpw6));  // ../RTL/cortexm0ds_logic.v(17595)
  AL_DFF Yzspw6_reg (
    .clk(HCLK),
    .d(Tivhu6),
    .reset(n5973),
    .set(1'b0),
    .q(Yzspw6));  // ../RTL/cortexm0ds_logic.v(17670)
  AL_DFF Z18bx6_reg (
    .clk(HCLK),
    .d(Ejqhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Z18bx6));  // ../RTL/cortexm0ds_logic.v(19789)
  AL_DFF Z1tpw6_reg (
    .clk(HCLK),
    .d(Sirhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Z1tpw6));  // ../RTL/cortexm0ds_logic.v(17672)
  AL_DFF Z2aax6_reg (
    .clk(DCLK),
    .d(P1whu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Z2aax6));  // ../RTL/cortexm0ds_logic.v(18178)
  AL_DFF Z38bx6_reg (
    .clk(HCLK),
    .d(Ljqhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Z38bx6));  // ../RTL/cortexm0ds_logic.v(19790)
  AL_DFF Z3spw6_reg (
    .clk(HCLK),
    .d(Xgshu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Z3spw6));  // ../RTL/cortexm0ds_logic.v(17640)
  AL_DFF Z3tpw6_reg (
    .clk(HCLK),
    .d(Zirhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Z3tpw6));  // ../RTL/cortexm0ds_logic.v(17673)
  AL_DFF Z47ax6_reg (
    .clk(HCLK),
    .d(Dmqhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Z47ax6));  // ../RTL/cortexm0ds_logic.v(18087)
  AL_DFF Z58bx6_reg (
    .clk(HCLK),
    .d(Sjqhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Z58bx6));  // ../RTL/cortexm0ds_logic.v(19791)
  AL_DFF Z5tpw6_reg (
    .clk(HCLK),
    .d(Bkrhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Z5tpw6));  // ../RTL/cortexm0ds_logic.v(17674)
  AL_DFF Z67ax6_reg (
    .clk(DCLK),
    .d(Taphu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Z67ax6));  // ../RTL/cortexm0ds_logic.v(18088)
  AL_DFF Z6qax6_reg (
    .clk(HCLK),
    .d(Upshu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Z6qax6));  // ../RTL/cortexm0ds_logic.v(18826)
  AL_DFF Z71bx6_reg (
    .clk(SCLK),
    .d(R2phu6),
    .reset(n5973),
    .set(1'b0),
    .q(Z71bx6));  // ../RTL/cortexm0ds_logic.v(19293)
  AL_DFF Z73qw6_reg (
    .clk(SWCLKTCK),
    .d(Psxhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Z73qw6));  // ../RTL/cortexm0ds_logic.v(18024)
  AL_DFF Z78bx6_reg (
    .clk(HCLK),
    .d(Zjqhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Z78bx6));  // ../RTL/cortexm0ds_logic.v(19792)
  AL_DFF Z7tpw6_reg (
    .clk(HCLK),
    .d(Pkrhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Z7tpw6));  // ../RTL/cortexm0ds_logic.v(17675)
  AL_DFF Z8jpw6_reg (
    .clk(SCLK),
    .d(N9uhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Z8jpw6));  // ../RTL/cortexm0ds_logic.v(17231)
  AL_DFF Z8zpw6_reg (
    .clk(HCLK),
    .d(Eashu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Z8zpw6));  // ../RTL/cortexm0ds_logic.v(17900)
  AL_DFF Z98bx6_reg (
    .clk(HCLK),
    .d(Gkqhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Z98bx6));  // ../RTL/cortexm0ds_logic.v(19793)
  AL_DFF Z9abx6_reg (
    .clk(HCLK),
    .d(Rxthu6),
    .reset(n5973),
    .set(1'b0),
    .q(Z9abx6));  // ../RTL/cortexm0ds_logic.v(19879)
  AL_DFF Z9opw6_reg (
    .clk(SCLK),
    .d(J4xhu6),
    .reset(n5973),
    .set(1'b0),
    .q(Z9opw6));  // ../RTL/cortexm0ds_logic.v(17500)
  AL_DFF Z9tpw6_reg (
    .clk(HCLK),
    .d(Dlrhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Z9tpw6));  // ../RTL/cortexm0ds_logic.v(17676)
  AL_DFF Zazpw6_reg (
    .clk(HCLK),
    .d(P5shu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Zazpw6));  // ../RTL/cortexm0ds_logic.v(17901)
  AL_DFF Zb8bx6_reg (
    .clk(HCLK),
    .d(Nkqhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Zb8bx6));  // ../RTL/cortexm0ds_logic.v(19794)
  AL_DFF Zbtpw6_reg (
    .clk(HCLK),
    .d(Tmrhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Zbtpw6));  // ../RTL/cortexm0ds_logic.v(17677)
  AL_DFF Zczpw6_reg (
    .clk(HCLK),
    .d(A1shu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Zczpw6));  // ../RTL/cortexm0ds_logic.v(17902)
  AL_DFF Zd8bx6_reg (
    .clk(HCLK),
    .d(Ukqhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Zd8bx6));  // ../RTL/cortexm0ds_logic.v(19795)
  AL_DFF Zdcbx6_reg (
    .clk(DCLK),
    .d(Mawhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Zdcbx6));  // ../RTL/cortexm0ds_logic.v(19949)
  AL_DFF Zdhax6_reg (
    .clk(HCLK),
    .d(Nmohu6),
    .reset(1'b0),
    .set(n5973),
    .q(Zdhax6));  // ../RTL/cortexm0ds_logic.v(18489)
  AL_DFF Zdiax6_reg (
    .clk(HCLK),
    .d(Tiohu6),
    .reset(n5973),
    .set(1'b0),
    .q(Zdiax6));  // ../RTL/cortexm0ds_logic.v(18583)
  AL_DFF Zdtpw6_reg (
    .clk(SCLK),
    .d(Qmthu6),
    .reset(n5973),
    .set(1'b0),
    .q(Zdtpw6));  // ../RTL/cortexm0ds_logic.v(17682)
  AL_DFF Zduax6_reg (
    .clk(HCLK),
    .d(Hmshu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Zduax6));  // ../RTL/cortexm0ds_logic.v(18902)
  AL_DFF Zezpw6_reg (
    .clk(HCLK),
    .d(Swrhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Zezpw6));  // ../RTL/cortexm0ds_logic.v(17903)
  AL_DFF Zf8bx6_reg (
    .clk(HCLK),
    .d(Blqhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Zf8bx6));  // ../RTL/cortexm0ds_logic.v(19796)
  AL_DFF Zgbax6_reg (
    .clk(DCLK),
    .d(Y2whu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Zgbax6));  // ../RTL/cortexm0ds_logic.v(18225)
  AL_DFF Zgfax6_reg (
    .clk(SWCLKTCK),
    .d(Dtxhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Zgfax6));  // ../RTL/cortexm0ds_logic.v(18358)
  AL_DFF Zgzpw6_reg (
    .clk(HCLK),
    .d(G3thu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Zgzpw6));  // ../RTL/cortexm0ds_logic.v(17904)
  AL_DFF Zh8bx6_reg (
    .clk(HCLK),
    .d(Ilqhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Zh8bx6));  // ../RTL/cortexm0ds_logic.v(19797)
  AL_DFF Zj8bx6_reg (
    .clk(HCLK),
    .d(Plqhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Zj8bx6));  // ../RTL/cortexm0ds_logic.v(19798)
  AL_DFF Zl8bx6_reg (
    .clk(HCLK),
    .d(Wlqhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Zl8bx6));  // ../RTL/cortexm0ds_logic.v(19799)
  AL_DFF Zl9bx6_reg (
    .clk(DCLK),
    .d(Itwhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Zl9bx6));  // ../RTL/cortexm0ds_logic.v(19818)
  AL_DFF Zm8ax6_reg (
    .clk(DCLK),
    .d(H3xhu6),
    .reset(n5974),
    .set(1'b0),
    .q(Zm8ax6));  // ../RTL/cortexm0ds_logic.v(18129)
  AL_DFF Zn8bx6_reg (
    .clk(HCLK),
    .d(T2qhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Zn8bx6));  // ../RTL/cortexm0ds_logic.v(19800)
  AL_DFF Zodbx6_reg (
    .clk(DCLK),
    .d(W8whu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Zodbx6));  // ../RTL/cortexm0ds_logic.v(19979)
  AL_DFF Zp8bx6_reg (
    .clk(HCLK),
    .d(A3qhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Zp8bx6));  // ../RTL/cortexm0ds_logic.v(19801)
  AL_DFF Zqiax6_reg (
    .clk(SCLK),
    .d(K3vhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Zqiax6));  // ../RTL/cortexm0ds_logic.v(18621)
  AL_DFF Zr7bx6_reg (
    .clk(HCLK),
    .d(Vhqhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Zr7bx6));  // ../RTL/cortexm0ds_logic.v(19784)
  AL_DFF Zr8bx6_reg (
    .clk(HCLK),
    .d(H3qhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Zr8bx6));  // ../RTL/cortexm0ds_logic.v(19802)
  AL_DFF Zrlax6_reg (
    .clk(HCLK),
    .d(Ehshu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Zrlax6));  // ../RTL/cortexm0ds_logic.v(18746)
  AL_DFF Zshax6_reg (
    .clk(HCLK),
    .d(Jkohu6),
    .reset(1'b0),
    .set(n5973),
    .q(Zshax6));  // ../RTL/cortexm0ds_logic.v(18537)
  AL_DFF Zslpw6_reg (
    .clk(SWCLKTCK),
    .d(Dvohu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Zslpw6));  // ../RTL/cortexm0ds_logic.v(17385)
  AL_DFF Zszax6_reg (
    .clk(HCLK),
    .d(Emuhu6),
    .reset(n5973),
    .set(1'b0),
    .q(Zszax6));  // ../RTL/cortexm0ds_logic.v(19143)
  AL_DFF Zt7bx6_reg (
    .clk(HCLK),
    .d(Ciqhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Zt7bx6));  // ../RTL/cortexm0ds_logic.v(19785)
  AL_DFF Ztgbx6_reg (
    .clk(HCLK),
    .d(Kavhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Ztgbx6));  // ../RTL/cortexm0ds_logic.v(20096)
  AL_DFF Ztupw6_reg (
    .clk(HCLK),
    .d(Fbvhu6),
    .reset(n5973),
    .set(1'b0),
    .q(Ztupw6));  // ../RTL/cortexm0ds_logic.v(17723)
  AL_DFF Zv7bx6_reg (
    .clk(HCLK),
    .d(Jiqhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Zv7bx6));  // ../RTL/cortexm0ds_logic.v(19786)
  AL_DFF Zvgbx6_reg (
    .clk(DCLK),
    .d(Yovhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Zvgbx6));  // ../RTL/cortexm0ds_logic.v(20097)
  AL_DFF Zvrpw6_reg (
    .clk(HCLK),
    .d(Ofshu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Zvrpw6));  // ../RTL/cortexm0ds_logic.v(17631)
  AL_DFF Zwnpw6_reg (
    .clk(SWCLKTCK),
    .d(A2yhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Zwnpw6));  // ../RTL/cortexm0ds_logic.v(17479)
  AL_DFF Zx7bx6_reg (
    .clk(HCLK),
    .d(Qiqhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Zx7bx6));  // ../RTL/cortexm0ds_logic.v(19787)
  AL_DFF Zx8ax6_reg (
    .clk(DCLK),
    .d(Z5xhu6),
    .reset(n5974),
    .set(1'b0),
    .q(Zx8ax6));  // ../RTL/cortexm0ds_logic.v(18145)
  AL_DFF Zycbx6_reg (
    .clk(DCLK),
    .d(Viwhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Zycbx6));  // ../RTL/cortexm0ds_logic.v(19965)
  AL_DFF Zz7bx6_reg (
    .clk(HCLK),
    .d(Xiqhu6),
    .reset(1'b0),
    .set(1'b0),
    .q(Zz7bx6));  // ../RTL/cortexm0ds_logic.v(19788)
  add_pu10_pu10_o10 add0 (
    .i0({Jshpw6[9:4],Tnhpw6}),
    .i1({7'b0000000,Aphpw6,E4yhu6}),
    .o(Vrkbx6[10:1]));  // ../RTL/cortexm0ds_logic.v(3108)
  add_pu31_pu31_o31 add1 (
    .i0(vis_pc_o),
    .i1(31'b0000000000000000000000000000001),
    .o(Zsfpw6));  // ../RTL/cortexm0ds_logic.v(3152)
  add_pu30_pu30_o30 add2 (
    .i0({vis_pc_o[30:2],R0ghu6}),
    .i1(30'b000000000000000000000000000001),
    .o({N5fpw6,open_n0}));  // ../RTL/cortexm0ds_logic.v(3153)
  add_pu33_pu33_o33 add3 (
    .i0({Qbehu6,Edehu6,Seehu6,Ggehu6,Uhehu6,Ijehu6,Wkehu6,Kmehu6,Ynehu6,Mpehu6,Arehu6,Osehu6,Cuehu6,Qvehu6,Exehu6,Syehu6,G0fhu6,U1fhu6,I3fhu6,W4fhu6,K6fhu6,Y7fhu6,M9fhu6,Abfhu6,Ocfhu6,Cefhu6,Qffhu6,Dhfhu6,Qifhu6,Dkfhu6,Qlfhu6,Dnfhu6,Qofhu6}),
    .i1({32'b00000000000000000000000000000000,Dqfhu6}),
    .o(Nxkbx6[33:1]));  // ../RTL/cortexm0ds_logic.v(3166)
  add_pu32_pu32_o33 add4 (
    .i0(Idfpw6),
    .i1({D5epw6,Qbfpw6[30:23],P4epw6,I4epw6,B4epw6,U3epw6,N3epw6,G3epw6,Z2epw6,L2epw6,X1epw6,Q1epw6,J1epw6,C1epw6,Qbfpw6[10],Q5phu6,W4epw6,S2epw6,E2epw6,Qbfpw6[5:0]}),
    .o(Ozkbx6[33:1]));  // ../RTL/cortexm0ds_logic.v(3171)
  eq_w32 eq0 (
    .i0({R9ohu6,Mzihu6,Eyihu6,Wwihu6,Ovihu6,Guihu6,Ysihu6,Qrihu6,Iqihu6,Apihu6,Snihu6,Kmihu6,Clihu6,Ujihu6,Miihu6,Ehihu6,Wfihu6,Oeihu6,Gdihu6,Ybihu6,Qaihu6,I9ihu6,A8ihu6,S6ihu6,K5ihu6,C4ihu6,U2ihu6,M1ihu6,E0ihu6,Wyhhu6,Oxhhu6,Gwhhu6}),
    .i1({E1hpw6,Edkhu6,Wbkhu6}),
    .o(Yuhhu6));  // ../RTL/cortexm0ds_logic.v(3114)
  eq_w32 eq1 (
    .i0({M9ohu6,Uilhu6,Nhlhu6,Gglhu6,Zelhu6,Sdlhu6,Lclhu6,Eblhu6,W9lhu6,O8lhu6,G7lhu6,Y5lhu6,Q4lhu6,I3lhu6,A2lhu6,S0lhu6,Kzkhu6,Cykhu6,Uwkhu6,Mvkhu6,Eukhu6,Wskhu6,Orkhu6,Gqkhu6,Yokhu6,Qnkhu6,Imkhu6,Alkhu6,Sjkhu6,Kikhu6,Chkhu6,Ufkhu6}),
    .i1({K7hpw6,Avmhu6,Ttmhu6}),
    .o(Mekhu6));  // ../RTL/cortexm0ds_logic.v(3128)
  eq_w27 eq2 (
    .i0({V0epw6,O0epw6,H0epw6,A0epw6,Tzdpw6,Mzdpw6,Fzdpw6,Yydpw6,Rydpw6,Kydpw6,Dydpw6,Wxdpw6,Pxdpw6,Tugpw6[13:11],Ixdpw6,Tugpw6[9:0]}),
    .i1(Togpw6),
    .o(Wphhu6));  // ../RTL/cortexm0ds_logic.v(3140)
  eq_w27 eq3 (
    .i0({V0epw6,O0epw6,H0epw6,A0epw6,Tzdpw6,Mzdpw6,Fzdpw6,Yydpw6,Rydpw6,Kydpw6,Dydpw6,Wxdpw6,Pxdpw6,Tugpw6[13:11],Ixdpw6,Tugpw6[9:0]}),
    .i1(Gqgpw6),
    .o(Drhhu6));  // ../RTL/cortexm0ds_logic.v(3143)
  eq_w27 eq4 (
    .i0({V0epw6,O0epw6,H0epw6,A0epw6,Tzdpw6,Mzdpw6,Fzdpw6,Yydpw6,Rydpw6,Kydpw6,Dydpw6,Wxdpw6,Pxdpw6,Tugpw6[13:11],Ixdpw6,Tugpw6[9:0]}),
    .i1(Trgpw6),
    .o(Kshhu6));  // ../RTL/cortexm0ds_logic.v(3146)
  eq_w27 eq5 (
    .i0({V0epw6,O0epw6,H0epw6,A0epw6,Tzdpw6,Mzdpw6,Fzdpw6,Yydpw6,Rydpw6,Kydpw6,Dydpw6,Wxdpw6,Pxdpw6,Tugpw6[13:11],Ixdpw6,Tugpw6[9:0]}),
    .i1(Gtgpw6),
    .o(Rthhu6));  // ../RTL/cortexm0ds_logic.v(3149)
  mult_u32_u32_o64 mult0 (
    .i0(Mifpw6),
    .i1(Tgfpw6),
    .o({open_n1,open_n2,open_n3,open_n4,open_n5,open_n6,open_n7,open_n8,open_n9,open_n10,open_n11,open_n12,open_n13,open_n14,open_n15,open_n16,open_n17,open_n18,open_n19,open_n20,open_n21,open_n22,open_n23,open_n24,open_n25,open_n26,open_n27,open_n28,open_n29,open_n30,open_n31,open_n32,Affpw6}));  // ../RTL/cortexm0ds_logic.v(3158)
  binary_mux_s1_w19 mux0 (
    .i0({Jshpw6[30],Jshpw6[28:11]}),
    .i1({Rx0iu6,V0epw6,O0epw6,H0epw6,A0epw6,Tzdpw6,Mzdpw6,Fzdpw6,Yydpw6,Rydpw6,Kydpw6,Dydpw6,Wxdpw6,Pxdpw6,Tugpw6[13:11],Ixdpw6,Tugpw6[9]}),
    .sel(Ze9iu6),
    .o({HADDR[30],HADDR[28:11]}));  // ../RTL/cortexm0ds_logic.v(15401)
  binary_mux_s1_w11 mux1 (
    .i0({Ef1iu6,Dx0iu6,Tugpw6[8:0]}),
    .i1({Jshpw6[31],Jshpw6[29],Jshpw6[10:4],I47iu6,P47iu6}),
    .sel(Xg6iu6),
    .o({HADDR[31],HADDR[29],HADDR[10:2]}));  // ../RTL/cortexm0ds_logic.v(15250)
  add_pu24_mu24_o24 sub0 (
    .i0(Tzfpw6),
    .i1(24'b000000000000000000000001),
    .o(L6gpw6));  // ../RTL/cortexm0ds_logic.v(3150)
  add_pu9_mu9_o9 sub1 (
    .i0({Vnfpw6,X5phu6}),
    .i1(9'b000000001),
    .o({Xlfpw6,open_n33}));  // ../RTL/cortexm0ds_logic.v(3151)
  buf u10 (TDO, 1'b0);  // ../RTL/cortexm0ds_logic.v(1733)
  buf u100 (E5ehu6, Fpnpw6);  // ../RTL/cortexm0ds_logic.v(1879)
  buf u1000 (R4gpw6[49], Wu3bx6);  // ../RTL/cortexm0ds_logic.v(2815)
  and u10000 (n2651, Jo4ju6, vis_r14_o[4]);  // ../RTL/cortexm0ds_logic.v(9404)
  not u10001 (Co4ju6, n2651);  // ../RTL/cortexm0ds_logic.v(9404)
  and u10002 (Vn4ju6, Qo4ju6, Xo4ju6);  // ../RTL/cortexm0ds_logic.v(9405)
  and u10003 (n2652, Ep4ju6, vis_psp_o[2]);  // ../RTL/cortexm0ds_logic.v(9406)
  not u10004 (Xo4ju6, n2652);  // ../RTL/cortexm0ds_logic.v(9406)
  and u10005 (n2653, Lp4ju6, vis_msp_o[2]);  // ../RTL/cortexm0ds_logic.v(9407)
  not u10006 (Qo4ju6, n2653);  // ../RTL/cortexm0ds_logic.v(9407)
  and u10007 (Hn4ju6, Sp4ju6, Zp4ju6);  // ../RTL/cortexm0ds_logic.v(9408)
  and u10008 (n2654, Gq4ju6, vis_r12_o[4]);  // ../RTL/cortexm0ds_logic.v(9409)
  not u10009 (Zp4ju6, n2654);  // ../RTL/cortexm0ds_logic.v(9409)
  buf u1001 (R4gpw6[50], Yw3bx6);  // ../RTL/cortexm0ds_logic.v(2815)
  and u10010 (n2655, Nq4ju6, vis_r11_o[4]);  // ../RTL/cortexm0ds_logic.v(9410)
  not u10011 (Sp4ju6, n2655);  // ../RTL/cortexm0ds_logic.v(9410)
  and u10012 (Tm4ju6, Uq4ju6, Br4ju6);  // ../RTL/cortexm0ds_logic.v(9411)
  and u10013 (Br4ju6, Ir4ju6, Pr4ju6);  // ../RTL/cortexm0ds_logic.v(9412)
  and u10014 (n2656, Wr4ju6, vis_r10_o[4]);  // ../RTL/cortexm0ds_logic.v(9413)
  not u10015 (Pr4ju6, n2656);  // ../RTL/cortexm0ds_logic.v(9413)
  and u10016 (n2657, Ds4ju6, vis_r9_o[4]);  // ../RTL/cortexm0ds_logic.v(9414)
  not u10017 (Ir4ju6, n2657);  // ../RTL/cortexm0ds_logic.v(9414)
  and u10018 (Uq4ju6, D50iu6, Ks4ju6);  // ../RTL/cortexm0ds_logic.v(9415)
  and u10019 (n2658, Rs4ju6, vis_r8_o[4]);  // ../RTL/cortexm0ds_logic.v(9416)
  buf u1002 (R4gpw6[51], Az3bx6);  // ../RTL/cortexm0ds_logic.v(2815)
  not u10020 (Ks4ju6, n2658);  // ../RTL/cortexm0ds_logic.v(9416)
  not u10021 (V3iiu6, Fkfpw6[4]);  // ../RTL/cortexm0ds_logic.v(9417)
  and u10022 (n2659, Ys4ju6, Qbfpw6[4]);  // ../RTL/cortexm0ds_logic.v(9418)
  not u10023 (Yl4ju6, n2659);  // ../RTL/cortexm0ds_logic.v(9418)
  or u10024 (n2660, Ft4ju6, Mt4ju6);  // ../RTL/cortexm0ds_logic.v(9419)
  not u10025 (Rl4ju6, n2660);  // ../RTL/cortexm0ds_logic.v(9419)
  AL_MUX u10026 (
    .i0(Ys4ju6),
    .i1(Tt4ju6),
    .sel(Qbfpw6[4]),
    .o(Ft4ju6));  // ../RTL/cortexm0ds_logic.v(9420)
  buf u10027 (Bagpw6[10], Tptpw6);  // ../RTL/cortexm0ds_logic.v(2680)
  buf u10028 (Bagpw6[17], Yjupw6);  // ../RTL/cortexm0ds_logic.v(2680)
  and u10029 (n2662, Ou4ju6, Vu4ju6);  // ../RTL/cortexm0ds_logic.v(9422)
  buf u1003 (R4gpw6[52], Jdgbx6);  // ../RTL/cortexm0ds_logic.v(2815)
  not u10030 (Au4ju6, n2662);  // ../RTL/cortexm0ds_logic.v(9422)
  and u10031 (Vu4ju6, Cv4ju6, Jv4ju6);  // ../RTL/cortexm0ds_logic.v(9423)
  or u10032 (Jv4ju6, B5kiu6, Qv4ju6);  // ../RTL/cortexm0ds_logic.v(9424)
  and u10033 (n2663, S8fpw6[4], Xv4ju6);  // ../RTL/cortexm0ds_logic.v(9425)
  not u10034 (Cv4ju6, n2663);  // ../RTL/cortexm0ds_logic.v(9425)
  and u10035 (Ou4ju6, Ew4ju6, Lw4ju6);  // ../RTL/cortexm0ds_logic.v(9426)
  and u10036 (n2664, Sw4ju6, Zw4ju6);  // ../RTL/cortexm0ds_logic.v(9427)
  not u10037 (Lw4ju6, n2664);  // ../RTL/cortexm0ds_logic.v(9427)
  or u10038 (Ew4ju6, V4aiu6, Gx4ju6);  // ../RTL/cortexm0ds_logic.v(9428)
  and u10039 (Dl4ju6, Nx4ju6, Ux4ju6);  // ../RTL/cortexm0ds_logic.v(9429)
  buf u1004 (R4gpw6[53], C14bx6);  // ../RTL/cortexm0ds_logic.v(2815)
  and u10040 (n2665, By4ju6, Eafpw6[4]);  // ../RTL/cortexm0ds_logic.v(9430)
  not u10041 (Ux4ju6, n2665);  // ../RTL/cortexm0ds_logic.v(9430)
  and u10042 (n2666, Iy4ju6, Zw4ju6);  // ../RTL/cortexm0ds_logic.v(9431)
  not u10043 (Nx4ju6, n2666);  // ../RTL/cortexm0ds_logic.v(9431)
  and u10044 (Ibliu6, Py4ju6, Wy4ju6);  // ../RTL/cortexm0ds_logic.v(9432)
  and u10045 (Wy4ju6, Dz4ju6, Kz4ju6);  // ../RTL/cortexm0ds_logic.v(9433)
  or u10046 (n2667, Affpw6[0], Wk4ju6);  // ../RTL/cortexm0ds_logic.v(9434)
  not u10047 (Kz4ju6, n2667);  // ../RTL/cortexm0ds_logic.v(9434)
  and u10048 (Dz4ju6, Rz4ju6, Yz4ju6);  // ../RTL/cortexm0ds_logic.v(9435)
  and u10049 (n2668, F05ju6, M05ju6);  // ../RTL/cortexm0ds_logic.v(9436)
  buf u1005 (R4gpw6[54], E34bx6);  // ../RTL/cortexm0ds_logic.v(2815)
  not u10050 (Yz4ju6, n2668);  // ../RTL/cortexm0ds_logic.v(9436)
  or u10051 (n2669, Qjoiu6, S8fpw6[2]);  // ../RTL/cortexm0ds_logic.v(9437)
  not u10052 (M05ju6, n2669);  // ../RTL/cortexm0ds_logic.v(9437)
  and u10053 (F05ju6, T05ju6, vis_primask_o);  // ../RTL/cortexm0ds_logic.v(9438)
  and u10054 (n2670, Pk4ju6, vis_ipsr_o[0]);  // ../RTL/cortexm0ds_logic.v(9439)
  not u10055 (Rz4ju6, n2670);  // ../RTL/cortexm0ds_logic.v(9439)
  and u10056 (Py4ju6, A15ju6, H15ju6);  // ../RTL/cortexm0ds_logic.v(9440)
  AL_MUX u10057 (
    .i0(O15ju6),
    .i1(V15ju6),
    .sel(Go0iu6),
    .o(H15ju6));  // ../RTL/cortexm0ds_logic.v(9441)
  or u10058 (n2671, C25ju6, Mt4ju6);  // ../RTL/cortexm0ds_logic.v(9442)
  not u10059 (V15ju6, n2671);  // ../RTL/cortexm0ds_logic.v(9442)
  buf u1006 (R4gpw6[55], G54bx6);  // ../RTL/cortexm0ds_logic.v(2815)
  AL_MUX u10060 (
    .i0(Ys4ju6),
    .i1(Tt4ju6),
    .sel(Qbfpw6[0]),
    .o(C25ju6));  // ../RTL/cortexm0ds_logic.v(9443)
  and u10061 (n2672, Ys4ju6, Qbfpw6[0]);  // ../RTL/cortexm0ds_logic.v(9444)
  not u10062 (O15ju6, n2672);  // ../RTL/cortexm0ds_logic.v(9444)
  buf u10063 (Bagpw6[14], Pdxax6);  // ../RTL/cortexm0ds_logic.v(2680)
  buf u10064 (Bagpw6[21], Rhkpw6);  // ../RTL/cortexm0ds_logic.v(2680)
  and u10065 (n2673, Q25ju6, X25ju6);  // ../RTL/cortexm0ds_logic.v(9446)
  not u10066 (J25ju6, n2673);  // ../RTL/cortexm0ds_logic.v(9446)
  and u10067 (n2674, S8fpw6[0], E35ju6);  // ../RTL/cortexm0ds_logic.v(9447)
  not u10068 (X25ju6, n2674);  // ../RTL/cortexm0ds_logic.v(9447)
  and u10069 (n2675, Sw4ju6, L35ju6);  // ../RTL/cortexm0ds_logic.v(9448)
  buf u1007 (R4gpw6[56], Pz9bx6);  // ../RTL/cortexm0ds_logic.v(2815)
  not u10070 (Q25ju6, n2675);  // ../RTL/cortexm0ds_logic.v(9448)
  and u10071 (A15ju6, S35ju6, Z35ju6);  // ../RTL/cortexm0ds_logic.v(9449)
  and u10072 (n2676, By4ju6, Eafpw6[0]);  // ../RTL/cortexm0ds_logic.v(9450)
  not u10073 (Z35ju6, n2676);  // ../RTL/cortexm0ds_logic.v(9450)
  and u10074 (n2677, Iy4ju6, L35ju6);  // ../RTL/cortexm0ds_logic.v(9451)
  not u10075 (S35ju6, n2677);  // ../RTL/cortexm0ds_logic.v(9451)
  and u10076 (Zi4ju6, K5liu6, Bbliu6);  // ../RTL/cortexm0ds_logic.v(9452)
  and u10077 (Bbliu6, G45ju6, N45ju6);  // ../RTL/cortexm0ds_logic.v(9453)
  and u10078 (N45ju6, U45ju6, B55ju6);  // ../RTL/cortexm0ds_logic.v(9454)
  and u10079 (n2678, vis_apsr_o[3], I55ju6);  // ../RTL/cortexm0ds_logic.v(9455)
  buf u1008 (R4gpw6[57], Sn4bx6);  // ../RTL/cortexm0ds_logic.v(2815)
  not u10080 (B55ju6, n2678);  // ../RTL/cortexm0ds_logic.v(9455)
  or u10081 (n2679, Affpw6[31], Wk4ju6);  // ../RTL/cortexm0ds_logic.v(9456)
  not u10082 (U45ju6, n2679);  // ../RTL/cortexm0ds_logic.v(9456)
  and u10083 (G45ju6, P55ju6, W55ju6);  // ../RTL/cortexm0ds_logic.v(9457)
  AL_MUX u10084 (
    .i0(D65ju6),
    .i1(K65ju6),
    .sel(To2ju6),
    .o(W55ju6));  // ../RTL/cortexm0ds_logic.v(9458)
  not u10085 (To2ju6, R65ju6);  // ../RTL/cortexm0ds_logic.v(9459)
  or u10086 (n2680, Y65ju6, Mt4ju6);  // ../RTL/cortexm0ds_logic.v(9460)
  not u10087 (K65ju6, n2680);  // ../RTL/cortexm0ds_logic.v(9460)
  AL_MUX u10088 (
    .i0(Tt4ju6),
    .i1(Ys4ju6),
    .sel(Nl2ju6),
    .o(Y65ju6));  // ../RTL/cortexm0ds_logic.v(9461)
  not u10089 (Nl2ju6, D5epw6);  // ../RTL/cortexm0ds_logic.v(9462)
  buf u1009 (R4gpw6[58], Up4bx6);  // ../RTL/cortexm0ds_logic.v(2815)
  and u10090 (n2681, Ys4ju6, D5epw6);  // ../RTL/cortexm0ds_logic.v(9463)
  not u10091 (D65ju6, n2681);  // ../RTL/cortexm0ds_logic.v(9463)
  or u10092 (D5epw6, F75ju6, M75ju6);  // ../RTL/cortexm0ds_logic.v(9464)
  AL_MUX u10093 (
    .i0(T75ju6),
    .i1(A85ju6),
    .sel(Aioiu6),
    .o(F75ju6));  // ../RTL/cortexm0ds_logic.v(9465)
  and u10094 (P55ju6, H85ju6, O85ju6);  // ../RTL/cortexm0ds_logic.v(9466)
  and u10095 (n2682, By4ju6, Eafpw6[31]);  // ../RTL/cortexm0ds_logic.v(9467)
  not u10096 (O85ju6, n2682);  // ../RTL/cortexm0ds_logic.v(9467)
  and u10097 (n2683, Iy4ju6, Aioiu6);  // ../RTL/cortexm0ds_logic.v(9468)
  not u10098 (H85ju6, n2683);  // ../RTL/cortexm0ds_logic.v(9468)
  and u10099 (K5liu6, V85ju6, C95ju6);  // ../RTL/cortexm0ds_logic.v(9469)
  buf u101 (Bagpw6[0], M6rpw6);  // ../RTL/cortexm0ds_logic.v(2680)
  buf u1010 (R4gpw6[59], Wr4bx6);  // ../RTL/cortexm0ds_logic.v(2815)
  and u10100 (C95ju6, J95ju6, Q95ju6);  // ../RTL/cortexm0ds_logic.v(9470)
  and u10101 (n2684, X95ju6, Sg0iu6);  // ../RTL/cortexm0ds_logic.v(9471)
  not u10102 (Q95ju6, n2684);  // ../RTL/cortexm0ds_logic.v(9471)
  and u10103 (X95ju6, Ys4ju6, Qbfpw6[30]);  // ../RTL/cortexm0ds_logic.v(9472)
  or u10104 (n2685, Affpw6[30], Ea5ju6);  // ../RTL/cortexm0ds_logic.v(9473)
  not u10105 (J95ju6, n2685);  // ../RTL/cortexm0ds_logic.v(9473)
  and u10106 (Ea5ju6, Iy4ju6, T6liu6);  // ../RTL/cortexm0ds_logic.v(9474)
  and u10107 (V85ju6, La5ju6, Sa5ju6);  // ../RTL/cortexm0ds_logic.v(9475)
  and u10108 (n2686, Za5ju6, Gb5ju6);  // ../RTL/cortexm0ds_logic.v(9476)
  not u10109 (Sa5ju6, n2686);  // ../RTL/cortexm0ds_logic.v(9476)
  buf u1011 (Odgpw6[0], U31bx6);  // ../RTL/cortexm0ds_logic.v(2789)
  or u10110 (Gb5ju6, Nb5ju6, Ub5ju6);  // ../RTL/cortexm0ds_logic.v(9477)
  or u10111 (Nb5ju6, Mt4ju6, Qbfpw6[30]);  // ../RTL/cortexm0ds_logic.v(9478)
  and u10112 (n2687, Bc5ju6, Ic5ju6);  // ../RTL/cortexm0ds_logic.v(9479)
  not u10113 (Za5ju6, n2687);  // ../RTL/cortexm0ds_logic.v(9479)
  or u10114 (Bc5ju6, Sg0iu6, Pc5ju6);  // ../RTL/cortexm0ds_logic.v(9480)
  and u10115 (Pc5ju6, Wc5ju6, Qbfpw6[30]);  // ../RTL/cortexm0ds_logic.v(9481)
  not u10116 (Idfpw6[1], n114[0]);  // ../RTL/cortexm0ds_logic.v(3453)
  AL_MUX u10117 (
    .i0(T75ju6),
    .i1(A85ju6),
    .sel(T6liu6),
    .o(Dd5ju6));  // ../RTL/cortexm0ds_logic.v(9483)
  and u10118 (La5ju6, Kd5ju6, Rd5ju6);  // ../RTL/cortexm0ds_logic.v(9484)
  and u10119 (n2688, vis_apsr_o[2], I55ju6);  // ../RTL/cortexm0ds_logic.v(9485)
  buf u1012 (Gmhpw6[0], Vrkbx6[1]);  // ../RTL/cortexm0ds_logic.v(3109)
  not u10120 (Rd5ju6, n2688);  // ../RTL/cortexm0ds_logic.v(9485)
  and u10121 (n2689, By4ju6, Eafpw6[30]);  // ../RTL/cortexm0ds_logic.v(9486)
  not u10122 (Kd5ju6, n2689);  // ../RTL/cortexm0ds_logic.v(9486)
  and u10123 (Li4ju6, Yd5ju6, Fe5ju6);  // ../RTL/cortexm0ds_logic.v(9487)
  and u10124 (Fe5ju6, Cgkiu6, Evkiu6);  // ../RTL/cortexm0ds_logic.v(9488)
  and u10125 (Evkiu6, Me5ju6, Te5ju6);  // ../RTL/cortexm0ds_logic.v(9489)
  and u10126 (Te5ju6, Af5ju6, Hf5ju6);  // ../RTL/cortexm0ds_logic.v(9490)
  and u10127 (n2690, By4ju6, Eafpw6[23]);  // ../RTL/cortexm0ds_logic.v(9491)
  not u10128 (Hf5ju6, n2690);  // ../RTL/cortexm0ds_logic.v(9491)
  or u10129 (n2691, Affpw6[23], Of5ju6);  // ../RTL/cortexm0ds_logic.v(9492)
  buf u1013 (A4khu6, Ntkbx6[0]);  // ../RTL/cortexm0ds_logic.v(3123)
  not u10130 (Af5ju6, n2691);  // ../RTL/cortexm0ds_logic.v(9492)
  or u10131 (n2692, Vf5ju6, Fk0iu6);  // ../RTL/cortexm0ds_logic.v(9493)
  not u10132 (Of5ju6, n2692);  // ../RTL/cortexm0ds_logic.v(9493)
  AL_MUX u10133 (
    .i0(Cg5ju6),
    .i1(Wc5ju6),
    .sel(Qbfpw6[23]),
    .o(Vf5ju6));  // ../RTL/cortexm0ds_logic.v(9494)
  and u10134 (Me5ju6, Jg5ju6, Qg5ju6);  // ../RTL/cortexm0ds_logic.v(9495)
  and u10135 (n2693, Iy4ju6, Xg5ju6);  // ../RTL/cortexm0ds_logic.v(9496)
  not u10136 (Qg5ju6, n2693);  // ../RTL/cortexm0ds_logic.v(9496)
  and u10137 (n2694, Ub5ju6, Eh5ju6);  // ../RTL/cortexm0ds_logic.v(9497)
  not u10138 (Jg5ju6, n2694);  // ../RTL/cortexm0ds_logic.v(9497)
  and u10139 (n2695, Lh5ju6, Ic5ju6);  // ../RTL/cortexm0ds_logic.v(9498)
  not u1014 (n6026, Knmhu6);  // ../RTL/cortexm0ds_logic.v(3132)
  not u10140 (Eh5ju6, n2695);  // ../RTL/cortexm0ds_logic.v(9498)
  and u10141 (n2696, Fk0iu6, Qbfpw6[23]);  // ../RTL/cortexm0ds_logic.v(9499)
  not u10142 (Lh5ju6, n2696);  // ../RTL/cortexm0ds_logic.v(9499)
  not u10143 (Qbfpw6[0], n2661[0]);  // ../RTL/cortexm0ds_logic.v(9500)
  and u10144 (Idfpw6[0], Go0iu6, Oe0iu6);  // ../RTL/cortexm0ds_logic.v(9222)
  or u10145 (Sh5ju6, Zh5ju6, Gi5ju6);  // ../RTL/cortexm0ds_logic.v(9501)
  AL_MUX u10146 (
    .i0(Ni5ju6),
    .i1(Ui5ju6),
    .sel(D7fpw6[13]),
    .o(Gi5ju6));  // ../RTL/cortexm0ds_logic.v(9502)
  or u10147 (Qbaju6, Gx4ju6, S8fpw6[11]);  // ../RTL/cortexm0ds_logic.v(9503)
  not u10148 (Ni5ju6, Qbaju6);  // ../RTL/cortexm0ds_logic.v(9503)
  and u10149 (n2697, Bj5ju6, Ij5ju6);  // ../RTL/cortexm0ds_logic.v(9504)
  buf u1015 (R4gpw6[33], H4zax6);  // ../RTL/cortexm0ds_logic.v(2815)
  not u10150 (Zh5ju6, n2697);  // ../RTL/cortexm0ds_logic.v(9504)
  and u10151 (n2698, Sw4ju6, Xg5ju6);  // ../RTL/cortexm0ds_logic.v(9505)
  not u10152 (Bj5ju6, n2698);  // ../RTL/cortexm0ds_logic.v(9505)
  and u10153 (Cgkiu6, Pj5ju6, Wj5ju6);  // ../RTL/cortexm0ds_logic.v(9506)
  and u10154 (Wj5ju6, Dk5ju6, Kk5ju6);  // ../RTL/cortexm0ds_logic.v(9507)
  or u10155 (n2699, Affpw6[2], Rk5ju6);  // ../RTL/cortexm0ds_logic.v(9508)
  not u10156 (Kk5ju6, n2699);  // ../RTL/cortexm0ds_logic.v(9508)
  and u10157 (Rk5ju6, Yk5ju6, L8ehu6);  // ../RTL/cortexm0ds_logic.v(9509)
  and u10158 (Yk5ju6, P8oiu6, H6ghu6);  // ../RTL/cortexm0ds_logic.v(9510)
  and u10159 (Dk5ju6, Fl5ju6, Ml5ju6);  // ../RTL/cortexm0ds_logic.v(9511)
  buf u1016 (Dmmhu6, Nvkbx6[0]);  // ../RTL/cortexm0ds_logic.v(3137)
  and u10160 (n2700, Pk4ju6, vis_ipsr_o[2]);  // ../RTL/cortexm0ds_logic.v(9512)
  not u10161 (Ml5ju6, n2700);  // ../RTL/cortexm0ds_logic.v(9512)
  and u10162 (n2701, By4ju6, Eafpw6[2]);  // ../RTL/cortexm0ds_logic.v(9513)
  not u10163 (Fl5ju6, n2701);  // ../RTL/cortexm0ds_logic.v(9513)
  and u10164 (Pj5ju6, Tl5ju6, Am5ju6);  // ../RTL/cortexm0ds_logic.v(9514)
  AL_MUX u10165 (
    .i0(Hm5ju6),
    .i1(Om5ju6),
    .sel(Gh0iu6),
    .o(Am5ju6));  // ../RTL/cortexm0ds_logic.v(9515)
  AL_MUX u10166 (
    .i0(Vm5ju6),
    .i1(Fkfpw6[2]),
    .sel(Cn5ju6),
    .o(Gh0iu6));  // ../RTL/cortexm0ds_logic.v(9516)
  and u10167 (n2702, Jn5ju6, Qn5ju6);  // ../RTL/cortexm0ds_logic.v(9517)
  not u10168 (Vm5ju6, n2702);  // ../RTL/cortexm0ds_logic.v(9517)
  and u10169 (Qn5ju6, Xn5ju6, Eo5ju6);  // ../RTL/cortexm0ds_logic.v(9518)
  buf u1017 (R4gpw6[32], V5abx6);  // ../RTL/cortexm0ds_logic.v(2815)
  and u10170 (Eo5ju6, Lo5ju6, So5ju6);  // ../RTL/cortexm0ds_logic.v(9519)
  and u10171 (n2703, Jo4ju6, vis_r14_o[2]);  // ../RTL/cortexm0ds_logic.v(9520)
  not u10172 (So5ju6, n2703);  // ../RTL/cortexm0ds_logic.v(9520)
  and u10173 (Lo5ju6, Zo5ju6, Gp5ju6);  // ../RTL/cortexm0ds_logic.v(9521)
  and u10174 (n2704, Ep4ju6, vis_psp_o[0]);  // ../RTL/cortexm0ds_logic.v(9522)
  not u10175 (Gp5ju6, n2704);  // ../RTL/cortexm0ds_logic.v(9522)
  and u10176 (n2705, Lp4ju6, vis_msp_o[0]);  // ../RTL/cortexm0ds_logic.v(9523)
  not u10177 (Zo5ju6, n2705);  // ../RTL/cortexm0ds_logic.v(9523)
  and u10178 (Xn5ju6, Np5ju6, Up5ju6);  // ../RTL/cortexm0ds_logic.v(9524)
  and u10179 (n2706, Gq4ju6, vis_r12_o[2]);  // ../RTL/cortexm0ds_logic.v(9525)
  buf u1018 (Eafpw6[0], Nxkbx6[1]);  // ../RTL/cortexm0ds_logic.v(3167)
  not u10180 (Up5ju6, n2706);  // ../RTL/cortexm0ds_logic.v(9525)
  and u10181 (n2707, Nq4ju6, vis_r11_o[2]);  // ../RTL/cortexm0ds_logic.v(9526)
  not u10182 (Np5ju6, n2707);  // ../RTL/cortexm0ds_logic.v(9526)
  and u10183 (Jn5ju6, Bq5ju6, Iq5ju6);  // ../RTL/cortexm0ds_logic.v(9527)
  and u10184 (Iq5ju6, Pq5ju6, Wq5ju6);  // ../RTL/cortexm0ds_logic.v(9528)
  and u10185 (n2708, Wr4ju6, vis_r10_o[2]);  // ../RTL/cortexm0ds_logic.v(9529)
  not u10186 (Wq5ju6, n2708);  // ../RTL/cortexm0ds_logic.v(9529)
  and u10187 (n2709, Ds4ju6, vis_r9_o[2]);  // ../RTL/cortexm0ds_logic.v(9530)
  not u10188 (Pq5ju6, n2709);  // ../RTL/cortexm0ds_logic.v(9530)
  and u10189 (Bq5ju6, F60iu6, Dr5ju6);  // ../RTL/cortexm0ds_logic.v(9531)
  and u1019 (n0, L4yhu6, S4yhu6);  // ../RTL/cortexm0ds_logic.v(3177)
  and u10190 (n2710, Rs4ju6, vis_r8_o[2]);  // ../RTL/cortexm0ds_logic.v(9532)
  not u10191 (Dr5ju6, n2710);  // ../RTL/cortexm0ds_logic.v(9532)
  or u10192 (n2711, Kr5ju6, Mt4ju6);  // ../RTL/cortexm0ds_logic.v(9533)
  not u10193 (Om5ju6, n2711);  // ../RTL/cortexm0ds_logic.v(9533)
  AL_MUX u10194 (
    .i0(Ys4ju6),
    .i1(Tt4ju6),
    .sel(Qbfpw6[2]),
    .o(Kr5ju6));  // ../RTL/cortexm0ds_logic.v(9534)
  and u10195 (n2712, Ys4ju6, Qbfpw6[2]);  // ../RTL/cortexm0ds_logic.v(9535)
  not u10196 (Hm5ju6, n2712);  // ../RTL/cortexm0ds_logic.v(9535)
  buf u10197 (Bagpw6[12], Tyipw6);  // ../RTL/cortexm0ds_logic.v(2680)
  buf u10198 (Bagpw6[19], Hhvpw6);  // ../RTL/cortexm0ds_logic.v(2680)
  and u10199 (n2713, Yr5ju6, Fs5ju6);  // ../RTL/cortexm0ds_logic.v(9537)
  buf u102 (vis_ipsr_o[0], Eliax6);  // ../RTL/cortexm0ds_logic.v(1815)
  not u1020 (I5nhu6, n0);  // ../RTL/cortexm0ds_logic.v(3177)
  not u10200 (Rr5ju6, n2713);  // ../RTL/cortexm0ds_logic.v(9537)
  and u10201 (Fs5ju6, Ms5ju6, Ts5ju6);  // ../RTL/cortexm0ds_logic.v(9538)
  and u10202 (n2714, S8fpw6[2], E35ju6);  // ../RTL/cortexm0ds_logic.v(9539)
  not u10203 (Ts5ju6, n2714);  // ../RTL/cortexm0ds_logic.v(9539)
  or u10204 (Ms5ju6, Je8iu6, Qv4ju6);  // ../RTL/cortexm0ds_logic.v(9540)
  and u10205 (Yr5ju6, At5ju6, Ht5ju6);  // ../RTL/cortexm0ds_logic.v(9541)
  and u10206 (n2715, Sw4ju6, Ot5ju6);  // ../RTL/cortexm0ds_logic.v(9542)
  not u10207 (Ht5ju6, n2715);  // ../RTL/cortexm0ds_logic.v(9542)
  or u10208 (At5ju6, Ccaiu6, Gx4ju6);  // ../RTL/cortexm0ds_logic.v(9543)
  and u10209 (Tl5ju6, Vt5ju6, Cu5ju6);  // ../RTL/cortexm0ds_logic.v(9544)
  and u1021 (n1, Z4yhu6, SWDOEN);  // ../RTL/cortexm0ds_logic.v(3178)
  and u10210 (n2716, Iy4ju6, Ot5ju6);  // ../RTL/cortexm0ds_logic.v(9545)
  not u10211 (Cu5ju6, n2716);  // ../RTL/cortexm0ds_logic.v(9545)
  and u10212 (n2717, vis_control_o, Wk4ju6);  // ../RTL/cortexm0ds_logic.v(9546)
  not u10213 (Vt5ju6, n2717);  // ../RTL/cortexm0ds_logic.v(9546)
  and u10214 (Yd5ju6, Lokiu6, Dkkiu6);  // ../RTL/cortexm0ds_logic.v(9547)
  and u10215 (Dkkiu6, Ju5ju6, Qu5ju6);  // ../RTL/cortexm0ds_logic.v(9548)
  and u10216 (Qu5ju6, Xu5ju6, Ev5ju6);  // ../RTL/cortexm0ds_logic.v(9549)
  and u10217 (n2718, By4ju6, Eafpw6[3]);  // ../RTL/cortexm0ds_logic.v(9550)
  not u10218 (Ev5ju6, n2718);  // ../RTL/cortexm0ds_logic.v(9550)
  or u10219 (n2719, Affpw6[3], Lv5ju6);  // ../RTL/cortexm0ds_logic.v(9551)
  not u1022 (S4yhu6, n1);  // ../RTL/cortexm0ds_logic.v(3178)
  not u10220 (Xu5ju6, n2719);  // ../RTL/cortexm0ds_logic.v(9551)
  and u10221 (Lv5ju6, Pk4ju6, vis_ipsr_o[3]);  // ../RTL/cortexm0ds_logic.v(9552)
  and u10222 (Ju5ju6, Sv5ju6, Zv5ju6);  // ../RTL/cortexm0ds_logic.v(9553)
  AL_MUX u10223 (
    .i0(Gw5ju6),
    .i1(Nw5ju6),
    .sel(Lg0iu6),
    .o(Zv5ju6));  // ../RTL/cortexm0ds_logic.v(9554)
  AL_MUX u10224 (
    .i0(Wjkiu6),
    .i1(Uw5ju6),
    .sel(Mm4ju6),
    .o(Lg0iu6));  // ../RTL/cortexm0ds_logic.v(9555)
  and u10225 (Uw5ju6, Bx5ju6, Ix5ju6);  // ../RTL/cortexm0ds_logic.v(9556)
  and u10226 (Ix5ju6, Px5ju6, Wx5ju6);  // ../RTL/cortexm0ds_logic.v(9557)
  and u10227 (Wx5ju6, Dy5ju6, Ky5ju6);  // ../RTL/cortexm0ds_logic.v(9558)
  and u10228 (n2720, Jo4ju6, vis_r14_o[3]);  // ../RTL/cortexm0ds_logic.v(9559)
  not u10229 (Ky5ju6, n2720);  // ../RTL/cortexm0ds_logic.v(9559)
  and u1023 (L4yhu6, G5yhu6, N5yhu6);  // ../RTL/cortexm0ds_logic.v(3179)
  and u10230 (Dy5ju6, Ry5ju6, Yy5ju6);  // ../RTL/cortexm0ds_logic.v(9560)
  and u10231 (n2721, Ep4ju6, vis_psp_o[1]);  // ../RTL/cortexm0ds_logic.v(9561)
  not u10232 (Yy5ju6, n2721);  // ../RTL/cortexm0ds_logic.v(9561)
  and u10233 (n2722, Lp4ju6, vis_msp_o[1]);  // ../RTL/cortexm0ds_logic.v(9562)
  not u10234 (Ry5ju6, n2722);  // ../RTL/cortexm0ds_logic.v(9562)
  and u10235 (Px5ju6, Fz5ju6, Mz5ju6);  // ../RTL/cortexm0ds_logic.v(9563)
  and u10236 (n2723, Gq4ju6, vis_r12_o[3]);  // ../RTL/cortexm0ds_logic.v(9564)
  not u10237 (Mz5ju6, n2723);  // ../RTL/cortexm0ds_logic.v(9564)
  and u10238 (n2724, Nq4ju6, vis_r11_o[3]);  // ../RTL/cortexm0ds_logic.v(9565)
  not u10239 (Fz5ju6, n2724);  // ../RTL/cortexm0ds_logic.v(9565)
  and u1024 (n2, U5yhu6, B6yhu6);  // ../RTL/cortexm0ds_logic.v(3180)
  and u10240 (Bx5ju6, Tz5ju6, A06ju6);  // ../RTL/cortexm0ds_logic.v(9566)
  and u10241 (A06ju6, H06ju6, O06ju6);  // ../RTL/cortexm0ds_logic.v(9567)
  and u10242 (n2725, Wr4ju6, vis_r10_o[3]);  // ../RTL/cortexm0ds_logic.v(9568)
  not u10243 (O06ju6, n2725);  // ../RTL/cortexm0ds_logic.v(9568)
  and u10244 (n2726, Ds4ju6, vis_r9_o[3]);  // ../RTL/cortexm0ds_logic.v(9569)
  not u10245 (H06ju6, n2726);  // ../RTL/cortexm0ds_logic.v(9569)
  and u10246 (Tz5ju6, K50iu6, V06ju6);  // ../RTL/cortexm0ds_logic.v(9570)
  and u10247 (n2727, Rs4ju6, vis_r8_o[3]);  // ../RTL/cortexm0ds_logic.v(9571)
  not u10248 (V06ju6, n2727);  // ../RTL/cortexm0ds_logic.v(9571)
  not u10249 (Wjkiu6, Fkfpw6[3]);  // ../RTL/cortexm0ds_logic.v(9572)
  not u1025 (G5yhu6, n2);  // ../RTL/cortexm0ds_logic.v(3180)
  and u10250 (n2728, Ys4ju6, Qbfpw6[3]);  // ../RTL/cortexm0ds_logic.v(9573)
  not u10251 (Nw5ju6, n2728);  // ../RTL/cortexm0ds_logic.v(9573)
  or u10252 (n2729, C16ju6, Mt4ju6);  // ../RTL/cortexm0ds_logic.v(9574)
  not u10253 (Gw5ju6, n2729);  // ../RTL/cortexm0ds_logic.v(9574)
  AL_MUX u10254 (
    .i0(Ys4ju6),
    .i1(Tt4ju6),
    .sel(Qbfpw6[3]),
    .o(C16ju6));  // ../RTL/cortexm0ds_logic.v(9575)
  buf u10255 (Bagpw6[11], Ofmpw6);  // ../RTL/cortexm0ds_logic.v(2680)
  buf u10256 (Bagpw6[18], Lywpw6);  // ../RTL/cortexm0ds_logic.v(2680)
  and u10257 (n2730, Q16ju6, X16ju6);  // ../RTL/cortexm0ds_logic.v(9577)
  not u10258 (J16ju6, n2730);  // ../RTL/cortexm0ds_logic.v(9577)
  and u10259 (X16ju6, E26ju6, L26ju6);  // ../RTL/cortexm0ds_logic.v(9578)
  and u1026 (n3, I6yhu6, P6yhu6);  // ../RTL/cortexm0ds_logic.v(3181)
  or u10260 (L26ju6, Y8biu6, Qv4ju6);  // ../RTL/cortexm0ds_logic.v(9579)
  and u10261 (n2731, S8fpw6[3], Xv4ju6);  // ../RTL/cortexm0ds_logic.v(9580)
  not u10262 (E26ju6, n2731);  // ../RTL/cortexm0ds_logic.v(9580)
  and u10263 (Q16ju6, S26ju6, Z26ju6);  // ../RTL/cortexm0ds_logic.v(9581)
  and u10264 (n2732, Sw4ju6, G36ju6);  // ../RTL/cortexm0ds_logic.v(9582)
  not u10265 (Z26ju6, n2732);  // ../RTL/cortexm0ds_logic.v(9582)
  or u10266 (S26ju6, Prjiu6, Gx4ju6);  // ../RTL/cortexm0ds_logic.v(9583)
  and u10267 (Sv5ju6, N36ju6, U36ju6);  // ../RTL/cortexm0ds_logic.v(9584)
  and u10268 (n2733, Iy4ju6, G36ju6);  // ../RTL/cortexm0ds_logic.v(9585)
  not u10269 (U36ju6, n2733);  // ../RTL/cortexm0ds_logic.v(9585)
  not u1027 (B6yhu6, n3);  // ../RTL/cortexm0ds_logic.v(3181)
  and u10270 (n2734, Hlliu6, Wk4ju6);  // ../RTL/cortexm0ds_logic.v(9586)
  not u10271 (N36ju6, n2734);  // ../RTL/cortexm0ds_logic.v(9586)
  and u10272 (Lokiu6, B46ju6, I46ju6);  // ../RTL/cortexm0ds_logic.v(9587)
  and u10273 (I46ju6, P46ju6, W46ju6);  // ../RTL/cortexm0ds_logic.v(9588)
  and u10274 (n2735, Pk4ju6, vis_ipsr_o[5]);  // ../RTL/cortexm0ds_logic.v(9589)
  not u10275 (W46ju6, n2735);  // ../RTL/cortexm0ds_logic.v(9589)
  or u10276 (n2736, Affpw6[5], Wk4ju6);  // ../RTL/cortexm0ds_logic.v(9590)
  not u10277 (P46ju6, n2736);  // ../RTL/cortexm0ds_logic.v(9590)
  and u10278 (B46ju6, D56ju6, K56ju6);  // ../RTL/cortexm0ds_logic.v(9591)
  AL_MUX u10279 (
    .i0(R56ju6),
    .i1(Y56ju6),
    .sel(Xf0iu6),
    .o(K56ju6));  // ../RTL/cortexm0ds_logic.v(9592)
  and u1028 (n4, W6yhu6, D7yhu6);  // ../RTL/cortexm0ds_logic.v(3182)
  AL_MUX u10280 (
    .i0(Eokiu6),
    .i1(F66ju6),
    .sel(Mm4ju6),
    .o(Xf0iu6));  // ../RTL/cortexm0ds_logic.v(9593)
  and u10281 (F66ju6, M66ju6, T66ju6);  // ../RTL/cortexm0ds_logic.v(9594)
  and u10282 (T66ju6, A76ju6, H76ju6);  // ../RTL/cortexm0ds_logic.v(9595)
  and u10283 (H76ju6, O76ju6, V76ju6);  // ../RTL/cortexm0ds_logic.v(9596)
  and u10284 (n2737, Jo4ju6, vis_r14_o[5]);  // ../RTL/cortexm0ds_logic.v(9597)
  not u10285 (V76ju6, n2737);  // ../RTL/cortexm0ds_logic.v(9597)
  and u10286 (O76ju6, C86ju6, J86ju6);  // ../RTL/cortexm0ds_logic.v(9598)
  and u10287 (n2738, Ep4ju6, vis_psp_o[3]);  // ../RTL/cortexm0ds_logic.v(9599)
  not u10288 (J86ju6, n2738);  // ../RTL/cortexm0ds_logic.v(9599)
  and u10289 (n2739, Lp4ju6, vis_msp_o[3]);  // ../RTL/cortexm0ds_logic.v(9600)
  not u1029 (P6yhu6, n4);  // ../RTL/cortexm0ds_logic.v(3182)
  not u10290 (C86ju6, n2739);  // ../RTL/cortexm0ds_logic.v(9600)
  and u10291 (A76ju6, Q86ju6, X86ju6);  // ../RTL/cortexm0ds_logic.v(9601)
  and u10292 (n2740, Gq4ju6, vis_r12_o[5]);  // ../RTL/cortexm0ds_logic.v(9602)
  not u10293 (X86ju6, n2740);  // ../RTL/cortexm0ds_logic.v(9602)
  and u10294 (n2741, Nq4ju6, vis_r11_o[5]);  // ../RTL/cortexm0ds_logic.v(9603)
  not u10295 (Q86ju6, n2741);  // ../RTL/cortexm0ds_logic.v(9603)
  and u10296 (M66ju6, E96ju6, L96ju6);  // ../RTL/cortexm0ds_logic.v(9604)
  and u10297 (L96ju6, S96ju6, Z96ju6);  // ../RTL/cortexm0ds_logic.v(9605)
  and u10298 (n2742, Wr4ju6, vis_r10_o[5]);  // ../RTL/cortexm0ds_logic.v(9606)
  not u10299 (Z96ju6, n2742);  // ../RTL/cortexm0ds_logic.v(9606)
  buf u103 (R4gpw6[34], J6zax6);  // ../RTL/cortexm0ds_logic.v(2815)
  or u1030 (n5, K7yhu6, Ighpw6[4]);  // ../RTL/cortexm0ds_logic.v(3183)
  and u10300 (n2743, Ds4ju6, vis_r9_o[5]);  // ../RTL/cortexm0ds_logic.v(9607)
  not u10301 (S96ju6, n2743);  // ../RTL/cortexm0ds_logic.v(9607)
  and u10302 (E96ju6, W40iu6, Ga6ju6);  // ../RTL/cortexm0ds_logic.v(9608)
  and u10303 (n2744, Rs4ju6, vis_r8_o[5]);  // ../RTL/cortexm0ds_logic.v(9609)
  not u10304 (Ga6ju6, n2744);  // ../RTL/cortexm0ds_logic.v(9609)
  not u10305 (Eokiu6, Fkfpw6[5]);  // ../RTL/cortexm0ds_logic.v(9610)
  and u10306 (n2745, Ys4ju6, Qbfpw6[5]);  // ../RTL/cortexm0ds_logic.v(9611)
  not u10307 (Y56ju6, n2745);  // ../RTL/cortexm0ds_logic.v(9611)
  or u10308 (n2746, Na6ju6, Mt4ju6);  // ../RTL/cortexm0ds_logic.v(9612)
  not u10309 (R56ju6, n2746);  // ../RTL/cortexm0ds_logic.v(9612)
  not u1031 (D7yhu6, n5);  // ../RTL/cortexm0ds_logic.v(3183)
  AL_MUX u10310 (
    .i0(Ys4ju6),
    .i1(Tt4ju6),
    .sel(Qbfpw6[5]),
    .o(Na6ju6));  // ../RTL/cortexm0ds_logic.v(9613)
  buf u10311 (Bagpw6[9], Tmjbx6);  // ../RTL/cortexm0ds_logic.v(2680)
  buf u10312 (Bagpw6[16], Ujspw6);  // ../RTL/cortexm0ds_logic.v(2680)
  and u10313 (n2747, Bb6ju6, Ib6ju6);  // ../RTL/cortexm0ds_logic.v(9615)
  not u10314 (Ua6ju6, n2747);  // ../RTL/cortexm0ds_logic.v(9615)
  and u10315 (Ib6ju6, Pb6ju6, Wb6ju6);  // ../RTL/cortexm0ds_logic.v(9616)
  or u10316 (Wb6ju6, Cajiu6, Qv4ju6);  // ../RTL/cortexm0ds_logic.v(9617)
  or u10317 (n2748, Dc6ju6, Kc6ju6);  // ../RTL/cortexm0ds_logic.v(9618)
  not u10318 (Qv4ju6, n2748);  // ../RTL/cortexm0ds_logic.v(9618)
  and u10319 (Dc6ju6, H6ghu6, Rc6ju6);  // ../RTL/cortexm0ds_logic.v(9619)
  or u1032 (n6, R7yhu6, Y7yhu6);  // ../RTL/cortexm0ds_logic.v(3184)
  and u10320 (n2749, Yc6ju6, Fd6ju6);  // ../RTL/cortexm0ds_logic.v(9620)
  not u10321 (Rc6ju6, n2749);  // ../RTL/cortexm0ds_logic.v(9620)
  and u10322 (Fd6ju6, Md6ju6, Fmjiu6);  // ../RTL/cortexm0ds_logic.v(9621)
  and u10323 (n2750, Td6ju6, Cyfpw6[7]);  // ../RTL/cortexm0ds_logic.v(9622)
  not u10324 (Md6ju6, n2750);  // ../RTL/cortexm0ds_logic.v(9622)
  and u10325 (Td6ju6, Ae6ju6, Jjhiu6);  // ../RTL/cortexm0ds_logic.v(9623)
  and u10326 (n2751, He6ju6, Oe6ju6);  // ../RTL/cortexm0ds_logic.v(9624)
  not u10327 (Ae6ju6, n2751);  // ../RTL/cortexm0ds_logic.v(9624)
  or u10328 (Oe6ju6, X5oiu6, Tfjiu6);  // ../RTL/cortexm0ds_logic.v(9625)
  and u10329 (Yc6ju6, Ve6ju6, Cf6ju6);  // ../RTL/cortexm0ds_logic.v(9626)
  not u1033 (W6yhu6, n6);  // ../RTL/cortexm0ds_logic.v(3184)
  and u10330 (n2752, Cyfpw6[0], F1jiu6);  // ../RTL/cortexm0ds_logic.v(9627)
  not u10331 (Cf6ju6, n2752);  // ../RTL/cortexm0ds_logic.v(9627)
  or u10332 (F1jiu6, Xzmiu6, Toaiu6);  // ../RTL/cortexm0ds_logic.v(9628)
  and u10333 (n2753, Jf6ju6, Oiaiu6);  // ../RTL/cortexm0ds_logic.v(9629)
  not u10334 (Ve6ju6, n2753);  // ../RTL/cortexm0ds_logic.v(9629)
  and u10335 (n2754, S8fpw6[5], Xv4ju6);  // ../RTL/cortexm0ds_logic.v(9630)
  not u10336 (Pb6ju6, n2754);  // ../RTL/cortexm0ds_logic.v(9630)
  and u10337 (Bb6ju6, Qf6ju6, Xf6ju6);  // ../RTL/cortexm0ds_logic.v(9631)
  and u10338 (n2755, Sw4ju6, Eg6ju6);  // ../RTL/cortexm0ds_logic.v(9632)
  not u10339 (Xf6ju6, n2755);  // ../RTL/cortexm0ds_logic.v(9632)
  buf u1034 (Qofhu6, Ozkbx6[1]);  // ../RTL/cortexm0ds_logic.v(3176)
  or u10340 (Qf6ju6, Gx4ju6, A1kiu6);  // ../RTL/cortexm0ds_logic.v(9633)
  and u10341 (D56ju6, Lg6ju6, Sg6ju6);  // ../RTL/cortexm0ds_logic.v(9634)
  and u10342 (n2756, By4ju6, Eafpw6[5]);  // ../RTL/cortexm0ds_logic.v(9635)
  not u10343 (Sg6ju6, n2756);  // ../RTL/cortexm0ds_logic.v(9635)
  and u10344 (n2757, Iy4ju6, Eg6ju6);  // ../RTL/cortexm0ds_logic.v(9636)
  not u10345 (Lg6ju6, n2757);  // ../RTL/cortexm0ds_logic.v(9636)
  and u10346 (Xh4ju6, Zg6ju6, Gh6ju6);  // ../RTL/cortexm0ds_logic.v(9637)
  and u10347 (Gh6ju6, Nh6ju6, Uh6ju6);  // ../RTL/cortexm0ds_logic.v(9638)
  or u10348 (n2758, Jukiu6, Pqkiu6);  // ../RTL/cortexm0ds_logic.v(9639)
  not u10349 (Uh6ju6, n2758);  // ../RTL/cortexm0ds_logic.v(9639)
  buf u1035 (Ighpw6[0], Bclpw6);  // ../RTL/cortexm0ds_logic.v(1840)
  and u10350 (n2759, Bi6ju6, Ii6ju6);  // ../RTL/cortexm0ds_logic.v(9640)
  not u10351 (Pqkiu6, n2759);  // ../RTL/cortexm0ds_logic.v(9640)
  and u10352 (Ii6ju6, Pi6ju6, Wi6ju6);  // ../RTL/cortexm0ds_logic.v(9641)
  and u10353 (n2760, By4ju6, Eafpw6[6]);  // ../RTL/cortexm0ds_logic.v(9642)
  not u10354 (Wi6ju6, n2760);  // ../RTL/cortexm0ds_logic.v(9642)
  or u10355 (n2761, Affpw6[6], Dj6ju6);  // ../RTL/cortexm0ds_logic.v(9643)
  not u10356 (Pi6ju6, n2761);  // ../RTL/cortexm0ds_logic.v(9643)
  and u10357 (Dj6ju6, Iy4ju6, Kj6ju6);  // ../RTL/cortexm0ds_logic.v(9644)
  and u10358 (Bi6ju6, Rj6ju6, Yj6ju6);  // ../RTL/cortexm0ds_logic.v(9645)
  or u10359 (Yj6ju6, Fk6ju6, Mk6ju6);  // ../RTL/cortexm0ds_logic.v(9646)
  and u1036 (n8, T8yhu6, Fnnhu6);  // ../RTL/cortexm0ds_logic.v(3186)
  AL_MUX u10360 (
    .i0(Cg5ju6),
    .i1(Wc5ju6),
    .sel(E2epw6),
    .o(Fk6ju6));  // ../RTL/cortexm0ds_logic.v(9647)
  and u10361 (n2762, Ub5ju6, Tk6ju6);  // ../RTL/cortexm0ds_logic.v(9648)
  not u10362 (Rj6ju6, n2762);  // ../RTL/cortexm0ds_logic.v(9648)
  and u10363 (n2763, Al6ju6, Ic5ju6);  // ../RTL/cortexm0ds_logic.v(9649)
  not u10364 (Tk6ju6, n2763);  // ../RTL/cortexm0ds_logic.v(9649)
  and u10365 (n2764, Mk6ju6, E2epw6);  // ../RTL/cortexm0ds_logic.v(9650)
  not u10366 (Al6ju6, n2764);  // ../RTL/cortexm0ds_logic.v(9650)
  xor u10367 (E2epw6, Hl6ju6, Ol6ju6);  // ../RTL/cortexm0ds_logic.v(9651)
  and u10368 (n2765, Vl6ju6, Cm6ju6);  // ../RTL/cortexm0ds_logic.v(9652)
  not u10369 (Hl6ju6, n2765);  // ../RTL/cortexm0ds_logic.v(9652)
  not u1037 (M8yhu6, n8);  // ../RTL/cortexm0ds_logic.v(3186)
  and u10370 (Cm6ju6, Jm6ju6, Qm6ju6);  // ../RTL/cortexm0ds_logic.v(9653)
  and u10371 (n2766, Kc6ju6, S8fpw6[4]);  // ../RTL/cortexm0ds_logic.v(9654)
  not u10372 (Qm6ju6, n2766);  // ../RTL/cortexm0ds_logic.v(9654)
  and u10373 (n2767, S8fpw6[6], Xv4ju6);  // ../RTL/cortexm0ds_logic.v(9655)
  not u10374 (Jm6ju6, n2767);  // ../RTL/cortexm0ds_logic.v(9655)
  and u10375 (Vl6ju6, Xm6ju6, En6ju6);  // ../RTL/cortexm0ds_logic.v(9656)
  and u10376 (n2768, Sw4ju6, Kj6ju6);  // ../RTL/cortexm0ds_logic.v(9657)
  not u10377 (En6ju6, n2768);  // ../RTL/cortexm0ds_logic.v(9657)
  or u10378 (Xm6ju6, Gx4ju6, Dzjiu6);  // ../RTL/cortexm0ds_logic.v(9658)
  not u10379 (Mk6ju6, Qf0iu6);  // ../RTL/cortexm0ds_logic.v(9659)
  and u1038 (F8yhu6, A9yhu6, H9yhu6);  // ../RTL/cortexm0ds_logic.v(3187)
  and u10380 (n2769, Ln6ju6, Sn6ju6);  // ../RTL/cortexm0ds_logic.v(9660)
  not u10381 (Jukiu6, n2769);  // ../RTL/cortexm0ds_logic.v(9660)
  and u10382 (Sn6ju6, Zn6ju6, Go6ju6);  // ../RTL/cortexm0ds_logic.v(9661)
  and u10383 (n2770, By4ju6, Eafpw6[7]);  // ../RTL/cortexm0ds_logic.v(9662)
  not u10384 (Go6ju6, n2770);  // ../RTL/cortexm0ds_logic.v(9662)
  or u10385 (n2771, Affpw6[7], No6ju6);  // ../RTL/cortexm0ds_logic.v(9663)
  not u10386 (Zn6ju6, n2771);  // ../RTL/cortexm0ds_logic.v(9663)
  and u10387 (No6ju6, Iy4ju6, Uo6ju6);  // ../RTL/cortexm0ds_logic.v(9664)
  and u10388 (Ln6ju6, Bp6ju6, Ip6ju6);  // ../RTL/cortexm0ds_logic.v(9665)
  and u10389 (n2772, Ub5ju6, Pp6ju6);  // ../RTL/cortexm0ds_logic.v(9666)
  and u1039 (n9, O9yhu6, V9yhu6);  // ../RTL/cortexm0ds_logic.v(3188)
  not u10390 (Ip6ju6, n2772);  // ../RTL/cortexm0ds_logic.v(9666)
  and u10391 (n2773, Wp6ju6, Ic5ju6);  // ../RTL/cortexm0ds_logic.v(9667)
  not u10392 (Pp6ju6, n2773);  // ../RTL/cortexm0ds_logic.v(9667)
  and u10393 (n2774, Jf0iu6, S2epw6);  // ../RTL/cortexm0ds_logic.v(9668)
  not u10394 (Wp6ju6, n2774);  // ../RTL/cortexm0ds_logic.v(9668)
  or u10395 (Bp6ju6, Dq6ju6, Jf0iu6);  // ../RTL/cortexm0ds_logic.v(9669)
  AL_MUX u10396 (
    .i0(Cukiu6),
    .i1(Kq6ju6),
    .sel(Mm4ju6),
    .o(Jf0iu6));  // ../RTL/cortexm0ds_logic.v(9670)
  and u10397 (Kq6ju6, Rq6ju6, Yq6ju6);  // ../RTL/cortexm0ds_logic.v(9671)
  and u10398 (Yq6ju6, Fr6ju6, Mr6ju6);  // ../RTL/cortexm0ds_logic.v(9672)
  and u10399 (Mr6ju6, Tr6ju6, As6ju6);  // ../RTL/cortexm0ds_logic.v(9673)
  and u104 (Vnfpw6[0], Ppfpw6[6], Ivfhu6);  // ../RTL/cortexm0ds_logic.v(3367)
  not u1040 (H9yhu6, n9);  // ../RTL/cortexm0ds_logic.v(3188)
  and u10400 (n2775, Jo4ju6, vis_r14_o[7]);  // ../RTL/cortexm0ds_logic.v(9674)
  not u10401 (As6ju6, n2775);  // ../RTL/cortexm0ds_logic.v(9674)
  and u10402 (Tr6ju6, Hs6ju6, Os6ju6);  // ../RTL/cortexm0ds_logic.v(9675)
  and u10403 (n2776, Ep4ju6, vis_psp_o[5]);  // ../RTL/cortexm0ds_logic.v(9676)
  not u10404 (Os6ju6, n2776);  // ../RTL/cortexm0ds_logic.v(9676)
  and u10405 (n2777, Lp4ju6, vis_msp_o[5]);  // ../RTL/cortexm0ds_logic.v(9677)
  not u10406 (Hs6ju6, n2777);  // ../RTL/cortexm0ds_logic.v(9677)
  and u10407 (Fr6ju6, Vs6ju6, Ct6ju6);  // ../RTL/cortexm0ds_logic.v(9678)
  and u10408 (n2778, Gq4ju6, vis_r12_o[7]);  // ../RTL/cortexm0ds_logic.v(9679)
  not u10409 (Ct6ju6, n2778);  // ../RTL/cortexm0ds_logic.v(9679)
  and u1041 (n10, Cayhu6, Jayhu6);  // ../RTL/cortexm0ds_logic.v(3189)
  and u10410 (n2779, Nq4ju6, vis_r11_o[7]);  // ../RTL/cortexm0ds_logic.v(9680)
  not u10411 (Vs6ju6, n2779);  // ../RTL/cortexm0ds_logic.v(9680)
  and u10412 (Rq6ju6, Jt6ju6, Qt6ju6);  // ../RTL/cortexm0ds_logic.v(9681)
  and u10413 (Qt6ju6, Xt6ju6, Eu6ju6);  // ../RTL/cortexm0ds_logic.v(9682)
  and u10414 (n2780, Wr4ju6, vis_r10_o[7]);  // ../RTL/cortexm0ds_logic.v(9683)
  not u10415 (Eu6ju6, n2780);  // ../RTL/cortexm0ds_logic.v(9683)
  and u10416 (n2781, Ds4ju6, vis_r9_o[7]);  // ../RTL/cortexm0ds_logic.v(9684)
  not u10417 (Xt6ju6, n2781);  // ../RTL/cortexm0ds_logic.v(9684)
  and u10418 (Jt6ju6, I40iu6, Lu6ju6);  // ../RTL/cortexm0ds_logic.v(9685)
  and u10419 (n2782, Rs4ju6, vis_r8_o[7]);  // ../RTL/cortexm0ds_logic.v(9686)
  not u1042 (V9yhu6, n10);  // ../RTL/cortexm0ds_logic.v(3189)
  not u10420 (Lu6ju6, n2782);  // ../RTL/cortexm0ds_logic.v(9686)
  not u10421 (Cukiu6, Fkfpw6[7]);  // ../RTL/cortexm0ds_logic.v(9687)
  AL_MUX u10422 (
    .i0(Cg5ju6),
    .i1(Wc5ju6),
    .sel(S2epw6),
    .o(Dq6ju6));  // ../RTL/cortexm0ds_logic.v(9688)
  xor u10423 (n2783, Su6ju6, Hu4ju6);  // ../RTL/cortexm0ds_logic.v(9689)
  not u10424 (S2epw6, n2783);  // ../RTL/cortexm0ds_logic.v(9689)
  and u10425 (n2784, Zu6ju6, Gv6ju6);  // ../RTL/cortexm0ds_logic.v(9690)
  not u10426 (Su6ju6, n2784);  // ../RTL/cortexm0ds_logic.v(9690)
  and u10427 (Gv6ju6, Nv6ju6, Uv6ju6);  // ../RTL/cortexm0ds_logic.v(9691)
  and u10428 (n2785, Kc6ju6, S8fpw6[5]);  // ../RTL/cortexm0ds_logic.v(9692)
  not u10429 (Uv6ju6, n2785);  // ../RTL/cortexm0ds_logic.v(9692)
  and u1043 (n11, U5yhu6, Qayhu6);  // ../RTL/cortexm0ds_logic.v(3190)
  and u10430 (n2786, S8fpw6[7], Xv4ju6);  // ../RTL/cortexm0ds_logic.v(9693)
  not u10431 (Nv6ju6, n2786);  // ../RTL/cortexm0ds_logic.v(9693)
  and u10432 (Zu6ju6, Bw6ju6, Iw6ju6);  // ../RTL/cortexm0ds_logic.v(9694)
  and u10433 (n2787, Sw4ju6, Uo6ju6);  // ../RTL/cortexm0ds_logic.v(9695)
  not u10434 (Iw6ju6, n2787);  // ../RTL/cortexm0ds_logic.v(9695)
  or u10435 (Bw6ju6, Gx4ju6, Ad8iu6);  // ../RTL/cortexm0ds_logic.v(9696)
  or u10436 (n2788, J1liu6, Yykiu6);  // ../RTL/cortexm0ds_logic.v(9697)
  not u10437 (Nh6ju6, n2788);  // ../RTL/cortexm0ds_logic.v(9697)
  and u10438 (n2789, Pw6ju6, Ww6ju6);  // ../RTL/cortexm0ds_logic.v(9698)
  not u10439 (Yykiu6, n2789);  // ../RTL/cortexm0ds_logic.v(9698)
  not u1044 (A9yhu6, n11);  // ../RTL/cortexm0ds_logic.v(3190)
  and u10440 (Ww6ju6, Dx6ju6, Kx6ju6);  // ../RTL/cortexm0ds_logic.v(9699)
  and u10441 (n2790, By4ju6, Eafpw6[24]);  // ../RTL/cortexm0ds_logic.v(9700)
  not u10442 (Kx6ju6, n2790);  // ../RTL/cortexm0ds_logic.v(9700)
  or u10443 (n2791, Affpw6[24], Wk4ju6);  // ../RTL/cortexm0ds_logic.v(9701)
  not u10444 (Dx6ju6, n2791);  // ../RTL/cortexm0ds_logic.v(9701)
  and u10445 (Pw6ju6, Rx6ju6, Yx6ju6);  // ../RTL/cortexm0ds_logic.v(9702)
  and u10446 (n2792, Iy4ju6, Fy6ju6);  // ../RTL/cortexm0ds_logic.v(9703)
  not u10447 (Yx6ju6, n2792);  // ../RTL/cortexm0ds_logic.v(9703)
  AL_MUX u10448 (
    .i0(My6ju6),
    .i1(Ty6ju6),
    .sel(Yj0iu6),
    .o(Rx6ju6));  // ../RTL/cortexm0ds_logic.v(9704)
  and u10449 (n2793, Ys4ju6, Qbfpw6[24]);  // ../RTL/cortexm0ds_logic.v(9705)
  and u1045 (n12, Xayhu6, Ebyhu6);  // ../RTL/cortexm0ds_logic.v(3191)
  not u10450 (Ty6ju6, n2793);  // ../RTL/cortexm0ds_logic.v(9705)
  or u10451 (n2794, Az6ju6, Mt4ju6);  // ../RTL/cortexm0ds_logic.v(9706)
  not u10452 (My6ju6, n2794);  // ../RTL/cortexm0ds_logic.v(9706)
  AL_MUX u10453 (
    .i0(Ys4ju6),
    .i1(Tt4ju6),
    .sel(Qbfpw6[24]),
    .o(Az6ju6));  // ../RTL/cortexm0ds_logic.v(9707)
  buf u10454 (vis_r2_o[4], Bxpax6);  // ../RTL/cortexm0ds_logic.v(2551)
  AL_MUX u10455 (
    .i0(T75ju6),
    .i1(A85ju6),
    .sel(Fy6ju6),
    .o(Hz6ju6));  // ../RTL/cortexm0ds_logic.v(9709)
  and u10456 (n2795, Oz6ju6, Vz6ju6);  // ../RTL/cortexm0ds_logic.v(9710)
  not u10457 (J1liu6, n2795);  // ../RTL/cortexm0ds_logic.v(9710)
  and u10458 (Vz6ju6, C07ju6, J07ju6);  // ../RTL/cortexm0ds_logic.v(9711)
  and u10459 (n2796, By4ju6, Eafpw6[26]);  // ../RTL/cortexm0ds_logic.v(9712)
  not u1046 (Qayhu6, n12);  // ../RTL/cortexm0ds_logic.v(3191)
  not u10460 (J07ju6, n2796);  // ../RTL/cortexm0ds_logic.v(9712)
  or u10461 (n2797, Affpw6[26], Q07ju6);  // ../RTL/cortexm0ds_logic.v(9713)
  not u10462 (C07ju6, n2797);  // ../RTL/cortexm0ds_logic.v(9713)
  or u10463 (n2798, X07ju6, E17ju6);  // ../RTL/cortexm0ds_logic.v(9714)
  not u10464 (Q07ju6, n2798);  // ../RTL/cortexm0ds_logic.v(9714)
  AL_MUX u10465 (
    .i0(Cg5ju6),
    .i1(Wc5ju6),
    .sel(Qbfpw6[26]),
    .o(X07ju6));  // ../RTL/cortexm0ds_logic.v(9715)
  and u10466 (Oz6ju6, L17ju6, S17ju6);  // ../RTL/cortexm0ds_logic.v(9716)
  and u10467 (n2799, Iy4ju6, Z17ju6);  // ../RTL/cortexm0ds_logic.v(9717)
  not u10468 (S17ju6, n2799);  // ../RTL/cortexm0ds_logic.v(9717)
  and u10469 (n2800, Ub5ju6, G27ju6);  // ../RTL/cortexm0ds_logic.v(9718)
  or u1047 (n13, Lbyhu6, Sbyhu6);  // ../RTL/cortexm0ds_logic.v(3192)
  not u10470 (L17ju6, n2800);  // ../RTL/cortexm0ds_logic.v(9718)
  and u10471 (n2801, N27ju6, Ic5ju6);  // ../RTL/cortexm0ds_logic.v(9719)
  not u10472 (G27ju6, n2801);  // ../RTL/cortexm0ds_logic.v(9719)
  and u10473 (n2802, E17ju6, Qbfpw6[26]);  // ../RTL/cortexm0ds_logic.v(9720)
  not u10474 (N27ju6, n2802);  // ../RTL/cortexm0ds_logic.v(9720)
  buf u10475 (vis_r2_o[2], Cvpax6);  // ../RTL/cortexm0ds_logic.v(2551)
  AL_MUX u10476 (
    .i0(T75ju6),
    .i1(A85ju6),
    .sel(Z17ju6),
    .o(U27ju6));  // ../RTL/cortexm0ds_logic.v(9722)
  not u10477 (E17ju6, Kj0iu6);  // ../RTL/cortexm0ds_logic.v(9723)
  and u10478 (Zg6ju6, B37ju6, I37ju6);  // ../RTL/cortexm0ds_logic.v(9724)
  or u10479 (n2803, W4liu6, B4liu6);  // ../RTL/cortexm0ds_logic.v(9725)
  not u1048 (Ebyhu6, n13);  // ../RTL/cortexm0ds_logic.v(3192)
  not u10480 (I37ju6, n2803);  // ../RTL/cortexm0ds_logic.v(9725)
  and u10481 (n2804, P37ju6, W37ju6);  // ../RTL/cortexm0ds_logic.v(9726)
  not u10482 (B4liu6, n2804);  // ../RTL/cortexm0ds_logic.v(9726)
  and u10483 (W37ju6, D47ju6, K47ju6);  // ../RTL/cortexm0ds_logic.v(9727)
  and u10484 (n2805, By4ju6, Eafpw6[27]);  // ../RTL/cortexm0ds_logic.v(9728)
  not u10485 (K47ju6, n2805);  // ../RTL/cortexm0ds_logic.v(9728)
  or u10486 (n2806, Affpw6[27], R47ju6);  // ../RTL/cortexm0ds_logic.v(9729)
  not u10487 (D47ju6, n2806);  // ../RTL/cortexm0ds_logic.v(9729)
  or u10488 (n2807, Y47ju6, F57ju6);  // ../RTL/cortexm0ds_logic.v(9730)
  not u10489 (R47ju6, n2807);  // ../RTL/cortexm0ds_logic.v(9730)
  and u1049 (Xayhu6, Zbyhu6, Gcyhu6);  // ../RTL/cortexm0ds_logic.v(3193)
  AL_MUX u10490 (
    .i0(Cg5ju6),
    .i1(Wc5ju6),
    .sel(Qbfpw6[27]),
    .o(Y47ju6));  // ../RTL/cortexm0ds_logic.v(9731)
  and u10491 (P37ju6, M57ju6, T57ju6);  // ../RTL/cortexm0ds_logic.v(9732)
  and u10492 (n2808, Iy4ju6, A67ju6);  // ../RTL/cortexm0ds_logic.v(9733)
  not u10493 (T57ju6, n2808);  // ../RTL/cortexm0ds_logic.v(9733)
  and u10494 (n2809, Ub5ju6, H67ju6);  // ../RTL/cortexm0ds_logic.v(9734)
  not u10495 (M57ju6, n2809);  // ../RTL/cortexm0ds_logic.v(9734)
  and u10496 (n2810, O67ju6, Ic5ju6);  // ../RTL/cortexm0ds_logic.v(9735)
  not u10497 (H67ju6, n2810);  // ../RTL/cortexm0ds_logic.v(9735)
  and u10498 (n2811, F57ju6, Qbfpw6[27]);  // ../RTL/cortexm0ds_logic.v(9736)
  not u10499 (O67ju6, n2811);  // ../RTL/cortexm0ds_logic.v(9736)
  not u105 (Vmdpw6, P13iu6);  // ../RTL/cortexm0ds_logic.v(1884)
  and u1050 (n14, Ighpw6[4], Ncyhu6);  // ../RTL/cortexm0ds_logic.v(3194)
  buf u10500 (vis_r2_o[1], Vmqax6);  // ../RTL/cortexm0ds_logic.v(2551)
  AL_MUX u10501 (
    .i0(T75ju6),
    .i1(A85ju6),
    .sel(A67ju6),
    .o(V67ju6));  // ../RTL/cortexm0ds_logic.v(9738)
  not u10502 (F57ju6, Dj0iu6);  // ../RTL/cortexm0ds_logic.v(9739)
  and u10503 (n2812, C77ju6, J77ju6);  // ../RTL/cortexm0ds_logic.v(9740)
  not u10504 (W4liu6, n2812);  // ../RTL/cortexm0ds_logic.v(9740)
  and u10505 (J77ju6, Q77ju6, X77ju6);  // ../RTL/cortexm0ds_logic.v(9741)
  and u10506 (n2813, I55ju6, vis_apsr_o[1]);  // ../RTL/cortexm0ds_logic.v(9742)
  not u10507 (X77ju6, n2813);  // ../RTL/cortexm0ds_logic.v(9742)
  or u10508 (n2814, Affpw6[29], Wk4ju6);  // ../RTL/cortexm0ds_logic.v(9743)
  not u10509 (Q77ju6, n2814);  // ../RTL/cortexm0ds_logic.v(9743)
  not u1051 (Gcyhu6, n14);  // ../RTL/cortexm0ds_logic.v(3194)
  and u10510 (C77ju6, E87ju6, L87ju6);  // ../RTL/cortexm0ds_logic.v(9744)
  AL_MUX u10511 (
    .i0(S87ju6),
    .i1(Z87ju6),
    .sel(Pi0iu6),
    .o(L87ju6));  // ../RTL/cortexm0ds_logic.v(9745)
  and u10512 (n2815, Ys4ju6, Qbfpw6[29]);  // ../RTL/cortexm0ds_logic.v(9746)
  not u10513 (Z87ju6, n2815);  // ../RTL/cortexm0ds_logic.v(9746)
  or u10514 (n2816, G97ju6, Mt4ju6);  // ../RTL/cortexm0ds_logic.v(9747)
  not u10515 (S87ju6, n2816);  // ../RTL/cortexm0ds_logic.v(9747)
  AL_MUX u10516 (
    .i0(Ys4ju6),
    .i1(Tt4ju6),
    .sel(Qbfpw6[29]),
    .o(G97ju6));  // ../RTL/cortexm0ds_logic.v(9748)
  buf u10517 (Bagpw6[22], D7gbx6);  // ../RTL/cortexm0ds_logic.v(2680)
  AL_MUX u10518 (
    .i0(T75ju6),
    .i1(A85ju6),
    .sel(Wh8iu6),
    .o(N97ju6));  // ../RTL/cortexm0ds_logic.v(9750)
  and u10519 (E87ju6, U97ju6, Ba7ju6);  // ../RTL/cortexm0ds_logic.v(9751)
  and u1052 (n15, Ucyhu6, Bdyhu6);  // ../RTL/cortexm0ds_logic.v(3195)
  and u10520 (n2817, By4ju6, Eafpw6[29]);  // ../RTL/cortexm0ds_logic.v(9752)
  not u10521 (Ba7ju6, n2817);  // ../RTL/cortexm0ds_logic.v(9752)
  and u10522 (n2818, Iy4ju6, Wh8iu6);  // ../RTL/cortexm0ds_logic.v(9753)
  not u10523 (U97ju6, n2818);  // ../RTL/cortexm0ds_logic.v(9753)
  and u10524 (B37ju6, Kgoiu6, Bpliu6);  // ../RTL/cortexm0ds_logic.v(9754)
  and u10525 (Bpliu6, Ia7ju6, Pa7ju6);  // ../RTL/cortexm0ds_logic.v(9755)
  and u10526 (Pa7ju6, Wa7ju6, Db7ju6);  // ../RTL/cortexm0ds_logic.v(9756)
  and u10527 (n2819, Pk4ju6, vis_ipsr_o[1]);  // ../RTL/cortexm0ds_logic.v(9757)
  not u10528 (Db7ju6, n2819);  // ../RTL/cortexm0ds_logic.v(9757)
  and u10529 (Pk4ju6, Kb7ju6, T05ju6);  // ../RTL/cortexm0ds_logic.v(9758)
  not u1053 (Ncyhu6, n15);  // ../RTL/cortexm0ds_logic.v(3195)
  or u10530 (n2820, Je8iu6, S8fpw6[4]);  // ../RTL/cortexm0ds_logic.v(9759)
  not u10531 (Kb7ju6, n2820);  // ../RTL/cortexm0ds_logic.v(9759)
  or u10532 (n2821, Affpw6[1], Rb7ju6);  // ../RTL/cortexm0ds_logic.v(9760)
  not u10533 (Wa7ju6, n2821);  // ../RTL/cortexm0ds_logic.v(9760)
  and u10534 (Rb7ju6, Yb7ju6, Fc7ju6);  // ../RTL/cortexm0ds_logic.v(9761)
  or u10535 (n2822, B5kiu6, Qjoiu6);  // ../RTL/cortexm0ds_logic.v(9762)
  not u10536 (Fc7ju6, n2822);  // ../RTL/cortexm0ds_logic.v(9762)
  and u10537 (Yb7ju6, vis_control_o, T05ju6);  // ../RTL/cortexm0ds_logic.v(9763)
  and u10538 (Ia7ju6, Mc7ju6, Tc7ju6);  // ../RTL/cortexm0ds_logic.v(9764)
  AL_MUX u10539 (
    .i0(Ad7ju6),
    .i1(Hd7ju6),
    .sel(Hl0iu6),
    .o(Tc7ju6));  // ../RTL/cortexm0ds_logic.v(9765)
  or u1054 (Bdyhu6, Ighpw6[1], Ighpw6[2]);  // ../RTL/cortexm0ds_logic.v(3196)
  and u10540 (n2823, Ys4ju6, Qbfpw6[1]);  // ../RTL/cortexm0ds_logic.v(9766)
  not u10541 (Hd7ju6, n2823);  // ../RTL/cortexm0ds_logic.v(9766)
  or u10542 (n2824, Od7ju6, Mt4ju6);  // ../RTL/cortexm0ds_logic.v(9767)
  not u10543 (Ad7ju6, n2824);  // ../RTL/cortexm0ds_logic.v(9767)
  AL_MUX u10544 (
    .i0(Ys4ju6),
    .i1(Tt4ju6),
    .sel(Qbfpw6[1]),
    .o(Od7ju6));  // ../RTL/cortexm0ds_logic.v(9768)
  buf u10545 (Bagpw6[13], R7kpw6);  // ../RTL/cortexm0ds_logic.v(2680)
  buf u10546 (Bagpw6[20], X6jpw6);  // ../RTL/cortexm0ds_logic.v(2680)
  and u10547 (n2825, Ce7ju6, Je7ju6);  // ../RTL/cortexm0ds_logic.v(9770)
  not u10548 (Vd7ju6, n2825);  // ../RTL/cortexm0ds_logic.v(9770)
  or u10549 (Je7ju6, Rb8iu6, Gx4ju6);  // ../RTL/cortexm0ds_logic.v(9771)
  and u1055 (Ucyhu6, Idyhu6, Pdyhu6);  // ../RTL/cortexm0ds_logic.v(3197)
  and u10550 (Ce7ju6, Qe7ju6, Xe7ju6);  // ../RTL/cortexm0ds_logic.v(9772)
  and u10551 (n2826, S8fpw6[1], E35ju6);  // ../RTL/cortexm0ds_logic.v(9773)
  not u10552 (Xe7ju6, n2826);  // ../RTL/cortexm0ds_logic.v(9773)
  or u10553 (E35ju6, Xv4ju6, Ef7ju6);  // ../RTL/cortexm0ds_logic.v(9774)
  and u10554 (Ef7ju6, Lf7ju6, Sf7ju6);  // ../RTL/cortexm0ds_logic.v(9775)
  and u10555 (Lf7ju6, H6ghu6, Cyfpw6[1]);  // ../RTL/cortexm0ds_logic.v(9776)
  or u10556 (Xv4ju6, Zf7ju6, Gg7ju6);  // ../RTL/cortexm0ds_logic.v(9777)
  and u10557 (Gg7ju6, H6ghu6, Ng7ju6);  // ../RTL/cortexm0ds_logic.v(9778)
  and u10558 (n2827, Ug7ju6, Bh7ju6);  // ../RTL/cortexm0ds_logic.v(9779)
  not u10559 (Ng7ju6, n2827);  // ../RTL/cortexm0ds_logic.v(9779)
  or u1056 (Idyhu6, Wdyhu6, Deyhu6);  // ../RTL/cortexm0ds_logic.v(3198)
  and u10560 (n2828, Ih7ju6, K9aiu6);  // ../RTL/cortexm0ds_logic.v(9780)
  not u10561 (Bh7ju6, n2828);  // ../RTL/cortexm0ds_logic.v(9780)
  and u10562 (n2829, Ph7ju6, Wh7ju6);  // ../RTL/cortexm0ds_logic.v(9781)
  not u10563 (Ih7ju6, n2829);  // ../RTL/cortexm0ds_logic.v(9781)
  or u10564 (Ph7ju6, M32ju6, Cyfpw6[6]);  // ../RTL/cortexm0ds_logic.v(9782)
  and u10565 (Ug7ju6, Di7ju6, Ki7ju6);  // ../RTL/cortexm0ds_logic.v(9783)
  and u10566 (n2830, Fd0iu6, Ri7ju6);  // ../RTL/cortexm0ds_logic.v(9784)
  not u10567 (Ki7ju6, n2830);  // ../RTL/cortexm0ds_logic.v(9784)
  or u10568 (Ri7ju6, Mo2ju6, Yi7ju6);  // ../RTL/cortexm0ds_logic.v(9785)
  and u10569 (n2831, C0ehu6, Fj7ju6);  // ../RTL/cortexm0ds_logic.v(9786)
  AL_MUX u1057 (
    .i0(Keyhu6),
    .i1(Reyhu6),
    .sel(Mdhpw6[3]),
    .o(Zbyhu6));  // ../RTL/cortexm0ds_logic.v(3199)
  not u10570 (Di7ju6, n2831);  // ../RTL/cortexm0ds_logic.v(9786)
  and u10571 (n2832, O60ju6, Mj7ju6);  // ../RTL/cortexm0ds_logic.v(9787)
  not u10572 (Fj7ju6, n2832);  // ../RTL/cortexm0ds_logic.v(9787)
  and u10573 (n2833, Jf6ju6, Cyfpw6[0]);  // ../RTL/cortexm0ds_logic.v(9788)
  not u10574 (Mj7ju6, n2833);  // ../RTL/cortexm0ds_logic.v(9788)
  and u10575 (n2834, Sw4ju6, Znliu6);  // ../RTL/cortexm0ds_logic.v(9789)
  not u10576 (Qe7ju6, n2834);  // ../RTL/cortexm0ds_logic.v(9789)
  and u10577 (Mc7ju6, Tj7ju6, Ak7ju6);  // ../RTL/cortexm0ds_logic.v(9790)
  and u10578 (n2835, By4ju6, Eafpw6[1]);  // ../RTL/cortexm0ds_logic.v(9791)
  not u10579 (Ak7ju6, n2835);  // ../RTL/cortexm0ds_logic.v(9791)
  and u1058 (Reyhu6, Yeyhu6, Ffyhu6);  // ../RTL/cortexm0ds_logic.v(3200)
  and u10580 (n2836, Iy4ju6, Znliu6);  // ../RTL/cortexm0ds_logic.v(9792)
  not u10581 (Tj7ju6, n2836);  // ../RTL/cortexm0ds_logic.v(9792)
  and u10582 (Kgoiu6, Hk7ju6, Ok7ju6);  // ../RTL/cortexm0ds_logic.v(9793)
  and u10583 (Ok7ju6, Vk7ju6, Cl7ju6);  // ../RTL/cortexm0ds_logic.v(9794)
  and u10584 (n2837, vis_apsr_o[0], I55ju6);  // ../RTL/cortexm0ds_logic.v(9795)
  not u10585 (Cl7ju6, n2837);  // ../RTL/cortexm0ds_logic.v(9795)
  and u10586 (I55ju6, Jl7ju6, T05ju6);  // ../RTL/cortexm0ds_logic.v(9796)
  and u10587 (T05ju6, Ql7ju6, Xl7ju6);  // ../RTL/cortexm0ds_logic.v(9797)
  or u10588 (n2838, Qxaiu6, C0ehu6);  // ../RTL/cortexm0ds_logic.v(9798)
  not u10589 (Xl7ju6, n2838);  // ../RTL/cortexm0ds_logic.v(9798)
  and u1059 (Yeyhu6, Mfyhu6, Tfyhu6);  // ../RTL/cortexm0ds_logic.v(3201)
  and u10590 (Ql7ju6, H6ghu6, D31ju6);  // ../RTL/cortexm0ds_logic.v(9799)
  or u10591 (n2839, S8fpw6[2], S8fpw6[4]);  // ../RTL/cortexm0ds_logic.v(9800)
  not u10592 (Jl7ju6, n2839);  // ../RTL/cortexm0ds_logic.v(9800)
  or u10593 (n2840, Affpw6[28], Wk4ju6);  // ../RTL/cortexm0ds_logic.v(9801)
  not u10594 (Vk7ju6, n2840);  // ../RTL/cortexm0ds_logic.v(9801)
  and u10595 (Hk7ju6, Em7ju6, Lm7ju6);  // ../RTL/cortexm0ds_logic.v(9802)
  AL_MUX u10596 (
    .i0(Sm7ju6),
    .i1(Zm7ju6),
    .sel(Wi0iu6),
    .o(Lm7ju6));  // ../RTL/cortexm0ds_logic.v(9803)
  and u10597 (n2841, Ys4ju6, Qbfpw6[28]);  // ../RTL/cortexm0ds_logic.v(9804)
  not u10598 (Zm7ju6, n2841);  // ../RTL/cortexm0ds_logic.v(9804)
  or u10599 (n2842, Gn7ju6, Mt4ju6);  // ../RTL/cortexm0ds_logic.v(9805)
  buf u106 (Fanhu6, I0opw6);  // ../RTL/cortexm0ds_logic.v(1885)
  or u1060 (n16, Agyhu6, Hgyhu6);  // ../RTL/cortexm0ds_logic.v(3202)
  not u10600 (Sm7ju6, n2842);  // ../RTL/cortexm0ds_logic.v(9805)
  AL_MUX u10601 (
    .i0(Ys4ju6),
    .i1(Tt4ju6),
    .sel(Qbfpw6[28]),
    .o(Gn7ju6));  // ../RTL/cortexm0ds_logic.v(9806)
  buf u10602 (Bagpw6[23], J7xax6);  // ../RTL/cortexm0ds_logic.v(2680)
  AL_MUX u10603 (
    .i0(A85ju6),
    .i1(T75ju6),
    .sel(Mbniu6),
    .o(Nn7ju6));  // ../RTL/cortexm0ds_logic.v(9808)
  and u10604 (Em7ju6, Un7ju6, Bo7ju6);  // ../RTL/cortexm0ds_logic.v(9809)
  and u10605 (n2843, By4ju6, Eafpw6[28]);  // ../RTL/cortexm0ds_logic.v(9810)
  not u10606 (Bo7ju6, n2843);  // ../RTL/cortexm0ds_logic.v(9810)
  or u10607 (Un7ju6, Io7ju6, Mbniu6);  // ../RTL/cortexm0ds_logic.v(9811)
  and u10608 (Jh4ju6, Wo7ju6, Dp7ju6);  // ../RTL/cortexm0ds_logic.v(9813)
  and u10609 (Dp7ju6, Kp7ju6, Rp7ju6);  // ../RTL/cortexm0ds_logic.v(9814)
  not u1061 (Keyhu6, n16);  // ../RTL/cortexm0ds_logic.v(3202)
  and u10610 (Rp7ju6, Yp7ju6, Fq7ju6);  // ../RTL/cortexm0ds_logic.v(9815)
  or u10611 (n2844, R3niu6, L7niu6);  // ../RTL/cortexm0ds_logic.v(9816)
  not u10612 (Fq7ju6, n2844);  // ../RTL/cortexm0ds_logic.v(9816)
  and u10613 (n2845, Mq7ju6, Tq7ju6);  // ../RTL/cortexm0ds_logic.v(9817)
  not u10614 (L7niu6, n2845);  // ../RTL/cortexm0ds_logic.v(9817)
  and u10615 (Tq7ju6, Ar7ju6, Hr7ju6);  // ../RTL/cortexm0ds_logic.v(9818)
  and u10616 (n2846, Or7ju6, Ub5ju6);  // ../RTL/cortexm0ds_logic.v(9819)
  not u10617 (Hr7ju6, n2846);  // ../RTL/cortexm0ds_logic.v(9819)
  and u10618 (n2847, Ic5ju6, Vr7ju6);  // ../RTL/cortexm0ds_logic.v(9820)
  not u10619 (Or7ju6, n2847);  // ../RTL/cortexm0ds_logic.v(9820)
  buf u1062 (vis_r5_o[4], O5ppw6);  // ../RTL/cortexm0ds_logic.v(1909)
  and u10620 (n2848, Ve0iu6, W4epw6);  // ../RTL/cortexm0ds_logic.v(9821)
  not u10621 (Vr7ju6, n2848);  // ../RTL/cortexm0ds_logic.v(9821)
  or u10622 (n2849, Affpw6[8], Cs7ju6);  // ../RTL/cortexm0ds_logic.v(9822)
  not u10623 (Ar7ju6, n2849);  // ../RTL/cortexm0ds_logic.v(9822)
  or u10624 (n2850, Js7ju6, Ve0iu6);  // ../RTL/cortexm0ds_logic.v(9823)
  not u10625 (Cs7ju6, n2850);  // ../RTL/cortexm0ds_logic.v(9823)
  AL_MUX u10626 (
    .i0(Q6niu6),
    .i1(Qs7ju6),
    .sel(Mm4ju6),
    .o(Ve0iu6));  // ../RTL/cortexm0ds_logic.v(9824)
  and u10627 (Qs7ju6, Xs7ju6, Et7ju6);  // ../RTL/cortexm0ds_logic.v(9825)
  and u10628 (Et7ju6, Lt7ju6, St7ju6);  // ../RTL/cortexm0ds_logic.v(9826)
  and u10629 (St7ju6, Zt7ju6, Gu7ju6);  // ../RTL/cortexm0ds_logic.v(9827)
  buf u1063 (vis_r5_o[10], Hsxpw6);  // ../RTL/cortexm0ds_logic.v(1909)
  and u10630 (n2851, Jo4ju6, vis_r14_o[8]);  // ../RTL/cortexm0ds_logic.v(9828)
  not u10631 (Gu7ju6, n2851);  // ../RTL/cortexm0ds_logic.v(9828)
  and u10632 (Zt7ju6, Nu7ju6, Uu7ju6);  // ../RTL/cortexm0ds_logic.v(9829)
  and u10633 (n2852, Ep4ju6, vis_psp_o[6]);  // ../RTL/cortexm0ds_logic.v(9830)
  not u10634 (Uu7ju6, n2852);  // ../RTL/cortexm0ds_logic.v(9830)
  and u10635 (n2853, Lp4ju6, vis_msp_o[6]);  // ../RTL/cortexm0ds_logic.v(9831)
  not u10636 (Nu7ju6, n2853);  // ../RTL/cortexm0ds_logic.v(9831)
  and u10637 (Lt7ju6, Bv7ju6, Iv7ju6);  // ../RTL/cortexm0ds_logic.v(9832)
  and u10638 (n2854, Gq4ju6, vis_r12_o[8]);  // ../RTL/cortexm0ds_logic.v(9833)
  not u10639 (Iv7ju6, n2854);  // ../RTL/cortexm0ds_logic.v(9833)
  and u1064 (n17, O9yhu6, Mdhpw6[3]);  // ../RTL/cortexm0ds_logic.v(3204)
  and u10640 (n2855, Nq4ju6, vis_r11_o[8]);  // ../RTL/cortexm0ds_logic.v(9834)
  not u10641 (Bv7ju6, n2855);  // ../RTL/cortexm0ds_logic.v(9834)
  and u10642 (Xs7ju6, Pv7ju6, Wv7ju6);  // ../RTL/cortexm0ds_logic.v(9835)
  and u10643 (Wv7ju6, Dw7ju6, Kw7ju6);  // ../RTL/cortexm0ds_logic.v(9836)
  and u10644 (n2856, Wr4ju6, vis_r10_o[8]);  // ../RTL/cortexm0ds_logic.v(9837)
  not u10645 (Kw7ju6, n2856);  // ../RTL/cortexm0ds_logic.v(9837)
  and u10646 (n2857, Ds4ju6, vis_r9_o[8]);  // ../RTL/cortexm0ds_logic.v(9838)
  not u10647 (Dw7ju6, n2857);  // ../RTL/cortexm0ds_logic.v(9838)
  and u10648 (Pv7ju6, B40iu6, Rw7ju6);  // ../RTL/cortexm0ds_logic.v(9839)
  and u10649 (n2858, Rs4ju6, vis_r8_o[8]);  // ../RTL/cortexm0ds_logic.v(9840)
  not u1065 (Vgyhu6, n17);  // ../RTL/cortexm0ds_logic.v(3204)
  not u10650 (Rw7ju6, n2858);  // ../RTL/cortexm0ds_logic.v(9840)
  not u10651 (Q6niu6, Fkfpw6[8]);  // ../RTL/cortexm0ds_logic.v(9841)
  AL_MUX u10652 (
    .i0(Cg5ju6),
    .i1(Wc5ju6),
    .sel(W4epw6),
    .o(Js7ju6));  // ../RTL/cortexm0ds_logic.v(9842)
  xor u10653 (n2859, Yw7ju6, Hu4ju6);  // ../RTL/cortexm0ds_logic.v(9843)
  not u10654 (W4epw6, n2859);  // ../RTL/cortexm0ds_logic.v(9843)
  and u10655 (n2860, Fx7ju6, Mx7ju6);  // ../RTL/cortexm0ds_logic.v(9844)
  not u10656 (Yw7ju6, n2860);  // ../RTL/cortexm0ds_logic.v(9844)
  and u10657 (Mx7ju6, Tx7ju6, Ay7ju6);  // ../RTL/cortexm0ds_logic.v(9845)
  and u10658 (n2861, Kc6ju6, S8fpw6[6]);  // ../RTL/cortexm0ds_logic.v(9846)
  not u10659 (Ay7ju6, n2861);  // ../RTL/cortexm0ds_logic.v(9846)
  and u1066 (Ogyhu6, Chyhu6, Jhyhu6);  // ../RTL/cortexm0ds_logic.v(3205)
  and u10660 (n2862, Zf7ju6, S8fpw6[8]);  // ../RTL/cortexm0ds_logic.v(9847)
  not u10661 (Tx7ju6, n2862);  // ../RTL/cortexm0ds_logic.v(9847)
  and u10662 (Fx7ju6, Hy7ju6, Oy7ju6);  // ../RTL/cortexm0ds_logic.v(9848)
  or u10663 (Oy7ju6, Vy7ju6, Cz7ju6);  // ../RTL/cortexm0ds_logic.v(9849)
  or u10664 (Hy7ju6, O95iu6, Gx4ju6);  // ../RTL/cortexm0ds_logic.v(9850)
  and u10665 (Mq7ju6, Jz7ju6, Qz7ju6);  // ../RTL/cortexm0ds_logic.v(9851)
  and u10666 (n2863, By4ju6, Eafpw6[8]);  // ../RTL/cortexm0ds_logic.v(9852)
  not u10667 (Qz7ju6, n2863);  // ../RTL/cortexm0ds_logic.v(9852)
  or u10668 (Jz7ju6, Io7ju6, Cz7ju6);  // ../RTL/cortexm0ds_logic.v(9853)
  and u10669 (n2864, Xz7ju6, E08ju6);  // ../RTL/cortexm0ds_logic.v(9854)
  and u1067 (n18, Qhyhu6, U5yhu6);  // ../RTL/cortexm0ds_logic.v(3206)
  not u10670 (R3niu6, n2864);  // ../RTL/cortexm0ds_logic.v(9854)
  and u10671 (E08ju6, L08ju6, S08ju6);  // ../RTL/cortexm0ds_logic.v(9855)
  and u10672 (n2865, By4ju6, Eafpw6[9]);  // ../RTL/cortexm0ds_logic.v(9856)
  not u10673 (S08ju6, n2865);  // ../RTL/cortexm0ds_logic.v(9856)
  or u10674 (n2866, Affpw6[9], Z08ju6);  // ../RTL/cortexm0ds_logic.v(9857)
  not u10675 (L08ju6, n2866);  // ../RTL/cortexm0ds_logic.v(9857)
  or u10676 (n2867, G18ju6, N18ju6);  // ../RTL/cortexm0ds_logic.v(9858)
  not u10677 (Z08ju6, n2867);  // ../RTL/cortexm0ds_logic.v(9858)
  AL_MUX u10678 (
    .i0(Cg5ju6),
    .i1(Wc5ju6),
    .sel(Q5phu6),
    .o(G18ju6));  // ../RTL/cortexm0ds_logic.v(9859)
  and u10679 (Xz7ju6, U18ju6, B28ju6);  // ../RTL/cortexm0ds_logic.v(9860)
  not u1068 (Jhyhu6, n18);  // ../RTL/cortexm0ds_logic.v(3206)
  or u10680 (B28ju6, Io7ju6, I28ju6);  // ../RTL/cortexm0ds_logic.v(9861)
  and u10681 (n2868, Ub5ju6, P28ju6);  // ../RTL/cortexm0ds_logic.v(9862)
  not u10682 (U18ju6, n2868);  // ../RTL/cortexm0ds_logic.v(9862)
  and u10683 (n2869, W28ju6, Ic5ju6);  // ../RTL/cortexm0ds_logic.v(9863)
  not u10684 (P28ju6, n2869);  // ../RTL/cortexm0ds_logic.v(9863)
  and u10685 (n2870, N18ju6, Q5phu6);  // ../RTL/cortexm0ds_logic.v(9864)
  not u10686 (W28ju6, n2870);  // ../RTL/cortexm0ds_logic.v(9864)
  xor u10687 (Q5phu6, D38ju6, Ol6ju6);  // ../RTL/cortexm0ds_logic.v(9865)
  and u10688 (n2871, K38ju6, R38ju6);  // ../RTL/cortexm0ds_logic.v(9866)
  not u10689 (D38ju6, n2871);  // ../RTL/cortexm0ds_logic.v(9866)
  and u1069 (Qhyhu6, Xhyhu6, Eiyhu6);  // ../RTL/cortexm0ds_logic.v(3207)
  and u10690 (R38ju6, Y38ju6, F48ju6);  // ../RTL/cortexm0ds_logic.v(9867)
  and u10691 (n2872, Kc6ju6, S8fpw6[7]);  // ../RTL/cortexm0ds_logic.v(9868)
  not u10692 (F48ju6, n2872);  // ../RTL/cortexm0ds_logic.v(9868)
  and u10693 (Kc6ju6, H6ghu6, M48ju6);  // ../RTL/cortexm0ds_logic.v(9869)
  and u10694 (n2873, T48ju6, A58ju6);  // ../RTL/cortexm0ds_logic.v(9870)
  not u10695 (M48ju6, n2873);  // ../RTL/cortexm0ds_logic.v(9870)
  AL_MUX u10696 (
    .i0(H58ju6),
    .i1(O58ju6),
    .sel(Cyfpw6[3]),
    .o(A58ju6));  // ../RTL/cortexm0ds_logic.v(9871)
  or u10697 (O58ju6, V58ju6, Jc2ju6);  // ../RTL/cortexm0ds_logic.v(9872)
  or u10698 (H58ju6, Szniu6, Knaiu6);  // ../RTL/cortexm0ds_logic.v(9873)
  and u10699 (T48ju6, C68ju6, J68ju6);  // ../RTL/cortexm0ds_logic.v(9874)
  buf u107 (vis_r14_o[15], Zh8bx6);  // ../RTL/cortexm0ds_logic.v(2497)
  and u1070 (n19, Liyhu6, Siyhu6);  // ../RTL/cortexm0ds_logic.v(3208)
  and u10700 (n2874, Y2aiu6, Vo3ju6);  // ../RTL/cortexm0ds_logic.v(9875)
  not u10701 (J68ju6, n2874);  // ../RTL/cortexm0ds_logic.v(9875)
  and u10702 (Y2aiu6, Q68ju6, Fd0iu6);  // ../RTL/cortexm0ds_logic.v(9876)
  or u10703 (n2875, As0iu6, C0ehu6);  // ../RTL/cortexm0ds_logic.v(9877)
  not u10704 (Q68ju6, n2875);  // ../RTL/cortexm0ds_logic.v(9877)
  and u10705 (n2876, D6kiu6, X68ju6);  // ../RTL/cortexm0ds_logic.v(9878)
  not u10706 (C68ju6, n2876);  // ../RTL/cortexm0ds_logic.v(9878)
  and u10707 (n2877, E78ju6, Jc2ju6);  // ../RTL/cortexm0ds_logic.v(9879)
  not u10708 (X68ju6, n2877);  // ../RTL/cortexm0ds_logic.v(9879)
  or u10709 (n2878, L78ju6, Cyfpw6[3]);  // ../RTL/cortexm0ds_logic.v(9880)
  not u1071 (Xhyhu6, n19);  // ../RTL/cortexm0ds_logic.v(3208)
  not u10710 (E78ju6, n2878);  // ../RTL/cortexm0ds_logic.v(9880)
  and u10711 (n2879, Zf7ju6, S8fpw6[9]);  // ../RTL/cortexm0ds_logic.v(9881)
  not u10712 (Y38ju6, n2879);  // ../RTL/cortexm0ds_logic.v(9881)
  and u10713 (K38ju6, S78ju6, Z78ju6);  // ../RTL/cortexm0ds_logic.v(9882)
  or u10714 (Z78ju6, Vy7ju6, I28ju6);  // ../RTL/cortexm0ds_logic.v(9883)
  or u10715 (S78ju6, Ndiiu6, Gx4ju6);  // ../RTL/cortexm0ds_logic.v(9884)
  not u10716 (N18ju6, He0iu6);  // ../RTL/cortexm0ds_logic.v(9885)
  or u10717 (n2880, Vsliu6, Vymiu6);  // ../RTL/cortexm0ds_logic.v(9886)
  not u10718 (Yp7ju6, n2880);  // ../RTL/cortexm0ds_logic.v(9886)
  and u10719 (n2881, G88ju6, N88ju6);  // ../RTL/cortexm0ds_logic.v(9887)
  and u1072 (n20, Ziyhu6, Mdhpw6[0]);  // ../RTL/cortexm0ds_logic.v(3209)
  not u10720 (Vymiu6, n2881);  // ../RTL/cortexm0ds_logic.v(9887)
  and u10721 (N88ju6, U88ju6, B98ju6);  // ../RTL/cortexm0ds_logic.v(9888)
  and u10722 (n2882, By4ju6, Eafpw6[10]);  // ../RTL/cortexm0ds_logic.v(9889)
  not u10723 (B98ju6, n2882);  // ../RTL/cortexm0ds_logic.v(9889)
  or u10724 (n2883, Affpw6[10], I98ju6);  // ../RTL/cortexm0ds_logic.v(9890)
  not u10725 (U88ju6, n2883);  // ../RTL/cortexm0ds_logic.v(9890)
  or u10726 (n2884, P98ju6, Zn0iu6);  // ../RTL/cortexm0ds_logic.v(9891)
  not u10727 (I98ju6, n2884);  // ../RTL/cortexm0ds_logic.v(9891)
  AL_MUX u10728 (
    .i0(Cg5ju6),
    .i1(Wc5ju6),
    .sel(Qbfpw6[10]),
    .o(P98ju6));  // ../RTL/cortexm0ds_logic.v(9892)
  and u10729 (G88ju6, W98ju6, Da8ju6);  // ../RTL/cortexm0ds_logic.v(9893)
  not u1073 (Siyhu6, n20);  // ../RTL/cortexm0ds_logic.v(3209)
  or u10730 (Da8ju6, Io7ju6, Ka8ju6);  // ../RTL/cortexm0ds_logic.v(9894)
  not u10731 (Io7ju6, Iy4ju6);  // ../RTL/cortexm0ds_logic.v(9895)
  and u10732 (n2885, Ub5ju6, Ra8ju6);  // ../RTL/cortexm0ds_logic.v(9896)
  not u10733 (W98ju6, n2885);  // ../RTL/cortexm0ds_logic.v(9896)
  and u10734 (n2886, Ya8ju6, Ic5ju6);  // ../RTL/cortexm0ds_logic.v(9897)
  not u10735 (Ra8ju6, n2886);  // ../RTL/cortexm0ds_logic.v(9897)
  and u10736 (n2887, Zn0iu6, Qbfpw6[10]);  // ../RTL/cortexm0ds_logic.v(9898)
  not u10737 (Ya8ju6, n2887);  // ../RTL/cortexm0ds_logic.v(9898)
  buf u10738 (Bagpw6[8], Rq0qw6);  // ../RTL/cortexm0ds_logic.v(2680)
  buf u10739 (Bagpw6[15], L9xax6);  // ../RTL/cortexm0ds_logic.v(2680)
  and u1074 (n21, Ighpw6[2], Gjyhu6);  // ../RTL/cortexm0ds_logic.v(3210)
  and u10740 (n2888, Mb8ju6, Tb8ju6);  // ../RTL/cortexm0ds_logic.v(9900)
  not u10741 (Fb8ju6, n2888);  // ../RTL/cortexm0ds_logic.v(9900)
  or u10742 (Tb8ju6, Tniiu6, Gx4ju6);  // ../RTL/cortexm0ds_logic.v(9901)
  and u10743 (Mb8ju6, Ac8ju6, Hc8ju6);  // ../RTL/cortexm0ds_logic.v(9902)
  and u10744 (n2889, Zf7ju6, S8fpw6[10]);  // ../RTL/cortexm0ds_logic.v(9903)
  not u10745 (Hc8ju6, n2889);  // ../RTL/cortexm0ds_logic.v(9903)
  or u10746 (Ac8ju6, Vy7ju6, Ka8ju6);  // ../RTL/cortexm0ds_logic.v(9904)
  AL_MUX u10747 (
    .i0(Oc8ju6),
    .i1(Aymiu6),
    .sel(Cn5ju6),
    .o(Zn0iu6));  // ../RTL/cortexm0ds_logic.v(9905)
  not u10748 (Aymiu6, Fkfpw6[10]);  // ../RTL/cortexm0ds_logic.v(9906)
  and u10749 (Oc8ju6, Vc8ju6, Cd8ju6);  // ../RTL/cortexm0ds_logic.v(9907)
  not u1075 (Liyhu6, n21);  // ../RTL/cortexm0ds_logic.v(3210)
  and u10750 (Cd8ju6, Jd8ju6, Qd8ju6);  // ../RTL/cortexm0ds_logic.v(9908)
  and u10751 (Qd8ju6, Xd8ju6, Ee8ju6);  // ../RTL/cortexm0ds_logic.v(9909)
  and u10752 (n2890, Jo4ju6, vis_r14_o[10]);  // ../RTL/cortexm0ds_logic.v(9910)
  not u10753 (Ee8ju6, n2890);  // ../RTL/cortexm0ds_logic.v(9910)
  and u10754 (Xd8ju6, Le8ju6, Se8ju6);  // ../RTL/cortexm0ds_logic.v(9911)
  and u10755 (n2891, Ep4ju6, vis_psp_o[8]);  // ../RTL/cortexm0ds_logic.v(9912)
  not u10756 (Se8ju6, n2891);  // ../RTL/cortexm0ds_logic.v(9912)
  and u10757 (n2892, Lp4ju6, vis_msp_o[8]);  // ../RTL/cortexm0ds_logic.v(9913)
  not u10758 (Le8ju6, n2892);  // ../RTL/cortexm0ds_logic.v(9913)
  and u10759 (Jd8ju6, Ze8ju6, Gf8ju6);  // ../RTL/cortexm0ds_logic.v(9914)
  and u1076 (n22, T8yhu6, Njyhu6);  // ../RTL/cortexm0ds_logic.v(3211)
  and u10760 (n2893, Gq4ju6, vis_r12_o[10]);  // ../RTL/cortexm0ds_logic.v(9915)
  not u10761 (Gf8ju6, n2893);  // ../RTL/cortexm0ds_logic.v(9915)
  and u10762 (n2894, Nq4ju6, vis_r11_o[10]);  // ../RTL/cortexm0ds_logic.v(9916)
  not u10763 (Ze8ju6, n2894);  // ../RTL/cortexm0ds_logic.v(9916)
  and u10764 (Vc8ju6, Nf8ju6, Uf8ju6);  // ../RTL/cortexm0ds_logic.v(9917)
  and u10765 (Uf8ju6, Bg8ju6, Ig8ju6);  // ../RTL/cortexm0ds_logic.v(9918)
  and u10766 (n2895, Wr4ju6, vis_r10_o[10]);  // ../RTL/cortexm0ds_logic.v(9919)
  not u10767 (Ig8ju6, n2895);  // ../RTL/cortexm0ds_logic.v(9919)
  and u10768 (n2896, Ds4ju6, vis_r9_o[10]);  // ../RTL/cortexm0ds_logic.v(9920)
  not u10769 (Bg8ju6, n2896);  // ../RTL/cortexm0ds_logic.v(9920)
  not u1077 (Chyhu6, n22);  // ../RTL/cortexm0ds_logic.v(3211)
  and u10770 (Nf8ju6, Wb0iu6, Pg8ju6);  // ../RTL/cortexm0ds_logic.v(9921)
  and u10771 (n2897, Rs4ju6, vis_r8_o[10]);  // ../RTL/cortexm0ds_logic.v(9922)
  not u10772 (Pg8ju6, n2897);  // ../RTL/cortexm0ds_logic.v(9922)
  and u10773 (n2898, Wg8ju6, Dh8ju6);  // ../RTL/cortexm0ds_logic.v(9923)
  not u10774 (Vsliu6, n2898);  // ../RTL/cortexm0ds_logic.v(9923)
  and u10775 (Dh8ju6, Kh8ju6, Rh8ju6);  // ../RTL/cortexm0ds_logic.v(9924)
  and u10776 (n2899, By4ju6, Eafpw6[25]);  // ../RTL/cortexm0ds_logic.v(9925)
  not u10777 (Rh8ju6, n2899);  // ../RTL/cortexm0ds_logic.v(9925)
  or u10778 (n2900, Affpw6[25], Yh8ju6);  // ../RTL/cortexm0ds_logic.v(9926)
  not u10779 (Kh8ju6, n2900);  // ../RTL/cortexm0ds_logic.v(9926)
  xor u1078 (n23, Ujyhu6, Bkyhu6);  // ../RTL/cortexm0ds_logic.v(3212)
  or u10780 (n2901, Fi8ju6, Mi8ju6);  // ../RTL/cortexm0ds_logic.v(9927)
  not u10781 (Yh8ju6, n2901);  // ../RTL/cortexm0ds_logic.v(9927)
  AL_MUX u10782 (
    .i0(Cg5ju6),
    .i1(Wc5ju6),
    .sel(Qbfpw6[25]),
    .o(Fi8ju6));  // ../RTL/cortexm0ds_logic.v(9928)
  and u10783 (Wg8ju6, Ti8ju6, Aj8ju6);  // ../RTL/cortexm0ds_logic.v(9929)
  and u10784 (n2902, Iy4ju6, Goliu6);  // ../RTL/cortexm0ds_logic.v(9930)
  not u10785 (Aj8ju6, n2902);  // ../RTL/cortexm0ds_logic.v(9930)
  and u10786 (n2903, Ub5ju6, Hj8ju6);  // ../RTL/cortexm0ds_logic.v(9931)
  not u10787 (Ti8ju6, n2903);  // ../RTL/cortexm0ds_logic.v(9931)
  and u10788 (n2904, Oj8ju6, Ic5ju6);  // ../RTL/cortexm0ds_logic.v(9932)
  not u10789 (Hj8ju6, n2904);  // ../RTL/cortexm0ds_logic.v(9932)
  not u1079 (Njyhu6, n23);  // ../RTL/cortexm0ds_logic.v(3212)
  and u10790 (n2905, Mi8ju6, Qbfpw6[25]);  // ../RTL/cortexm0ds_logic.v(9933)
  not u10791 (Oj8ju6, n2905);  // ../RTL/cortexm0ds_logic.v(9933)
  buf u10792 (vis_r2_o[3], Z6qax6);  // ../RTL/cortexm0ds_logic.v(2551)
  and u10793 (n2906, Ck8ju6, Jk8ju6);  // ../RTL/cortexm0ds_logic.v(9935)
  not u10794 (M75ju6, n2906);  // ../RTL/cortexm0ds_logic.v(9935)
  and u10795 (n2907, T75ju6, Vy7ju6);  // ../RTL/cortexm0ds_logic.v(9936)
  not u10796 (Jk8ju6, n2907);  // ../RTL/cortexm0ds_logic.v(9936)
  and u10797 (n2908, Hu4ju6, Qk8ju6);  // ../RTL/cortexm0ds_logic.v(9937)
  not u10798 (Ck8ju6, n2908);  // ../RTL/cortexm0ds_logic.v(9937)
  and u10799 (El8ju6, Xk8ju6, Ij5ju6);  // ../RTL/cortexm0ds_logic.v(9938)
  buf u108 (vis_r8_o[24], Yxspw6);  // ../RTL/cortexm0ds_logic.v(2579)
  and u1080 (Bkyhu6, Ikyhu6, Pkyhu6);  // ../RTL/cortexm0ds_logic.v(3213)
  not u10800 (Qk8ju6, El8ju6);  // ../RTL/cortexm0ds_logic.v(9938)
  AL_MUX u10801 (
    .i0(T75ju6),
    .i1(A85ju6),
    .sel(Goliu6),
    .o(Vj8ju6));  // ../RTL/cortexm0ds_logic.v(9939)
  or u10802 (n2909, Vy7ju6, Ol6ju6);  // ../RTL/cortexm0ds_logic.v(9940)
  not u10803 (A85ju6, n2909);  // ../RTL/cortexm0ds_logic.v(9940)
  and u10804 (T75ju6, El8ju6, Ol6ju6);  // ../RTL/cortexm0ds_logic.v(9941)
  buf u10805 (Exehu6, Ozkbx6[19]);  // ../RTL/cortexm0ds_logic.v(3176)
  not u10806 (Mi8ju6, Rj0iu6);  // ../RTL/cortexm0ds_logic.v(9944)
  and u10807 (Kp7ju6, Ll8ju6, Sl8ju6);  // ../RTL/cortexm0ds_logic.v(9945)
  or u10808 (n2910, Pomiu6, Bvmiu6);  // ../RTL/cortexm0ds_logic.v(9946)
  not u10809 (Sl8ju6, n2910);  // ../RTL/cortexm0ds_logic.v(9946)
  or u1081 (n24, Eiyhu6, Wdyhu6);  // ../RTL/cortexm0ds_logic.v(3214)
  and u10810 (n2911, Zl8ju6, Gm8ju6);  // ../RTL/cortexm0ds_logic.v(9947)
  not u10811 (Bvmiu6, n2911);  // ../RTL/cortexm0ds_logic.v(9947)
  and u10812 (Gm8ju6, Nm8ju6, Um8ju6);  // ../RTL/cortexm0ds_logic.v(9948)
  and u10813 (n2912, By4ju6, Eafpw6[11]);  // ../RTL/cortexm0ds_logic.v(9949)
  not u10814 (Um8ju6, n2912);  // ../RTL/cortexm0ds_logic.v(9949)
  or u10815 (n2913, Affpw6[11], Bn8ju6);  // ../RTL/cortexm0ds_logic.v(9950)
  not u10816 (Nm8ju6, n2913);  // ../RTL/cortexm0ds_logic.v(9950)
  and u10817 (Bn8ju6, Iy4ju6, In8ju6);  // ../RTL/cortexm0ds_logic.v(9951)
  and u10818 (Zl8ju6, Pn8ju6, Wn8ju6);  // ../RTL/cortexm0ds_logic.v(9952)
  and u10819 (n2914, Ub5ju6, Do8ju6);  // ../RTL/cortexm0ds_logic.v(9953)
  not u1082 (Ikyhu6, n24);  // ../RTL/cortexm0ds_logic.v(3214)
  not u10820 (Wn8ju6, n2914);  // ../RTL/cortexm0ds_logic.v(9953)
  and u10821 (n2915, Ko8ju6, Ic5ju6);  // ../RTL/cortexm0ds_logic.v(9954)
  not u10822 (Do8ju6, n2915);  // ../RTL/cortexm0ds_logic.v(9954)
  and u10823 (n2916, Sn0iu6, C1epw6);  // ../RTL/cortexm0ds_logic.v(9955)
  not u10824 (Ko8ju6, n2916);  // ../RTL/cortexm0ds_logic.v(9955)
  or u10825 (Pn8ju6, Ro8ju6, Sn0iu6);  // ../RTL/cortexm0ds_logic.v(9956)
  AL_MUX u10826 (
    .i0(Yo8ju6),
    .i1(Ormiu6),
    .sel(Cn5ju6),
    .o(Sn0iu6));  // ../RTL/cortexm0ds_logic.v(9957)
  not u10827 (Ormiu6, Fkfpw6[11]);  // ../RTL/cortexm0ds_logic.v(9958)
  and u10828 (Yo8ju6, Fp8ju6, Mp8ju6);  // ../RTL/cortexm0ds_logic.v(9959)
  and u10829 (Mp8ju6, Tp8ju6, Aq8ju6);  // ../RTL/cortexm0ds_logic.v(9960)
  buf u1083 (vis_r5_o[5], Mdppw6);  // ../RTL/cortexm0ds_logic.v(1909)
  and u10830 (Aq8ju6, Hq8ju6, Oq8ju6);  // ../RTL/cortexm0ds_logic.v(9961)
  and u10831 (n2917, Jo4ju6, vis_r14_o[11]);  // ../RTL/cortexm0ds_logic.v(9962)
  not u10832 (Oq8ju6, n2917);  // ../RTL/cortexm0ds_logic.v(9962)
  and u10833 (Hq8ju6, Vq8ju6, Cr8ju6);  // ../RTL/cortexm0ds_logic.v(9963)
  and u10834 (n2918, Ep4ju6, vis_psp_o[9]);  // ../RTL/cortexm0ds_logic.v(9964)
  not u10835 (Cr8ju6, n2918);  // ../RTL/cortexm0ds_logic.v(9964)
  and u10836 (n2919, Lp4ju6, vis_msp_o[9]);  // ../RTL/cortexm0ds_logic.v(9965)
  not u10837 (Vq8ju6, n2919);  // ../RTL/cortexm0ds_logic.v(9965)
  and u10838 (Tp8ju6, Jr8ju6, Qr8ju6);  // ../RTL/cortexm0ds_logic.v(9966)
  and u10839 (n2920, Gq4ju6, vis_r12_o[11]);  // ../RTL/cortexm0ds_logic.v(9967)
  buf u1084 (vis_r5_o[11], Ck7bx6);  // ../RTL/cortexm0ds_logic.v(1909)
  not u10840 (Qr8ju6, n2920);  // ../RTL/cortexm0ds_logic.v(9967)
  and u10841 (n2921, Nq4ju6, vis_r11_o[11]);  // ../RTL/cortexm0ds_logic.v(9968)
  not u10842 (Jr8ju6, n2921);  // ../RTL/cortexm0ds_logic.v(9968)
  and u10843 (Fp8ju6, Xr8ju6, Es8ju6);  // ../RTL/cortexm0ds_logic.v(9969)
  and u10844 (Es8ju6, Ls8ju6, Ss8ju6);  // ../RTL/cortexm0ds_logic.v(9970)
  and u10845 (n2922, Wr4ju6, vis_r10_o[11]);  // ../RTL/cortexm0ds_logic.v(9971)
  not u10846 (Ss8ju6, n2922);  // ../RTL/cortexm0ds_logic.v(9971)
  and u10847 (n2923, Ds4ju6, vis_r9_o[11]);  // ../RTL/cortexm0ds_logic.v(9972)
  not u10848 (Ls8ju6, n2923);  // ../RTL/cortexm0ds_logic.v(9972)
  and u10849 (Xr8ju6, Pb0iu6, Zs8ju6);  // ../RTL/cortexm0ds_logic.v(9973)
  and u1085 (Dlyhu6, Klyhu6, Rlyhu6);  // ../RTL/cortexm0ds_logic.v(3216)
  and u10850 (n2924, Rs4ju6, vis_r8_o[11]);  // ../RTL/cortexm0ds_logic.v(9974)
  not u10851 (Zs8ju6, n2924);  // ../RTL/cortexm0ds_logic.v(9974)
  AL_MUX u10852 (
    .i0(Cg5ju6),
    .i1(Wc5ju6),
    .sel(C1epw6),
    .o(Ro8ju6));  // ../RTL/cortexm0ds_logic.v(9975)
  xor u10853 (n2925, Gt8ju6, Hu4ju6);  // ../RTL/cortexm0ds_logic.v(9976)
  not u10854 (C1epw6, n2925);  // ../RTL/cortexm0ds_logic.v(9976)
  and u10855 (n2926, Nt8ju6, Ut8ju6);  // ../RTL/cortexm0ds_logic.v(9977)
  not u10856 (Gt8ju6, n2926);  // ../RTL/cortexm0ds_logic.v(9977)
  or u10857 (Ut8ju6, I6jiu6, Gx4ju6);  // ../RTL/cortexm0ds_logic.v(9978)
  and u10858 (Nt8ju6, Bu8ju6, Ij5ju6);  // ../RTL/cortexm0ds_logic.v(9979)
  and u10859 (n2927, Sw4ju6, In8ju6);  // ../RTL/cortexm0ds_logic.v(9980)
  and u1086 (n25, Ylyhu6, Fmyhu6);  // ../RTL/cortexm0ds_logic.v(3217)
  not u10860 (Bu8ju6, n2927);  // ../RTL/cortexm0ds_logic.v(9980)
  and u10861 (n2928, Iu8ju6, Pu8ju6);  // ../RTL/cortexm0ds_logic.v(9981)
  not u10862 (Pomiu6, n2928);  // ../RTL/cortexm0ds_logic.v(9981)
  and u10863 (Pu8ju6, Wu8ju6, Dv8ju6);  // ../RTL/cortexm0ds_logic.v(9982)
  and u10864 (n2929, By4ju6, Eafpw6[12]);  // ../RTL/cortexm0ds_logic.v(9983)
  not u10865 (Dv8ju6, n2929);  // ../RTL/cortexm0ds_logic.v(9983)
  or u10866 (n2930, Affpw6[12], Kv8ju6);  // ../RTL/cortexm0ds_logic.v(9984)
  not u10867 (Wu8ju6, n2930);  // ../RTL/cortexm0ds_logic.v(9984)
  and u10868 (Kv8ju6, Iy4ju6, Rv8ju6);  // ../RTL/cortexm0ds_logic.v(9985)
  and u10869 (Iu8ju6, Yv8ju6, Fw8ju6);  // ../RTL/cortexm0ds_logic.v(9986)
  not u1087 (Klyhu6, n25);  // ../RTL/cortexm0ds_logic.v(3217)
  and u10870 (n2931, Ub5ju6, Mw8ju6);  // ../RTL/cortexm0ds_logic.v(9987)
  not u10871 (Fw8ju6, n2931);  // ../RTL/cortexm0ds_logic.v(9987)
  and u10872 (n2932, Tw8ju6, Ic5ju6);  // ../RTL/cortexm0ds_logic.v(9988)
  not u10873 (Mw8ju6, n2932);  // ../RTL/cortexm0ds_logic.v(9988)
  and u10874 (n2933, Ln0iu6, J1epw6);  // ../RTL/cortexm0ds_logic.v(9989)
  not u10875 (Tw8ju6, n2933);  // ../RTL/cortexm0ds_logic.v(9989)
  or u10876 (Yv8ju6, Ax8ju6, Ln0iu6);  // ../RTL/cortexm0ds_logic.v(9990)
  AL_MUX u10877 (
    .i0(Cg5ju6),
    .i1(Wc5ju6),
    .sel(J1epw6),
    .o(Ax8ju6));  // ../RTL/cortexm0ds_logic.v(9991)
  xor u10878 (n2934, Hx8ju6, Hu4ju6);  // ../RTL/cortexm0ds_logic.v(9992)
  not u10879 (J1epw6, n2934);  // ../RTL/cortexm0ds_logic.v(9992)
  or u1088 (n26, Mmyhu6, B7nhu6);  // ../RTL/cortexm0ds_logic.v(3218)
  and u10880 (n2935, Ox8ju6, Vx8ju6);  // ../RTL/cortexm0ds_logic.v(9993)
  not u10881 (Hx8ju6, n2935);  // ../RTL/cortexm0ds_logic.v(9993)
  or u10882 (Vx8ju6, Y8biu6, Gx4ju6);  // ../RTL/cortexm0ds_logic.v(9994)
  and u10883 (Ox8ju6, Cy8ju6, Ij5ju6);  // ../RTL/cortexm0ds_logic.v(9995)
  and u10884 (n2936, Sw4ju6, Rv8ju6);  // ../RTL/cortexm0ds_logic.v(9996)
  not u10885 (Cy8ju6, n2936);  // ../RTL/cortexm0ds_logic.v(9996)
  or u10886 (n2937, Fjmiu6, Xlmiu6);  // ../RTL/cortexm0ds_logic.v(9997)
  not u10887 (Ll8ju6, n2937);  // ../RTL/cortexm0ds_logic.v(9997)
  and u10888 (n2938, Jy8ju6, Qy8ju6);  // ../RTL/cortexm0ds_logic.v(9998)
  not u10889 (Xlmiu6, n2938);  // ../RTL/cortexm0ds_logic.v(9998)
  not u1089 (Ylyhu6, n26);  // ../RTL/cortexm0ds_logic.v(3218)
  and u10890 (Qy8ju6, Xy8ju6, Ez8ju6);  // ../RTL/cortexm0ds_logic.v(9999)
  and u10891 (n2939, By4ju6, Eafpw6[13]);  // ../RTL/cortexm0ds_logic.v(10000)
  not u10892 (Ez8ju6, n2939);  // ../RTL/cortexm0ds_logic.v(10000)
  or u10893 (n2940, Affpw6[13], Lz8ju6);  // ../RTL/cortexm0ds_logic.v(10001)
  not u10894 (Xy8ju6, n2940);  // ../RTL/cortexm0ds_logic.v(10001)
  and u10895 (Lz8ju6, Iy4ju6, Sz8ju6);  // ../RTL/cortexm0ds_logic.v(10002)
  and u10896 (Jy8ju6, Zz8ju6, G09ju6);  // ../RTL/cortexm0ds_logic.v(10003)
  and u10897 (n2941, Ub5ju6, N09ju6);  // ../RTL/cortexm0ds_logic.v(10004)
  not u10898 (G09ju6, n2941);  // ../RTL/cortexm0ds_logic.v(10004)
  and u10899 (n2942, U09ju6, Ic5ju6);  // ../RTL/cortexm0ds_logic.v(10005)
  buf u109 (Uthpw6[15], Z67ax6);  // ../RTL/cortexm0ds_logic.v(1882)
  and u1090 (Wkyhu6, Tmyhu6, Anyhu6);  // ../RTL/cortexm0ds_logic.v(3219)
  not u10900 (N09ju6, n2942);  // ../RTL/cortexm0ds_logic.v(10005)
  and u10901 (n2943, En0iu6, Q1epw6);  // ../RTL/cortexm0ds_logic.v(10006)
  not u10902 (U09ju6, n2943);  // ../RTL/cortexm0ds_logic.v(10006)
  or u10903 (Zz8ju6, B19ju6, En0iu6);  // ../RTL/cortexm0ds_logic.v(10007)
  AL_MUX u10904 (
    .i0(Cg5ju6),
    .i1(Wc5ju6),
    .sel(Q1epw6),
    .o(B19ju6));  // ../RTL/cortexm0ds_logic.v(10008)
  xor u10905 (n2944, I19ju6, Hu4ju6);  // ../RTL/cortexm0ds_logic.v(10009)
  not u10906 (Q1epw6, n2944);  // ../RTL/cortexm0ds_logic.v(10009)
  and u10907 (n2945, P19ju6, W19ju6);  // ../RTL/cortexm0ds_logic.v(10010)
  not u10908 (I19ju6, n2945);  // ../RTL/cortexm0ds_logic.v(10010)
  or u10909 (W19ju6, B5kiu6, Gx4ju6);  // ../RTL/cortexm0ds_logic.v(10011)
  and u1091 (n27, U5yhu6, Hnyhu6);  // ../RTL/cortexm0ds_logic.v(3220)
  and u10910 (P19ju6, D29ju6, Ij5ju6);  // ../RTL/cortexm0ds_logic.v(10012)
  and u10911 (n2946, Sw4ju6, Sz8ju6);  // ../RTL/cortexm0ds_logic.v(10013)
  not u10912 (D29ju6, n2946);  // ../RTL/cortexm0ds_logic.v(10013)
  and u10913 (n2947, K29ju6, R29ju6);  // ../RTL/cortexm0ds_logic.v(10014)
  not u10914 (Fjmiu6, n2947);  // ../RTL/cortexm0ds_logic.v(10014)
  and u10915 (R29ju6, Y29ju6, F39ju6);  // ../RTL/cortexm0ds_logic.v(10015)
  and u10916 (n2948, By4ju6, Eafpw6[14]);  // ../RTL/cortexm0ds_logic.v(10016)
  not u10917 (F39ju6, n2948);  // ../RTL/cortexm0ds_logic.v(10016)
  or u10918 (n2949, Affpw6[14], M39ju6);  // ../RTL/cortexm0ds_logic.v(10017)
  not u10919 (Y29ju6, n2949);  // ../RTL/cortexm0ds_logic.v(10017)
  not u1092 (Anyhu6, n27);  // ../RTL/cortexm0ds_logic.v(3220)
  and u10920 (M39ju6, Iy4ju6, T39ju6);  // ../RTL/cortexm0ds_logic.v(10018)
  and u10921 (K29ju6, A49ju6, H49ju6);  // ../RTL/cortexm0ds_logic.v(10019)
  and u10922 (n2950, Ub5ju6, O49ju6);  // ../RTL/cortexm0ds_logic.v(10020)
  not u10923 (H49ju6, n2950);  // ../RTL/cortexm0ds_logic.v(10020)
  and u10924 (n2951, V49ju6, Ic5ju6);  // ../RTL/cortexm0ds_logic.v(10021)
  not u10925 (O49ju6, n2951);  // ../RTL/cortexm0ds_logic.v(10021)
  and u10926 (n2952, Xm0iu6, X1epw6);  // ../RTL/cortexm0ds_logic.v(10022)
  not u10927 (V49ju6, n2952);  // ../RTL/cortexm0ds_logic.v(10022)
  or u10928 (A49ju6, C59ju6, Xm0iu6);  // ../RTL/cortexm0ds_logic.v(10023)
  AL_MUX u10929 (
    .i0(Cg5ju6),
    .i1(Wc5ju6),
    .sel(X1epw6),
    .o(C59ju6));  // ../RTL/cortexm0ds_logic.v(10024)
  or u1093 (Hnyhu6, Onyhu6, Vnyhu6);  // ../RTL/cortexm0ds_logic.v(3221)
  xor u10930 (n2953, J59ju6, Hu4ju6);  // ../RTL/cortexm0ds_logic.v(10025)
  not u10931 (X1epw6, n2953);  // ../RTL/cortexm0ds_logic.v(10025)
  and u10932 (n2954, Q59ju6, X59ju6);  // ../RTL/cortexm0ds_logic.v(10026)
  not u10933 (J59ju6, n2954);  // ../RTL/cortexm0ds_logic.v(10026)
  or u10934 (X59ju6, Gx4ju6, Cajiu6);  // ../RTL/cortexm0ds_logic.v(10027)
  and u10935 (Q59ju6, E69ju6, Ij5ju6);  // ../RTL/cortexm0ds_logic.v(10028)
  and u10936 (n2955, Sw4ju6, T39ju6);  // ../RTL/cortexm0ds_logic.v(10029)
  not u10937 (E69ju6, n2955);  // ../RTL/cortexm0ds_logic.v(10029)
  and u10938 (Wo7ju6, L69ju6, S69ju6);  // ../RTL/cortexm0ds_logic.v(10030)
  and u10939 (S69ju6, Z69ju6, G79ju6);  // ../RTL/cortexm0ds_logic.v(10031)
  and u1094 (n28, Coyhu6, Joyhu6);  // ../RTL/cortexm0ds_logic.v(3222)
  and u10940 (G79ju6, Vdmiu6, Ngmiu6);  // ../RTL/cortexm0ds_logic.v(10032)
  and u10941 (Ngmiu6, N79ju6, U79ju6);  // ../RTL/cortexm0ds_logic.v(10033)
  and u10942 (U79ju6, B89ju6, I89ju6);  // ../RTL/cortexm0ds_logic.v(10034)
  and u10943 (n2956, By4ju6, Eafpw6[15]);  // ../RTL/cortexm0ds_logic.v(10035)
  not u10944 (I89ju6, n2956);  // ../RTL/cortexm0ds_logic.v(10035)
  or u10945 (n2957, Affpw6[15], P89ju6);  // ../RTL/cortexm0ds_logic.v(10036)
  not u10946 (B89ju6, n2957);  // ../RTL/cortexm0ds_logic.v(10036)
  and u10947 (P89ju6, Iy4ju6, W89ju6);  // ../RTL/cortexm0ds_logic.v(10037)
  and u10948 (N79ju6, D99ju6, K99ju6);  // ../RTL/cortexm0ds_logic.v(10038)
  and u10949 (n2958, Ub5ju6, R99ju6);  // ../RTL/cortexm0ds_logic.v(10039)
  not u1095 (Onyhu6, n28);  // ../RTL/cortexm0ds_logic.v(3222)
  not u10950 (K99ju6, n2958);  // ../RTL/cortexm0ds_logic.v(10039)
  and u10951 (n2959, Y99ju6, Ic5ju6);  // ../RTL/cortexm0ds_logic.v(10040)
  not u10952 (R99ju6, n2959);  // ../RTL/cortexm0ds_logic.v(10040)
  and u10953 (n2960, Qm0iu6, L2epw6);  // ../RTL/cortexm0ds_logic.v(10041)
  not u10954 (Y99ju6, n2960);  // ../RTL/cortexm0ds_logic.v(10041)
  or u10955 (D99ju6, Fa9ju6, Qm0iu6);  // ../RTL/cortexm0ds_logic.v(10042)
  AL_MUX u10956 (
    .i0(Cg5ju6),
    .i1(Wc5ju6),
    .sel(L2epw6),
    .o(Fa9ju6));  // ../RTL/cortexm0ds_logic.v(10043)
  xor u10957 (n2961, Ma9ju6, Hu4ju6);  // ../RTL/cortexm0ds_logic.v(10044)
  not u10958 (L2epw6, n2961);  // ../RTL/cortexm0ds_logic.v(10044)
  and u10959 (n2962, Ta9ju6, Ab9ju6);  // ../RTL/cortexm0ds_logic.v(10045)
  or u1096 (Coyhu6, Eiyhu6, I6yhu6);  // ../RTL/cortexm0ds_logic.v(3223)
  not u10960 (Ma9ju6, n2962);  // ../RTL/cortexm0ds_logic.v(10045)
  or u10961 (Ab9ju6, Gx4ju6, Qjoiu6);  // ../RTL/cortexm0ds_logic.v(10046)
  and u10962 (Ta9ju6, Hb9ju6, Ij5ju6);  // ../RTL/cortexm0ds_logic.v(10047)
  and u10963 (n2963, Sw4ju6, W89ju6);  // ../RTL/cortexm0ds_logic.v(10048)
  not u10964 (Hb9ju6, n2963);  // ../RTL/cortexm0ds_logic.v(10048)
  and u10965 (Vdmiu6, Ob9ju6, Vb9ju6);  // ../RTL/cortexm0ds_logic.v(10049)
  and u10966 (Vb9ju6, Cc9ju6, Jc9ju6);  // ../RTL/cortexm0ds_logic.v(10050)
  and u10967 (n2964, By4ju6, Eafpw6[16]);  // ../RTL/cortexm0ds_logic.v(10051)
  not u10968 (Jc9ju6, n2964);  // ../RTL/cortexm0ds_logic.v(10051)
  or u10969 (n2965, Affpw6[16], Qc9ju6);  // ../RTL/cortexm0ds_logic.v(10052)
  and u1097 (n29, T8yhu6, Qoyhu6);  // ../RTL/cortexm0ds_logic.v(3224)
  not u10970 (Cc9ju6, n2965);  // ../RTL/cortexm0ds_logic.v(10052)
  and u10971 (Qc9ju6, Iy4ju6, Xc9ju6);  // ../RTL/cortexm0ds_logic.v(10053)
  and u10972 (Ob9ju6, Ed9ju6, Ld9ju6);  // ../RTL/cortexm0ds_logic.v(10054)
  and u10973 (n2966, Ub5ju6, Sd9ju6);  // ../RTL/cortexm0ds_logic.v(10055)
  not u10974 (Ld9ju6, n2966);  // ../RTL/cortexm0ds_logic.v(10055)
  and u10975 (n2967, Zd9ju6, Ic5ju6);  // ../RTL/cortexm0ds_logic.v(10056)
  not u10976 (Sd9ju6, n2967);  // ../RTL/cortexm0ds_logic.v(10056)
  and u10977 (n2968, Jm0iu6, Z2epw6);  // ../RTL/cortexm0ds_logic.v(10057)
  not u10978 (Zd9ju6, n2968);  // ../RTL/cortexm0ds_logic.v(10057)
  or u10979 (Ed9ju6, Ge9ju6, Jm0iu6);  // ../RTL/cortexm0ds_logic.v(10058)
  not u1098 (Tmyhu6, n29);  // ../RTL/cortexm0ds_logic.v(3224)
  AL_MUX u10980 (
    .i0(Cg5ju6),
    .i1(Wc5ju6),
    .sel(Z2epw6),
    .o(Ge9ju6));  // ../RTL/cortexm0ds_logic.v(10059)
  xor u10981 (n2969, Ne9ju6, Hu4ju6);  // ../RTL/cortexm0ds_logic.v(10060)
  not u10982 (Z2epw6, n2969);  // ../RTL/cortexm0ds_logic.v(10060)
  and u10983 (n2970, Ue9ju6, Bf9ju6);  // ../RTL/cortexm0ds_logic.v(10061)
  not u10984 (Ne9ju6, n2970);  // ../RTL/cortexm0ds_logic.v(10061)
  and u10985 (n2971, If9ju6, S8fpw6[5]);  // ../RTL/cortexm0ds_logic.v(10062)
  not u10986 (Bf9ju6, n2971);  // ../RTL/cortexm0ds_logic.v(10062)
  and u10987 (Ue9ju6, Pf9ju6, Ij5ju6);  // ../RTL/cortexm0ds_logic.v(10063)
  and u10988 (n2972, Sw4ju6, Xc9ju6);  // ../RTL/cortexm0ds_logic.v(10064)
  not u10989 (Pf9ju6, n2972);  // ../RTL/cortexm0ds_logic.v(10064)
  or u1099 (Qoyhu6, Xoyhu6, Epyhu6);  // ../RTL/cortexm0ds_logic.v(3225)
  and u10990 (Z69ju6, X7miu6, Wamiu6);  // ../RTL/cortexm0ds_logic.v(10065)
  and u10991 (Wamiu6, Wf9ju6, Dg9ju6);  // ../RTL/cortexm0ds_logic.v(10066)
  and u10992 (Dg9ju6, Kg9ju6, Rg9ju6);  // ../RTL/cortexm0ds_logic.v(10067)
  and u10993 (n2973, By4ju6, Eafpw6[17]);  // ../RTL/cortexm0ds_logic.v(10068)
  not u10994 (Rg9ju6, n2973);  // ../RTL/cortexm0ds_logic.v(10068)
  or u10995 (n2974, Affpw6[17], Yg9ju6);  // ../RTL/cortexm0ds_logic.v(10069)
  not u10996 (Kg9ju6, n2974);  // ../RTL/cortexm0ds_logic.v(10069)
  and u10997 (Yg9ju6, Iy4ju6, Fh9ju6);  // ../RTL/cortexm0ds_logic.v(10070)
  and u10998 (Wf9ju6, Mh9ju6, Th9ju6);  // ../RTL/cortexm0ds_logic.v(10071)
  and u10999 (n2975, Ub5ju6, Ai9ju6);  // ../RTL/cortexm0ds_logic.v(10072)
  not u11 (HPROT[0], n5200[0]);  // ../RTL/cortexm0ds_logic.v(15247)
  buf u110 (E1hpw6[3], Ftaax6);  // ../RTL/cortexm0ds_logic.v(2367)
  AL_MUX u1100 (
    .i0(Ighpw6[4]),
    .i1(Lpyhu6),
    .sel(Pkyhu6),
    .o(Xoyhu6));  // ../RTL/cortexm0ds_logic.v(3226)
  not u11000 (Th9ju6, n2975);  // ../RTL/cortexm0ds_logic.v(10072)
  and u11001 (n2976, Hi9ju6, Ic5ju6);  // ../RTL/cortexm0ds_logic.v(10073)
  not u11002 (Ai9ju6, n2976);  // ../RTL/cortexm0ds_logic.v(10073)
  and u11003 (n2977, Cm0iu6, G3epw6);  // ../RTL/cortexm0ds_logic.v(10074)
  not u11004 (Hi9ju6, n2977);  // ../RTL/cortexm0ds_logic.v(10074)
  or u11005 (Mh9ju6, Oi9ju6, Cm0iu6);  // ../RTL/cortexm0ds_logic.v(10075)
  AL_MUX u11006 (
    .i0(Cg5ju6),
    .i1(Wc5ju6),
    .sel(G3epw6),
    .o(Oi9ju6));  // ../RTL/cortexm0ds_logic.v(10076)
  xor u11007 (n2978, Vi9ju6, Hu4ju6);  // ../RTL/cortexm0ds_logic.v(10077)
  not u11008 (G3epw6, n2978);  // ../RTL/cortexm0ds_logic.v(10077)
  and u11009 (n2979, Cj9ju6, Jj9ju6);  // ../RTL/cortexm0ds_logic.v(10078)
  or u1101 (n30, Wdyhu6, Ighpw6[4]);  // ../RTL/cortexm0ds_logic.v(3227)
  not u11010 (Vi9ju6, n2979);  // ../RTL/cortexm0ds_logic.v(10078)
  and u11011 (n2980, If9ju6, S8fpw6[6]);  // ../RTL/cortexm0ds_logic.v(10079)
  not u11012 (Jj9ju6, n2980);  // ../RTL/cortexm0ds_logic.v(10079)
  and u11013 (Cj9ju6, Qj9ju6, Ij5ju6);  // ../RTL/cortexm0ds_logic.v(10080)
  and u11014 (n2981, Sw4ju6, Fh9ju6);  // ../RTL/cortexm0ds_logic.v(10081)
  not u11015 (Qj9ju6, n2981);  // ../RTL/cortexm0ds_logic.v(10081)
  and u11016 (X7miu6, Xj9ju6, Ek9ju6);  // ../RTL/cortexm0ds_logic.v(10082)
  and u11017 (Ek9ju6, Lk9ju6, Sk9ju6);  // ../RTL/cortexm0ds_logic.v(10083)
  and u11018 (n2982, By4ju6, Eafpw6[18]);  // ../RTL/cortexm0ds_logic.v(10084)
  not u11019 (Sk9ju6, n2982);  // ../RTL/cortexm0ds_logic.v(10084)
  not u1102 (Lpyhu6, n30);  // ../RTL/cortexm0ds_logic.v(3227)
  or u11020 (n2983, Affpw6[18], Zk9ju6);  // ../RTL/cortexm0ds_logic.v(10085)
  not u11021 (Lk9ju6, n2983);  // ../RTL/cortexm0ds_logic.v(10085)
  and u11022 (Zk9ju6, Iy4ju6, Gl9ju6);  // ../RTL/cortexm0ds_logic.v(10086)
  and u11023 (Xj9ju6, Nl9ju6, Ul9ju6);  // ../RTL/cortexm0ds_logic.v(10087)
  and u11024 (n2984, Ub5ju6, Bm9ju6);  // ../RTL/cortexm0ds_logic.v(10088)
  not u11025 (Ul9ju6, n2984);  // ../RTL/cortexm0ds_logic.v(10088)
  and u11026 (n2985, Im9ju6, Ic5ju6);  // ../RTL/cortexm0ds_logic.v(10089)
  not u11027 (Bm9ju6, n2985);  // ../RTL/cortexm0ds_logic.v(10089)
  and u11028 (n2986, Vl0iu6, N3epw6);  // ../RTL/cortexm0ds_logic.v(10090)
  not u11029 (Im9ju6, n2986);  // ../RTL/cortexm0ds_logic.v(10090)
  buf u1103 (vis_r5_o[6], X7spw6);  // ../RTL/cortexm0ds_logic.v(1909)
  or u11030 (Nl9ju6, Pm9ju6, Vl0iu6);  // ../RTL/cortexm0ds_logic.v(10091)
  AL_MUX u11031 (
    .i0(Cg5ju6),
    .i1(Wc5ju6),
    .sel(N3epw6),
    .o(Pm9ju6));  // ../RTL/cortexm0ds_logic.v(10092)
  xor u11032 (n2987, Wm9ju6, Hu4ju6);  // ../RTL/cortexm0ds_logic.v(10093)
  not u11033 (N3epw6, n2987);  // ../RTL/cortexm0ds_logic.v(10093)
  and u11034 (n2988, Dn9ju6, Kn9ju6);  // ../RTL/cortexm0ds_logic.v(10094)
  not u11035 (Wm9ju6, n2988);  // ../RTL/cortexm0ds_logic.v(10094)
  and u11036 (n2989, If9ju6, S8fpw6[7]);  // ../RTL/cortexm0ds_logic.v(10095)
  not u11037 (Kn9ju6, n2989);  // ../RTL/cortexm0ds_logic.v(10095)
  and u11038 (Dn9ju6, Rn9ju6, Ij5ju6);  // ../RTL/cortexm0ds_logic.v(10096)
  and u11039 (n2990, Sw4ju6, Gl9ju6);  // ../RTL/cortexm0ds_logic.v(10097)
  buf u1104 (vis_r5_o[12], Lpppw6);  // ../RTL/cortexm0ds_logic.v(1909)
  not u11040 (Rn9ju6, n2990);  // ../RTL/cortexm0ds_logic.v(10097)
  and u11041 (L69ju6, Yn9ju6, Fo9ju6);  // ../RTL/cortexm0ds_logic.v(10098)
  and u11042 (Fo9ju6, Z1miu6, Y4miu6);  // ../RTL/cortexm0ds_logic.v(10099)
  and u11043 (Y4miu6, Mo9ju6, To9ju6);  // ../RTL/cortexm0ds_logic.v(10100)
  and u11044 (To9ju6, Ap9ju6, Hp9ju6);  // ../RTL/cortexm0ds_logic.v(10101)
  and u11045 (n2991, By4ju6, Eafpw6[19]);  // ../RTL/cortexm0ds_logic.v(10102)
  not u11046 (Hp9ju6, n2991);  // ../RTL/cortexm0ds_logic.v(10102)
  or u11047 (n2992, Affpw6[19], Op9ju6);  // ../RTL/cortexm0ds_logic.v(10103)
  not u11048 (Ap9ju6, n2992);  // ../RTL/cortexm0ds_logic.v(10103)
  and u11049 (Op9ju6, Iy4ju6, Vp9ju6);  // ../RTL/cortexm0ds_logic.v(10104)
  and u1105 (n31, U5yhu6, Gqyhu6);  // ../RTL/cortexm0ds_logic.v(3229)
  and u11050 (Mo9ju6, Cq9ju6, Jq9ju6);  // ../RTL/cortexm0ds_logic.v(10105)
  and u11051 (n2993, Ub5ju6, Qq9ju6);  // ../RTL/cortexm0ds_logic.v(10106)
  not u11052 (Jq9ju6, n2993);  // ../RTL/cortexm0ds_logic.v(10106)
  and u11053 (n2994, Xq9ju6, Ic5ju6);  // ../RTL/cortexm0ds_logic.v(10107)
  not u11054 (Qq9ju6, n2994);  // ../RTL/cortexm0ds_logic.v(10107)
  and u11055 (n2995, Ol0iu6, U3epw6);  // ../RTL/cortexm0ds_logic.v(10108)
  not u11056 (Xq9ju6, n2995);  // ../RTL/cortexm0ds_logic.v(10108)
  or u11057 (Cq9ju6, Er9ju6, Ol0iu6);  // ../RTL/cortexm0ds_logic.v(10109)
  AL_MUX u11058 (
    .i0(Cg5ju6),
    .i1(Wc5ju6),
    .sel(U3epw6),
    .o(Er9ju6));  // ../RTL/cortexm0ds_logic.v(10110)
  xor u11059 (n2996, Lr9ju6, Hu4ju6);  // ../RTL/cortexm0ds_logic.v(10111)
  not u1106 (Zpyhu6, n31);  // ../RTL/cortexm0ds_logic.v(3229)
  not u11060 (U3epw6, n2996);  // ../RTL/cortexm0ds_logic.v(10111)
  and u11061 (n2997, Sr9ju6, Zr9ju6);  // ../RTL/cortexm0ds_logic.v(10112)
  not u11062 (Lr9ju6, n2997);  // ../RTL/cortexm0ds_logic.v(10112)
  or u11063 (Zr9ju6, Gx4ju6, I65iu6);  // ../RTL/cortexm0ds_logic.v(10113)
  and u11064 (Sr9ju6, Gs9ju6, Ij5ju6);  // ../RTL/cortexm0ds_logic.v(10114)
  and u11065 (n2998, Sw4ju6, Vp9ju6);  // ../RTL/cortexm0ds_logic.v(10115)
  not u11066 (Gs9ju6, n2998);  // ../RTL/cortexm0ds_logic.v(10115)
  and u11067 (Z1miu6, Ns9ju6, Us9ju6);  // ../RTL/cortexm0ds_logic.v(10116)
  and u11068 (Us9ju6, Bt9ju6, It9ju6);  // ../RTL/cortexm0ds_logic.v(10117)
  and u11069 (n2999, By4ju6, Eafpw6[20]);  // ../RTL/cortexm0ds_logic.v(10118)
  and u1107 (n32, Nqyhu6, Uqyhu6);  // ../RTL/cortexm0ds_logic.v(3230)
  not u11070 (It9ju6, n2999);  // ../RTL/cortexm0ds_logic.v(10118)
  or u11071 (n3000, Affpw6[20], Pt9ju6);  // ../RTL/cortexm0ds_logic.v(10119)
  not u11072 (Bt9ju6, n3000);  // ../RTL/cortexm0ds_logic.v(10119)
  and u11073 (Pt9ju6, Iy4ju6, Wt9ju6);  // ../RTL/cortexm0ds_logic.v(10120)
  and u11074 (Ns9ju6, Du9ju6, Ku9ju6);  // ../RTL/cortexm0ds_logic.v(10121)
  and u11075 (n3001, Ub5ju6, Ru9ju6);  // ../RTL/cortexm0ds_logic.v(10122)
  not u11076 (Ku9ju6, n3001);  // ../RTL/cortexm0ds_logic.v(10122)
  and u11077 (n3002, Yu9ju6, Ic5ju6);  // ../RTL/cortexm0ds_logic.v(10123)
  not u11078 (Ru9ju6, n3002);  // ../RTL/cortexm0ds_logic.v(10123)
  and u11079 (n3003, Al0iu6, B4epw6);  // ../RTL/cortexm0ds_logic.v(10124)
  not u1108 (Gqyhu6, n32);  // ../RTL/cortexm0ds_logic.v(3230)
  not u11080 (Yu9ju6, n3003);  // ../RTL/cortexm0ds_logic.v(10124)
  or u11081 (Du9ju6, Fv9ju6, Al0iu6);  // ../RTL/cortexm0ds_logic.v(10125)
  AL_MUX u11082 (
    .i0(Cg5ju6),
    .i1(Wc5ju6),
    .sel(B4epw6),
    .o(Fv9ju6));  // ../RTL/cortexm0ds_logic.v(10126)
  xor u11083 (n3004, Mv9ju6, Hu4ju6);  // ../RTL/cortexm0ds_logic.v(10127)
  not u11084 (B4epw6, n3004);  // ../RTL/cortexm0ds_logic.v(10127)
  and u11085 (n3005, Tv9ju6, Aw9ju6);  // ../RTL/cortexm0ds_logic.v(10128)
  not u11086 (Mv9ju6, n3005);  // ../RTL/cortexm0ds_logic.v(10128)
  or u11087 (Aw9ju6, Gx4ju6, P65iu6);  // ../RTL/cortexm0ds_logic.v(10129)
  and u11088 (Tv9ju6, Hw9ju6, Ij5ju6);  // ../RTL/cortexm0ds_logic.v(10130)
  and u11089 (n3006, Sw4ju6, Wt9ju6);  // ../RTL/cortexm0ds_logic.v(10131)
  and u1109 (Uqyhu6, Bryhu6, Iryhu6);  // ../RTL/cortexm0ds_logic.v(3231)
  not u11090 (Hw9ju6, n3006);  // ../RTL/cortexm0ds_logic.v(10131)
  and u11091 (Yn9ju6, Uvliu6, Azliu6);  // ../RTL/cortexm0ds_logic.v(10132)
  and u11092 (Azliu6, Ow9ju6, Vw9ju6);  // ../RTL/cortexm0ds_logic.v(10133)
  and u11093 (Vw9ju6, Cx9ju6, Jx9ju6);  // ../RTL/cortexm0ds_logic.v(10134)
  and u11094 (n3007, By4ju6, Eafpw6[21]);  // ../RTL/cortexm0ds_logic.v(10135)
  not u11095 (Jx9ju6, n3007);  // ../RTL/cortexm0ds_logic.v(10135)
  or u11096 (n3008, Affpw6[21], Qx9ju6);  // ../RTL/cortexm0ds_logic.v(10136)
  not u11097 (Cx9ju6, n3008);  // ../RTL/cortexm0ds_logic.v(10136)
  and u11098 (Qx9ju6, Iy4ju6, Xx9ju6);  // ../RTL/cortexm0ds_logic.v(10137)
  and u11099 (Ow9ju6, Ey9ju6, Ly9ju6);  // ../RTL/cortexm0ds_logic.v(10138)
  buf u111 (Fsdhu6, Z9opw6);  // ../RTL/cortexm0ds_logic.v(1890)
  or u1110 (Bryhu6, Ffyhu6, Mdhpw6[3]);  // ../RTL/cortexm0ds_logic.v(3232)
  and u11100 (n3009, Ub5ju6, Sy9ju6);  // ../RTL/cortexm0ds_logic.v(10139)
  not u11101 (Ly9ju6, n3009);  // ../RTL/cortexm0ds_logic.v(10139)
  and u11102 (n3010, Zy9ju6, Ic5ju6);  // ../RTL/cortexm0ds_logic.v(10140)
  not u11103 (Sy9ju6, n3010);  // ../RTL/cortexm0ds_logic.v(10140)
  and u11104 (n3011, Tk0iu6, I4epw6);  // ../RTL/cortexm0ds_logic.v(10141)
  not u11105 (Zy9ju6, n3011);  // ../RTL/cortexm0ds_logic.v(10141)
  or u11106 (Ey9ju6, Gz9ju6, Tk0iu6);  // ../RTL/cortexm0ds_logic.v(10142)
  AL_MUX u11107 (
    .i0(Cg5ju6),
    .i1(Wc5ju6),
    .sel(I4epw6),
    .o(Gz9ju6));  // ../RTL/cortexm0ds_logic.v(10143)
  xor u11108 (n3012, Nz9ju6, Hu4ju6);  // ../RTL/cortexm0ds_logic.v(10144)
  not u11109 (I4epw6, n3012);  // ../RTL/cortexm0ds_logic.v(10144)
  and u1111 (Ffyhu6, Pryhu6, Wryhu6);  // ../RTL/cortexm0ds_logic.v(3233)
  and u11110 (n3013, Uz9ju6, B0aju6);  // ../RTL/cortexm0ds_logic.v(10145)
  not u11111 (Nz9ju6, n3013);  // ../RTL/cortexm0ds_logic.v(10145)
  and u11112 (n3014, If9ju6, S8fpw6[10]);  // ../RTL/cortexm0ds_logic.v(10146)
  not u11113 (B0aju6, n3014);  // ../RTL/cortexm0ds_logic.v(10146)
  and u11114 (Uz9ju6, I0aju6, Ij5ju6);  // ../RTL/cortexm0ds_logic.v(10147)
  and u11115 (n3015, Sw4ju6, Xx9ju6);  // ../RTL/cortexm0ds_logic.v(10148)
  not u11116 (I0aju6, n3015);  // ../RTL/cortexm0ds_logic.v(10148)
  and u11117 (Uvliu6, P0aju6, W0aju6);  // ../RTL/cortexm0ds_logic.v(10149)
  and u11118 (W0aju6, D1aju6, K1aju6);  // ../RTL/cortexm0ds_logic.v(10150)
  and u11119 (n3016, By4ju6, Eafpw6[22]);  // ../RTL/cortexm0ds_logic.v(10151)
  or u1112 (n33, Dsyhu6, Ksyhu6);  // ../RTL/cortexm0ds_logic.v(3234)
  not u11120 (K1aju6, n3016);  // ../RTL/cortexm0ds_logic.v(10151)
  and u11121 (By4ju6, H6ghu6, R1aju6);  // ../RTL/cortexm0ds_logic.v(10152)
  or u11122 (R1aju6, Y1aju6, Pt2ju6);  // ../RTL/cortexm0ds_logic.v(10153)
  AL_MUX u11123 (
    .i0(F2aju6),
    .i1(Difiu6),
    .sel(Cyfpw6[4]),
    .o(Y1aju6));  // ../RTL/cortexm0ds_logic.v(10154)
  and u11124 (n3017, M2aju6, T2aju6);  // ../RTL/cortexm0ds_logic.v(10155)
  not u11125 (F2aju6, n3017);  // ../RTL/cortexm0ds_logic.v(10155)
  or u11126 (T2aju6, Qcoiu6, H4ghu6);  // ../RTL/cortexm0ds_logic.v(10156)
  or u11127 (n3018, A3aju6, H3aju6);  // ../RTL/cortexm0ds_logic.v(10157)
  not u11128 (M2aju6, n3018);  // ../RTL/cortexm0ds_logic.v(10157)
  or u11129 (n3019, Affpw6[22], O3aju6);  // ../RTL/cortexm0ds_logic.v(10158)
  not u1113 (Nqyhu6, n33);  // ../RTL/cortexm0ds_logic.v(3234)
  not u11130 (D1aju6, n3019);  // ../RTL/cortexm0ds_logic.v(10158)
  and u11131 (O3aju6, Iy4ju6, V3aju6);  // ../RTL/cortexm0ds_logic.v(10159)
  and u11132 (Iy4ju6, H6ghu6, C4aju6);  // ../RTL/cortexm0ds_logic.v(10160)
  or u11133 (C4aju6, J4aju6, S6aiu6);  // ../RTL/cortexm0ds_logic.v(10161)
  and u11134 (P0aju6, Q4aju6, X4aju6);  // ../RTL/cortexm0ds_logic.v(10162)
  and u11135 (n3020, Ub5ju6, E5aju6);  // ../RTL/cortexm0ds_logic.v(10163)
  not u11136 (X4aju6, n3020);  // ../RTL/cortexm0ds_logic.v(10163)
  and u11137 (n3021, L5aju6, Ic5ju6);  // ../RTL/cortexm0ds_logic.v(10164)
  not u11138 (E5aju6, n3021);  // ../RTL/cortexm0ds_logic.v(10164)
  and u11139 (n3022, Mk0iu6, P4epw6);  // ../RTL/cortexm0ds_logic.v(10165)
  AL_MUX u1114 (
    .i0(Rsyhu6),
    .i1(Ysyhu6),
    .sel(Ighpw6[3]),
    .o(Dsyhu6));  // ../RTL/cortexm0ds_logic.v(3235)
  not u11140 (L5aju6, n3022);  // ../RTL/cortexm0ds_logic.v(10165)
  or u11141 (Ub5ju6, Wk4ju6, Ys4ju6);  // ../RTL/cortexm0ds_logic.v(10166)
  and u11142 (Wk4ju6, S5aju6, H6ghu6);  // ../RTL/cortexm0ds_logic.v(10168)
  not u11143 (Ic5ju6, Wk4ju6);  // ../RTL/cortexm0ds_logic.v(10168)
  and u11144 (S5aju6, Md0iu6, H4ghu6);  // ../RTL/cortexm0ds_logic.v(10169)
  or u11145 (Q4aju6, Z5aju6, Mk0iu6);  // ../RTL/cortexm0ds_logic.v(10170)
  AL_MUX u11146 (
    .i0(Cg5ju6),
    .i1(Wc5ju6),
    .sel(P4epw6),
    .o(Z5aju6));  // ../RTL/cortexm0ds_logic.v(10171)
  xor u11147 (n3023, G6aju6, Hu4ju6);  // ../RTL/cortexm0ds_logic.v(10172)
  not u11148 (P4epw6, n3023);  // ../RTL/cortexm0ds_logic.v(10172)
  and u11149 (Ol6ju6, H6ghu6, N6aju6);  // ../RTL/cortexm0ds_logic.v(10173)
  not u1115 (n6019, Ypmhu6);  // ../RTL/cortexm0ds_logic.v(3132)
  not u11150 (Hu4ju6, Ol6ju6);  // ../RTL/cortexm0ds_logic.v(10173)
  and u11151 (n3024, U6aju6, B7aju6);  // ../RTL/cortexm0ds_logic.v(10174)
  not u11152 (N6aju6, n3024);  // ../RTL/cortexm0ds_logic.v(10174)
  and u11153 (B7aju6, I7aju6, P7aju6);  // ../RTL/cortexm0ds_logic.v(10175)
  and u11154 (n3025, W7aju6, Cyfpw6[4]);  // ../RTL/cortexm0ds_logic.v(10176)
  not u11155 (P7aju6, n3025);  // ../RTL/cortexm0ds_logic.v(10176)
  and u11156 (W7aju6, D8aju6, Hs0iu6);  // ../RTL/cortexm0ds_logic.v(10177)
  and u11157 (n3026, Wfoiu6, K8aju6);  // ../RTL/cortexm0ds_logic.v(10178)
  not u11158 (D8aju6, n3026);  // ../RTL/cortexm0ds_logic.v(10178)
  buf u11159 (Syehu6, Ozkbx6[18]);  // ../RTL/cortexm0ds_logic.v(3176)
  or u1116 (n34, Pdyhu6, Ighpw6[4]);  // ../RTL/cortexm0ds_logic.v(3237)
  and u11160 (I7aju6, R8aju6, Zu0iu6);  // ../RTL/cortexm0ds_logic.v(10180)
  and u11161 (n3027, Y8aju6, F9aju6);  // ../RTL/cortexm0ds_logic.v(10181)
  not u11162 (Zu0iu6, n3027);  // ../RTL/cortexm0ds_logic.v(10181)
  and u11163 (n3028, M9aju6, A3aju6);  // ../RTL/cortexm0ds_logic.v(10182)
  not u11164 (R8aju6, n3028);  // ../RTL/cortexm0ds_logic.v(10182)
  and u11165 (M9aju6, S2ziu6, C0ehu6);  // ../RTL/cortexm0ds_logic.v(10183)
  and u11166 (U6aju6, Lu0iu6, T9aju6);  // ../RTL/cortexm0ds_logic.v(10184)
  and u11167 (n3029, Bi0iu6, Tfjiu6);  // ../RTL/cortexm0ds_logic.v(10185)
  not u11168 (T9aju6, n3029);  // ../RTL/cortexm0ds_logic.v(10185)
  and u11169 (Lu0iu6, Aaaju6, Haaju6);  // ../RTL/cortexm0ds_logic.v(10186)
  not u1117 (Rsyhu6, n34);  // ../RTL/cortexm0ds_logic.v(3237)
  or u11170 (Haaju6, Ey2ju6, Ezniu6);  // ../RTL/cortexm0ds_logic.v(10187)
  not u11171 (Ezniu6, F23ju6);  // ../RTL/cortexm0ds_logic.v(10188)
  and u11172 (Aaaju6, Oaaju6, Vaaju6);  // ../RTL/cortexm0ds_logic.v(10189)
  and u11173 (n3030, Mo2ju6, C0ehu6);  // ../RTL/cortexm0ds_logic.v(10190)
  not u11174 (Vaaju6, n3030);  // ../RTL/cortexm0ds_logic.v(10190)
  and u11175 (n3031, L78ju6, D6kiu6);  // ../RTL/cortexm0ds_logic.v(10191)
  not u11176 (Oaaju6, n3031);  // ../RTL/cortexm0ds_logic.v(10191)
  and u11177 (n3032, Cbaju6, Jbaju6);  // ../RTL/cortexm0ds_logic.v(10192)
  not u11178 (G6aju6, n3032);  // ../RTL/cortexm0ds_logic.v(10192)
  AL_MUX u11179 (
    .i0(Qbaju6),
    .i1(Xk8ju6),
    .sel(D7fpw6[11]),
    .o(Jbaju6));  // ../RTL/cortexm0ds_logic.v(10193)
  and u1118 (Spyhu6, Mtyhu6, N5yhu6);  // ../RTL/cortexm0ds_logic.v(3238)
  not u11180 (Xk8ju6, Ui5ju6);  // ../RTL/cortexm0ds_logic.v(10194)
  and u11181 (Ui5ju6, If9ju6, S8fpw6[11]);  // ../RTL/cortexm0ds_logic.v(10195)
  buf u11182 (G0fhu6, Ozkbx6[17]);  // ../RTL/cortexm0ds_logic.v(3176)
  not u11183 (Gx4ju6, If9ju6);  // ../RTL/cortexm0ds_logic.v(10197)
  and u11184 (If9ju6, Xbaju6, Sy2ju6);  // ../RTL/cortexm0ds_logic.v(10198)
  and u11185 (Xbaju6, H6ghu6, Fd0iu6);  // ../RTL/cortexm0ds_logic.v(10199)
  and u11186 (Cbaju6, Ecaju6, Ij5ju6);  // ../RTL/cortexm0ds_logic.v(10200)
  and u11187 (n3033, Zf7ju6, S8fpw6[11]);  // ../RTL/cortexm0ds_logic.v(10201)
  not u11188 (Ij5ju6, n3033);  // ../RTL/cortexm0ds_logic.v(10201)
  and u11189 (Zf7ju6, Lcaju6, H6ghu6);  // ../RTL/cortexm0ds_logic.v(10202)
  and u1119 (n35, T8yhu6, Ttyhu6);  // ../RTL/cortexm0ds_logic.v(3239)
  and u11190 (Lcaju6, Pt2ju6, Hzziu6);  // ../RTL/cortexm0ds_logic.v(10203)
  and u11191 (n3034, Sw4ju6, V3aju6);  // ../RTL/cortexm0ds_logic.v(10204)
  not u11192 (Ecaju6, n3034);  // ../RTL/cortexm0ds_logic.v(10204)
  and u11193 (Sw4ju6, H6ghu6, Scaju6);  // ../RTL/cortexm0ds_logic.v(10206)
  not u11194 (Vy7ju6, Sw4ju6);  // ../RTL/cortexm0ds_logic.v(10206)
  and u11195 (n3035, Zcaju6, Gdaju6);  // ../RTL/cortexm0ds_logic.v(10207)
  not u11196 (Scaju6, n3035);  // ../RTL/cortexm0ds_logic.v(10207)
  and u11197 (Gdaju6, Ndaju6, Udaju6);  // ../RTL/cortexm0ds_logic.v(10208)
  and u11198 (n3036, H4ghu6, Beaju6);  // ../RTL/cortexm0ds_logic.v(10209)
  not u11199 (Udaju6, n3036);  // ../RTL/cortexm0ds_logic.v(10209)
  buf u112 (SLEEPHOLDACKn, Xbopw6);  // ../RTL/cortexm0ds_logic.v(1891)
  not u1120 (Mtyhu6, n35);  // ../RTL/cortexm0ds_logic.v(3239)
  and u11200 (n3037, Ieaju6, Peaju6);  // ../RTL/cortexm0ds_logic.v(10210)
  not u11201 (Beaju6, n3037);  // ../RTL/cortexm0ds_logic.v(10210)
  or u11202 (n3038, Owoiu6, Kfiiu6);  // ../RTL/cortexm0ds_logic.v(10211)
  not u11203 (Peaju6, n3038);  // ../RTL/cortexm0ds_logic.v(10211)
  and u11204 (Ieaju6, Weaju6, Dfaju6);  // ../RTL/cortexm0ds_logic.v(10212)
  or u11205 (Dfaju6, Wfoiu6, Vwaiu6);  // ../RTL/cortexm0ds_logic.v(10213)
  or u11206 (Weaju6, Y2oiu6, Ii0iu6);  // ../RTL/cortexm0ds_logic.v(10214)
  and u11207 (Ndaju6, Kfaju6, Rfaju6);  // ../RTL/cortexm0ds_logic.v(10215)
  and u11208 (n3039, Yfaju6, Whfiu6);  // ../RTL/cortexm0ds_logic.v(10216)
  not u11209 (Rfaju6, n3039);  // ../RTL/cortexm0ds_logic.v(10216)
  xor u1121 (n36, Wdyhu6, Pkyhu6);  // ../RTL/cortexm0ds_logic.v(3240)
  and u11210 (Yfaju6, Oiaiu6, Sq3ju6);  // ../RTL/cortexm0ds_logic.v(10217)
  and u11211 (n3040, Cyfpw6[3], Fgaju6);  // ../RTL/cortexm0ds_logic.v(10218)
  not u11212 (Kfaju6, n3040);  // ../RTL/cortexm0ds_logic.v(10218)
  and u11213 (n3041, Yn2ju6, Mgaju6);  // ../RTL/cortexm0ds_logic.v(10219)
  not u11214 (Fgaju6, n3041);  // ../RTL/cortexm0ds_logic.v(10219)
  or u11215 (Mgaju6, Z6oiu6, Wfoiu6);  // ../RTL/cortexm0ds_logic.v(10220)
  and u11216 (Zcaju6, Tgaju6, Ahaju6);  // ../RTL/cortexm0ds_logic.v(10221)
  and u11217 (n3042, Pt2ju6, Pthiu6);  // ../RTL/cortexm0ds_logic.v(10222)
  not u11218 (Ahaju6, n3042);  // ../RTL/cortexm0ds_logic.v(10222)
  or u11219 (Tgaju6, Y2oiu6, Cyfpw6[7]);  // ../RTL/cortexm0ds_logic.v(10223)
  not u1122 (Ttyhu6, n36);  // ../RTL/cortexm0ds_logic.v(3240)
  or u11220 (n3043, Tt4ju6, Mt4ju6);  // ../RTL/cortexm0ds_logic.v(10224)
  not u11221 (Wc5ju6, n3043);  // ../RTL/cortexm0ds_logic.v(10224)
  and u11222 (n3044, Hhaju6, Ohaju6);  // ../RTL/cortexm0ds_logic.v(10225)
  not u11223 (Tt4ju6, n3044);  // ../RTL/cortexm0ds_logic.v(10225)
  and u11224 (n3045, Vhaju6, H4ghu6);  // ../RTL/cortexm0ds_logic.v(10226)
  not u11225 (Ohaju6, n3045);  // ../RTL/cortexm0ds_logic.v(10226)
  and u11226 (Vhaju6, Ciaju6, Tr0iu6);  // ../RTL/cortexm0ds_logic.v(10227)
  or u11227 (Ciaju6, Hs0iu6, Kfiiu6);  // ../RTL/cortexm0ds_logic.v(10228)
  or u11228 (Hhaju6, Szniu6, Wfoiu6);  // ../RTL/cortexm0ds_logic.v(10229)
  or u11229 (n3046, Ys4ju6, Mt4ju6);  // ../RTL/cortexm0ds_logic.v(10230)
  buf u1123 (vis_r5_o[7], Aurpw6);  // ../RTL/cortexm0ds_logic.v(1909)
  not u11230 (Cg5ju6, n3046);  // ../RTL/cortexm0ds_logic.v(10230)
  and u11231 (Mt4ju6, H6ghu6, Jiaju6);  // ../RTL/cortexm0ds_logic.v(10231)
  and u11232 (n3047, Qiaju6, Xiaju6);  // ../RTL/cortexm0ds_logic.v(10232)
  not u11233 (Jiaju6, n3047);  // ../RTL/cortexm0ds_logic.v(10232)
  and u11234 (Qiaju6, Ejaju6, Ljaju6);  // ../RTL/cortexm0ds_logic.v(10233)
  and u11235 (n3048, Ae0iu6, N3ziu6);  // ../RTL/cortexm0ds_logic.v(10234)
  not u11236 (Ljaju6, n3048);  // ../RTL/cortexm0ds_logic.v(10234)
  AL_MUX u11237 (
    .i0(Sjaju6),
    .i1(Zjaju6),
    .sel(Cyfpw6[6]),
    .o(Ejaju6));  // ../RTL/cortexm0ds_logic.v(10235)
  or u11238 (Zjaju6, Y2oiu6, R75iu6);  // ../RTL/cortexm0ds_logic.v(10236)
  or u11239 (Sjaju6, Yn2ju6, Cyfpw6[4]);  // ../RTL/cortexm0ds_logic.v(10237)
  buf u1124 (vis_r5_o[13], Lnppw6);  // ../RTL/cortexm0ds_logic.v(1909)
  and u11240 (Ys4ju6, Gkaju6, Nkaju6);  // ../RTL/cortexm0ds_logic.v(10238)
  buf u11241 (U1fhu6, Ozkbx6[16]);  // ../RTL/cortexm0ds_logic.v(3176)
  not u11242 (Nkaju6, Tgaju6);  // ../RTL/cortexm0ds_logic.v(10239)
  and u11243 (Gkaju6, H6ghu6, Qyniu6);  // ../RTL/cortexm0ds_logic.v(10240)
  not u11244 (Xe0ju6, Nzoiu6);  // ../RTL/cortexm0ds_logic.v(10241)
  and u11245 (Nzoiu6, I6jiu6, Oviiu6);  // ../RTL/cortexm0ds_logic.v(10242)
  not u11246 (Utohu6, Ukaju6);  // ../RTL/cortexm0ds_logic.v(10243)
  AL_MUX u11247 (
    .i0(Ii0iu6),
    .i1(Blaju6),
    .sel(HREADY),
    .o(Ukaju6));  // ../RTL/cortexm0ds_logic.v(10244)
  and u11248 (Blaju6, Ilaju6, Plaju6);  // ../RTL/cortexm0ds_logic.v(10245)
  and u11249 (Plaju6, Wlaju6, Dmaju6);  // ../RTL/cortexm0ds_logic.v(10246)
  and u1125 (n37, T8yhu6, Ouyhu6);  // ../RTL/cortexm0ds_logic.v(3242)
  and u11250 (Dmaju6, Kmaju6, Rmaju6);  // ../RTL/cortexm0ds_logic.v(10247)
  and u11251 (n3049, Ymaju6, Eoyiu6);  // ../RTL/cortexm0ds_logic.v(10248)
  not u11252 (Rmaju6, n3049);  // ../RTL/cortexm0ds_logic.v(10248)
  or u11253 (n3050, H3piu6, Lkaiu6);  // ../RTL/cortexm0ds_logic.v(10249)
  not u11254 (Ymaju6, n3050);  // ../RTL/cortexm0ds_logic.v(10249)
  and u11255 (Kmaju6, Fnaju6, Mnaju6);  // ../RTL/cortexm0ds_logic.v(10250)
  and u11256 (n3051, Tnaju6, W8aiu6);  // ../RTL/cortexm0ds_logic.v(10251)
  not u11257 (Mnaju6, n3051);  // ../RTL/cortexm0ds_logic.v(10251)
  and u11258 (Tnaju6, Cyfpw6[3], Aoaju6);  // ../RTL/cortexm0ds_logic.v(10252)
  and u11259 (n3052, Hoaju6, Ooaju6);  // ../RTL/cortexm0ds_logic.v(10253)
  not u1126 (Huyhu6, n37);  // ../RTL/cortexm0ds_logic.v(3242)
  not u11260 (Aoaju6, n3052);  // ../RTL/cortexm0ds_logic.v(10253)
  and u11261 (Ooaju6, Voaju6, T0hhu6);  // ../RTL/cortexm0ds_logic.v(10254)
  or u11262 (n3053, Ftjiu6, D7fpw6[3]);  // ../RTL/cortexm0ds_logic.v(10255)
  not u11263 (Voaju6, n3053);  // ../RTL/cortexm0ds_logic.v(10255)
  or u11264 (n3054, Rg2ju6, Q5aiu6);  // ../RTL/cortexm0ds_logic.v(10256)
  not u11265 (Hoaju6, n3054);  // ../RTL/cortexm0ds_logic.v(10256)
  and u11266 (n3055, Cpaju6, Jpaju6);  // ../RTL/cortexm0ds_logic.v(10257)
  not u11267 (Fnaju6, n3055);  // ../RTL/cortexm0ds_logic.v(10257)
  or u11268 (n3056, Qpaju6, D7fpw6[10]);  // ../RTL/cortexm0ds_logic.v(10258)
  not u11269 (Jpaju6, n3056);  // ../RTL/cortexm0ds_logic.v(10258)
  xor u1127 (n38, Vuyhu6, Cvyhu6);  // ../RTL/cortexm0ds_logic.v(3243)
  and u11270 (Cpaju6, D7fpw6[8], J9kiu6);  // ../RTL/cortexm0ds_logic.v(10259)
  and u11271 (Wlaju6, Xpaju6, Eqaju6);  // ../RTL/cortexm0ds_logic.v(10260)
  and u11272 (n3057, Wwziu6, Lqaju6);  // ../RTL/cortexm0ds_logic.v(10261)
  not u11273 (Eqaju6, n3057);  // ../RTL/cortexm0ds_logic.v(10261)
  and u11274 (n3058, Y2oiu6, Sqaju6);  // ../RTL/cortexm0ds_logic.v(10262)
  not u11275 (Lqaju6, n3058);  // ../RTL/cortexm0ds_logic.v(10262)
  or u11276 (Sqaju6, Zqaju6, Cyfpw6[5]);  // ../RTL/cortexm0ds_logic.v(10263)
  and u11277 (Xpaju6, Graju6, Nraju6);  // ../RTL/cortexm0ds_logic.v(10264)
  and u11278 (n3059, Btoiu6, Uraju6);  // ../RTL/cortexm0ds_logic.v(10265)
  not u11279 (Nraju6, n3059);  // ../RTL/cortexm0ds_logic.v(10265)
  not u1128 (Ouyhu6, n38);  // ../RTL/cortexm0ds_logic.v(3243)
  and u11280 (n3060, Ctziu6, Bsaju6);  // ../RTL/cortexm0ds_logic.v(10266)
  not u11281 (Uraju6, n3060);  // ../RTL/cortexm0ds_logic.v(10266)
  and u11282 (n3061, U98iu6, Xe8iu6);  // ../RTL/cortexm0ds_logic.v(10267)
  not u11283 (Bsaju6, n3061);  // ../RTL/cortexm0ds_logic.v(10267)
  or u11284 (n3062, Cyfpw6[1], H4ghu6);  // ../RTL/cortexm0ds_logic.v(10268)
  not u11285 (Btoiu6, n3062);  // ../RTL/cortexm0ds_logic.v(10268)
  and u11286 (n3063, Isaju6, F23ju6);  // ../RTL/cortexm0ds_logic.v(10269)
  not u11287 (Graju6, n3063);  // ../RTL/cortexm0ds_logic.v(10269)
  and u11288 (Isaju6, Frziu6, Qe8iu6);  // ../RTL/cortexm0ds_logic.v(10270)
  and u11289 (Ilaju6, Psaju6, Wsaju6);  // ../RTL/cortexm0ds_logic.v(10271)
  and u1129 (n39, U5yhu6, Jvyhu6);  // ../RTL/cortexm0ds_logic.v(3244)
  and u11290 (Wsaju6, Dtaju6, K76ow6);  // ../RTL/cortexm0ds_logic.v(10272)
  or u11291 (K76ow6, P5kiu6, Sijiu6);  // ../RTL/cortexm0ds_logic.v(10273)
  and u11292 (Dtaju6, R76ow6, Y76ow6);  // ../RTL/cortexm0ds_logic.v(10274)
  or u11293 (Y76ow6, Ctziu6, V58ju6);  // ../RTL/cortexm0ds_logic.v(10275)
  or u11294 (Ctziu6, Jcaiu6, R75iu6);  // ../RTL/cortexm0ds_logic.v(10277)
  and u11295 (n3064, M86ow6, Tfjiu6);  // ../RTL/cortexm0ds_logic.v(10278)
  not u11296 (R76ow6, n3064);  // ../RTL/cortexm0ds_logic.v(10278)
  and u11297 (n3065, T86ow6, A96ow6);  // ../RTL/cortexm0ds_logic.v(10279)
  not u11298 (M86ow6, n3065);  // ../RTL/cortexm0ds_logic.v(10279)
  and u11299 (n3066, H96ow6, W8aiu6);  // ../RTL/cortexm0ds_logic.v(10280)
  not u113 (E6phu6, Xbopw6);  // ../RTL/cortexm0ds_logic.v(1892)
  not u1130 (Auyhu6, n39);  // ../RTL/cortexm0ds_logic.v(3244)
  not u11300 (A96ow6, n3066);  // ../RTL/cortexm0ds_logic.v(10280)
  or u11301 (n3067, O96ow6, Cyfpw6[5]);  // ../RTL/cortexm0ds_logic.v(10281)
  not u11302 (H96ow6, n3067);  // ../RTL/cortexm0ds_logic.v(10281)
  and u11303 (T86ow6, V96ow6, P5kiu6);  // ../RTL/cortexm0ds_logic.v(10282)
  not u11304 (P5kiu6, Lijiu6);  // ../RTL/cortexm0ds_logic.v(10283)
  and u11305 (Lijiu6, Whfiu6, Y7ghu6);  // ../RTL/cortexm0ds_logic.v(10284)
  and u11306 (n3068, Ca6ow6, Ae0iu6);  // ../RTL/cortexm0ds_logic.v(10285)
  not u11307 (V96ow6, n3068);  // ../RTL/cortexm0ds_logic.v(10285)
  and u11308 (Ca6ow6, U4kiu6, I30ju6);  // ../RTL/cortexm0ds_logic.v(10286)
  and u11309 (Psaju6, Ja6ow6, Qa6ow6);  // ../RTL/cortexm0ds_logic.v(10287)
  and u1131 (n40, Qvyhu6, Xvyhu6);  // ../RTL/cortexm0ds_logic.v(3245)
  or u11310 (Qa6ow6, Xa6ow6, Jcaiu6);  // ../RTL/cortexm0ds_logic.v(10288)
  and u11311 (n3069, Eb6ow6, Zraiu6);  // ../RTL/cortexm0ds_logic.v(10289)
  not u11312 (Ja6ow6, n3069);  // ../RTL/cortexm0ds_logic.v(10289)
  and u11313 (n3070, Lb6ow6, Sb6ow6);  // ../RTL/cortexm0ds_logic.v(10290)
  not u11314 (Eb6ow6, n3070);  // ../RTL/cortexm0ds_logic.v(10290)
  and u11315 (Sb6ow6, Zb6ow6, Gc6ow6);  // ../RTL/cortexm0ds_logic.v(10291)
  and u11316 (Gc6ow6, Nc6ow6, Kb0ju6);  // ../RTL/cortexm0ds_logic.v(10292)
  and u11317 (n3071, Nyiiu6, Mtjiu6);  // ../RTL/cortexm0ds_logic.v(10293)
  not u11318 (Kb0ju6, n3071);  // ../RTL/cortexm0ds_logic.v(10293)
  and u11319 (Nc6ow6, Xs0ju6, Xl0ju6);  // ../RTL/cortexm0ds_logic.v(10294)
  not u1132 (Jvyhu6, n40);  // ../RTL/cortexm0ds_logic.v(3245)
  and u11320 (Zb6ow6, Uc6ow6, Bd6ow6);  // ../RTL/cortexm0ds_logic.v(10295)
  and u11321 (n3072, Dxziu6, Id6ow6);  // ../RTL/cortexm0ds_logic.v(10296)
  not u11322 (Bd6ow6, n3072);  // ../RTL/cortexm0ds_logic.v(10296)
  and u11323 (n3073, Pd6ow6, Wd6ow6);  // ../RTL/cortexm0ds_logic.v(10297)
  not u11324 (Id6ow6, n3073);  // ../RTL/cortexm0ds_logic.v(10297)
  and u11325 (n3074, De6ow6, Frziu6);  // ../RTL/cortexm0ds_logic.v(10298)
  not u11326 (Wd6ow6, n3074);  // ../RTL/cortexm0ds_logic.v(10298)
  and u11327 (Uc6ow6, Ke6ow6, Re6ow6);  // ../RTL/cortexm0ds_logic.v(10299)
  and u11328 (n3075, Ye6ow6, Cyfpw6[0]);  // ../RTL/cortexm0ds_logic.v(10300)
  not u11329 (Ke6ow6, n3075);  // ../RTL/cortexm0ds_logic.v(10300)
  and u1133 (Xvyhu6, Ewyhu6, Lwyhu6);  // ../RTL/cortexm0ds_logic.v(3246)
  and u11330 (Ye6ow6, Omyiu6, Ff6ow6);  // ../RTL/cortexm0ds_logic.v(10301)
  or u11331 (Ff6ow6, Tr0iu6, D31ju6);  // ../RTL/cortexm0ds_logic.v(10302)
  and u11332 (Lb6ow6, Mf6ow6, Tf6ow6);  // ../RTL/cortexm0ds_logic.v(10303)
  and u11333 (Tf6ow6, Ag6ow6, Hg6ow6);  // ../RTL/cortexm0ds_logic.v(10304)
  and u11334 (n3076, Il3ju6, A95iu6);  // ../RTL/cortexm0ds_logic.v(10305)
  not u11335 (Hg6ow6, n3076);  // ../RTL/cortexm0ds_logic.v(10305)
  and u11336 (Ag6ow6, Og6ow6, Vg6ow6);  // ../RTL/cortexm0ds_logic.v(10306)
  and u11337 (n3077, Evyiu6, D7fpw6[15]);  // ../RTL/cortexm0ds_logic.v(10307)
  not u11338 (Vg6ow6, n3077);  // ../RTL/cortexm0ds_logic.v(10307)
  and u11339 (n3078, N3ziu6, Xzmiu6);  // ../RTL/cortexm0ds_logic.v(10308)
  and u1134 (n41, Swyhu6, Zwyhu6);  // ../RTL/cortexm0ds_logic.v(3247)
  not u11340 (Og6ow6, n3078);  // ../RTL/cortexm0ds_logic.v(10308)
  and u11341 (Mf6ow6, Ch6ow6, Jh6ow6);  // ../RTL/cortexm0ds_logic.v(10309)
  AL_MUX u11342 (
    .i0(Qh6ow6),
    .i1(Xh6ow6),
    .sel(C0ehu6),
    .o(Jh6ow6));  // ../RTL/cortexm0ds_logic.v(10310)
  and u11343 (Xh6ow6, Ei6ow6, Li6ow6);  // ../RTL/cortexm0ds_logic.v(10311)
  and u11344 (Li6ow6, Si6ow6, Zi6ow6);  // ../RTL/cortexm0ds_logic.v(10312)
  and u11345 (Zi6ow6, Gj6ow6, Geaiu6);  // ../RTL/cortexm0ds_logic.v(10313)
  or u11346 (Gj6ow6, Nj6ow6, D7fpw6[11]);  // ../RTL/cortexm0ds_logic.v(10314)
  and u11347 (Si6ow6, Uj6ow6, Bk6ow6);  // ../RTL/cortexm0ds_logic.v(10315)
  and u11348 (n3079, Ik6ow6, D7fpw6[9]);  // ../RTL/cortexm0ds_logic.v(10316)
  not u11349 (Bk6ow6, n3079);  // ../RTL/cortexm0ds_logic.v(10316)
  not u1135 (Lwyhu6, n41);  // ../RTL/cortexm0ds_logic.v(3247)
  AL_MUX u11350 (
    .i0(Pk6ow6),
    .i1(Wk6ow6),
    .sel(D7fpw6[7]),
    .o(Ik6ow6));  // ../RTL/cortexm0ds_logic.v(10317)
  and u11351 (n3080, Dl6ow6, Kl6ow6);  // ../RTL/cortexm0ds_logic.v(10318)
  not u11352 (Wk6ow6, n3080);  // ../RTL/cortexm0ds_logic.v(10318)
  and u11353 (n3081, Y40ju6, D7fpw6[6]);  // ../RTL/cortexm0ds_logic.v(10319)
  not u11354 (Kl6ow6, n3081);  // ../RTL/cortexm0ds_logic.v(10319)
  or u11355 (Dl6ow6, Oviiu6, Gaziu6);  // ../RTL/cortexm0ds_logic.v(10320)
  or u11356 (n3082, Gkiiu6, D7fpw6[6]);  // ../RTL/cortexm0ds_logic.v(10321)
  not u11357 (Pk6ow6, n3082);  // ../RTL/cortexm0ds_logic.v(10321)
  and u11358 (n3083, Rl6ow6, Ftjiu6);  // ../RTL/cortexm0ds_logic.v(10322)
  not u11359 (Uj6ow6, n3083);  // ../RTL/cortexm0ds_logic.v(10322)
  and u1136 (Ewyhu6, Gxyhu6, Ftyhu6);  // ../RTL/cortexm0ds_logic.v(3248)
  or u11360 (Rl6ow6, Yl6ow6, Fm6ow6);  // ../RTL/cortexm0ds_logic.v(10323)
  or u11361 (n3084, O7ziu6, X1ziu6);  // ../RTL/cortexm0ds_logic.v(10324)
  not u11362 (Fm6ow6, n3084);  // ../RTL/cortexm0ds_logic.v(10324)
  AL_MUX u11363 (
    .i0(Mm6ow6),
    .i1(D7fpw6[12]),
    .sel(D7fpw6[13]),
    .o(Yl6ow6));  // ../RTL/cortexm0ds_logic.v(10325)
  and u11364 (n3085, Tm6ow6, An6ow6);  // ../RTL/cortexm0ds_logic.v(10326)
  not u11365 (Mm6ow6, n3085);  // ../RTL/cortexm0ds_logic.v(10326)
  or u11366 (n3086, X8ziu6, Jwiiu6);  // ../RTL/cortexm0ds_logic.v(10327)
  not u11367 (Tm6ow6, n3086);  // ../RTL/cortexm0ds_logic.v(10327)
  and u11368 (Ei6ow6, Hn6ow6, Y31ju6);  // ../RTL/cortexm0ds_logic.v(10328)
  and u11369 (Hn6ow6, On6ow6, Vn6ow6);  // ../RTL/cortexm0ds_logic.v(10329)
  and u1137 (n42, Mdhpw6[3], Nxyhu6);  // ../RTL/cortexm0ds_logic.v(3249)
  or u11370 (Vn6ow6, Co6ow6, Xuyiu6);  // ../RTL/cortexm0ds_logic.v(10330)
  or u11371 (n3087, Jo6ow6, Qo6ow6);  // ../RTL/cortexm0ds_logic.v(10331)
  not u11372 (Xuyiu6, n3087);  // ../RTL/cortexm0ds_logic.v(10331)
  AL_MUX u11373 (
    .i0(Kcziu6),
    .i1(Xo6ow6),
    .sel(D7fpw6[5]),
    .o(Qo6ow6));  // ../RTL/cortexm0ds_logic.v(10332)
  or u11374 (Xo6ow6, O95iu6, Ad8iu6);  // ../RTL/cortexm0ds_logic.v(10333)
  and u11375 (n3088, D7fpw6[8], D7fpw6[9]);  // ../RTL/cortexm0ds_logic.v(10334)
  not u11376 (Jo6ow6, n3088);  // ../RTL/cortexm0ds_logic.v(10334)
  and u11377 (n3089, Qxoiu6, D7fpw6[12]);  // ../RTL/cortexm0ds_logic.v(10335)
  not u11378 (On6ow6, n3089);  // ../RTL/cortexm0ds_logic.v(10335)
  and u11379 (n3090, Ep6ow6, F23ju6);  // ../RTL/cortexm0ds_logic.v(10336)
  not u1138 (Gxyhu6, n42);  // ../RTL/cortexm0ds_logic.v(3249)
  not u11380 (Qh6ow6, n3090);  // ../RTL/cortexm0ds_logic.v(10336)
  and u11381 (Ch6ow6, Lp6ow6, Sp6ow6);  // ../RTL/cortexm0ds_logic.v(10337)
  and u11382 (n3091, Pthiu6, S6aiu6);  // ../RTL/cortexm0ds_logic.v(10338)
  not u11383 (Sp6ow6, n3091);  // ../RTL/cortexm0ds_logic.v(10338)
  or u11384 (Lp6ow6, H95iu6, D7fpw6[11]);  // ../RTL/cortexm0ds_logic.v(10339)
  AL_MUX u11385 (
    .i0(Zp6ow6),
    .i1(H2fpw6[0]),
    .sel(G81ju6),
    .o(Ntohu6));  // ../RTL/cortexm0ds_logic.v(10340)
  and u11386 (n3092, Gq6ow6, Nq6ow6);  // ../RTL/cortexm0ds_logic.v(10341)
  not u11387 (Zp6ow6, n3092);  // ../RTL/cortexm0ds_logic.v(10341)
  and u11388 (Nq6ow6, Uq6ow6, Br6ow6);  // ../RTL/cortexm0ds_logic.v(10342)
  and u11389 (n3093, Fb1ju6, D7fpw6[8]);  // ../RTL/cortexm0ds_logic.v(10343)
  and u1139 (n43, Uxyhu6, Byyhu6);  // ../RTL/cortexm0ds_logic.v(3250)
  not u11390 (Br6ow6, n3093);  // ../RTL/cortexm0ds_logic.v(10343)
  and u11391 (n3094, P91ju6, D7fpw6[3]);  // ../RTL/cortexm0ds_logic.v(10344)
  not u11392 (Uq6ow6, n3094);  // ../RTL/cortexm0ds_logic.v(10344)
  and u11393 (Gq6ow6, Ir6ow6, Pr6ow6);  // ../RTL/cortexm0ds_logic.v(10345)
  and u11394 (n3095, D7fpw6[0], Ac1ju6);  // ../RTL/cortexm0ds_logic.v(10346)
  not u11395 (Pr6ow6, n3095);  // ../RTL/cortexm0ds_logic.v(10346)
  and u11396 (n3096, Wr6ow6, Ds6ow6);  // ../RTL/cortexm0ds_logic.v(10347)
  not u11397 (Gtohu6, n3096);  // ../RTL/cortexm0ds_logic.v(10347)
  and u11398 (Ds6ow6, Ks6ow6, Rs6ow6);  // ../RTL/cortexm0ds_logic.v(10348)
  and u11399 (n3097, Egziu6, Eafpw6[1]);  // ../RTL/cortexm0ds_logic.v(10349)
  buf u114 (C0ehu6, Ydopw6);  // ../RTL/cortexm0ds_logic.v(1893)
  not u1140 (Nxyhu6, n43);  // ../RTL/cortexm0ds_logic.v(3250)
  not u11400 (Rs6ow6, n3097);  // ../RTL/cortexm0ds_logic.v(10349)
  and u11401 (Ks6ow6, Ys6ow6, Sgziu6);  // ../RTL/cortexm0ds_logic.v(10350)
  or u11402 (Ys6ow6, Ft6ow6, Njciu6);  // ../RTL/cortexm0ds_logic.v(10351)
  and u11403 (Njciu6, Mt6ow6, Tt6ow6);  // ../RTL/cortexm0ds_logic.v(10352)
  and u11404 (Tt6ow6, Au6ow6, Hu6ow6);  // ../RTL/cortexm0ds_logic.v(10353)
  or u11405 (Hu6ow6, Cfliu6, Ou6ow6);  // ../RTL/cortexm0ds_logic.v(10354)
  and u11406 (Au6ow6, Vu6ow6, Mdliu6);  // ../RTL/cortexm0ds_logic.v(10355)
  and u11407 (n3098, Qfliu6, Cv6ow6);  // ../RTL/cortexm0ds_logic.v(10356)
  not u11408 (Vu6ow6, n3098);  // ../RTL/cortexm0ds_logic.v(10356)
  and u11409 (Mt6ow6, Jv6ow6, Qv6ow6);  // ../RTL/cortexm0ds_logic.v(10357)
  and u1141 (n44, Iyyhu6, Cvyhu6);  // ../RTL/cortexm0ds_logic.v(3251)
  or u11410 (Qv6ow6, Ycliu6, Xv6ow6);  // ../RTL/cortexm0ds_logic.v(10358)
  and u11411 (n3099, Aeliu6, Ew6ow6);  // ../RTL/cortexm0ds_logic.v(10359)
  not u11412 (Jv6ow6, n3099);  // ../RTL/cortexm0ds_logic.v(10359)
  and u11413 (Wr6ow6, Lw6ow6, Sw6ow6);  // ../RTL/cortexm0ds_logic.v(10360)
  and u11414 (n3100, Zsfpw6[0], Cmziu6);  // ../RTL/cortexm0ds_logic.v(10361)
  not u11415 (Sw6ow6, n3100);  // ../RTL/cortexm0ds_logic.v(10361)
  or u11416 (Lw6ow6, Zkhiu6, Ar8iu6);  // ../RTL/cortexm0ds_logic.v(10362)
  not u11417 (Zkhiu6, vis_pc_o[0]);  // ../RTL/cortexm0ds_logic.v(10363)
  not u11418 (Zsohu6, Zw6ow6);  // ../RTL/cortexm0ds_logic.v(10364)
  AL_MUX u11419 (
    .i0(Mr0iu6),
    .i1(Gx6ow6),
    .sel(HREADY),
    .o(Zw6ow6));  // ../RTL/cortexm0ds_logic.v(10365)
  not u1142 (Byyhu6, n44);  // ../RTL/cortexm0ds_logic.v(3251)
  and u11420 (Gx6ow6, Nx6ow6, Ux6ow6);  // ../RTL/cortexm0ds_logic.v(10366)
  and u11421 (Ux6ow6, By6ow6, Iy6ow6);  // ../RTL/cortexm0ds_logic.v(10367)
  and u11422 (Iy6ow6, Py6ow6, Wy6ow6);  // ../RTL/cortexm0ds_logic.v(10368)
  and u11423 (Wy6ow6, Dz6ow6, X5aiu6);  // ../RTL/cortexm0ds_logic.v(10369)
  and u11424 (Py6ow6, Kz6ow6, Rz6ow6);  // ../RTL/cortexm0ds_logic.v(10370)
  and u11425 (By6ow6, Yz6ow6, F07ow6);  // ../RTL/cortexm0ds_logic.v(10371)
  and u11426 (F07ow6, B1aiu6, Uloiu6);  // ../RTL/cortexm0ds_logic.v(10372)
  and u11427 (Yz6ow6, M07ow6, T07ow6);  // ../RTL/cortexm0ds_logic.v(10373)
  and u11428 (n3101, A17ow6, Cyfpw6[4]);  // ../RTL/cortexm0ds_logic.v(10374)
  not u11429 (T07ow6, n3101);  // ../RTL/cortexm0ds_logic.v(10374)
  and u1143 (n45, Pyyhu6, Wyyhu6);  // ../RTL/cortexm0ds_logic.v(3252)
  and u11430 (A17ow6, Cyfpw6[5], H17ow6);  // ../RTL/cortexm0ds_logic.v(10375)
  and u11431 (n3102, R2aiu6, O17ow6);  // ../RTL/cortexm0ds_logic.v(10376)
  not u11432 (H17ow6, n3102);  // ../RTL/cortexm0ds_logic.v(10376)
  and u11433 (n3103, Ae0iu6, D6kiu6);  // ../RTL/cortexm0ds_logic.v(10377)
  not u11434 (O17ow6, n3103);  // ../RTL/cortexm0ds_logic.v(10377)
  and u11435 (n3104, V17ow6, Htyiu6);  // ../RTL/cortexm0ds_logic.v(10378)
  not u11436 (M07ow6, n3104);  // ../RTL/cortexm0ds_logic.v(10378)
  or u11437 (n3105, C27ow6, D7fpw6[14]);  // ../RTL/cortexm0ds_logic.v(10379)
  not u11438 (V17ow6, n3105);  // ../RTL/cortexm0ds_logic.v(10379)
  and u11439 (Nx6ow6, J27ow6, Q27ow6);  // ../RTL/cortexm0ds_logic.v(10380)
  not u1144 (Uxyhu6, n45);  // ../RTL/cortexm0ds_logic.v(3252)
  and u11440 (Q27ow6, X27ow6, E37ow6);  // ../RTL/cortexm0ds_logic.v(10381)
  and u11441 (E37ow6, L37ow6, S37ow6);  // ../RTL/cortexm0ds_logic.v(10382)
  and u11442 (n3106, Z37ow6, K2aiu6);  // ../RTL/cortexm0ds_logic.v(10383)
  not u11443 (S37ow6, n3106);  // ../RTL/cortexm0ds_logic.v(10383)
  or u11444 (n3107, Sijiu6, Kq0iu6);  // ../RTL/cortexm0ds_logic.v(10384)
  not u11445 (Z37ow6, n3107);  // ../RTL/cortexm0ds_logic.v(10384)
  or u11446 (L37ow6, Jojiu6, E62ju6);  // ../RTL/cortexm0ds_logic.v(10385)
  not u11447 (E62ju6, G47ow6);  // ../RTL/cortexm0ds_logic.v(10386)
  and u11448 (X27ow6, N47ow6, U47ow6);  // ../RTL/cortexm0ds_logic.v(10387)
  and u11449 (n3108, B57ow6, Ii0iu6);  // ../RTL/cortexm0ds_logic.v(10388)
  and u1145 (n46, Dzyhu6, Kzyhu6);  // ../RTL/cortexm0ds_logic.v(3253)
  not u11450 (U47ow6, n3108);  // ../RTL/cortexm0ds_logic.v(10388)
  and u11451 (n3109, I57ow6, P57ow6);  // ../RTL/cortexm0ds_logic.v(10389)
  not u11452 (B57ow6, n3109);  // ../RTL/cortexm0ds_logic.v(10389)
  or u11453 (P57ow6, Yn2ju6, K9aiu6);  // ../RTL/cortexm0ds_logic.v(10390)
  and u11454 (I57ow6, W57ow6, D67ow6);  // ../RTL/cortexm0ds_logic.v(10391)
  and u11455 (n3110, K67ow6, Ae0iu6);  // ../RTL/cortexm0ds_logic.v(10392)
  not u11456 (D67ow6, n3110);  // ../RTL/cortexm0ds_logic.v(10392)
  and u11457 (K67ow6, I30ju6, Y2oiu6);  // ../RTL/cortexm0ds_logic.v(10393)
  or u11458 (W57ow6, E45iu6, L62ju6);  // ../RTL/cortexm0ds_logic.v(10394)
  and u11459 (n3111, R67ow6, Geaiu6);  // ../RTL/cortexm0ds_logic.v(10395)
  not u1146 (Wyyhu6, n46);  // ../RTL/cortexm0ds_logic.v(3253)
  not u11460 (N47ow6, n3111);  // ../RTL/cortexm0ds_logic.v(10395)
  and u11461 (n3112, Y67ow6, F77ow6);  // ../RTL/cortexm0ds_logic.v(10396)
  not u11462 (R67ow6, n3112);  // ../RTL/cortexm0ds_logic.v(10396)
  and u11463 (F77ow6, M77ow6, T77ow6);  // ../RTL/cortexm0ds_logic.v(10397)
  and u11464 (T77ow6, A87ow6, H87ow6);  // ../RTL/cortexm0ds_logic.v(10398)
  and u11465 (n3113, O87ow6, V87ow6);  // ../RTL/cortexm0ds_logic.v(10399)
  not u11466 (H87ow6, n3113);  // ../RTL/cortexm0ds_logic.v(10399)
  or u11467 (n3114, Q1ziu6, Gaziu6);  // ../RTL/cortexm0ds_logic.v(10400)
  not u11468 (V87ow6, n3114);  // ../RTL/cortexm0ds_logic.v(10400)
  not u11469 (Q1ziu6, Y31ju6);  // ../RTL/cortexm0ds_logic.v(10401)
  and u1147 (n47, Lbyhu6, Mdhpw6[0]);  // ../RTL/cortexm0ds_logic.v(3254)
  and u11470 (O87ow6, Nyiiu6, Evyiu6);  // ../RTL/cortexm0ds_logic.v(10402)
  and u11471 (n3115, Ipziu6, S6aiu6);  // ../RTL/cortexm0ds_logic.v(10403)
  not u11472 (A87ow6, n3115);  // ../RTL/cortexm0ds_logic.v(10403)
  or u11473 (n3116, Lkaiu6, Dxziu6);  // ../RTL/cortexm0ds_logic.v(10404)
  not u11474 (Ipziu6, n3116);  // ../RTL/cortexm0ds_logic.v(10404)
  and u11475 (M77ow6, C97ow6, J97ow6);  // ../RTL/cortexm0ds_logic.v(10405)
  and u11476 (n3117, Q97ow6, X97ow6);  // ../RTL/cortexm0ds_logic.v(10406)
  not u11477 (J97ow6, n3117);  // ../RTL/cortexm0ds_logic.v(10406)
  and u11478 (n3118, Vviiu6, Ea7ow6);  // ../RTL/cortexm0ds_logic.v(10407)
  not u11479 (C97ow6, n3118);  // ../RTL/cortexm0ds_logic.v(10407)
  not u1148 (Kzyhu6, n47);  // ../RTL/cortexm0ds_logic.v(3254)
  and u11480 (n3119, Nj6ow6, La7ow6);  // ../RTL/cortexm0ds_logic.v(10408)
  not u11481 (Ea7ow6, n3119);  // ../RTL/cortexm0ds_logic.v(10408)
  and u11482 (n3120, Y40ju6, Db0ju6);  // ../RTL/cortexm0ds_logic.v(10409)
  not u11483 (La7ow6, n3120);  // ../RTL/cortexm0ds_logic.v(10409)
  and u11484 (Y67ow6, Sa7ow6, Za7ow6);  // ../RTL/cortexm0ds_logic.v(10410)
  or u11485 (Za7ow6, Kgaiu6, Wthiu6);  // ../RTL/cortexm0ds_logic.v(10411)
  not u11486 (Wthiu6, K2aiu6);  // ../RTL/cortexm0ds_logic.v(10412)
  and u11487 (Sa7ow6, Gb7ow6, Nb7ow6);  // ../RTL/cortexm0ds_logic.v(10413)
  and u11488 (n3121, Ub7ow6, Q5aiu6);  // ../RTL/cortexm0ds_logic.v(10414)
  not u11489 (Nb7ow6, n3121);  // ../RTL/cortexm0ds_logic.v(10414)
  or u1149 (Dzyhu6, Pryhu6, Rzyhu6);  // ../RTL/cortexm0ds_logic.v(3255)
  and u11490 (n3122, Bc7ow6, Ic7ow6);  // ../RTL/cortexm0ds_logic.v(10415)
  not u11491 (Ub7ow6, n3122);  // ../RTL/cortexm0ds_logic.v(10415)
  and u11492 (n3123, Pc7ow6, Wc7ow6);  // ../RTL/cortexm0ds_logic.v(10416)
  not u11493 (Ic7ow6, n3123);  // ../RTL/cortexm0ds_logic.v(10416)
  or u11494 (n3124, H95iu6, Oviiu6);  // ../RTL/cortexm0ds_logic.v(10417)
  not u11495 (Wc7ow6, n3124);  // ../RTL/cortexm0ds_logic.v(10417)
  and u11496 (Pc7ow6, Dmiiu6, Jwiiu6);  // ../RTL/cortexm0ds_logic.v(10418)
  and u11497 (n3125, Dd7ow6, J8ziu6);  // ../RTL/cortexm0ds_logic.v(10419)
  not u11498 (Bc7ow6, n3125);  // ../RTL/cortexm0ds_logic.v(10419)
  and u11499 (J8ziu6, Kd7ow6, Wh0ju6);  // ../RTL/cortexm0ds_logic.v(10420)
  buf u115 (E1hpw6[12], Biaax6);  // ../RTL/cortexm0ds_logic.v(2367)
  or u1150 (n48, Ksyhu6, Vnyhu6);  // ../RTL/cortexm0ds_logic.v(3256)
  or u11500 (n3126, Ph0ju6, D7fpw6[5]);  // ../RTL/cortexm0ds_logic.v(10421)
  not u11501 (Kd7ow6, n3126);  // ../RTL/cortexm0ds_logic.v(10421)
  or u11502 (Ph0ju6, Aq1ju6, D7fpw6[7]);  // ../RTL/cortexm0ds_logic.v(10422)
  and u11503 (n3127, Uyiiu6, Rd7ow6);  // ../RTL/cortexm0ds_logic.v(10423)
  not u11504 (Gb7ow6, n3127);  // ../RTL/cortexm0ds_logic.v(10423)
  and u11505 (n3128, Yd7ow6, Fe7ow6);  // ../RTL/cortexm0ds_logic.v(10424)
  not u11506 (Rd7ow6, n3128);  // ../RTL/cortexm0ds_logic.v(10424)
  and u11507 (n3129, Wliiu6, Me7ow6);  // ../RTL/cortexm0ds_logic.v(10425)
  not u11508 (Fe7ow6, n3129);  // ../RTL/cortexm0ds_logic.v(10425)
  and u11509 (n3130, Ftjiu6, Te7ow6);  // ../RTL/cortexm0ds_logic.v(10426)
  not u1151 (Qvyhu6, n48);  // ../RTL/cortexm0ds_logic.v(3256)
  not u11510 (Me7ow6, n3130);  // ../RTL/cortexm0ds_logic.v(10426)
  and u11511 (n3131, Af7ow6, Uriiu6);  // ../RTL/cortexm0ds_logic.v(10427)
  not u11512 (Te7ow6, n3131);  // ../RTL/cortexm0ds_logic.v(10427)
  and u11513 (n3132, Hf7ow6, Of7ow6);  // ../RTL/cortexm0ds_logic.v(10428)
  not u11514 (Af7ow6, n3132);  // ../RTL/cortexm0ds_logic.v(10428)
  and u11515 (Of7ow6, Vf7ow6, Cg7ow6);  // ../RTL/cortexm0ds_logic.v(10429)
  or u11516 (Cg7ow6, Ar0ju6, D7fpw6[10]);  // ../RTL/cortexm0ds_logic.v(10430)
  or u11517 (Vf7ow6, Hk0ju6, Kcziu6);  // ../RTL/cortexm0ds_logic.v(10431)
  and u11518 (Hf7ow6, Qz0ju6, D7fpw6[14]);  // ../RTL/cortexm0ds_logic.v(10432)
  and u11519 (Qz0ju6, Jg7ow6, Qg7ow6);  // ../RTL/cortexm0ds_logic.v(10433)
  AL_MUX u1152 (
    .i0(Yzyhu6),
    .i1(Hgyhu6),
    .sel(Mdhpw6[3]),
    .o(Vnyhu6));  // ../RTL/cortexm0ds_logic.v(3257)
  and u11520 (n3133, Xg7ow6, D7fpw6[7]);  // ../RTL/cortexm0ds_logic.v(10434)
  not u11521 (Qg7ow6, n3133);  // ../RTL/cortexm0ds_logic.v(10434)
  and u11522 (n3134, D7fpw6[10], Eh7ow6);  // ../RTL/cortexm0ds_logic.v(10435)
  not u11523 (Jg7ow6, n3134);  // ../RTL/cortexm0ds_logic.v(10435)
  or u11524 (Eh7ow6, D7fpw6[8], Qe0ju6);  // ../RTL/cortexm0ds_logic.v(10436)
  and u11525 (n3135, Dmiiu6, Lh7ow6);  // ../RTL/cortexm0ds_logic.v(10438)
  not u11526 (Yd7ow6, n3135);  // ../RTL/cortexm0ds_logic.v(10438)
  and u11527 (n3136, Sh7ow6, Zh7ow6);  // ../RTL/cortexm0ds_logic.v(10439)
  not u11528 (Lh7ow6, n3136);  // ../RTL/cortexm0ds_logic.v(10439)
  or u11529 (Zh7ow6, H95iu6, D7fpw6[9]);  // ../RTL/cortexm0ds_logic.v(10440)
  buf u1153 (Ggehu6, Ozkbx6[30]);  // ../RTL/cortexm0ds_logic.v(3176)
  and u11530 (Sh7ow6, Z01ju6, Gi7ow6);  // ../RTL/cortexm0ds_logic.v(10441)
  or u11531 (Gi7ow6, Wiliu6, Gaziu6);  // ../RTL/cortexm0ds_logic.v(10442)
  and u11532 (n3137, Qxoiu6, Nbkiu6);  // ../RTL/cortexm0ds_logic.v(10443)
  not u11533 (Z01ju6, n3137);  // ../RTL/cortexm0ds_logic.v(10443)
  and u11534 (J27ow6, Ni7ow6, K0jiu6);  // ../RTL/cortexm0ds_logic.v(10444)
  and u11535 (Ni7ow6, Ui7ow6, Bj7ow6);  // ../RTL/cortexm0ds_logic.v(10445)
  and u11536 (n3138, Moaiu6, Us2ju6);  // ../RTL/cortexm0ds_logic.v(10446)
  not u11537 (Bj7ow6, n3138);  // ../RTL/cortexm0ds_logic.v(10446)
  or u11538 (Ui7ow6, Qojiu6, Cyfpw6[7]);  // ../RTL/cortexm0ds_logic.v(10447)
  or u11539 (Ssohu6, Ij7ow6, Pj7ow6);  // ../RTL/cortexm0ds_logic.v(10448)
  not u1154 (Yzyhu6, Yeyhu6);  // ../RTL/cortexm0ds_logic.v(3258)
  or u11540 (n3139, Wj7ow6, Dk7ow6);  // ../RTL/cortexm0ds_logic.v(10449)
  not u11541 (Pj7ow6, n3139);  // ../RTL/cortexm0ds_logic.v(10449)
  AL_MUX u11542 (
    .i0(Kk7ow6),
    .i1(S8fpw6[5]),
    .sel(Rk7ow6),
    .o(Ij7ow6));  // ../RTL/cortexm0ds_logic.v(10450)
  and u11543 (n3140, Yk7ow6, Fl7ow6);  // ../RTL/cortexm0ds_logic.v(10451)
  not u11544 (Kk7ow6, n3140);  // ../RTL/cortexm0ds_logic.v(10451)
  and u11545 (Fl7ow6, Ml7ow6, Tl7ow6);  // ../RTL/cortexm0ds_logic.v(10452)
  and u11546 (n3141, Am7ow6, Ppfpw6[5]);  // ../RTL/cortexm0ds_logic.v(10453)
  not u11547 (Tl7ow6, n3141);  // ../RTL/cortexm0ds_logic.v(10453)
  or u11548 (Ml7ow6, Dzjiu6, Hm7ow6);  // ../RTL/cortexm0ds_logic.v(10454)
  and u11549 (Yk7ow6, Om7ow6, Vm7ow6);  // ../RTL/cortexm0ds_logic.v(10455)
  and u1155 (n49, I6yhu6, F0zhu6);  // ../RTL/cortexm0ds_logic.v(3259)
  and u11550 (n3142, Cbbiu6, D7fpw6[10]);  // ../RTL/cortexm0ds_logic.v(10456)
  not u11551 (Vm7ow6, n3142);  // ../RTL/cortexm0ds_logic.v(10456)
  or u11552 (Om7ow6, A1kiu6, Cn7ow6);  // ../RTL/cortexm0ds_logic.v(10457)
  AL_MUX u11553 (
    .i0(Jn7ow6),
    .i1(X3fpw6[0]),
    .sel(O25iu6),
    .o(Lsohu6));  // ../RTL/cortexm0ds_logic.v(10458)
  and u11554 (n3143, HREADY, Qn7ow6);  // ../RTL/cortexm0ds_logic.v(10459)
  not u11555 (O25iu6, n3143);  // ../RTL/cortexm0ds_logic.v(10459)
  and u11556 (n3144, Xn7ow6, Eo7ow6);  // ../RTL/cortexm0ds_logic.v(10460)
  not u11557 (Qn7ow6, n3144);  // ../RTL/cortexm0ds_logic.v(10460)
  and u11558 (Eo7ow6, Lo7ow6, So7ow6);  // ../RTL/cortexm0ds_logic.v(10461)
  or u11559 (n3145, Zo7ow6, Ujjiu6);  // ../RTL/cortexm0ds_logic.v(10462)
  not u1156 (Ksyhu6, n49);  // ../RTL/cortexm0ds_logic.v(3259)
  not u11560 (So7ow6, n3145);  // ../RTL/cortexm0ds_logic.v(10462)
  and u11561 (n3146, Isiiu6, Dz6ow6);  // ../RTL/cortexm0ds_logic.v(10463)
  not u11562 (Zo7ow6, n3146);  // ../RTL/cortexm0ds_logic.v(10463)
  and u11563 (n3147, Gp7ow6, Np7ow6);  // ../RTL/cortexm0ds_logic.v(10464)
  not u11564 (Isiiu6, n3147);  // ../RTL/cortexm0ds_logic.v(10464)
  buf u11565 (I3fhu6, Ozkbx6[15]);  // ../RTL/cortexm0ds_logic.v(3176)
  not u11566 (Np7ow6, Qq2ju6);  // ../RTL/cortexm0ds_logic.v(10465)
  or u11567 (n3148, R2aiu6, Xojiu6);  // ../RTL/cortexm0ds_logic.v(10466)
  not u11568 (Gp7ow6, n3148);  // ../RTL/cortexm0ds_logic.v(10466)
  and u11569 (Lo7ow6, Up7ow6, Bq7ow6);  // ../RTL/cortexm0ds_logic.v(10467)
  and u1157 (n50, M0zhu6, Ziyhu6);  // ../RTL/cortexm0ds_logic.v(3260)
  and u11570 (n3149, Iq7ow6, Cyfpw6[0]);  // ../RTL/cortexm0ds_logic.v(10468)
  not u11571 (Bq7ow6, n3149);  // ../RTL/cortexm0ds_logic.v(10468)
  or u11572 (n3150, Kq0iu6, Cyfpw6[3]);  // ../RTL/cortexm0ds_logic.v(10469)
  not u11573 (Iq7ow6, n3150);  // ../RTL/cortexm0ds_logic.v(10469)
  and u11574 (Up7ow6, Pq7ow6, Wq7ow6);  // ../RTL/cortexm0ds_logic.v(10470)
  and u11575 (n3151, Dr7ow6, Kr7ow6);  // ../RTL/cortexm0ds_logic.v(10471)
  not u11576 (Wq7ow6, n3151);  // ../RTL/cortexm0ds_logic.v(10471)
  and u11577 (Dr7ow6, L45iu6, Zraiu6);  // ../RTL/cortexm0ds_logic.v(10472)
  and u11578 (n3152, Rr7ow6, Y31ju6);  // ../RTL/cortexm0ds_logic.v(10473)
  not u11579 (Pq7ow6, n3152);  // ../RTL/cortexm0ds_logic.v(10473)
  not u1158 (F0zhu6, n50);  // ../RTL/cortexm0ds_logic.v(3260)
  and u11580 (Rr7ow6, M7kiu6, Yr7ow6);  // ../RTL/cortexm0ds_logic.v(10474)
  or u11581 (Yr7ow6, D7fpw6[14], Fs7ow6);  // ../RTL/cortexm0ds_logic.v(10475)
  and u11582 (Xn7ow6, Ms7ow6, Ts7ow6);  // ../RTL/cortexm0ds_logic.v(10476)
  and u11583 (Ts7ow6, At7ow6, Ht7ow6);  // ../RTL/cortexm0ds_logic.v(10477)
  and u11584 (n3153, Ot7ow6, D7fpw6[3]);  // ../RTL/cortexm0ds_logic.v(10478)
  not u11585 (Ht7ow6, n3153);  // ../RTL/cortexm0ds_logic.v(10478)
  and u11586 (At7ow6, Vt7ow6, Cu7ow6);  // ../RTL/cortexm0ds_logic.v(10479)
  and u11587 (n3154, Zzniu6, Ju7ow6);  // ../RTL/cortexm0ds_logic.v(10480)
  not u11588 (Cu7ow6, n3154);  // ../RTL/cortexm0ds_logic.v(10480)
  or u11589 (Ju7ow6, Qu7ow6, Ae0iu6);  // ../RTL/cortexm0ds_logic.v(10481)
  or u1159 (n51, Mdhpw6[0], Ighpw6[4]);  // ../RTL/cortexm0ds_logic.v(3261)
  and u11590 (n3155, U98iu6, Xu7ow6);  // ../RTL/cortexm0ds_logic.v(10482)
  not u11591 (Vt7ow6, n3155);  // ../RTL/cortexm0ds_logic.v(10482)
  or u11592 (Xu7ow6, Mo2ju6, Us2ju6);  // ../RTL/cortexm0ds_logic.v(10483)
  and u11593 (Ms7ow6, Ev7ow6, Lv7ow6);  // ../RTL/cortexm0ds_logic.v(10484)
  and u11594 (Ev7ow6, Sv7ow6, Zv7ow6);  // ../RTL/cortexm0ds_logic.v(10485)
  and u11595 (n3156, Uyiiu6, Gw7ow6);  // ../RTL/cortexm0ds_logic.v(10486)
  not u11596 (Zv7ow6, n3156);  // ../RTL/cortexm0ds_logic.v(10486)
  and u11597 (n3157, Nw7ow6, Uw7ow6);  // ../RTL/cortexm0ds_logic.v(10487)
  not u11598 (Gw7ow6, n3157);  // ../RTL/cortexm0ds_logic.v(10487)
  and u11599 (n3158, Bx7ow6, Dmiiu6);  // ../RTL/cortexm0ds_logic.v(10488)
  buf u116 (vis_r1_o[5], Jvppw6);  // ../RTL/cortexm0ds_logic.v(1876)
  not u1160 (M0zhu6, n51);  // ../RTL/cortexm0ds_logic.v(3261)
  not u11600 (Uw7ow6, n3158);  // ../RTL/cortexm0ds_logic.v(10488)
  and u11601 (Bx7ow6, Nbkiu6, Zraiu6);  // ../RTL/cortexm0ds_logic.v(10489)
  and u11602 (Nw7ow6, Ix7ow6, Px7ow6);  // ../RTL/cortexm0ds_logic.v(10490)
  and u11603 (n3159, Wx7ow6, Dy7ow6);  // ../RTL/cortexm0ds_logic.v(10491)
  not u11604 (Px7ow6, n3159);  // ../RTL/cortexm0ds_logic.v(10491)
  and u11605 (Dy7ow6, Ky7ow6, Ry7ow6);  // ../RTL/cortexm0ds_logic.v(10492)
  and u11606 (Ky7ow6, L88iu6, Dzjiu6);  // ../RTL/cortexm0ds_logic.v(10493)
  or u11607 (n3160, Ndiiu6, Gkiiu6);  // ../RTL/cortexm0ds_logic.v(10494)
  not u11608 (L88iu6, n3160);  // ../RTL/cortexm0ds_logic.v(10494)
  or u11609 (n3161, Kcziu6, U5jiu6);  // ../RTL/cortexm0ds_logic.v(10495)
  or u1161 (n52, T0zhu6, A1zhu6);  // ../RTL/cortexm0ds_logic.v(3262)
  not u11610 (Wx7ow6, n3161);  // ../RTL/cortexm0ds_logic.v(10495)
  and u11611 (n3162, Yy7ow6, Fz7ow6);  // ../RTL/cortexm0ds_logic.v(10496)
  not u11612 (Ix7ow6, n3162);  // ../RTL/cortexm0ds_logic.v(10496)
  and u11613 (Fz7ow6, Th2ju6, Ak0ju6);  // ../RTL/cortexm0ds_logic.v(10497)
  and u11614 (Yy7ow6, Cwiiu6, Aujiu6);  // ../RTL/cortexm0ds_logic.v(10498)
  and u11615 (n3163, Y0jiu6, Gwyiu6);  // ../RTL/cortexm0ds_logic.v(10499)
  not u11616 (Sv7ow6, n3163);  // ../RTL/cortexm0ds_logic.v(10499)
  and u11617 (n3164, Mz7ow6, Tz7ow6);  // ../RTL/cortexm0ds_logic.v(10500)
  not u11618 (Jn7ow6, n3164);  // ../RTL/cortexm0ds_logic.v(10500)
  and u11619 (Tz7ow6, A08ow6, H08ow6);  // ../RTL/cortexm0ds_logic.v(10501)
  not u1162 (I6yhu6, n52);  // ../RTL/cortexm0ds_logic.v(3262)
  or u11620 (H08ow6, R75iu6, I65iu6);  // ../RTL/cortexm0ds_logic.v(10502)
  not u11621 (I65iu6, S8fpw6[8]);  // ../RTL/cortexm0ds_logic.v(10503)
  and u11622 (A08ow6, O08ow6, V08ow6);  // ../RTL/cortexm0ds_logic.v(10504)
  and u11623 (n3165, L45iu6, C18ow6);  // ../RTL/cortexm0ds_logic.v(10505)
  not u11624 (V08ow6, n3165);  // ../RTL/cortexm0ds_logic.v(10505)
  and u11625 (n3166, J18ow6, Q18ow6);  // ../RTL/cortexm0ds_logic.v(10506)
  not u11626 (C18ow6, n3166);  // ../RTL/cortexm0ds_logic.v(10506)
  and u11627 (Q18ow6, X18ow6, E28ow6);  // ../RTL/cortexm0ds_logic.v(10507)
  or u11628 (E28ow6, L28ow6, Eoyiu6);  // ../RTL/cortexm0ds_logic.v(10508)
  and u11629 (n3167, Zoyiu6, G55iu6);  // ../RTL/cortexm0ds_logic.v(10509)
  buf u1163 (vis_r5_o[8], P21qw6);  // ../RTL/cortexm0ds_logic.v(1909)
  not u11630 (X18ow6, n3167);  // ../RTL/cortexm0ds_logic.v(10509)
  and u11631 (J18ow6, S28ow6, Z28ow6);  // ../RTL/cortexm0ds_logic.v(10510)
  or u11632 (Z28ow6, B65iu6, N55iu6);  // ../RTL/cortexm0ds_logic.v(10511)
  or u11633 (S28ow6, P65iu6, S8fpw6[8]);  // ../RTL/cortexm0ds_logic.v(10512)
  not u11634 (P65iu6, S8fpw6[9]);  // ../RTL/cortexm0ds_logic.v(10513)
  and u11635 (n3168, D7fpw6[3], K75iu6);  // ../RTL/cortexm0ds_logic.v(10514)
  not u11636 (O08ow6, n3168);  // ../RTL/cortexm0ds_logic.v(10514)
  and u11637 (n3169, Wiliu6, G38ow6);  // ../RTL/cortexm0ds_logic.v(10515)
  not u11638 (K75iu6, n3169);  // ../RTL/cortexm0ds_logic.v(10515)
  or u11639 (G38ow6, N38ow6, I6jiu6);  // ../RTL/cortexm0ds_logic.v(10516)
  buf u1164 (vis_r5_o[14], S58ax6);  // ../RTL/cortexm0ds_logic.v(1909)
  and u11640 (Mz7ow6, U38ow6, Gpyiu6);  // ../RTL/cortexm0ds_logic.v(10517)
  and u11641 (Gpyiu6, B48ow6, F85iu6);  // ../RTL/cortexm0ds_logic.v(10518)
  and u11642 (F85iu6, K0jiu6, Twniu6);  // ../RTL/cortexm0ds_logic.v(10519)
  or u11643 (K0jiu6, R2aiu6, Tr0iu6);  // ../RTL/cortexm0ds_logic.v(10520)
  or u11644 (n3170, N20ju6, Hzziu6);  // ../RTL/cortexm0ds_logic.v(10521)
  not u11645 (B48ow6, n3170);  // ../RTL/cortexm0ds_logic.v(10521)
  and u11646 (U38ow6, I48ow6, P48ow6);  // ../RTL/cortexm0ds_logic.v(10522)
  and u11647 (n3171, A95iu6, D7fpw6[0]);  // ../RTL/cortexm0ds_logic.v(10523)
  not u11648 (P48ow6, n3171);  // ../RTL/cortexm0ds_logic.v(10523)
  or u11649 (I48ow6, H95iu6, Ad8iu6);  // ../RTL/cortexm0ds_logic.v(10524)
  and u1165 (n53, U5yhu6, V1zhu6);  // ../RTL/cortexm0ds_logic.v(3264)
  and u11650 (n3172, W48ow6, D58ow6);  // ../RTL/cortexm0ds_logic.v(10525)
  not u11651 (Esohu6, n3172);  // ../RTL/cortexm0ds_logic.v(10525)
  and u11652 (D58ow6, K58ow6, R58ow6);  // ../RTL/cortexm0ds_logic.v(10526)
  and u11653 (n3173, Egziu6, Eafpw6[7]);  // ../RTL/cortexm0ds_logic.v(10527)
  not u11654 (R58ow6, n3173);  // ../RTL/cortexm0ds_logic.v(10527)
  and u11655 (K58ow6, Y58ow6, Sgziu6);  // ../RTL/cortexm0ds_logic.v(10528)
  and u11656 (n3174, Zgziu6, Qukiu6);  // ../RTL/cortexm0ds_logic.v(10529)
  not u11657 (Y58ow6, n3174);  // ../RTL/cortexm0ds_logic.v(10529)
  and u11658 (n3175, F68ow6, M68ow6);  // ../RTL/cortexm0ds_logic.v(10530)
  not u11659 (Qukiu6, n3175);  // ../RTL/cortexm0ds_logic.v(10530)
  not u1166 (O1zhu6, n53);  // ../RTL/cortexm0ds_logic.v(3264)
  and u11660 (M68ow6, T68ow6, A78ow6);  // ../RTL/cortexm0ds_logic.v(10531)
  or u11661 (A78ow6, Cfliu6, H78ow6);  // ../RTL/cortexm0ds_logic.v(10532)
  and u11662 (T68ow6, O78ow6, Mdliu6);  // ../RTL/cortexm0ds_logic.v(10533)
  and u11663 (n3176, Qfliu6, V78ow6);  // ../RTL/cortexm0ds_logic.v(10534)
  not u11664 (O78ow6, n3176);  // ../RTL/cortexm0ds_logic.v(10534)
  and u11665 (F68ow6, C88ow6, J88ow6);  // ../RTL/cortexm0ds_logic.v(10535)
  or u11666 (J88ow6, Ycliu6, Q88ow6);  // ../RTL/cortexm0ds_logic.v(10536)
  and u11667 (n3177, Aeliu6, X88ow6);  // ../RTL/cortexm0ds_logic.v(10537)
  not u11668 (C88ow6, n3177);  // ../RTL/cortexm0ds_logic.v(10537)
  and u11669 (W48ow6, E98ow6, L98ow6);  // ../RTL/cortexm0ds_logic.v(10538)
  and u1167 (n54, C2zhu6, J2zhu6);  // ../RTL/cortexm0ds_logic.v(3265)
  and u11670 (n3178, Zsfpw6[6], Cmziu6);  // ../RTL/cortexm0ds_logic.v(10539)
  not u11671 (L98ow6, n3178);  // ../RTL/cortexm0ds_logic.v(10539)
  and u11672 (n3179, vis_pc_o[6], Jmziu6);  // ../RTL/cortexm0ds_logic.v(10540)
  not u11673 (E98ow6, n3179);  // ../RTL/cortexm0ds_logic.v(10540)
  and u11674 (n3180, S98ow6, Z98ow6);  // ../RTL/cortexm0ds_logic.v(10541)
  not u11675 (Xrohu6, n3180);  // ../RTL/cortexm0ds_logic.v(10541)
  and u11676 (Z98ow6, Ga8ow6, Na8ow6);  // ../RTL/cortexm0ds_logic.v(10542)
  and u11677 (n3181, Egziu6, Eafpw6[31]);  // ../RTL/cortexm0ds_logic.v(10543)
  not u11678 (Na8ow6, n3181);  // ../RTL/cortexm0ds_logic.v(10543)
  and u11679 (Ga8ow6, Ua8ow6, Sgziu6);  // ../RTL/cortexm0ds_logic.v(10544)
  not u1168 (V1zhu6, n54);  // ../RTL/cortexm0ds_logic.v(3265)
  or u11680 (Ua8ow6, Ft6ow6, Ualiu6);  // ../RTL/cortexm0ds_logic.v(10545)
  and u11681 (Ualiu6, Bb8ow6, Ib8ow6);  // ../RTL/cortexm0ds_logic.v(10546)
  and u11682 (Ib8ow6, Pb8ow6, Wb8ow6);  // ../RTL/cortexm0ds_logic.v(10547)
  and u11683 (n3182, Dc8ow6, X88ow6);  // ../RTL/cortexm0ds_logic.v(10548)
  not u11684 (Wb8ow6, n3182);  // ../RTL/cortexm0ds_logic.v(10548)
  and u11685 (Pb8ow6, Kc8ow6, Djziu6);  // ../RTL/cortexm0ds_logic.v(10549)
  and u11686 (n3183, Rc8ow6, V78ow6);  // ../RTL/cortexm0ds_logic.v(10550)
  not u11687 (Kc8ow6, n3183);  // ../RTL/cortexm0ds_logic.v(10550)
  and u11688 (Bb8ow6, Yc8ow6, Fd8ow6);  // ../RTL/cortexm0ds_logic.v(10551)
  or u11689 (Fd8ow6, Mkziu6, Q88ow6);  // ../RTL/cortexm0ds_logic.v(10552)
  and u1169 (J2zhu6, Q2zhu6, X2zhu6);  // ../RTL/cortexm0ds_logic.v(3266)
  or u11690 (Yc8ow6, Hlziu6, H78ow6);  // ../RTL/cortexm0ds_logic.v(10553)
  and u11691 (S98ow6, Md8ow6, Td8ow6);  // ../RTL/cortexm0ds_logic.v(10554)
  and u11692 (n3184, Zsfpw6[30], Cmziu6);  // ../RTL/cortexm0ds_logic.v(10555)
  not u11693 (Td8ow6, n3184);  // ../RTL/cortexm0ds_logic.v(10555)
  and u11694 (n3185, vis_pc_o[30], Jmziu6);  // ../RTL/cortexm0ds_logic.v(10556)
  not u11695 (Md8ow6, n3185);  // ../RTL/cortexm0ds_logic.v(10556)
  or u11696 (Qrohu6, Ae8ow6, He8ow6);  // ../RTL/cortexm0ds_logic.v(10557)
  or u11697 (U7iow6, Oe8ow6, Cyfpw6[6]);  // ../RTL/cortexm0ds_logic.v(10558)
  not u11698 (He8ow6, U7iow6);  // ../RTL/cortexm0ds_logic.v(10558)
  AL_MUX u11699 (
    .i0(Cyfpw6[1]),
    .i1(Ve8ow6),
    .sel(HREADY),
    .o(Ae8ow6));  // ../RTL/cortexm0ds_logic.v(10559)
  buf u117 (Zbhpw6[26], Hpcbx6);  // ../RTL/cortexm0ds_logic.v(2147)
  and u1170 (n55, E3zhu6, Ighpw6[0]);  // ../RTL/cortexm0ds_logic.v(3267)
  and u11700 (n3186, Cf8ow6, Jf8ow6);  // ../RTL/cortexm0ds_logic.v(10560)
  not u11701 (Ve8ow6, n3186);  // ../RTL/cortexm0ds_logic.v(10560)
  and u11702 (Jf8ow6, Qf8ow6, Xf8ow6);  // ../RTL/cortexm0ds_logic.v(10561)
  and u11703 (Xf8ow6, Eg8ow6, Lg8ow6);  // ../RTL/cortexm0ds_logic.v(10562)
  and u11704 (n3187, Sg8ow6, Neoiu6);  // ../RTL/cortexm0ds_logic.v(10563)
  not u11705 (Lg8ow6, n3187);  // ../RTL/cortexm0ds_logic.v(10563)
  and u11706 (Sg8ow6, Zg8ow6, Mr0iu6);  // ../RTL/cortexm0ds_logic.v(10564)
  and u11707 (n3188, E4jiu6, Gh8ow6);  // ../RTL/cortexm0ds_logic.v(10565)
  not u11708 (Zg8ow6, n3188);  // ../RTL/cortexm0ds_logic.v(10565)
  and u11709 (n3189, Nh8ow6, Pthiu6);  // ../RTL/cortexm0ds_logic.v(10566)
  not u1171 (X2zhu6, n55);  // ../RTL/cortexm0ds_logic.v(3267)
  not u11710 (Gh8ow6, n3189);  // ../RTL/cortexm0ds_logic.v(10566)
  or u11711 (n3190, R75iu6, Cyfpw6[5]);  // ../RTL/cortexm0ds_logic.v(10567)
  not u11712 (Nh8ow6, n3190);  // ../RTL/cortexm0ds_logic.v(10567)
  and u11713 (n3191, Uh8ow6, Hiaiu6);  // ../RTL/cortexm0ds_logic.v(10568)
  not u11714 (Eg8ow6, n3191);  // ../RTL/cortexm0ds_logic.v(10568)
  and u11715 (Uh8ow6, Bi8ow6, Q5aiu6);  // ../RTL/cortexm0ds_logic.v(10569)
  and u11716 (n3192, Ii8ow6, Pi8ow6);  // ../RTL/cortexm0ds_logic.v(10570)
  not u11717 (Bi8ow6, n3192);  // ../RTL/cortexm0ds_logic.v(10570)
  and u11718 (Pi8ow6, Wi8ow6, Dj8ow6);  // ../RTL/cortexm0ds_logic.v(10571)
  and u11719 (n3193, J9kiu6, Kj8ow6);  // ../RTL/cortexm0ds_logic.v(10572)
  and u1172 (E3zhu6, L3zhu6, Eiyhu6);  // ../RTL/cortexm0ds_logic.v(3268)
  not u11720 (Dj8ow6, n3193);  // ../RTL/cortexm0ds_logic.v(10572)
  and u11721 (n3194, Rj8ow6, Yj8ow6);  // ../RTL/cortexm0ds_logic.v(10573)
  not u11722 (Kj8ow6, n3194);  // ../RTL/cortexm0ds_logic.v(10573)
  and u11723 (Yj8ow6, Fk8ow6, S01ju6);  // ../RTL/cortexm0ds_logic.v(10574)
  not u11724 (S01ju6, Fs7ow6);  // ../RTL/cortexm0ds_logic.v(10575)
  and u11725 (Fs7ow6, D7fpw6[11], I6jiu6);  // ../RTL/cortexm0ds_logic.v(10576)
  and u11726 (n3195, Mk8ow6, X1ziu6);  // ../RTL/cortexm0ds_logic.v(10577)
  not u11727 (Fk8ow6, n3195);  // ../RTL/cortexm0ds_logic.v(10577)
  or u11728 (Mk8ow6, Zwciu6, D7fpw6[8]);  // ../RTL/cortexm0ds_logic.v(10578)
  not u11729 (Zwciu6, Jehhu6);  // ../RTL/cortexm0ds_logic.v(10579)
  and u1173 (n56, S3zhu6, Z3zhu6);  // ../RTL/cortexm0ds_logic.v(3269)
  and u11730 (Rj8ow6, Tk8ow6, Al8ow6);  // ../RTL/cortexm0ds_logic.v(10580)
  or u11731 (Al8ow6, Hl8ow6, D7fpw6[11]);  // ../RTL/cortexm0ds_logic.v(10581)
  or u11732 (Tk8ow6, D7fpw6[13], D7fpw6[8]);  // ../RTL/cortexm0ds_logic.v(10582)
  and u11733 (Wi8ow6, Ol8ow6, Vl8ow6);  // ../RTL/cortexm0ds_logic.v(10583)
  and u11734 (n3196, Cm8ow6, Jm8ow6);  // ../RTL/cortexm0ds_logic.v(10584)
  not u11735 (Vl8ow6, n3196);  // ../RTL/cortexm0ds_logic.v(10584)
  or u11736 (n3197, I6jiu6, Jjhiu6);  // ../RTL/cortexm0ds_logic.v(10585)
  not u11737 (Jm8ow6, n3197);  // ../RTL/cortexm0ds_logic.v(10585)
  and u11738 (Cm8ow6, Y40ju6, Nyiiu6);  // ../RTL/cortexm0ds_logic.v(10586)
  and u11739 (Nyiiu6, D7fpw6[11], Ftjiu6);  // ../RTL/cortexm0ds_logic.v(10587)
  not u1174 (L3zhu6, n56);  // ../RTL/cortexm0ds_logic.v(3269)
  and u11740 (n3198, Qm8ow6, Evyiu6);  // ../RTL/cortexm0ds_logic.v(10588)
  not u11741 (Ol8ow6, n3198);  // ../RTL/cortexm0ds_logic.v(10588)
  buf u11742 (W4fhu6, Ozkbx6[14]);  // ../RTL/cortexm0ds_logic.v(3176)
  not u11743 (Qm8ow6, Dl6ow6);  // ../RTL/cortexm0ds_logic.v(10589)
  or u11744 (n3199, Xm8ow6, En8ow6);  // ../RTL/cortexm0ds_logic.v(10590)
  not u11745 (Ii8ow6, n3199);  // ../RTL/cortexm0ds_logic.v(10590)
  and u11746 (En8ow6, Ejiiu6, Dmiiu6);  // ../RTL/cortexm0ds_logic.v(10591)
  and u11747 (Dmiiu6, Jiiiu6, D7fpw6[14]);  // ../RTL/cortexm0ds_logic.v(10592)
  AL_MUX u11748 (
    .i0(Ln8ow6),
    .i1(Sn8ow6),
    .sel(S1ehu6),
    .o(Xm8ow6));  // ../RTL/cortexm0ds_logic.v(10593)
  and u11749 (n3200, Zn8ow6, Go8ow6);  // ../RTL/cortexm0ds_logic.v(10594)
  or u1175 (Z3zhu6, Y7yhu6, Mdhpw6[0]);  // ../RTL/cortexm0ds_logic.v(3270)
  not u11750 (Ln8ow6, n3200);  // ../RTL/cortexm0ds_logic.v(10594)
  or u11751 (Go8ow6, No8ow6, Lroiu6);  // ../RTL/cortexm0ds_logic.v(10595)
  not u11752 (Lroiu6, Ejiiu6);  // ../RTL/cortexm0ds_logic.v(10596)
  not u11753 (No8ow6, Il3ju6);  // ../RTL/cortexm0ds_logic.v(10597)
  and u11754 (Zn8ow6, Uo8ow6, Xs0ju6);  // ../RTL/cortexm0ds_logic.v(10598)
  or u11755 (Xs0ju6, Wiliu6, Co6ow6);  // ../RTL/cortexm0ds_logic.v(10599)
  not u11756 (Wiliu6, Mtjiu6);  // ../RTL/cortexm0ds_logic.v(10600)
  and u11757 (n3201, Bp8ow6, Mtjiu6);  // ../RTL/cortexm0ds_logic.v(10601)
  not u11758 (Uo8ow6, n3201);  // ../RTL/cortexm0ds_logic.v(10601)
  and u11759 (Bp8ow6, D7fpw6[14], Ip8ow6);  // ../RTL/cortexm0ds_logic.v(10602)
  or u1176 (S3zhu6, Ighpw6[1], Ighpw6[3]);  // ../RTL/cortexm0ds_logic.v(3271)
  and u11760 (n3202, Pp8ow6, Wp8ow6);  // ../RTL/cortexm0ds_logic.v(10603)
  not u11761 (Ip8ow6, n3202);  // ../RTL/cortexm0ds_logic.v(10603)
  AL_MUX u11762 (
    .i0(D7fpw6[9]),
    .i1(Dq8ow6),
    .sel(Aq1ju6),
    .o(Wp8ow6));  // ../RTL/cortexm0ds_logic.v(10604)
  and u11763 (n3203, D7fpw6[8], Ad8iu6);  // ../RTL/cortexm0ds_logic.v(10605)
  not u11764 (Aq1ju6, n3203);  // ../RTL/cortexm0ds_logic.v(10605)
  or u11765 (Dq8ow6, U5jiu6, O95iu6);  // ../RTL/cortexm0ds_logic.v(10606)
  and u11766 (Pp8ow6, Kq8ow6, Oviiu6);  // ../RTL/cortexm0ds_logic.v(10607)
  and u11767 (n3204, D7fpw6[8], Rq8ow6);  // ../RTL/cortexm0ds_logic.v(10608)
  not u11768 (Kq8ow6, n3204);  // ../RTL/cortexm0ds_logic.v(10608)
  and u11769 (n3205, Yq8ow6, Fr8ow6);  // ../RTL/cortexm0ds_logic.v(10609)
  and u1177 (Q2zhu6, G4zhu6, Joyhu6);  // ../RTL/cortexm0ds_logic.v(3272)
  not u11770 (Rq8ow6, n3205);  // ../RTL/cortexm0ds_logic.v(10609)
  or u11771 (Fr8ow6, I6jiu6, D7fpw6[7]);  // ../RTL/cortexm0ds_logic.v(10610)
  or u11772 (n3206, Db0ju6, Dcziu6);  // ../RTL/cortexm0ds_logic.v(10611)
  not u11773 (Yq8ow6, n3206);  // ../RTL/cortexm0ds_logic.v(10611)
  and u11774 (Qf8ow6, Mr8ow6, Tr8ow6);  // ../RTL/cortexm0ds_logic.v(10612)
  and u11775 (n3207, As8ow6, Hs8ow6);  // ../RTL/cortexm0ds_logic.v(10613)
  not u11776 (Tr8ow6, n3207);  // ../RTL/cortexm0ds_logic.v(10613)
  and u11777 (As8ow6, Frziu6, Hzziu6);  // ../RTL/cortexm0ds_logic.v(10614)
  and u11778 (n3208, Os8ow6, Geaiu6);  // ../RTL/cortexm0ds_logic.v(10615)
  not u11779 (Mr8ow6, n3208);  // ../RTL/cortexm0ds_logic.v(10615)
  and u1178 (n57, N4zhu6, U4zhu6);  // ../RTL/cortexm0ds_logic.v(3273)
  and u11780 (n3209, Vs8ow6, Ct8ow6);  // ../RTL/cortexm0ds_logic.v(10616)
  not u11781 (Os8ow6, n3209);  // ../RTL/cortexm0ds_logic.v(10616)
  and u11782 (n3210, Jt8ow6, Vs0iu6);  // ../RTL/cortexm0ds_logic.v(10617)
  not u11783 (Ct8ow6, n3210);  // ../RTL/cortexm0ds_logic.v(10617)
  and u11784 (Vs0iu6, F86ow6, Cyfpw6[0]);  // ../RTL/cortexm0ds_logic.v(10618)
  or u11785 (V58ju6, Knaiu6, Tfjiu6);  // ../RTL/cortexm0ds_logic.v(10619)
  not u11786 (F86ow6, V58ju6);  // ../RTL/cortexm0ds_logic.v(10619)
  and u11787 (Jt8ow6, Qe8iu6, Gwyiu6);  // ../RTL/cortexm0ds_logic.v(10620)
  and u11788 (n3211, Qt8ow6, D7fpw6[11]);  // ../RTL/cortexm0ds_logic.v(10621)
  not u11789 (Vs8ow6, n3211);  // ../RTL/cortexm0ds_logic.v(10621)
  not u1179 (G4zhu6, n57);  // ../RTL/cortexm0ds_logic.v(3273)
  and u11790 (Qt8ow6, Xt8ow6, Q5aiu6);  // ../RTL/cortexm0ds_logic.v(10622)
  or u11791 (Xt8ow6, Ry7ow6, Zakiu6);  // ../RTL/cortexm0ds_logic.v(10623)
  and u11792 (Zakiu6, Th2ju6, I6jiu6);  // ../RTL/cortexm0ds_logic.v(10624)
  and u11793 (Cf8ow6, Eu8ow6, Lu8ow6);  // ../RTL/cortexm0ds_logic.v(10626)
  and u11794 (Lu8ow6, Su8ow6, Zu8ow6);  // ../RTL/cortexm0ds_logic.v(10627)
  and u11795 (n3212, Gv8ow6, Zraiu6);  // ../RTL/cortexm0ds_logic.v(10628)
  not u11796 (Zu8ow6, n3212);  // ../RTL/cortexm0ds_logic.v(10628)
  and u11797 (n3213, Nv8ow6, Uv8ow6);  // ../RTL/cortexm0ds_logic.v(10629)
  not u11798 (Gv8ow6, n3213);  // ../RTL/cortexm0ds_logic.v(10629)
  and u11799 (Uv8ow6, Bw8ow6, Td0iu6);  // ../RTL/cortexm0ds_logic.v(10630)
  buf u118 (vis_r10_o[0], Cmlax6);  // ../RTL/cortexm0ds_logic.v(2469)
  and u1180 (N4zhu6, Hknhu6, B5zhu6);  // ../RTL/cortexm0ds_logic.v(3274)
  and u11800 (Bw8ow6, Re6ow6, Iw8ow6);  // ../RTL/cortexm0ds_logic.v(10631)
  and u11801 (n3214, Pw8ow6, Ww8ow6);  // ../RTL/cortexm0ds_logic.v(10632)
  not u11802 (Re6ow6, n3214);  // ../RTL/cortexm0ds_logic.v(10632)
  or u11803 (n3215, Iuniu6, Xmliu6);  // ../RTL/cortexm0ds_logic.v(10633)
  not u11804 (Pw8ow6, n3215);  // ../RTL/cortexm0ds_logic.v(10633)
  and u11805 (Nv8ow6, Dx8ow6, Kx8ow6);  // ../RTL/cortexm0ds_logic.v(10634)
  and u11806 (n3216, U0aiu6, Rx8ow6);  // ../RTL/cortexm0ds_logic.v(10635)
  not u11807 (Kx8ow6, n3216);  // ../RTL/cortexm0ds_logic.v(10635)
  or u11808 (Rx8ow6, Tfjiu6, X97ow6);  // ../RTL/cortexm0ds_logic.v(10636)
  and u11809 (n3217, S6aiu6, Yx8ow6);  // ../RTL/cortexm0ds_logic.v(10637)
  and u1181 (n58, Pyyhu6, I5zhu6);  // ../RTL/cortexm0ds_logic.v(3275)
  not u11810 (Dx8ow6, n3217);  // ../RTL/cortexm0ds_logic.v(10637)
  or u11811 (Yx8ow6, Geoiu6, Ly2ju6);  // ../RTL/cortexm0ds_logic.v(10638)
  and u11812 (Ly2ju6, Vo3ju6, Tr0iu6);  // ../RTL/cortexm0ds_logic.v(10639)
  and u11813 (Eu8ow6, Fy8ow6, My8ow6);  // ../RTL/cortexm0ds_logic.v(10640)
  or u11814 (My8ow6, Ty8ow6, Xe8iu6);  // ../RTL/cortexm0ds_logic.v(10641)
  AL_MUX u11815 (
    .i0(Az8ow6),
    .i1(Hz8ow6),
    .sel(Dxziu6),
    .o(Fy8ow6));  // ../RTL/cortexm0ds_logic.v(10642)
  and u11816 (n3218, Oz8ow6, Moaiu6);  // ../RTL/cortexm0ds_logic.v(10643)
  not u11817 (Hz8ow6, n3218);  // ../RTL/cortexm0ds_logic.v(10643)
  and u11818 (Oz8ow6, Toaiu6, Cyfpw6[7]);  // ../RTL/cortexm0ds_logic.v(10644)
  and u11819 (n3219, Vz8ow6, F9aju6);  // ../RTL/cortexm0ds_logic.v(10645)
  not u1182 (B5zhu6, n58);  // ../RTL/cortexm0ds_logic.v(3275)
  not u11820 (Az8ow6, n3219);  // ../RTL/cortexm0ds_logic.v(10645)
  and u11821 (Vz8ow6, Ls1ju6, Sq3ju6);  // ../RTL/cortexm0ds_logic.v(10646)
  and u11822 (Jrohu6, C09ow6, J09ow6);  // ../RTL/cortexm0ds_logic.v(10647)
  and u11823 (n3220, Q09ow6, X09ow6);  // ../RTL/cortexm0ds_logic.v(10648)
  not u11824 (J09ow6, n3220);  // ../RTL/cortexm0ds_logic.v(10648)
  and u11825 (X09ow6, E19ow6, L19ow6);  // ../RTL/cortexm0ds_logic.v(10649)
  and u11826 (L19ow6, S19ow6, Z19ow6);  // ../RTL/cortexm0ds_logic.v(10650)
  and u11827 (Z19ow6, G29ow6, Yryiu6);  // ../RTL/cortexm0ds_logic.v(10651)
  and u11828 (n3221, Ujjiu6, Bkjiu6);  // ../RTL/cortexm0ds_logic.v(10652)
  not u11829 (Yryiu6, n3221);  // ../RTL/cortexm0ds_logic.v(10652)
  or u1183 (I5zhu6, P5zhu6, R7yhu6);  // ../RTL/cortexm0ds_logic.v(3276)
  and u11830 (n3222, N29ow6, Cyfpw6[0]);  // ../RTL/cortexm0ds_logic.v(10653)
  not u11831 (G29ow6, n3222);  // ../RTL/cortexm0ds_logic.v(10653)
  and u11832 (N29ow6, U29ow6, B39ow6);  // ../RTL/cortexm0ds_logic.v(10654)
  and u11833 (n3223, I39ow6, R75iu6);  // ../RTL/cortexm0ds_logic.v(10655)
  not u11834 (B39ow6, n3223);  // ../RTL/cortexm0ds_logic.v(10655)
  and u11835 (n3224, P39ow6, Yljiu6);  // ../RTL/cortexm0ds_logic.v(10656)
  not u11836 (I39ow6, n3224);  // ../RTL/cortexm0ds_logic.v(10656)
  or u11837 (n3225, Hs0iu6, Dxziu6);  // ../RTL/cortexm0ds_logic.v(10657)
  not u11838 (P39ow6, n3225);  // ../RTL/cortexm0ds_logic.v(10657)
  or u11839 (U29ow6, Difiu6, Pugiu6);  // ../RTL/cortexm0ds_logic.v(10658)
  and u1184 (C2zhu6, W5zhu6, D6zhu6);  // ../RTL/cortexm0ds_logic.v(3277)
  and u11840 (Difiu6, Cyfpw6[6], Ii0iu6);  // ../RTL/cortexm0ds_logic.v(10659)
  and u11841 (S19ow6, W39ow6, D49ow6);  // ../RTL/cortexm0ds_logic.v(10660)
  and u11842 (n3226, K49ow6, T23ju6);  // ../RTL/cortexm0ds_logic.v(10661)
  not u11843 (D49ow6, n3226);  // ../RTL/cortexm0ds_logic.v(10661)
  or u11844 (n3227, C0ehu6, Cyfpw6[7]);  // ../RTL/cortexm0ds_logic.v(10662)
  not u11845 (K49ow6, n3227);  // ../RTL/cortexm0ds_logic.v(10662)
  and u11846 (n3228, R49ow6, W0piu6);  // ../RTL/cortexm0ds_logic.v(10663)
  not u11847 (W39ow6, n3228);  // ../RTL/cortexm0ds_logic.v(10663)
  and u11848 (R49ow6, D7fpw6[11], Y49ow6);  // ../RTL/cortexm0ds_logic.v(10664)
  and u11849 (n3229, C27ow6, F59ow6);  // ../RTL/cortexm0ds_logic.v(10665)
  AL_MUX u1185 (
    .i0(K6zhu6),
    .i1(R6zhu6),
    .sel(Mdhpw6[3]),
    .o(D6zhu6));  // ../RTL/cortexm0ds_logic.v(3278)
  not u11850 (Y49ow6, n3229);  // ../RTL/cortexm0ds_logic.v(10665)
  and u11851 (n3230, M59ow6, C0ehu6);  // ../RTL/cortexm0ds_logic.v(10666)
  not u11852 (F59ow6, n3230);  // ../RTL/cortexm0ds_logic.v(10666)
  or u11853 (n3231, X1ziu6, D7fpw6[10]);  // ../RTL/cortexm0ds_logic.v(10667)
  not u11854 (M59ow6, n3231);  // ../RTL/cortexm0ds_logic.v(10667)
  and u11855 (E19ow6, T59ow6, A69ow6);  // ../RTL/cortexm0ds_logic.v(10668)
  and u11856 (A69ow6, H69ow6, O69ow6);  // ../RTL/cortexm0ds_logic.v(10669)
  and u11857 (n3232, V69ow6, Hzziu6);  // ../RTL/cortexm0ds_logic.v(10670)
  not u11858 (O69ow6, n3232);  // ../RTL/cortexm0ds_logic.v(10670)
  or u11859 (n3233, Yp8iu6, Y7ghu6);  // ../RTL/cortexm0ds_logic.v(10671)
  and u1186 (R6zhu6, Mfyhu6, Y6zhu6);  // ../RTL/cortexm0ds_logic.v(3279)
  not u11860 (V69ow6, n3233);  // ../RTL/cortexm0ds_logic.v(10671)
  and u11861 (n3234, C79ow6, J79ow6);  // ../RTL/cortexm0ds_logic.v(10672)
  not u11862 (H69ow6, n3234);  // ../RTL/cortexm0ds_logic.v(10672)
  and u11863 (C79ow6, Yljiu6, Taaiu6);  // ../RTL/cortexm0ds_logic.v(10673)
  and u11864 (T59ow6, Q79ow6, X79ow6);  // ../RTL/cortexm0ds_logic.v(10674)
  and u11865 (n3235, Hwaiu6, A3aju6);  // ../RTL/cortexm0ds_logic.v(10675)
  not u11866 (X79ow6, n3235);  // ../RTL/cortexm0ds_logic.v(10675)
  or u11867 (n3236, R75iu6, Knaiu6);  // ../RTL/cortexm0ds_logic.v(10676)
  not u11868 (Hwaiu6, n3236);  // ../RTL/cortexm0ds_logic.v(10676)
  and u11869 (n3237, Dxziu6, E89ow6);  // ../RTL/cortexm0ds_logic.v(10677)
  and u1187 (n59, F7zhu6, Lbyhu6);  // ../RTL/cortexm0ds_logic.v(3280)
  not u11870 (Q79ow6, n3237);  // ../RTL/cortexm0ds_logic.v(10677)
  and u11871 (n3238, L89ow6, S89ow6);  // ../RTL/cortexm0ds_logic.v(10678)
  not u11872 (E89ow6, n3238);  // ../RTL/cortexm0ds_logic.v(10678)
  and u11873 (n3239, Z89ow6, X97ow6);  // ../RTL/cortexm0ds_logic.v(10679)
  not u11874 (S89ow6, n3239);  // ../RTL/cortexm0ds_logic.v(10679)
  and u11875 (Z89ow6, D1piu6, Tfjiu6);  // ../RTL/cortexm0ds_logic.v(10680)
  and u11876 (n3240, Jf6ju6, N3ziu6);  // ../RTL/cortexm0ds_logic.v(10681)
  not u11877 (L89ow6, n3240);  // ../RTL/cortexm0ds_logic.v(10681)
  and u11878 (Q09ow6, G99ow6, N99ow6);  // ../RTL/cortexm0ds_logic.v(10682)
  and u11879 (N99ow6, U99ow6, Ba9ow6);  // ../RTL/cortexm0ds_logic.v(10683)
  not u1188 (Y6zhu6, n59);  // ../RTL/cortexm0ds_logic.v(3280)
  and u11880 (Ba9ow6, Ia9ow6, Pa9ow6);  // ../RTL/cortexm0ds_logic.v(10684)
  and u11881 (n3241, Uyiiu6, Wa9ow6);  // ../RTL/cortexm0ds_logic.v(10685)
  not u11882 (Pa9ow6, n3241);  // ../RTL/cortexm0ds_logic.v(10685)
  and u11883 (n3242, Xl0ju6, Db9ow6);  // ../RTL/cortexm0ds_logic.v(10686)
  not u11884 (Wa9ow6, n3242);  // ../RTL/cortexm0ds_logic.v(10686)
  and u11885 (n3243, Kb9ow6, Ftjiu6);  // ../RTL/cortexm0ds_logic.v(10687)
  not u11886 (Db9ow6, n3243);  // ../RTL/cortexm0ds_logic.v(10687)
  and u11887 (n3244, Biliu6, Rb9ow6);  // ../RTL/cortexm0ds_logic.v(10688)
  not u11888 (Kb9ow6, n3244);  // ../RTL/cortexm0ds_logic.v(10688)
  or u11889 (Rb9ow6, Yb9ow6, I6jiu6);  // ../RTL/cortexm0ds_logic.v(10689)
  and u1189 (Lbyhu6, M7zhu6, T7zhu6);  // ../RTL/cortexm0ds_logic.v(3281)
  not u11890 (Biliu6, Sn8ow6);  // ../RTL/cortexm0ds_logic.v(10690)
  and u11891 (Sn8ow6, C0ehu6, X1ziu6);  // ../RTL/cortexm0ds_logic.v(10691)
  or u11892 (Ia9ow6, Thaiu6, Cyfpw6[5]);  // ../RTL/cortexm0ds_logic.v(10692)
  and u11893 (U99ow6, Fc9ow6, Mc9ow6);  // ../RTL/cortexm0ds_logic.v(10693)
  and u11894 (n3245, De6ow6, Vxniu6);  // ../RTL/cortexm0ds_logic.v(10694)
  not u11895 (Mc9ow6, n3245);  // ../RTL/cortexm0ds_logic.v(10694)
  or u11896 (Fc9ow6, Iw8ow6, Ae0iu6);  // ../RTL/cortexm0ds_logic.v(10695)
  and u11897 (G99ow6, Tc9ow6, Ad9ow6);  // ../RTL/cortexm0ds_logic.v(10696)
  and u11898 (Ad9ow6, Hd9ow6, Od9ow6);  // ../RTL/cortexm0ds_logic.v(10697)
  and u11899 (n3246, S6aiu6, Vd9ow6);  // ../RTL/cortexm0ds_logic.v(10698)
  buf u119 (K7hpw6[29], Wahbx6);  // ../RTL/cortexm0ds_logic.v(2366)
  and u1190 (F7zhu6, Mdhpw6[2], A8zhu6);  // ../RTL/cortexm0ds_logic.v(3282)
  not u11900 (Od9ow6, n3246);  // ../RTL/cortexm0ds_logic.v(10698)
  and u11901 (n3247, Ce9ow6, Je9ow6);  // ../RTL/cortexm0ds_logic.v(10699)
  not u11902 (Vd9ow6, n3247);  // ../RTL/cortexm0ds_logic.v(10699)
  AL_MUX u11903 (
    .i0(Cyfpw6[1]),
    .i1(Ey2ju6),
    .sel(Nlaiu6),
    .o(Je9ow6));  // ../RTL/cortexm0ds_logic.v(10700)
  or u11904 (n3248, Qe9ow6, Ep6ow6);  // ../RTL/cortexm0ds_logic.v(10701)
  not u11905 (Ce9ow6, n3248);  // ../RTL/cortexm0ds_logic.v(10701)
  or u11906 (n3249, Lkaiu6, Eoyiu6);  // ../RTL/cortexm0ds_logic.v(10702)
  not u11907 (Qe9ow6, n3249);  // ../RTL/cortexm0ds_logic.v(10702)
  or u11908 (Hd9ow6, Xe9ow6, Wxyiu6);  // ../RTL/cortexm0ds_logic.v(10703)
  and u11909 (Wxyiu6, L62ju6, Zraiu6);  // ../RTL/cortexm0ds_logic.v(10704)
  and u1191 (n60, H8zhu6, Mdhpw6[0]);  // ../RTL/cortexm0ds_logic.v(3283)
  and u11910 (Tc9ow6, T41ju6, Ef9ow6);  // ../RTL/cortexm0ds_logic.v(10706)
  and u11911 (n3250, Lf9ow6, Q5aiu6);  // ../RTL/cortexm0ds_logic.v(10707)
  not u11912 (Ef9ow6, n3250);  // ../RTL/cortexm0ds_logic.v(10707)
  and u11913 (n3251, Sf9ow6, Zf9ow6);  // ../RTL/cortexm0ds_logic.v(10708)
  not u11914 (Lf9ow6, n3251);  // ../RTL/cortexm0ds_logic.v(10708)
  and u11915 (Zf9ow6, Gg9ow6, Ng9ow6);  // ../RTL/cortexm0ds_logic.v(10709)
  and u11916 (n3252, Ug9ow6, Vboiu6);  // ../RTL/cortexm0ds_logic.v(10710)
  not u11917 (Ng9ow6, n3252);  // ../RTL/cortexm0ds_logic.v(10710)
  or u11918 (n3253, R75iu6, H4ghu6);  // ../RTL/cortexm0ds_logic.v(10711)
  not u11919 (Ug9ow6, n3253);  // ../RTL/cortexm0ds_logic.v(10711)
  not u1192 (A8zhu6, n60);  // ../RTL/cortexm0ds_logic.v(3283)
  and u11920 (Gg9ow6, Bh9ow6, Ih9ow6);  // ../RTL/cortexm0ds_logic.v(10712)
  and u11921 (n3254, Ph9ow6, P0piu6);  // ../RTL/cortexm0ds_logic.v(10713)
  not u11922 (Ih9ow6, n3254);  // ../RTL/cortexm0ds_logic.v(10713)
  and u11923 (Ph9ow6, Wh9ow6, Ftjiu6);  // ../RTL/cortexm0ds_logic.v(10714)
  or u11924 (Wh9ow6, Di9ow6, Ki9ow6);  // ../RTL/cortexm0ds_logic.v(10715)
  AL_MUX u11925 (
    .i0(Ad8iu6),
    .i1(Dcziu6),
    .sel(Tniiu6),
    .o(Ki9ow6));  // ../RTL/cortexm0ds_logic.v(10716)
  and u11926 (n3255, Ri9ow6, Ar0ju6);  // ../RTL/cortexm0ds_logic.v(10717)
  not u11927 (Di9ow6, n3255);  // ../RTL/cortexm0ds_logic.v(10717)
  not u11928 (Ar0ju6, Jz0ju6);  // ../RTL/cortexm0ds_logic.v(10718)
  or u11929 (Ri9ow6, Ndiiu6, O95iu6);  // ../RTL/cortexm0ds_logic.v(10719)
  or u1193 (n61, O8zhu6, Ulnhu6);  // ../RTL/cortexm0ds_logic.v(3284)
  and u11930 (n3256, Yi9ow6, Db0ju6);  // ../RTL/cortexm0ds_logic.v(10720)
  not u11931 (Bh9ow6, n3256);  // ../RTL/cortexm0ds_logic.v(10720)
  or u11932 (n3257, H95iu6, X1ziu6);  // ../RTL/cortexm0ds_logic.v(10721)
  not u11933 (Yi9ow6, n3257);  // ../RTL/cortexm0ds_logic.v(10721)
  not u11934 (H95iu6, Ozziu6);  // ../RTL/cortexm0ds_logic.v(10722)
  and u11935 (Sf9ow6, Fj9ow6, Mj9ow6);  // ../RTL/cortexm0ds_logic.v(10723)
  and u11936 (n3258, Xiiiu6, Tj9ow6);  // ../RTL/cortexm0ds_logic.v(10724)
  not u11937 (Mj9ow6, n3258);  // ../RTL/cortexm0ds_logic.v(10724)
  and u11938 (n3259, Ak9ow6, Hk9ow6);  // ../RTL/cortexm0ds_logic.v(10725)
  not u11939 (Tj9ow6, n3259);  // ../RTL/cortexm0ds_logic.v(10725)
  not u1194 (H8zhu6, n61);  // ../RTL/cortexm0ds_logic.v(3284)
  and u11940 (n3260, Aujiu6, U5jiu6);  // ../RTL/cortexm0ds_logic.v(10726)
  not u11941 (Hk9ow6, n3260);  // ../RTL/cortexm0ds_logic.v(10726)
  not u11942 (U5jiu6, Jwiiu6);  // ../RTL/cortexm0ds_logic.v(10727)
  or u11943 (n3261, Ok9ow6, Vk9ow6);  // ../RTL/cortexm0ds_logic.v(10728)
  not u11944 (Ak9ow6, n3261);  // ../RTL/cortexm0ds_logic.v(10728)
  and u11945 (Ok9ow6, Y40ju6, Cl9ow6);  // ../RTL/cortexm0ds_logic.v(10729)
  and u11946 (n3262, Jl9ow6, Ql9ow6);  // ../RTL/cortexm0ds_logic.v(10730)
  not u11947 (Cl9ow6, n3262);  // ../RTL/cortexm0ds_logic.v(10730)
  or u11948 (Ql9ow6, Oviiu6, D7fpw6[6]);  // ../RTL/cortexm0ds_logic.v(10731)
  or u11949 (n3263, Dcziu6, D7fpw6[8]);  // ../RTL/cortexm0ds_logic.v(10732)
  and u1195 (n62, V8zhu6, Epyhu6);  // ../RTL/cortexm0ds_logic.v(3285)
  not u11950 (Jl9ow6, n3263);  // ../RTL/cortexm0ds_logic.v(10732)
  and u11951 (Fj9ow6, Xl9ow6, Em9ow6);  // ../RTL/cortexm0ds_logic.v(10733)
  and u11952 (n3264, Hl8ow6, Lm9ow6);  // ../RTL/cortexm0ds_logic.v(10734)
  not u11953 (Em9ow6, n3264);  // ../RTL/cortexm0ds_logic.v(10734)
  and u11954 (n3265, S80ju6, Sm9ow6);  // ../RTL/cortexm0ds_logic.v(10735)
  not u11955 (Lm9ow6, n3265);  // ../RTL/cortexm0ds_logic.v(10735)
  and u11956 (n3266, J9kiu6, Zm9ow6);  // ../RTL/cortexm0ds_logic.v(10736)
  not u11957 (Sm9ow6, n3266);  // ../RTL/cortexm0ds_logic.v(10736)
  and u11958 (n3267, Gn9ow6, Nn9ow6);  // ../RTL/cortexm0ds_logic.v(10737)
  not u11959 (Zm9ow6, n3267);  // ../RTL/cortexm0ds_logic.v(10737)
  not u1196 (Mfyhu6, n62);  // ../RTL/cortexm0ds_logic.v(3285)
  and u11960 (Nn9ow6, Un9ow6, I6jiu6);  // ../RTL/cortexm0ds_logic.v(10738)
  buf u11961 (K6fhu6, Ozkbx6[13]);  // ../RTL/cortexm0ds_logic.v(3176)
  or u11962 (n3268, O95iu6, Dzjiu6);  // ../RTL/cortexm0ds_logic.v(10740)
  not u11963 (Gn9ow6, n3268);  // ../RTL/cortexm0ds_logic.v(10740)
  and u11964 (n3269, C0ehu6, Bo9ow6);  // ../RTL/cortexm0ds_logic.v(10741)
  not u11965 (Xl9ow6, n3269);  // ../RTL/cortexm0ds_logic.v(10741)
  and u11966 (n3270, Io9ow6, Po9ow6);  // ../RTL/cortexm0ds_logic.v(10742)
  not u11967 (Bo9ow6, n3270);  // ../RTL/cortexm0ds_logic.v(10742)
  and u11968 (n3271, Wo9ow6, Aujiu6);  // ../RTL/cortexm0ds_logic.v(10743)
  not u11969 (Po9ow6, n3271);  // ../RTL/cortexm0ds_logic.v(10743)
  or u1197 (n63, C9zhu6, Ighpw6[2]);  // ../RTL/cortexm0ds_logic.v(3286)
  or u11970 (n3272, X1ziu6, D7fpw6[8]);  // ../RTL/cortexm0ds_logic.v(10744)
  not u11971 (Wo9ow6, n3272);  // ../RTL/cortexm0ds_logic.v(10744)
  and u11972 (Io9ow6, Dp9ow6, Uriiu6);  // ../RTL/cortexm0ds_logic.v(10745)
  and u11973 (n3273, Kp9ow6, Y40ju6);  // ../RTL/cortexm0ds_logic.v(10746)
  not u11974 (Dp9ow6, n3273);  // ../RTL/cortexm0ds_logic.v(10746)
  or u11975 (n3274, Jwiiu6, D7fpw6[15]);  // ../RTL/cortexm0ds_logic.v(10747)
  not u11976 (Kp9ow6, n3274);  // ../RTL/cortexm0ds_logic.v(10747)
  and u11977 (T41ju6, Rp9ow6, Yp9ow6);  // ../RTL/cortexm0ds_logic.v(10748)
  and u11978 (Yp9ow6, Fq9ow6, B1aiu6);  // ../RTL/cortexm0ds_logic.v(10749)
  and u11979 (n3275, Mq9ow6, Cyfpw6[4]);  // ../RTL/cortexm0ds_logic.v(10750)
  not u1198 (V8zhu6, n63);  // ../RTL/cortexm0ds_logic.v(3286)
  not u11980 (Fq9ow6, n3275);  // ../RTL/cortexm0ds_logic.v(10750)
  or u11981 (n3276, Geaiu6, Cyfpw6[5]);  // ../RTL/cortexm0ds_logic.v(10751)
  not u11982 (Mq9ow6, n3276);  // ../RTL/cortexm0ds_logic.v(10751)
  and u11983 (Rp9ow6, HREADY, Tq9ow6);  // ../RTL/cortexm0ds_logic.v(10752)
  or u11984 (C09ow6, Cyfpw6[0], HREADY);  // ../RTL/cortexm0ds_logic.v(10753)
  and u11985 (Crohu6, Ar9ow6, Hr9ow6);  // ../RTL/cortexm0ds_logic.v(10754)
  and u11986 (n3277, Or9ow6, Vr9ow6);  // ../RTL/cortexm0ds_logic.v(10755)
  not u11987 (Hr9ow6, n3277);  // ../RTL/cortexm0ds_logic.v(10755)
  and u11988 (Vr9ow6, Cs9ow6, Js9ow6);  // ../RTL/cortexm0ds_logic.v(10756)
  and u11989 (Js9ow6, Qs9ow6, Xs9ow6);  // ../RTL/cortexm0ds_logic.v(10757)
  and u1199 (K6zhu6, Pryhu6, Tfyhu6);  // ../RTL/cortexm0ds_logic.v(3287)
  and u11990 (Xs9ow6, Et9ow6, A42ju6);  // ../RTL/cortexm0ds_logic.v(10758)
  and u11991 (n3278, Lt9ow6, Htyiu6);  // ../RTL/cortexm0ds_logic.v(10759)
  not u11992 (A42ju6, n3278);  // ../RTL/cortexm0ds_logic.v(10759)
  and u11993 (Lt9ow6, Th2ju6, St9ow6);  // ../RTL/cortexm0ds_logic.v(10760)
  and u11994 (n3279, D7fpw6[12], Zt9ow6);  // ../RTL/cortexm0ds_logic.v(10761)
  not u11995 (St9ow6, n3279);  // ../RTL/cortexm0ds_logic.v(10761)
  or u11996 (n3280, Ujjiu6, Ot7ow6);  // ../RTL/cortexm0ds_logic.v(10762)
  not u11997 (Et9ow6, n3280);  // ../RTL/cortexm0ds_logic.v(10762)
  and u11998 (Ot7ow6, Gu9ow6, Nu9ow6);  // ../RTL/cortexm0ds_logic.v(10763)
  or u11999 (n3281, Jcaiu6, Cyfpw6[0]);  // ../RTL/cortexm0ds_logic.v(10764)
  buf u12 (WAKEUP, 1'b0);  // ../RTL/cortexm0ds_logic.v(1768)
  buf u120 (R4gpw6[62], Aw4bx6);  // ../RTL/cortexm0ds_logic.v(2815)
  and u1200 (W5zhu6, J9zhu6, Q9zhu6);  // ../RTL/cortexm0ds_logic.v(3288)
  not u12000 (Gu9ow6, n3281);  // ../RTL/cortexm0ds_logic.v(10764)
  and u12001 (Ujjiu6, Uu9ow6, D7fpw6[15]);  // ../RTL/cortexm0ds_logic.v(10765)
  and u12002 (Qs9ow6, Bv9ow6, Iv9ow6);  // ../RTL/cortexm0ds_logic.v(10766)
  and u12003 (n3282, Pv9ow6, Wv9ow6);  // ../RTL/cortexm0ds_logic.v(10767)
  not u12004 (Iv9ow6, n3282);  // ../RTL/cortexm0ds_logic.v(10767)
  and u12005 (Wv9ow6, D7fpw6[11], Dw9ow6);  // ../RTL/cortexm0ds_logic.v(10768)
  or u12006 (Dw9ow6, Gkiiu6, Fp1ju6);  // ../RTL/cortexm0ds_logic.v(10769)
  buf u12007 (Y7fhu6, Ozkbx6[12]);  // ../RTL/cortexm0ds_logic.v(3176)
  and u12008 (n3283, Kw9ow6, Rw9ow6);  // ../RTL/cortexm0ds_logic.v(10771)
  not u12009 (Bv9ow6, n3283);  // ../RTL/cortexm0ds_logic.v(10771)
  and u1201 (n64, X9zhu6, R7yhu6);  // ../RTL/cortexm0ds_logic.v(3289)
  or u12010 (n3284, D7fpw6[5], D7fpw6[7]);  // ../RTL/cortexm0ds_logic.v(10772)
  not u12011 (Rw9ow6, n3284);  // ../RTL/cortexm0ds_logic.v(10772)
  or u12012 (n3285, P82ju6, Yw9ow6);  // ../RTL/cortexm0ds_logic.v(10773)
  not u12013 (Kw9ow6, n3285);  // ../RTL/cortexm0ds_logic.v(10773)
  and u12014 (Yw9ow6, D7fpw6[4], D7fpw6[6]);  // ../RTL/cortexm0ds_logic.v(10774)
  and u12015 (Cs9ow6, Fx9ow6, Mx9ow6);  // ../RTL/cortexm0ds_logic.v(10775)
  and u12016 (Mx9ow6, Tx9ow6, Ay9ow6);  // ../RTL/cortexm0ds_logic.v(10776)
  and u12017 (n3286, Hy9ow6, Vviiu6);  // ../RTL/cortexm0ds_logic.v(10777)
  not u12018 (Ay9ow6, n3286);  // ../RTL/cortexm0ds_logic.v(10777)
  and u12019 (Hy9ow6, Hiaiu6, Oy9ow6);  // ../RTL/cortexm0ds_logic.v(10778)
  not u1202 (Q9zhu6, n64);  // ../RTL/cortexm0ds_logic.v(3289)
  and u12020 (n3287, Vy9ow6, Cz9ow6);  // ../RTL/cortexm0ds_logic.v(10779)
  not u12021 (Oy9ow6, n3287);  // ../RTL/cortexm0ds_logic.v(10779)
  or u12022 (Cz9ow6, Jz9ow6, Gaziu6);  // ../RTL/cortexm0ds_logic.v(10780)
  or u12023 (Vy9ow6, X1ziu6, Gkiiu6);  // ../RTL/cortexm0ds_logic.v(10781)
  and u12024 (n3288, Qz9ow6, Htyiu6);  // ../RTL/cortexm0ds_logic.v(10782)
  not u12025 (Tx9ow6, n3288);  // ../RTL/cortexm0ds_logic.v(10782)
  and u12026 (Qz9ow6, Xz9ow6, Zraiu6);  // ../RTL/cortexm0ds_logic.v(10783)
  and u12027 (n3289, E0aow6, L0aow6);  // ../RTL/cortexm0ds_logic.v(10784)
  not u12028 (Xz9ow6, n3289);  // ../RTL/cortexm0ds_logic.v(10784)
  and u12029 (n3290, X8ziu6, A95iu6);  // ../RTL/cortexm0ds_logic.v(10785)
  and u1203 (H1zhu6, Eazhu6, Rlyhu6);  // ../RTL/cortexm0ds_logic.v(3290)
  not u12030 (L0aow6, n3290);  // ../RTL/cortexm0ds_logic.v(10785)
  or u12031 (n3291, D7fpw6[11], D7fpw6[8]);  // ../RTL/cortexm0ds_logic.v(10786)
  not u12032 (X8ziu6, n3291);  // ../RTL/cortexm0ds_logic.v(10786)
  or u12033 (E0aow6, S80ju6, Gaziu6);  // ../RTL/cortexm0ds_logic.v(10787)
  and u12034 (Fx9ow6, S0aow6, Z0aow6);  // ../RTL/cortexm0ds_logic.v(10788)
  and u12035 (n3292, G1aow6, K2aiu6);  // ../RTL/cortexm0ds_logic.v(10789)
  not u12036 (Z0aow6, n3292);  // ../RTL/cortexm0ds_logic.v(10789)
  and u12037 (G1aow6, N1aow6, Y2oiu6);  // ../RTL/cortexm0ds_logic.v(10790)
  and u12038 (n3293, U1aow6, Neoiu6);  // ../RTL/cortexm0ds_logic.v(10791)
  not u12039 (S0aow6, n3293);  // ../RTL/cortexm0ds_logic.v(10791)
  and u1204 (n65, O9yhu6, Cayhu6);  // ../RTL/cortexm0ds_logic.v(3291)
  and u12040 (U1aow6, Omyiu6, B2aow6);  // ../RTL/cortexm0ds_logic.v(10792)
  and u12041 (n3294, I2aow6, P2aow6);  // ../RTL/cortexm0ds_logic.v(10793)
  not u12042 (B2aow6, n3294);  // ../RTL/cortexm0ds_logic.v(10793)
  or u12043 (P2aow6, Vwaiu6, Mr0iu6);  // ../RTL/cortexm0ds_logic.v(10794)
  or u12044 (n3295, G47ow6, W2aow6);  // ../RTL/cortexm0ds_logic.v(10795)
  not u12045 (I2aow6, n3295);  // ../RTL/cortexm0ds_logic.v(10795)
  and u12046 (Or9ow6, D3aow6, K3aow6);  // ../RTL/cortexm0ds_logic.v(10796)
  and u12047 (K3aow6, R3aow6, Y3aow6);  // ../RTL/cortexm0ds_logic.v(10797)
  and u12048 (Y3aow6, F4aow6, M4aow6);  // ../RTL/cortexm0ds_logic.v(10798)
  or u12049 (M4aow6, Tdziu6, Qpaju6);  // ../RTL/cortexm0ds_logic.v(10799)
  not u1205 (Rlyhu6, n65);  // ../RTL/cortexm0ds_logic.v(3291)
  and u12050 (n3296, Q97ow6, T4aow6);  // ../RTL/cortexm0ds_logic.v(10800)
  not u12051 (Tdziu6, n3296);  // ../RTL/cortexm0ds_logic.v(10800)
  or u12052 (n3297, E4jiu6, Cyfpw6[0]);  // ../RTL/cortexm0ds_logic.v(10801)
  not u12053 (Q97ow6, n3297);  // ../RTL/cortexm0ds_logic.v(10801)
  and u12054 (F4aow6, A5aow6, H5aow6);  // ../RTL/cortexm0ds_logic.v(10802)
  and u12055 (n3298, O5aow6, Yo1ju6);  // ../RTL/cortexm0ds_logic.v(10803)
  not u12056 (H5aow6, n3298);  // ../RTL/cortexm0ds_logic.v(10803)
  and u12057 (O5aow6, D7fpw6[14], V5aow6);  // ../RTL/cortexm0ds_logic.v(10804)
  or u12058 (V5aow6, C6aow6, J6aow6);  // ../RTL/cortexm0ds_logic.v(10805)
  AL_MUX u12059 (
    .i0(Q6aow6),
    .i1(X6aow6),
    .sel(D7fpw6[7]),
    .o(J6aow6));  // ../RTL/cortexm0ds_logic.v(10806)
  and u1206 (n66, T8yhu6, Lazhu6);  // ../RTL/cortexm0ds_logic.v(3292)
  or u12060 (n3299, Jz0ju6, D7fpw6[10]);  // ../RTL/cortexm0ds_logic.v(10807)
  not u12061 (X6aow6, n3299);  // ../RTL/cortexm0ds_logic.v(10807)
  and u12062 (Jz0ju6, Ad8iu6, Ndiiu6);  // ../RTL/cortexm0ds_logic.v(10808)
  and u12063 (n3300, E7aow6, Hk0ju6);  // ../RTL/cortexm0ds_logic.v(10809)
  not u12064 (C6aow6, n3300);  // ../RTL/cortexm0ds_logic.v(10809)
  not u12065 (Hk0ju6, Fp1ju6);  // ../RTL/cortexm0ds_logic.v(10810)
  and u12066 (Fp1ju6, I6jiu6, Tniiu6);  // ../RTL/cortexm0ds_logic.v(10811)
  or u12067 (E7aow6, L7aow6, D7fpw6[9]);  // ../RTL/cortexm0ds_logic.v(10812)
  and u12068 (n3301, Pthiu6, S7aow6);  // ../RTL/cortexm0ds_logic.v(10813)
  not u12069 (A5aow6, n3301);  // ../RTL/cortexm0ds_logic.v(10813)
  not u1207 (Eazhu6, n66);  // ../RTL/cortexm0ds_logic.v(3292)
  and u12070 (n3302, Z7aow6, G8aow6);  // ../RTL/cortexm0ds_logic.v(10814)
  not u12071 (S7aow6, n3302);  // ../RTL/cortexm0ds_logic.v(10814)
  or u12072 (G8aow6, Jojiu6, Y2oiu6);  // ../RTL/cortexm0ds_logic.v(10815)
  and u12073 (n3303, Ls1ju6, Cyfpw6[5]);  // ../RTL/cortexm0ds_logic.v(10816)
  not u12074 (Z7aow6, n3303);  // ../RTL/cortexm0ds_logic.v(10816)
  and u12075 (R3aow6, N8aow6, U8aow6);  // ../RTL/cortexm0ds_logic.v(10817)
  and u12076 (n3304, B9aow6, Geaiu6);  // ../RTL/cortexm0ds_logic.v(10818)
  not u12077 (U8aow6, n3304);  // ../RTL/cortexm0ds_logic.v(10818)
  and u12078 (n3305, I9aow6, P9aow6);  // ../RTL/cortexm0ds_logic.v(10819)
  not u12079 (B9aow6, n3305);  // ../RTL/cortexm0ds_logic.v(10819)
  and u1208 (n67, Deyhu6, Sazhu6);  // ../RTL/cortexm0ds_logic.v(3293)
  or u12080 (P9aow6, R2aiu6, Y2oiu6);  // ../RTL/cortexm0ds_logic.v(10820)
  and u12081 (I9aow6, W9aow6, Daaow6);  // ../RTL/cortexm0ds_logic.v(10821)
  and u12082 (n3306, Kaaow6, Raaow6);  // ../RTL/cortexm0ds_logic.v(10822)
  not u12083 (Daaow6, n3306);  // ../RTL/cortexm0ds_logic.v(10822)
  and u12084 (Kaaow6, M7kiu6, X1ziu6);  // ../RTL/cortexm0ds_logic.v(10823)
  and u12085 (M7kiu6, Yaaow6, Ozziu6);  // ../RTL/cortexm0ds_logic.v(10824)
  or u12086 (n3307, Ae0iu6, D7fpw6[15]);  // ../RTL/cortexm0ds_logic.v(10825)
  not u12087 (Yaaow6, n3307);  // ../RTL/cortexm0ds_logic.v(10825)
  or u12088 (W9aow6, Jxoiu6, Ak0ju6);  // ../RTL/cortexm0ds_logic.v(10826)
  and u12089 (Ak0ju6, Qxoiu6, Ndiiu6);  // ../RTL/cortexm0ds_logic.v(10827)
  not u1209 (Lazhu6, n67);  // ../RTL/cortexm0ds_logic.v(3293)
  and u12090 (n3308, Fbaow6, R7jiu6);  // ../RTL/cortexm0ds_logic.v(10828)
  not u12091 (Jxoiu6, n3308);  // ../RTL/cortexm0ds_logic.v(10828)
  and u12092 (Fbaow6, Ia8iu6, Q5aiu6);  // ../RTL/cortexm0ds_logic.v(10829)
  and u12093 (n3309, Dxziu6, Mbaow6);  // ../RTL/cortexm0ds_logic.v(10830)
  not u12094 (N8aow6, n3309);  // ../RTL/cortexm0ds_logic.v(10830)
  and u12095 (n3310, Tbaow6, Acaow6);  // ../RTL/cortexm0ds_logic.v(10831)
  not u12096 (Mbaow6, n3310);  // ../RTL/cortexm0ds_logic.v(10831)
  and u12097 (n3311, Ls1ju6, Hcaow6);  // ../RTL/cortexm0ds_logic.v(10832)
  not u12098 (Acaow6, n3311);  // ../RTL/cortexm0ds_logic.v(10832)
  or u12099 (Hcaow6, Rljiu6, Ocaow6);  // ../RTL/cortexm0ds_logic.v(10833)
  buf u121 (vis_r5_o[23], Gt6ax6);  // ../RTL/cortexm0ds_logic.v(1909)
  or u1210 (Sazhu6, Zazhu6, Ighpw6[1]);  // ../RTL/cortexm0ds_logic.v(3294)
  or u12100 (n3312, Qjaiu6, Cyfpw6[0]);  // ../RTL/cortexm0ds_logic.v(10834)
  not u12101 (Ocaow6, n3312);  // ../RTL/cortexm0ds_logic.v(10834)
  and u12102 (Tbaow6, Vcaow6, Cdaow6);  // ../RTL/cortexm0ds_logic.v(10835)
  and u12103 (n3313, Jdaow6, Qdaow6);  // ../RTL/cortexm0ds_logic.v(10836)
  not u12104 (Cdaow6, n3313);  // ../RTL/cortexm0ds_logic.v(10836)
  buf u12105 (M9fhu6, Ozkbx6[11]);  // ../RTL/cortexm0ds_logic.v(3176)
  and u12106 (Jdaow6, Eoyiu6, Geoiu6);  // ../RTL/cortexm0ds_logic.v(10838)
  and u12107 (Geoiu6, Wp0iu6, Ii0iu6);  // ../RTL/cortexm0ds_logic.v(10839)
  or u12108 (n3314, L28ow6, S8fpw6[7]);  // ../RTL/cortexm0ds_logic.v(10840)
  not u12109 (Eoyiu6, n3314);  // ../RTL/cortexm0ds_logic.v(10840)
  buf u1211 (vis_r5_o[9], Fx1qw6);  // ../RTL/cortexm0ds_logic.v(1909)
  and u12110 (n3315, Xdaow6, Vxniu6);  // ../RTL/cortexm0ds_logic.v(10841)
  not u12111 (Vcaow6, n3315);  // ../RTL/cortexm0ds_logic.v(10841)
  and u12112 (Xdaow6, D1piu6, Zraiu6);  // ../RTL/cortexm0ds_logic.v(10842)
  and u12113 (D3aow6, Eeaow6, Leaow6);  // ../RTL/cortexm0ds_logic.v(10843)
  and u12114 (Leaow6, Seaow6, Zeaow6);  // ../RTL/cortexm0ds_logic.v(10844)
  and u12115 (n3316, Hs8ow6, Nriiu6);  // ../RTL/cortexm0ds_logic.v(10845)
  not u12116 (Zeaow6, n3316);  // ../RTL/cortexm0ds_logic.v(10845)
  or u12117 (Seaow6, Qojiu6, M32ju6);  // ../RTL/cortexm0ds_logic.v(10846)
  not u12118 (Qojiu6, M2piu6);  // ../RTL/cortexm0ds_logic.v(10847)
  and u12119 (Eeaow6, Ez1ju6, Oeziu6);  // ../RTL/cortexm0ds_logic.v(10848)
  buf u1212 (vis_r5_o[15], Z98bx6);  // ../RTL/cortexm0ds_logic.v(1909)
  and u12120 (Oeziu6, Gfaow6, HREADY);  // ../RTL/cortexm0ds_logic.v(10849)
  and u12121 (Gfaow6, Thaiu6, Dz6ow6);  // ../RTL/cortexm0ds_logic.v(10850)
  or u12122 (Thaiu6, E45iu6, Y2oiu6);  // ../RTL/cortexm0ds_logic.v(10851)
  and u12123 (Ez1ju6, Nfaow6, J5aiu6);  // ../RTL/cortexm0ds_logic.v(10852)
  or u12124 (J5aiu6, Qp3ju6, Jojiu6);  // ../RTL/cortexm0ds_logic.v(10853)
  not u12125 (Qp3ju6, J79ow6);  // ../RTL/cortexm0ds_logic.v(10854)
  and u12126 (Nfaow6, Ufaow6, Bgaow6);  // ../RTL/cortexm0ds_logic.v(10855)
  or u12127 (Ufaow6, H3piu6, Cyfpw6[6]);  // ../RTL/cortexm0ds_logic.v(10856)
  not u12128 (H3piu6, C78iu6);  // ../RTL/cortexm0ds_logic.v(10857)
  and u12129 (C78iu6, S6aiu6, Neoiu6);  // ../RTL/cortexm0ds_logic.v(10858)
  and u1213 (n68, T8yhu6, Zazhu6);  // ../RTL/cortexm0ds_logic.v(3296)
  or u12130 (Ar9ow6, Cyfpw6[4], HREADY);  // ../RTL/cortexm0ds_logic.v(10859)
  not u12131 (Vqohu6, Igaow6);  // ../RTL/cortexm0ds_logic.v(10860)
  AL_MUX u12132 (
    .i0(Xe8iu6),
    .i1(Pgaow6),
    .sel(HREADY),
    .o(Igaow6));  // ../RTL/cortexm0ds_logic.v(10861)
  and u12133 (Pgaow6, Wgaow6, Dhaow6);  // ../RTL/cortexm0ds_logic.v(10862)
  and u12134 (Dhaow6, Khaow6, Rhaow6);  // ../RTL/cortexm0ds_logic.v(10863)
  and u12135 (Rhaow6, Yhaow6, Fiaow6);  // ../RTL/cortexm0ds_logic.v(10864)
  and u12136 (Fiaow6, Miaow6, Tiaow6);  // ../RTL/cortexm0ds_logic.v(10865)
  and u12137 (n3317, Ajaow6, Hjaow6);  // ../RTL/cortexm0ds_logic.v(10866)
  not u12138 (Tiaow6, n3317);  // ../RTL/cortexm0ds_logic.v(10866)
  or u12139 (n3318, Qpaju6, D7fpw6[13]);  // ../RTL/cortexm0ds_logic.v(10867)
  not u1214 (Nbzhu6, n68);  // ../RTL/cortexm0ds_logic.v(3296)
  not u12140 (Hjaow6, n3318);  // ../RTL/cortexm0ds_logic.v(10867)
  and u12141 (Ajaow6, Raaow6, Imaiu6);  // ../RTL/cortexm0ds_logic.v(10868)
  and u12142 (Miaow6, Imoiu6, Dz6ow6);  // ../RTL/cortexm0ds_logic.v(10869)
  and u12143 (n3319, Ojaow6, N20ju6);  // ../RTL/cortexm0ds_logic.v(10870)
  not u12144 (Dz6ow6, n3319);  // ../RTL/cortexm0ds_logic.v(10870)
  or u12145 (n3320, Ii0iu6, Lraiu6);  // ../RTL/cortexm0ds_logic.v(10871)
  not u12146 (Ojaow6, n3320);  // ../RTL/cortexm0ds_logic.v(10871)
  and u12147 (n3321, Pfoiu6, Pu1ju6);  // ../RTL/cortexm0ds_logic.v(10872)
  not u12148 (Imoiu6, n3321);  // ../RTL/cortexm0ds_logic.v(10872)
  and u12149 (Yhaow6, Vjaow6, Ckaow6);  // ../RTL/cortexm0ds_logic.v(10873)
  or u1215 (n69, O9yhu6, U5yhu6);  // ../RTL/cortexm0ds_logic.v(3297)
  and u12150 (n3322, Jkaow6, Qkaow6);  // ../RTL/cortexm0ds_logic.v(10874)
  not u12151 (Ckaow6, n3322);  // ../RTL/cortexm0ds_logic.v(10874)
  and u12152 (Qkaow6, L45iu6, Oiaiu6);  // ../RTL/cortexm0ds_logic.v(10875)
  or u12153 (n3323, Wfoiu6, Xkaow6);  // ../RTL/cortexm0ds_logic.v(10876)
  not u12154 (Jkaow6, n3323);  // ../RTL/cortexm0ds_logic.v(10876)
  and u12155 (n3324, Elaow6, J79ow6);  // ../RTL/cortexm0ds_logic.v(10877)
  not u12156 (Vjaow6, n3324);  // ../RTL/cortexm0ds_logic.v(10877)
  and u12157 (Elaow6, U98iu6, Taaiu6);  // ../RTL/cortexm0ds_logic.v(10878)
  and u12158 (U98iu6, Llaow6, Jjhiu6);  // ../RTL/cortexm0ds_logic.v(10879)
  and u12159 (Khaow6, Slaow6, Zlaow6);  // ../RTL/cortexm0ds_logic.v(10880)
  not u1216 (T8yhu6, n69);  // ../RTL/cortexm0ds_logic.v(3297)
  and u12160 (Zlaow6, Gmaow6, Nmaow6);  // ../RTL/cortexm0ds_logic.v(10881)
  and u12161 (n3325, Llaow6, Umaow6);  // ../RTL/cortexm0ds_logic.v(10882)
  not u12162 (Nmaow6, n3325);  // ../RTL/cortexm0ds_logic.v(10882)
  and u12163 (n3326, Bnaow6, Inaow6);  // ../RTL/cortexm0ds_logic.v(10883)
  not u12164 (Umaow6, n3326);  // ../RTL/cortexm0ds_logic.v(10883)
  and u12165 (n3327, Pnaow6, Ruaiu6);  // ../RTL/cortexm0ds_logic.v(10884)
  not u12166 (Inaow6, n3327);  // ../RTL/cortexm0ds_logic.v(10884)
  and u12167 (n3328, Wnaow6, Doaow6);  // ../RTL/cortexm0ds_logic.v(10885)
  not u12168 (Pnaow6, n3328);  // ../RTL/cortexm0ds_logic.v(10885)
  and u12169 (Doaow6, Koaow6, Xa6ow6);  // ../RTL/cortexm0ds_logic.v(10886)
  and u1217 (O9yhu6, Fnnhu6, Ubzhu6);  // ../RTL/cortexm0ds_logic.v(3298)
  and u12170 (n3329, Roaow6, Cyfpw6[7]);  // ../RTL/cortexm0ds_logic.v(10887)
  not u12171 (Xa6ow6, n3329);  // ../RTL/cortexm0ds_logic.v(10887)
  or u12172 (n3330, Geaiu6, Cyfpw6[3]);  // ../RTL/cortexm0ds_logic.v(10888)
  not u12173 (Roaow6, n3330);  // ../RTL/cortexm0ds_logic.v(10888)
  and u12174 (n3331, Yoaow6, Hzziu6);  // ../RTL/cortexm0ds_logic.v(10889)
  not u12175 (Koaow6, n3331);  // ../RTL/cortexm0ds_logic.v(10889)
  and u12176 (Yoaow6, Fpaow6, Mr0iu6);  // ../RTL/cortexm0ds_logic.v(10890)
  and u12177 (n3332, Mpaow6, Tpaow6);  // ../RTL/cortexm0ds_logic.v(10891)
  not u12178 (Fpaow6, n3332);  // ../RTL/cortexm0ds_logic.v(10891)
  or u12179 (Tpaow6, X1ziu6, S1ehu6);  // ../RTL/cortexm0ds_logic.v(10892)
  or u1218 (Ubzhu6, Jayhu6, Cayhu6);  // ../RTL/cortexm0ds_logic.v(3299)
  and u12180 (Wnaow6, Aqaow6, Hqaow6);  // ../RTL/cortexm0ds_logic.v(10893)
  or u12181 (Hqaow6, Z6oiu6, Geaiu6);  // ../RTL/cortexm0ds_logic.v(10894)
  or u12182 (Aqaow6, R75iu6, Cyfpw6[6]);  // ../RTL/cortexm0ds_logic.v(10895)
  and u12183 (n3333, Nu9ow6, V4aiu6);  // ../RTL/cortexm0ds_logic.v(10896)
  not u12184 (Bnaow6, n3333);  // ../RTL/cortexm0ds_logic.v(10896)
  and u12185 (Gmaow6, Oqaow6, Vqaow6);  // ../RTL/cortexm0ds_logic.v(10897)
  and u12186 (n3334, Yi7ju6, Pu1ju6);  // ../RTL/cortexm0ds_logic.v(10898)
  not u12187 (Vqaow6, n3334);  // ../RTL/cortexm0ds_logic.v(10898)
  or u12188 (n3335, Ii0iu6, Cyfpw6[6]);  // ../RTL/cortexm0ds_logic.v(10899)
  not u12189 (Yi7ju6, n3335);  // ../RTL/cortexm0ds_logic.v(10899)
  and u1219 (Cayhu6, Bczhu6, Ighpw6[4]);  // ../RTL/cortexm0ds_logic.v(3300)
  and u12190 (n3336, Yo1ju6, Craow6);  // ../RTL/cortexm0ds_logic.v(10900)
  not u12191 (Oqaow6, n3336);  // ../RTL/cortexm0ds_logic.v(10900)
  and u12192 (n3337, Jraow6, Qraow6);  // ../RTL/cortexm0ds_logic.v(10901)
  not u12193 (Craow6, n3337);  // ../RTL/cortexm0ds_logic.v(10901)
  or u12194 (Qraow6, L7aow6, O7ziu6);  // ../RTL/cortexm0ds_logic.v(10902)
  and u12195 (n3338, D7fpw6[8], Xraow6);  // ../RTL/cortexm0ds_logic.v(10903)
  not u12196 (Jraow6, n3338);  // ../RTL/cortexm0ds_logic.v(10903)
  and u12197 (n3339, Esaow6, Lsaow6);  // ../RTL/cortexm0ds_logic.v(10904)
  not u12198 (Xraow6, n3339);  // ../RTL/cortexm0ds_logic.v(10904)
  and u12199 (n3340, D7fpw6[9], Dcziu6);  // ../RTL/cortexm0ds_logic.v(10905)
  buf u122 (vis_r5_o[19], Jrvpw6);  // ../RTL/cortexm0ds_logic.v(1909)
  or u1220 (n70, Ujyhu6, Zwyhu6);  // ../RTL/cortexm0ds_logic.v(3301)
  not u12200 (Lsaow6, n3340);  // ../RTL/cortexm0ds_logic.v(10905)
  and u12201 (n3341, Qxoiu6, O95iu6);  // ../RTL/cortexm0ds_logic.v(10906)
  not u12202 (Esaow6, n3341);  // ../RTL/cortexm0ds_logic.v(10906)
  and u12203 (Yo1ju6, Ba8iu6, Ssaow6);  // ../RTL/cortexm0ds_logic.v(10907)
  or u12204 (n3342, S80ju6, D7fpw6[13]);  // ../RTL/cortexm0ds_logic.v(10908)
  not u12205 (Ba8iu6, n3342);  // ../RTL/cortexm0ds_logic.v(10908)
  and u12206 (Slaow6, Zsaow6, Gtaow6);  // ../RTL/cortexm0ds_logic.v(10909)
  and u12207 (n3343, Ntaow6, Zraiu6);  // ../RTL/cortexm0ds_logic.v(10910)
  not u12208 (Gtaow6, n3343);  // ../RTL/cortexm0ds_logic.v(10910)
  and u12209 (n3344, Rz6ow6, Utaow6);  // ../RTL/cortexm0ds_logic.v(10911)
  not u1221 (Bczhu6, n70);  // ../RTL/cortexm0ds_logic.v(3301)
  not u12210 (Ntaow6, n3344);  // ../RTL/cortexm0ds_logic.v(10911)
  or u12211 (Utaow6, Gtgiu6, Iuniu6);  // ../RTL/cortexm0ds_logic.v(10912)
  not u12212 (Gtgiu6, Buaow6);  // ../RTL/cortexm0ds_logic.v(10913)
  and u12213 (n3345, Iuaow6, Nu9ow6);  // ../RTL/cortexm0ds_logic.v(10914)
  not u12214 (Rz6ow6, n3345);  // ../RTL/cortexm0ds_logic.v(10914)
  or u12215 (n3346, Nlaiu6, H4ghu6);  // ../RTL/cortexm0ds_logic.v(10915)
  not u12216 (Iuaow6, n3346);  // ../RTL/cortexm0ds_logic.v(10915)
  and u12217 (n3347, Rljiu6, It2ju6);  // ../RTL/cortexm0ds_logic.v(10916)
  not u12218 (Zsaow6, n3347);  // ../RTL/cortexm0ds_logic.v(10916)
  and u12219 (Rljiu6, Xzmiu6, Cyfpw6[5]);  // ../RTL/cortexm0ds_logic.v(10917)
  and u1222 (n71, U5yhu6, Iczhu6);  // ../RTL/cortexm0ds_logic.v(3302)
  and u12220 (Wgaow6, Puaow6, Wuaow6);  // ../RTL/cortexm0ds_logic.v(10918)
  and u12221 (Wuaow6, Dvaow6, Kvaow6);  // ../RTL/cortexm0ds_logic.v(10919)
  and u12222 (Kvaow6, Rvaow6, Yvaow6);  // ../RTL/cortexm0ds_logic.v(10920)
  or u12223 (Yvaow6, Rb0ju6, Fwaow6);  // ../RTL/cortexm0ds_logic.v(10921)
  and u12224 (n3348, Bziiu6, Oviiu6);  // ../RTL/cortexm0ds_logic.v(10922)
  not u12225 (Rb0ju6, n3348);  // ../RTL/cortexm0ds_logic.v(10922)
  and u12226 (Rvaow6, Mwaow6, Twaow6);  // ../RTL/cortexm0ds_logic.v(10923)
  and u12227 (n3349, D7fpw6[12], Axaow6);  // ../RTL/cortexm0ds_logic.v(10924)
  not u12228 (Twaow6, n3349);  // ../RTL/cortexm0ds_logic.v(10924)
  and u12229 (n3350, Hxaow6, Oxaow6);  // ../RTL/cortexm0ds_logic.v(10925)
  not u1223 (Gbzhu6, n71);  // ../RTL/cortexm0ds_logic.v(3302)
  not u12230 (Axaow6, n3350);  // ../RTL/cortexm0ds_logic.v(10925)
  or u12231 (Oxaow6, Fwaow6, N38ow6);  // ../RTL/cortexm0ds_logic.v(10926)
  not u12232 (Fwaow6, Ssaow6);  // ../RTL/cortexm0ds_logic.v(10927)
  and u12233 (Hxaow6, Vxaow6, Cyaow6);  // ../RTL/cortexm0ds_logic.v(10928)
  and u12234 (n3351, Jyaow6, Qyaow6);  // ../RTL/cortexm0ds_logic.v(10929)
  not u12235 (Cyaow6, n3351);  // ../RTL/cortexm0ds_logic.v(10929)
  and u12236 (Qyaow6, Xyaow6, Geaiu6);  // ../RTL/cortexm0ds_logic.v(10930)
  and u12237 (n3352, Jz9ow6, Ezaow6);  // ../RTL/cortexm0ds_logic.v(10931)
  not u12238 (Xyaow6, n3352);  // ../RTL/cortexm0ds_logic.v(10931)
  or u12239 (Ezaow6, O7ziu6, Ndiiu6);  // ../RTL/cortexm0ds_logic.v(10932)
  and u1224 (n72, Pczhu6, Wczhu6);  // ../RTL/cortexm0ds_logic.v(3303)
  and u12240 (n3353, Xg7ow6, Cwiiu6);  // ../RTL/cortexm0ds_logic.v(10933)
  not u12241 (Jz9ow6, n3353);  // ../RTL/cortexm0ds_logic.v(10933)
  or u12242 (n3354, Tniiu6, D7fpw6[8]);  // ../RTL/cortexm0ds_logic.v(10934)
  not u12243 (Xg7ow6, n3354);  // ../RTL/cortexm0ds_logic.v(10934)
  and u12244 (Jyaow6, Vviiu6, Kxziu6);  // ../RTL/cortexm0ds_logic.v(10935)
  and u12245 (n3355, Lzaow6, W82ju6);  // ../RTL/cortexm0ds_logic.v(10936)
  not u12246 (Vxaow6, n3355);  // ../RTL/cortexm0ds_logic.v(10936)
  and u12247 (W82ju6, Szaow6, D7fpw6[5]);  // ../RTL/cortexm0ds_logic.v(10937)
  or u12248 (n3356, D7fpw6[6], D7fpw6[7]);  // ../RTL/cortexm0ds_logic.v(10938)
  not u12249 (Szaow6, n3356);  // ../RTL/cortexm0ds_logic.v(10938)
  not u1225 (Iczhu6, n72);  // ../RTL/cortexm0ds_logic.v(3303)
  or u12250 (n3357, P82ju6, A1kiu6);  // ../RTL/cortexm0ds_logic.v(10939)
  not u12251 (Lzaow6, n3357);  // ../RTL/cortexm0ds_logic.v(10939)
  and u12252 (n3358, Zzaow6, G0bow6);  // ../RTL/cortexm0ds_logic.v(10940)
  not u12253 (P82ju6, n3358);  // ../RTL/cortexm0ds_logic.v(10940)
  and u12254 (G0bow6, Rmiiu6, D7fpw6[8]);  // ../RTL/cortexm0ds_logic.v(10941)
  and u12255 (Rmiiu6, F6ziu6, Th2ju6);  // ../RTL/cortexm0ds_logic.v(10942)
  and u12256 (Zzaow6, Wh0ju6, Htyiu6);  // ../RTL/cortexm0ds_logic.v(10943)
  and u12257 (n3359, Hzziu6, N0bow6);  // ../RTL/cortexm0ds_logic.v(10944)
  not u12258 (Mwaow6, n3359);  // ../RTL/cortexm0ds_logic.v(10944)
  and u12259 (n3360, U0bow6, B1bow6);  // ../RTL/cortexm0ds_logic.v(10945)
  and u1226 (Wczhu6, Ddzhu6, Kdzhu6);  // ../RTL/cortexm0ds_logic.v(3304)
  not u12260 (N0bow6, n3360);  // ../RTL/cortexm0ds_logic.v(10945)
  and u12261 (n3361, Oxniu6, Tfjiu6);  // ../RTL/cortexm0ds_logic.v(10946)
  not u12262 (B1bow6, n3361);  // ../RTL/cortexm0ds_logic.v(10946)
  and u12263 (U0bow6, I1bow6, P1bow6);  // ../RTL/cortexm0ds_logic.v(10947)
  and u12264 (n3362, W1bow6, Ia8iu6);  // ../RTL/cortexm0ds_logic.v(10948)
  not u12265 (I1bow6, n3362);  // ../RTL/cortexm0ds_logic.v(10948)
  and u12266 (W1bow6, Aujiu6, Frziu6);  // ../RTL/cortexm0ds_logic.v(10949)
  and u12267 (Dvaow6, D2bow6, K2bow6);  // ../RTL/cortexm0ds_logic.v(10950)
  and u12268 (n3363, Qe8iu6, R2bow6);  // ../RTL/cortexm0ds_logic.v(10951)
  not u12269 (K2bow6, n3363);  // ../RTL/cortexm0ds_logic.v(10951)
  or u1227 (n73, X9zhu6, A1zhu6);  // ../RTL/cortexm0ds_logic.v(3305)
  and u12270 (n3364, Y2bow6, F3bow6);  // ../RTL/cortexm0ds_logic.v(10952)
  not u12271 (R2bow6, n3364);  // ../RTL/cortexm0ds_logic.v(10952)
  or u12272 (n3365, J79ow6, D31ju6);  // ../RTL/cortexm0ds_logic.v(10953)
  not u12273 (F3bow6, n3365);  // ../RTL/cortexm0ds_logic.v(10953)
  and u12274 (Y2bow6, M3bow6, T3bow6);  // ../RTL/cortexm0ds_logic.v(10954)
  or u12275 (T3bow6, Jc2ju6, Knaiu6);  // ../RTL/cortexm0ds_logic.v(10955)
  and u12276 (n3366, Frziu6, K2aiu6);  // ../RTL/cortexm0ds_logic.v(10956)
  not u12277 (M3bow6, n3366);  // ../RTL/cortexm0ds_logic.v(10956)
  and u12278 (n3367, D7fpw6[11], A4bow6);  // ../RTL/cortexm0ds_logic.v(10957)
  not u12279 (D2bow6, n3367);  // ../RTL/cortexm0ds_logic.v(10957)
  not u1228 (Kdzhu6, n73);  // ../RTL/cortexm0ds_logic.v(3305)
  and u12280 (n3368, H4bow6, O4bow6);  // ../RTL/cortexm0ds_logic.v(10958)
  not u12281 (A4bow6, n3368);  // ../RTL/cortexm0ds_logic.v(10958)
  and u12282 (O4bow6, V4bow6, C5bow6);  // ../RTL/cortexm0ds_logic.v(10959)
  and u12283 (n3369, J5bow6, Yv1ju6);  // ../RTL/cortexm0ds_logic.v(10960)
  not u12284 (C5bow6, n3369);  // ../RTL/cortexm0ds_logic.v(10960)
  and u12285 (Yv1ju6, Ssaow6, X1ziu6);  // ../RTL/cortexm0ds_logic.v(10961)
  or u12286 (n3370, Tniiu6, Jjhiu6);  // ../RTL/cortexm0ds_logic.v(10962)
  not u12287 (J5bow6, n3370);  // ../RTL/cortexm0ds_logic.v(10962)
  and u12288 (n3371, Q5bow6, Htyiu6);  // ../RTL/cortexm0ds_logic.v(10963)
  not u12289 (V4bow6, n3371);  // ../RTL/cortexm0ds_logic.v(10963)
  and u1229 (X9zhu6, Rdzhu6, Iyyhu6);  // ../RTL/cortexm0ds_logic.v(3306)
  or u12290 (n3372, C27ow6, Ae0iu6);  // ../RTL/cortexm0ds_logic.v(10964)
  not u12291 (Q5bow6, n3372);  // ../RTL/cortexm0ds_logic.v(10964)
  and u12292 (H4bow6, X5bow6, E6bow6);  // ../RTL/cortexm0ds_logic.v(10965)
  and u12293 (n3373, Ssaow6, Evyiu6);  // ../RTL/cortexm0ds_logic.v(10966)
  not u12294 (E6bow6, n3373);  // ../RTL/cortexm0ds_logic.v(10966)
  and u12295 (Ssaow6, L6bow6, Y31ju6);  // ../RTL/cortexm0ds_logic.v(10967)
  or u12296 (n3374, Xkaow6, D7fpw6[15]);  // ../RTL/cortexm0ds_logic.v(10968)
  not u12297 (L6bow6, n3374);  // ../RTL/cortexm0ds_logic.v(10968)
  or u12298 (X5bow6, Ax1ju6, Ad8iu6);  // ../RTL/cortexm0ds_logic.v(10969)
  and u12299 (Puaow6, S6bow6, Z6bow6);  // ../RTL/cortexm0ds_logic.v(10970)
  buf u123 (Punhu6, Cjqpw6);  // ../RTL/cortexm0ds_logic.v(1932)
  or u1230 (n74, Sbyhu6, Ighpw6[0]);  // ../RTL/cortexm0ds_logic.v(3307)
  and u12300 (Z6bow6, G7bow6, N7bow6);  // ../RTL/cortexm0ds_logic.v(10971)
  and u12301 (n3375, Omyiu6, U7bow6);  // ../RTL/cortexm0ds_logic.v(10972)
  not u12302 (N7bow6, n3375);  // ../RTL/cortexm0ds_logic.v(10972)
  and u12303 (n3376, B8bow6, I8bow6);  // ../RTL/cortexm0ds_logic.v(10973)
  not u12304 (U7bow6, n3376);  // ../RTL/cortexm0ds_logic.v(10973)
  and u12305 (I8bow6, P8bow6, W8bow6);  // ../RTL/cortexm0ds_logic.v(10974)
  and u12306 (n3377, Apaiu6, D9bow6);  // ../RTL/cortexm0ds_logic.v(10975)
  not u12307 (W8bow6, n3377);  // ../RTL/cortexm0ds_logic.v(10975)
  and u12308 (n3378, K9bow6, R9bow6);  // ../RTL/cortexm0ds_logic.v(10976)
  not u12309 (D9bow6, n3378);  // ../RTL/cortexm0ds_logic.v(10976)
  not u1231 (Rdzhu6, n74);  // ../RTL/cortexm0ds_logic.v(3307)
  and u12310 (n3379, Y9bow6, Tfjiu6);  // ../RTL/cortexm0ds_logic.v(10977)
  not u12311 (R9bow6, n3379);  // ../RTL/cortexm0ds_logic.v(10977)
  or u12312 (Y9bow6, Y2oiu6, P0biu6);  // ../RTL/cortexm0ds_logic.v(10978)
  and u12313 (P8bow6, Fabow6, Mabow6);  // ../RTL/cortexm0ds_logic.v(10979)
  and u12314 (n3380, Tabow6, T4aow6);  // ../RTL/cortexm0ds_logic.v(10980)
  not u12315 (Mabow6, n3380);  // ../RTL/cortexm0ds_logic.v(10980)
  and u12316 (T4aow6, Abbow6, Hbbow6);  // ../RTL/cortexm0ds_logic.v(10981)
  and u12317 (Abbow6, Ya1ju6, Frziu6);  // ../RTL/cortexm0ds_logic.v(10982)
  or u12318 (n3381, G7oiu6, Qpaju6);  // ../RTL/cortexm0ds_logic.v(10983)
  not u12319 (Tabow6, n3381);  // ../RTL/cortexm0ds_logic.v(10983)
  and u1232 (Sbyhu6, Ydzhu6, Fezhu6);  // ../RTL/cortexm0ds_logic.v(3308)
  and u12320 (n3382, Obbow6, Vbbow6);  // ../RTL/cortexm0ds_logic.v(10984)
  not u12321 (Fabow6, n3382);  // ../RTL/cortexm0ds_logic.v(10984)
  or u12322 (Vbbow6, Wp0iu6, Ep6ow6);  // ../RTL/cortexm0ds_logic.v(10985)
  and u12323 (Ep6ow6, Taaiu6, Tr0iu6);  // ../RTL/cortexm0ds_logic.v(10986)
  and u12324 (B8bow6, Ccbow6, Jcbow6);  // ../RTL/cortexm0ds_logic.v(10987)
  and u12325 (n3383, Qcbow6, Ruaiu6);  // ../RTL/cortexm0ds_logic.v(10988)
  not u12326 (Jcbow6, n3383);  // ../RTL/cortexm0ds_logic.v(10988)
  and u12327 (n3384, Xcbow6, Edbow6);  // ../RTL/cortexm0ds_logic.v(10989)
  not u12328 (Qcbow6, n3384);  // ../RTL/cortexm0ds_logic.v(10989)
  and u12329 (n3385, Sy2ju6, Kxziu6);  // ../RTL/cortexm0ds_logic.v(10990)
  and u1233 (Fezhu6, Mdhpw6[1], Mezhu6);  // ../RTL/cortexm0ds_logic.v(3309)
  not u12330 (Edbow6, n3385);  // ../RTL/cortexm0ds_logic.v(10990)
  and u12331 (Sy2ju6, Cyfpw6[4], Mr0iu6);  // ../RTL/cortexm0ds_logic.v(10991)
  or u12332 (Xcbow6, P1bow6, Knaiu6);  // ../RTL/cortexm0ds_logic.v(10992)
  and u12333 (n3386, Oxniu6, Pugiu6);  // ../RTL/cortexm0ds_logic.v(10993)
  not u12334 (Ccbow6, n3386);  // ../RTL/cortexm0ds_logic.v(10993)
  and u12335 (Oxniu6, Cyfpw6[0], Zraiu6);  // ../RTL/cortexm0ds_logic.v(10994)
  or u12336 (G7bow6, Ax1ju6, D7fpw6[7]);  // ../RTL/cortexm0ds_logic.v(10995)
  and u12337 (n3387, Ldbow6, Z4jiu6);  // ../RTL/cortexm0ds_logic.v(10996)
  not u12338 (Ax1ju6, n3387);  // ../RTL/cortexm0ds_logic.v(10996)
  or u12339 (n3388, Hujiu6, Gkiiu6);  // ../RTL/cortexm0ds_logic.v(10997)
  or u1234 (Mezhu6, Iahpw6[8], Iahpw6[7]);  // ../RTL/cortexm0ds_logic.v(3310)
  not u12340 (Z4jiu6, n3388);  // ../RTL/cortexm0ds_logic.v(10997)
  and u12341 (Ldbow6, Htyiu6, Sdbow6);  // ../RTL/cortexm0ds_logic.v(10998)
  and u12342 (Htyiu6, W0piu6, Geaiu6);  // ../RTL/cortexm0ds_logic.v(10999)
  or u12343 (n3389, Zdbow6, Gebow6);  // ../RTL/cortexm0ds_logic.v(11000)
  not u12344 (S6bow6, n3389);  // ../RTL/cortexm0ds_logic.v(11000)
  or u12345 (n3390, R2aiu6, Lkaiu6);  // ../RTL/cortexm0ds_logic.v(11001)
  not u12346 (Gebow6, n3390);  // ../RTL/cortexm0ds_logic.v(11001)
  AL_MUX u12347 (
    .i0(Mfjiu6),
    .i1(Nebow6),
    .sel(Cyfpw6[7]),
    .o(Zdbow6));  // ../RTL/cortexm0ds_logic.v(11002)
  and u12348 (n3391, Uebow6, Bfbow6);  // ../RTL/cortexm0ds_logic.v(11003)
  not u12349 (Nebow6, n3391);  // ../RTL/cortexm0ds_logic.v(11003)
  and u1235 (Ydzhu6, Tezhu6, Pinhu6);  // ../RTL/cortexm0ds_logic.v(3311)
  and u12350 (n3392, D6kiu6, Pugiu6);  // ../RTL/cortexm0ds_logic.v(11004)
  not u12351 (Bfbow6, n3392);  // ../RTL/cortexm0ds_logic.v(11004)
  and u12352 (Uebow6, Ifbow6, Pfbow6);  // ../RTL/cortexm0ds_logic.v(11005)
  and u12353 (n3393, I82ju6, Xojiu6);  // ../RTL/cortexm0ds_logic.v(11006)
  not u12354 (Pfbow6, n3393);  // ../RTL/cortexm0ds_logic.v(11006)
  and u12355 (n3394, Jf6ju6, It2ju6);  // ../RTL/cortexm0ds_logic.v(11007)
  not u12356 (Ifbow6, n3394);  // ../RTL/cortexm0ds_logic.v(11007)
  and u12357 (n3395, Wfbow6, Dgbow6);  // ../RTL/cortexm0ds_logic.v(11008)
  not u12358 (Oqohu6, n3395);  // ../RTL/cortexm0ds_logic.v(11008)
  and u12359 (n3396, Y7ghu6, Kgbow6);  // ../RTL/cortexm0ds_logic.v(11009)
  and u1236 (Ddzhu6, Afzhu6, Iryhu6);  // ../RTL/cortexm0ds_logic.v(3312)
  not u12360 (Dgbow6, n3396);  // ../RTL/cortexm0ds_logic.v(11009)
  or u12361 (Kgbow6, Eh6iu6, J79ow6);  // ../RTL/cortexm0ds_logic.v(11010)
  and u12362 (J79ow6, Ii0iu6, Hs0iu6);  // ../RTL/cortexm0ds_logic.v(11011)
  and u12363 (n3397, HREADY, Rgbow6);  // ../RTL/cortexm0ds_logic.v(11012)
  not u12364 (Wfbow6, n3397);  // ../RTL/cortexm0ds_logic.v(11012)
  and u12365 (n3398, Ygbow6, Fhbow6);  // ../RTL/cortexm0ds_logic.v(11013)
  not u12366 (Rgbow6, n3398);  // ../RTL/cortexm0ds_logic.v(11013)
  and u12367 (Fhbow6, Mhbow6, Thbow6);  // ../RTL/cortexm0ds_logic.v(11014)
  and u12368 (Thbow6, Aibow6, Hibow6);  // ../RTL/cortexm0ds_logic.v(11015)
  and u12369 (n3399, Oibow6, Vibow6);  // ../RTL/cortexm0ds_logic.v(11016)
  and u1237 (n75, Hfzhu6, M7zhu6);  // ../RTL/cortexm0ds_logic.v(3313)
  not u12370 (Hibow6, n3399);  // ../RTL/cortexm0ds_logic.v(11016)
  or u12371 (n3400, D7fpw6[8], Sbghu6);  // ../RTL/cortexm0ds_logic.v(11017)
  not u12372 (Vibow6, n3400);  // ../RTL/cortexm0ds_logic.v(11017)
  and u12373 (Oibow6, Dd7ow6, Jehhu6);  // ../RTL/cortexm0ds_logic.v(11018)
  and u12374 (Dd7ow6, Cjbow6, Jjbow6);  // ../RTL/cortexm0ds_logic.v(11019)
  and u12375 (Jjbow6, J9kiu6, D7fpw6[13]);  // ../RTL/cortexm0ds_logic.v(11020)
  and u12376 (Cjbow6, Y40ju6, F6ziu6);  // ../RTL/cortexm0ds_logic.v(11021)
  and u12377 (n3401, Imaiu6, Qjbow6);  // ../RTL/cortexm0ds_logic.v(11022)
  not u12378 (Aibow6, n3401);  // ../RTL/cortexm0ds_logic.v(11022)
  or u12379 (Qjbow6, Lraiu6, Xjbow6);  // ../RTL/cortexm0ds_logic.v(11023)
  not u1238 (Iryhu6, n75);  // ../RTL/cortexm0ds_logic.v(3313)
  and u12380 (Mhbow6, Vx1ju6, Ekbow6);  // ../RTL/cortexm0ds_logic.v(11024)
  and u12381 (n3402, Lkbow6, Xe8iu6);  // ../RTL/cortexm0ds_logic.v(11025)
  not u12382 (Ekbow6, n3402);  // ../RTL/cortexm0ds_logic.v(11025)
  and u12383 (n3403, Skbow6, Zkbow6);  // ../RTL/cortexm0ds_logic.v(11026)
  not u12384 (Lkbow6, n3403);  // ../RTL/cortexm0ds_logic.v(11026)
  or u12385 (Zkbow6, K9aiu6, Sbghu6);  // ../RTL/cortexm0ds_logic.v(11027)
  and u12386 (Skbow6, Glbow6, Nlbow6);  // ../RTL/cortexm0ds_logic.v(11028)
  and u12387 (n3404, Ulbow6, Xjbow6);  // ../RTL/cortexm0ds_logic.v(11029)
  not u12388 (Nlbow6, n3404);  // ../RTL/cortexm0ds_logic.v(11029)
  buf u12389 (Abfhu6, Ozkbx6[10]);  // ../RTL/cortexm0ds_logic.v(3176)
  and u1239 (Hfzhu6, Ofzhu6, Vfzhu6);  // ../RTL/cortexm0ds_logic.v(3315)
  not u12390 (Ulbow6, Hhaju6);  // ../RTL/cortexm0ds_logic.v(11030)
  not u12391 (Szniu6, Kfiiu6);  // ../RTL/cortexm0ds_logic.v(11031)
  and u12392 (Kfiiu6, Cyfpw6[4], K9aiu6);  // ../RTL/cortexm0ds_logic.v(11032)
  and u12393 (n3405, Bmbow6, E6oiu6);  // ../RTL/cortexm0ds_logic.v(11033)
  not u12394 (Glbow6, n3405);  // ../RTL/cortexm0ds_logic.v(11033)
  or u12395 (n3406, Q5aiu6, As0iu6);  // ../RTL/cortexm0ds_logic.v(11034)
  not u12396 (Bmbow6, n3406);  // ../RTL/cortexm0ds_logic.v(11034)
  or u12397 (Vx1ju6, Jojiu6, Mjfiu6);  // ../RTL/cortexm0ds_logic.v(11035)
  and u12398 (Ygbow6, Imbow6, Pmbow6);  // ../RTL/cortexm0ds_logic.v(11036)
  and u12399 (Imbow6, Wmbow6, Dnbow6);  // ../RTL/cortexm0ds_logic.v(11037)
  buf u124 (CDBGPWRUPREQ, Xkqpw6);  // ../RTL/cortexm0ds_logic.v(1933)
  not u1240 (T7zhu6, Hfzhu6);  // ../RTL/cortexm0ds_logic.v(3315)
  or u12400 (Dnbow6, Kq0iu6, W2aow6);  // ../RTL/cortexm0ds_logic.v(11038)
  or u12401 (Wmbow6, Zraiu6, Lkaiu6);  // ../RTL/cortexm0ds_logic.v(11039)
  AL_MUX u12402 (
    .i0(V9ghu6),
    .i1(B0biu6),
    .sel(F2biu6),
    .o(Hqohu6));  // ../RTL/cortexm0ds_logic.v(11040)
  not u12403 (B0biu6, Knbow6);  // ../RTL/cortexm0ds_logic.v(11041)
  AL_MUX u12404 (
    .i0(Rnbow6),
    .i1(H2fpw6[2]),
    .sel(G81ju6),
    .o(Aqohu6));  // ../RTL/cortexm0ds_logic.v(11042)
  and u12405 (n3407, Ynbow6, Fobow6);  // ../RTL/cortexm0ds_logic.v(11043)
  not u12406 (Rnbow6, n3407);  // ../RTL/cortexm0ds_logic.v(11043)
  and u12407 (Fobow6, Mobow6, Tobow6);  // ../RTL/cortexm0ds_logic.v(11044)
  and u12408 (n3408, Fb1ju6, D7fpw6[10]);  // ../RTL/cortexm0ds_logic.v(11045)
  not u12409 (Tobow6, n3408);  // ../RTL/cortexm0ds_logic.v(11045)
  and u1241 (n76, Cgzhu6, Jgzhu6);  // ../RTL/cortexm0ds_logic.v(3316)
  and u12410 (Fb1ju6, Llaow6, Apbow6);  // ../RTL/cortexm0ds_logic.v(11046)
  and u12411 (n3409, Hpbow6, Opbow6);  // ../RTL/cortexm0ds_logic.v(11047)
  not u12412 (Apbow6, n3409);  // ../RTL/cortexm0ds_logic.v(11047)
  and u12413 (n3410, Vk9ow6, D7fpw6[13]);  // ../RTL/cortexm0ds_logic.v(11048)
  not u12414 (Opbow6, n3410);  // ../RTL/cortexm0ds_logic.v(11048)
  or u12415 (Hpbow6, Ftjiu6, X1ziu6);  // ../RTL/cortexm0ds_logic.v(11049)
  and u12416 (n3411, P91ju6, D7fpw6[5]);  // ../RTL/cortexm0ds_logic.v(11050)
  not u12417 (Mobow6, n3411);  // ../RTL/cortexm0ds_logic.v(11050)
  and u12418 (P91ju6, Llaow6, Vpbow6);  // ../RTL/cortexm0ds_logic.v(11051)
  and u12419 (n3412, Cqbow6, Jqbow6);  // ../RTL/cortexm0ds_logic.v(11052)
  not u1242 (Vfzhu6, n76);  // ../RTL/cortexm0ds_logic.v(3316)
  not u12420 (Vpbow6, n3412);  // ../RTL/cortexm0ds_logic.v(11052)
  AL_MUX u12421 (
    .i0(Qqbow6),
    .i1(Xqbow6),
    .sel(D7fpw6[13]),
    .o(Jqbow6));  // ../RTL/cortexm0ds_logic.v(11053)
  and u12422 (n3413, Aujiu6, D7fpw6[9]);  // ../RTL/cortexm0ds_logic.v(11054)
  not u12423 (Xqbow6, n3413);  // ../RTL/cortexm0ds_logic.v(11054)
  or u12424 (Qqbow6, Gkiiu6, D7fpw6[15]);  // ../RTL/cortexm0ds_logic.v(11055)
  and u12425 (Cqbow6, Erbow6, Co6ow6);  // ../RTL/cortexm0ds_logic.v(11056)
  or u12426 (Erbow6, Nj6ow6, D7fpw6[12]);  // ../RTL/cortexm0ds_logic.v(11057)
  or u12427 (Nj6ow6, D7fpw6[13], D7fpw6[14]);  // ../RTL/cortexm0ds_logic.v(11058)
  and u12428 (Ynbow6, Ir6ow6, Lrbow6);  // ../RTL/cortexm0ds_logic.v(11059)
  and u12429 (n3414, D7fpw6[2], Ac1ju6);  // ../RTL/cortexm0ds_logic.v(11060)
  or u1243 (n77, Ulnhu6, Mdhpw6[1]);  // ../RTL/cortexm0ds_logic.v(3317)
  not u12430 (Lrbow6, n3414);  // ../RTL/cortexm0ds_logic.v(11060)
  or u12431 (Ac1ju6, Srbow6, Zrbow6);  // ../RTL/cortexm0ds_logic.v(11061)
  and u12432 (Zrbow6, Gsbow6, V4aiu6);  // ../RTL/cortexm0ds_logic.v(11062)
  and u12433 (n3415, Nsbow6, Usbow6);  // ../RTL/cortexm0ds_logic.v(11063)
  not u12434 (Tpohu6, n3415);  // ../RTL/cortexm0ds_logic.v(11063)
  or u12435 (Usbow6, Btbow6, Dk7ow6);  // ../RTL/cortexm0ds_logic.v(11064)
  AL_MUX u12436 (
    .i0(Itbow6),
    .i1(Qjoiu6),
    .sel(Rk7ow6),
    .o(Nsbow6));  // ../RTL/cortexm0ds_logic.v(11065)
  and u12437 (Itbow6, Ptbow6, Wtbow6);  // ../RTL/cortexm0ds_logic.v(11066)
  and u12438 (Wtbow6, Dubow6, Kubow6);  // ../RTL/cortexm0ds_logic.v(11067)
  and u12439 (Kubow6, W6jiu6, Faaiu6);  // ../RTL/cortexm0ds_logic.v(11068)
  not u1244 (Jgzhu6, n77);  // ../RTL/cortexm0ds_logic.v(3317)
  or u12440 (W6jiu6, Jc2ju6, K9aiu6);  // ../RTL/cortexm0ds_logic.v(11069)
  and u12441 (Dubow6, Rubow6, Yubow6);  // ../RTL/cortexm0ds_logic.v(11070)
  and u12442 (n3416, Fvbow6, D7fpw6[10]);  // ../RTL/cortexm0ds_logic.v(11071)
  not u12443 (Yubow6, n3416);  // ../RTL/cortexm0ds_logic.v(11071)
  and u12444 (Fvbow6, Mvbow6, Ftjiu6);  // ../RTL/cortexm0ds_logic.v(11072)
  and u12445 (n3417, O8kiu6, Tvbow6);  // ../RTL/cortexm0ds_logic.v(11073)
  not u12446 (Mvbow6, n3417);  // ../RTL/cortexm0ds_logic.v(11073)
  or u12447 (Tvbow6, Yb9ow6, Qpaju6);  // ../RTL/cortexm0ds_logic.v(11074)
  and u12448 (n3418, Bziiu6, Zraiu6);  // ../RTL/cortexm0ds_logic.v(11075)
  not u12449 (O8kiu6, n3418);  // ../RTL/cortexm0ds_logic.v(11075)
  or u1245 (n78, Qgzhu6, R7yhu6);  // ../RTL/cortexm0ds_logic.v(3318)
  or u12450 (n3419, Co6ow6, Jjhiu6);  // ../RTL/cortexm0ds_logic.v(11076)
  not u12451 (Bziiu6, n3419);  // ../RTL/cortexm0ds_logic.v(11076)
  and u12452 (n3420, Am7ow6, Ppfpw6[4]);  // ../RTL/cortexm0ds_logic.v(11077)
  not u12453 (Rubow6, n3420);  // ../RTL/cortexm0ds_logic.v(11077)
  and u12454 (Am7ow6, Ivfhu6, Awbow6);  // ../RTL/cortexm0ds_logic.v(11078)
  and u12455 (n3421, Hwbow6, Twniu6);  // ../RTL/cortexm0ds_logic.v(11079)
  not u12456 (Awbow6, n3421);  // ../RTL/cortexm0ds_logic.v(11079)
  and u12457 (n3422, D6kiu6, Cyfpw6[1]);  // ../RTL/cortexm0ds_logic.v(11080)
  not u12458 (Twniu6, n3422);  // ../RTL/cortexm0ds_logic.v(11080)
  or u12459 (n3423, Mfjiu6, Gsbow6);  // ../RTL/cortexm0ds_logic.v(11081)
  not u1246 (Cgzhu6, n78);  // ../RTL/cortexm0ds_logic.v(3318)
  not u12460 (Hwbow6, n3423);  // ../RTL/cortexm0ds_logic.v(11081)
  and u12461 (Ptbow6, Owbow6, Vwbow6);  // ../RTL/cortexm0ds_logic.v(11082)
  or u12462 (Vwbow6, V4aiu6, Cn7ow6);  // ../RTL/cortexm0ds_logic.v(11083)
  not u12463 (V4aiu6, D7fpw6[3]);  // ../RTL/cortexm0ds_logic.v(11084)
  and u12464 (Owbow6, Cxbow6, Jxbow6);  // ../RTL/cortexm0ds_logic.v(11085)
  or u12465 (Jxbow6, A1kiu6, Hm7ow6);  // ../RTL/cortexm0ds_logic.v(11086)
  and u12466 (n3424, Cbbiu6, D7fpw6[9]);  // ../RTL/cortexm0ds_logic.v(11087)
  not u12467 (Cxbow6, n3424);  // ../RTL/cortexm0ds_logic.v(11087)
  or u12468 (n3425, Vhiiu6, Ftjiu6);  // ../RTL/cortexm0ds_logic.v(11088)
  not u12469 (Cbbiu6, n3425);  // ../RTL/cortexm0ds_logic.v(11088)
  and u1247 (n79, Ziyhu6, Ighpw6[4]);  // ../RTL/cortexm0ds_logic.v(3319)
  or u12470 (Vhiiu6, C27ow6, Qpaju6);  // ../RTL/cortexm0ds_logic.v(11089)
  and u12471 (n3426, Qxbow6, Xxbow6);  // ../RTL/cortexm0ds_logic.v(11090)
  not u12472 (Mpohu6, n3426);  // ../RTL/cortexm0ds_logic.v(11090)
  and u12473 (Xxbow6, Eybow6, Lybow6);  // ../RTL/cortexm0ds_logic.v(11091)
  and u12474 (n3427, Egziu6, Eafpw6[28]);  // ../RTL/cortexm0ds_logic.v(11092)
  not u12475 (Lybow6, n3427);  // ../RTL/cortexm0ds_logic.v(11092)
  and u12476 (Eybow6, Sybow6, Sgziu6);  // ../RTL/cortexm0ds_logic.v(11093)
  or u12477 (Sybow6, Ft6ow6, Acniu6);  // ../RTL/cortexm0ds_logic.v(11094)
  and u12478 (Acniu6, Zybow6, Gzbow6);  // ../RTL/cortexm0ds_logic.v(11095)
  and u12479 (Gzbow6, Nzbow6, Uzbow6);  // ../RTL/cortexm0ds_logic.v(11096)
  not u1248 (Afzhu6, n79);  // ../RTL/cortexm0ds_logic.v(3319)
  or u12480 (Uzbow6, Iiziu6, B0cow6);  // ../RTL/cortexm0ds_logic.v(11097)
  and u12481 (Nzbow6, I0cow6, Djziu6);  // ../RTL/cortexm0ds_logic.v(11098)
  or u12482 (I0cow6, Kjziu6, P0cow6);  // ../RTL/cortexm0ds_logic.v(11099)
  and u12483 (Zybow6, W0cow6, D1cow6);  // ../RTL/cortexm0ds_logic.v(11100)
  or u12484 (D1cow6, K1cow6, Hlziu6);  // ../RTL/cortexm0ds_logic.v(11101)
  or u12485 (W0cow6, Mkziu6, R1cow6);  // ../RTL/cortexm0ds_logic.v(11102)
  and u12486 (Qxbow6, Y1cow6, F2cow6);  // ../RTL/cortexm0ds_logic.v(11103)
  and u12487 (n3428, Zsfpw6[27], Cmziu6);  // ../RTL/cortexm0ds_logic.v(11104)
  not u12488 (F2cow6, n3428);  // ../RTL/cortexm0ds_logic.v(11104)
  and u12489 (n3429, vis_pc_o[27], Jmziu6);  // ../RTL/cortexm0ds_logic.v(11105)
  or u1249 (n80, Y7yhu6, Zazhu6);  // ../RTL/cortexm0ds_logic.v(3320)
  not u12490 (Y1cow6, n3429);  // ../RTL/cortexm0ds_logic.v(11105)
  and u12491 (n3430, M2cow6, T2cow6);  // ../RTL/cortexm0ds_logic.v(11106)
  not u12492 (Fpohu6, n3430);  // ../RTL/cortexm0ds_logic.v(11106)
  and u12493 (T2cow6, A3cow6, H3cow6);  // ../RTL/cortexm0ds_logic.v(11107)
  and u12494 (n3431, Egziu6, Eafpw6[30]);  // ../RTL/cortexm0ds_logic.v(11108)
  not u12495 (H3cow6, n3431);  // ../RTL/cortexm0ds_logic.v(11108)
  and u12496 (A3cow6, O3cow6, Sgziu6);  // ../RTL/cortexm0ds_logic.v(11109)
  or u12497 (O3cow6, Ft6ow6, D5liu6);  // ../RTL/cortexm0ds_logic.v(11110)
  and u12498 (D5liu6, V3cow6, C4cow6);  // ../RTL/cortexm0ds_logic.v(11111)
  and u12499 (C4cow6, J4cow6, Q4cow6);  // ../RTL/cortexm0ds_logic.v(11112)
  not u125 (W9ohu6, Xkqpw6);  // ../RTL/cortexm0ds_logic.v(1934)
  not u1250 (Ziyhu6, n80);  // ../RTL/cortexm0ds_logic.v(3320)
  and u12500 (n3432, X4cow6, Rc8ow6);  // ../RTL/cortexm0ds_logic.v(11113)
  not u12501 (Q4cow6, n3432);  // ../RTL/cortexm0ds_logic.v(11113)
  and u12502 (J4cow6, E5cow6, Djziu6);  // ../RTL/cortexm0ds_logic.v(11114)
  or u12503 (E5cow6, Mkziu6, L5cow6);  // ../RTL/cortexm0ds_logic.v(11115)
  and u12504 (V3cow6, S5cow6, Z5cow6);  // ../RTL/cortexm0ds_logic.v(11116)
  or u12505 (Z5cow6, Hlziu6, G6cow6);  // ../RTL/cortexm0ds_logic.v(11117)
  and u12506 (n3433, N6cow6, Dc8ow6);  // ../RTL/cortexm0ds_logic.v(11118)
  not u12507 (S5cow6, n3433);  // ../RTL/cortexm0ds_logic.v(11118)
  and u12508 (M2cow6, U6cow6, B7cow6);  // ../RTL/cortexm0ds_logic.v(11119)
  and u12509 (n3434, Zsfpw6[29], Cmziu6);  // ../RTL/cortexm0ds_logic.v(11120)
  and u1251 (Pczhu6, Xgzhu6, J9zhu6);  // ../RTL/cortexm0ds_logic.v(3321)
  not u12510 (B7cow6, n3434);  // ../RTL/cortexm0ds_logic.v(11120)
  and u12511 (n3435, vis_pc_o[29], Jmziu6);  // ../RTL/cortexm0ds_logic.v(11121)
  not u12512 (U6cow6, n3435);  // ../RTL/cortexm0ds_logic.v(11121)
  AL_MUX u12513 (
    .i0(I7cow6),
    .i1(Yyfhu6),
    .sel(n3436),
    .o(Yoohu6));  // ../RTL/cortexm0ds_logic.v(11122)
  or u12514 (n3436, Q08iu6, Eh6iu6);  // ../RTL/cortexm0ds_logic.v(11123)
  buf u12515 (Eafpw6[1], Nxkbx6[2]);  // ../RTL/cortexm0ds_logic.v(3167)
  not u12516 (Q08iu6, W7cow6);  // ../RTL/cortexm0ds_logic.v(11124)
  and u12517 (n3437, D8cow6, K8cow6);  // ../RTL/cortexm0ds_logic.v(11125)
  not u12518 (Roohu6, n3437);  // ../RTL/cortexm0ds_logic.v(11125)
  and u12519 (K8cow6, R8cow6, Y8cow6);  // ../RTL/cortexm0ds_logic.v(11126)
  and u1252 (J9zhu6, Ehzhu6, Lhzhu6);  // ../RTL/cortexm0ds_logic.v(3322)
  and u12520 (n3438, Zsfpw6[22], Cmziu6);  // ../RTL/cortexm0ds_logic.v(11127)
  not u12521 (Y8cow6, n3438);  // ../RTL/cortexm0ds_logic.v(11127)
  and u12522 (R8cow6, F9cow6, M9cow6);  // ../RTL/cortexm0ds_logic.v(11128)
  or u12523 (M9cow6, Ft6ow6, Lvkiu6);  // ../RTL/cortexm0ds_logic.v(11129)
  and u12524 (Lvkiu6, T9cow6, Aacow6);  // ../RTL/cortexm0ds_logic.v(11130)
  and u12525 (Aacow6, Hacow6, Oacow6);  // ../RTL/cortexm0ds_logic.v(11131)
  or u12526 (Oacow6, Vacow6, Q88ow6);  // ../RTL/cortexm0ds_logic.v(11132)
  and u12527 (n3439, Cbcow6, V78ow6);  // ../RTL/cortexm0ds_logic.v(11133)
  not u12528 (Hacow6, n3439);  // ../RTL/cortexm0ds_logic.v(11133)
  and u12529 (T9cow6, Jbcow6, Qbcow6);  // ../RTL/cortexm0ds_logic.v(11134)
  and u1253 (n81, Mdhpw6[3], Agyhu6);  // ../RTL/cortexm0ds_logic.v(3323)
  and u12530 (n3440, Xbcow6, X88ow6);  // ../RTL/cortexm0ds_logic.v(11135)
  not u12531 (Qbcow6, n3440);  // ../RTL/cortexm0ds_logic.v(11135)
  or u12532 (Jbcow6, H78ow6, Eccow6);  // ../RTL/cortexm0ds_logic.v(11136)
  and u12533 (n3441, Egziu6, Eafpw6[23]);  // ../RTL/cortexm0ds_logic.v(11137)
  not u12534 (F9cow6, n3441);  // ../RTL/cortexm0ds_logic.v(11137)
  and u12535 (D8cow6, Lccow6, Sccow6);  // ../RTL/cortexm0ds_logic.v(11138)
  and u12536 (n3442, vis_pc_o[22], Jmziu6);  // ../RTL/cortexm0ds_logic.v(11139)
  not u12537 (Sccow6, n3442);  // ../RTL/cortexm0ds_logic.v(11139)
  and u12538 (n3443, Zccow6, Gdcow6);  // ../RTL/cortexm0ds_logic.v(11140)
  not u12539 (Koohu6, n3443);  // ../RTL/cortexm0ds_logic.v(11140)
  not u1254 (Lhzhu6, n81);  // ../RTL/cortexm0ds_logic.v(3323)
  and u12540 (Gdcow6, Ndcow6, Udcow6);  // ../RTL/cortexm0ds_logic.v(11141)
  and u12541 (n3444, Egziu6, Eafpw6[27]);  // ../RTL/cortexm0ds_logic.v(11142)
  not u12542 (Udcow6, n3444);  // ../RTL/cortexm0ds_logic.v(11142)
  and u12543 (Ndcow6, Becow6, Sgziu6);  // ../RTL/cortexm0ds_logic.v(11143)
  and u12544 (n3445, Zgziu6, I4liu6);  // ../RTL/cortexm0ds_logic.v(11144)
  not u12545 (Becow6, n3445);  // ../RTL/cortexm0ds_logic.v(11144)
  and u12546 (n3446, Iecow6, Pecow6);  // ../RTL/cortexm0ds_logic.v(11145)
  not u12547 (I4liu6, n3446);  // ../RTL/cortexm0ds_logic.v(11145)
  and u12548 (Pecow6, Wecow6, Dfcow6);  // ../RTL/cortexm0ds_logic.v(11146)
  or u12549 (Dfcow6, Iiziu6, Kfcow6);  // ../RTL/cortexm0ds_logic.v(11147)
  and u1255 (Ehzhu6, Shzhu6, Ftyhu6);  // ../RTL/cortexm0ds_logic.v(3324)
  and u12550 (Wecow6, Rfcow6, Djziu6);  // ../RTL/cortexm0ds_logic.v(11148)
  or u12551 (Rfcow6, Kjziu6, Yfcow6);  // ../RTL/cortexm0ds_logic.v(11149)
  and u12552 (Iecow6, Fgcow6, Mgcow6);  // ../RTL/cortexm0ds_logic.v(11150)
  or u12553 (Mgcow6, Mkziu6, Tgcow6);  // ../RTL/cortexm0ds_logic.v(11151)
  or u12554 (Fgcow6, Ahcow6, Hlziu6);  // ../RTL/cortexm0ds_logic.v(11152)
  and u12555 (Zccow6, Hhcow6, Ohcow6);  // ../RTL/cortexm0ds_logic.v(11153)
  and u12556 (n3447, Zsfpw6[26], Cmziu6);  // ../RTL/cortexm0ds_logic.v(11154)
  not u12557 (Ohcow6, n3447);  // ../RTL/cortexm0ds_logic.v(11154)
  and u12558 (n3448, vis_pc_o[26], Jmziu6);  // ../RTL/cortexm0ds_logic.v(11155)
  not u12559 (Hhcow6, n3448);  // ../RTL/cortexm0ds_logic.v(11155)
  and u1256 (Ysyhu6, Zhzhu6, Ighpw6[2]);  // ../RTL/cortexm0ds_logic.v(3325)
  and u12560 (n3449, Vhcow6, Cicow6);  // ../RTL/cortexm0ds_logic.v(11156)
  not u12561 (Doohu6, n3449);  // ../RTL/cortexm0ds_logic.v(11156)
  and u12562 (Cicow6, Jicow6, Qicow6);  // ../RTL/cortexm0ds_logic.v(11157)
  and u12563 (n3450, Egziu6, Eafpw6[26]);  // ../RTL/cortexm0ds_logic.v(11158)
  not u12564 (Qicow6, n3450);  // ../RTL/cortexm0ds_logic.v(11158)
  and u12565 (Jicow6, Xicow6, Sgziu6);  // ../RTL/cortexm0ds_logic.v(11159)
  and u12566 (n3451, Zgziu6, Q1liu6);  // ../RTL/cortexm0ds_logic.v(11160)
  not u12567 (Xicow6, n3451);  // ../RTL/cortexm0ds_logic.v(11160)
  and u12568 (n3452, Ejcow6, Ljcow6);  // ../RTL/cortexm0ds_logic.v(11161)
  not u12569 (Q1liu6, n3452);  // ../RTL/cortexm0ds_logic.v(11161)
  not u1257 (Ftyhu6, Ysyhu6);  // ../RTL/cortexm0ds_logic.v(3325)
  and u12570 (Ljcow6, Sjcow6, Zjcow6);  // ../RTL/cortexm0ds_logic.v(11162)
  or u12571 (Zjcow6, Iiziu6, Gkcow6);  // ../RTL/cortexm0ds_logic.v(11163)
  and u12572 (Sjcow6, Nkcow6, Djziu6);  // ../RTL/cortexm0ds_logic.v(11165)
  or u12573 (Nkcow6, Kjziu6, Ukcow6);  // ../RTL/cortexm0ds_logic.v(11166)
  not u12574 (Kjziu6, Rc8ow6);  // ../RTL/cortexm0ds_logic.v(11167)
  and u12575 (Ejcow6, Blcow6, Ilcow6);  // ../RTL/cortexm0ds_logic.v(11168)
  or u12576 (Ilcow6, Mkziu6, Plcow6);  // ../RTL/cortexm0ds_logic.v(11169)
  or u12577 (Blcow6, Hlziu6, Wlcow6);  // ../RTL/cortexm0ds_logic.v(11170)
  and u12578 (Vhcow6, Dmcow6, Kmcow6);  // ../RTL/cortexm0ds_logic.v(11171)
  and u12579 (n3453, Zsfpw6[25], Cmziu6);  // ../RTL/cortexm0ds_logic.v(11172)
  or u1258 (n82, Deyhu6, Ighpw6[4]);  // ../RTL/cortexm0ds_logic.v(3326)
  not u12580 (Kmcow6, n3453);  // ../RTL/cortexm0ds_logic.v(11172)
  and u12581 (n3454, vis_pc_o[25], Jmziu6);  // ../RTL/cortexm0ds_logic.v(11173)
  not u12582 (Dmcow6, n3454);  // ../RTL/cortexm0ds_logic.v(11173)
  and u12583 (n3455, Rmcow6, Ymcow6);  // ../RTL/cortexm0ds_logic.v(11174)
  not u12584 (Wnohu6, n3455);  // ../RTL/cortexm0ds_logic.v(11174)
  and u12585 (Ymcow6, Fncow6, Mncow6);  // ../RTL/cortexm0ds_logic.v(11175)
  and u12586 (n3456, Egziu6, Eafpw6[25]);  // ../RTL/cortexm0ds_logic.v(11176)
  not u12587 (Mncow6, n3456);  // ../RTL/cortexm0ds_logic.v(11176)
  and u12588 (Fncow6, Tncow6, Sgziu6);  // ../RTL/cortexm0ds_logic.v(11177)
  and u12589 (n3457, Zgziu6, Osliu6);  // ../RTL/cortexm0ds_logic.v(11178)
  not u1259 (Zhzhu6, n82);  // ../RTL/cortexm0ds_logic.v(3326)
  not u12590 (Tncow6, n3457);  // ../RTL/cortexm0ds_logic.v(11178)
  and u12591 (n3458, Aocow6, Hocow6);  // ../RTL/cortexm0ds_logic.v(11179)
  not u12592 (Osliu6, n3458);  // ../RTL/cortexm0ds_logic.v(11179)
  and u12593 (Hocow6, Oocow6, Vocow6);  // ../RTL/cortexm0ds_logic.v(11180)
  and u12594 (n3459, Dc8ow6, Ew6ow6);  // ../RTL/cortexm0ds_logic.v(11181)
  not u12595 (Vocow6, n3459);  // ../RTL/cortexm0ds_logic.v(11181)
  and u12596 (Oocow6, Cpcow6, Djziu6);  // ../RTL/cortexm0ds_logic.v(11182)
  and u12597 (n3460, Rc8ow6, Cv6ow6);  // ../RTL/cortexm0ds_logic.v(11183)
  not u12598 (Cpcow6, n3460);  // ../RTL/cortexm0ds_logic.v(11183)
  and u12599 (Aocow6, Jpcow6, Qpcow6);  // ../RTL/cortexm0ds_logic.v(11184)
  buf u126 (Iqnhu6, Gnqpw6);  // ../RTL/cortexm0ds_logic.v(1935)
  and u1260 (n83, Iyyhu6, Gizhu6);  // ../RTL/cortexm0ds_logic.v(3327)
  or u12600 (Qpcow6, Mkziu6, Xv6ow6);  // ../RTL/cortexm0ds_logic.v(11185)
  or u12601 (Jpcow6, Ou6ow6, Hlziu6);  // ../RTL/cortexm0ds_logic.v(11186)
  and u12602 (Rmcow6, Xpcow6, Eqcow6);  // ../RTL/cortexm0ds_logic.v(11187)
  and u12603 (n3461, Zsfpw6[24], Cmziu6);  // ../RTL/cortexm0ds_logic.v(11188)
  not u12604 (Eqcow6, n3461);  // ../RTL/cortexm0ds_logic.v(11188)
  and u12605 (n3462, vis_pc_o[24], Jmziu6);  // ../RTL/cortexm0ds_logic.v(11189)
  not u12606 (Xpcow6, n3462);  // ../RTL/cortexm0ds_logic.v(11189)
  and u12607 (n3463, Lqcow6, Sqcow6);  // ../RTL/cortexm0ds_logic.v(11190)
  not u12608 (Pnohu6, n3463);  // ../RTL/cortexm0ds_logic.v(11190)
  and u12609 (Sqcow6, Zqcow6, Grcow6);  // ../RTL/cortexm0ds_logic.v(11191)
  not u1261 (Shzhu6, n83);  // ../RTL/cortexm0ds_logic.v(3327)
  and u12610 (n3464, Egziu6, Eafpw6[24]);  // ../RTL/cortexm0ds_logic.v(11192)
  not u12611 (Grcow6, n3464);  // ../RTL/cortexm0ds_logic.v(11192)
  and u12612 (Zqcow6, Nrcow6, Sgziu6);  // ../RTL/cortexm0ds_logic.v(11193)
  and u12613 (n3465, Zgziu6, Nu8iu6);  // ../RTL/cortexm0ds_logic.v(11194)
  not u12614 (Nrcow6, n3465);  // ../RTL/cortexm0ds_logic.v(11194)
  and u12615 (n3466, Urcow6, Bscow6);  // ../RTL/cortexm0ds_logic.v(11195)
  not u12616 (Nu8iu6, n3466);  // ../RTL/cortexm0ds_logic.v(11195)
  and u12617 (Bscow6, Iscow6, Pscow6);  // ../RTL/cortexm0ds_logic.v(11196)
  and u12618 (n3467, Dc8ow6, Tdliu6);  // ../RTL/cortexm0ds_logic.v(11197)
  not u12619 (Pscow6, n3467);  // ../RTL/cortexm0ds_logic.v(11197)
  and u1262 (n84, Deyhu6, Nizhu6);  // ../RTL/cortexm0ds_logic.v(3328)
  and u12620 (Iiziu6, Wscow6, Dtcow6);  // ../RTL/cortexm0ds_logic.v(11198)
  not u12621 (Dc8ow6, Iiziu6);  // ../RTL/cortexm0ds_logic.v(11198)
  or u12622 (Wscow6, Ah3ju6, Ktcow6);  // ../RTL/cortexm0ds_logic.v(11199)
  and u12623 (Iscow6, Rtcow6, Djziu6);  // ../RTL/cortexm0ds_logic.v(11200)
  and u12624 (n3468, Ytcow6, Fucow6);  // ../RTL/cortexm0ds_logic.v(11201)
  not u12625 (Djziu6, n3468);  // ../RTL/cortexm0ds_logic.v(11201)
  and u12626 (n3469, Mucow6, Tucow6);  // ../RTL/cortexm0ds_logic.v(11202)
  not u12627 (Fucow6, n3469);  // ../RTL/cortexm0ds_logic.v(11202)
  and u12628 (n3470, Fg3ju6, Ah3ju6);  // ../RTL/cortexm0ds_logic.v(11203)
  not u12629 (Mucow6, n3470);  // ../RTL/cortexm0ds_logic.v(11203)
  not u1263 (Gizhu6, n84);  // ../RTL/cortexm0ds_logic.v(3328)
  or u12630 (Ah3ju6, Avcow6, Df3ju6);  // ../RTL/cortexm0ds_logic.v(11204)
  and u12631 (n3471, Rc8ow6, Jfliu6);  // ../RTL/cortexm0ds_logic.v(11205)
  not u12632 (Rtcow6, n3471);  // ../RTL/cortexm0ds_logic.v(11205)
  or u12633 (Rc8ow6, Hvcow6, Ovcow6);  // ../RTL/cortexm0ds_logic.v(11206)
  or u12634 (n3472, Fg3ju6, Ktcow6);  // ../RTL/cortexm0ds_logic.v(11207)
  not u12635 (Hvcow6, n3472);  // ../RTL/cortexm0ds_logic.v(11207)
  and u12636 (Urcow6, Vvcow6, Cwcow6);  // ../RTL/cortexm0ds_logic.v(11208)
  or u12637 (Cwcow6, Mkziu6, Rcliu6);  // ../RTL/cortexm0ds_logic.v(11209)
  or u12638 (Vvcow6, Veliu6, Hlziu6);  // ../RTL/cortexm0ds_logic.v(11210)
  and u12639 (Lqcow6, Jwcow6, Qwcow6);  // ../RTL/cortexm0ds_logic.v(11211)
  or u1264 (Nizhu6, C9zhu6, Mdhpw6[3]);  // ../RTL/cortexm0ds_logic.v(3329)
  and u12640 (n3473, Zsfpw6[23], Cmziu6);  // ../RTL/cortexm0ds_logic.v(11212)
  not u12641 (Qwcow6, n3473);  // ../RTL/cortexm0ds_logic.v(11212)
  and u12642 (n3474, vis_pc_o[23], Jmziu6);  // ../RTL/cortexm0ds_logic.v(11213)
  not u12643 (Jwcow6, n3474);  // ../RTL/cortexm0ds_logic.v(11213)
  and u12644 (n3475, Xwcow6, Excow6);  // ../RTL/cortexm0ds_logic.v(11214)
  not u12645 (Inohu6, n3475);  // ../RTL/cortexm0ds_logic.v(11214)
  and u12646 (Excow6, Lxcow6, Sxcow6);  // ../RTL/cortexm0ds_logic.v(11215)
  and u12647 (n3476, Zsfpw6[20], Cmziu6);  // ../RTL/cortexm0ds_logic.v(11216)
  not u12648 (Sxcow6, n3476);  // ../RTL/cortexm0ds_logic.v(11216)
  and u12649 (Lxcow6, Zxcow6, Gycow6);  // ../RTL/cortexm0ds_logic.v(11217)
  and u1265 (Xgzhu6, Uizhu6, Bjzhu6);  // ../RTL/cortexm0ds_logic.v(3330)
  or u12650 (Gycow6, Ft6ow6, Tyliu6);  // ../RTL/cortexm0ds_logic.v(11218)
  and u12651 (Tyliu6, Nycow6, Uycow6);  // ../RTL/cortexm0ds_logic.v(11219)
  and u12652 (Uycow6, Bzcow6, Izcow6);  // ../RTL/cortexm0ds_logic.v(11220)
  or u12653 (Izcow6, Tkziu6, Vacow6);  // ../RTL/cortexm0ds_logic.v(11221)
  or u12654 (Bzcow6, Rjziu6, Pzcow6);  // ../RTL/cortexm0ds_logic.v(11222)
  and u12655 (Nycow6, Wzcow6, D0dow6);  // ../RTL/cortexm0ds_logic.v(11223)
  or u12656 (D0dow6, Alziu6, Eccow6);  // ../RTL/cortexm0ds_logic.v(11224)
  or u12657 (Wzcow6, Mkziu6, Piziu6);  // ../RTL/cortexm0ds_logic.v(11225)
  and u12658 (n3477, Egziu6, Eafpw6[21]);  // ../RTL/cortexm0ds_logic.v(11226)
  not u12659 (Zxcow6, n3477);  // ../RTL/cortexm0ds_logic.v(11226)
  and u1266 (n85, Swyhu6, Zazhu6);  // ../RTL/cortexm0ds_logic.v(3331)
  and u12660 (Xwcow6, Lccow6, K0dow6);  // ../RTL/cortexm0ds_logic.v(11227)
  and u12661 (n3478, vis_pc_o[20], Jmziu6);  // ../RTL/cortexm0ds_logic.v(11228)
  not u12662 (K0dow6, n3478);  // ../RTL/cortexm0ds_logic.v(11228)
  and u12663 (n3479, R0dow6, Y0dow6);  // ../RTL/cortexm0ds_logic.v(11229)
  not u12664 (Bnohu6, n3479);  // ../RTL/cortexm0ds_logic.v(11229)
  and u12665 (Y0dow6, F1dow6, M1dow6);  // ../RTL/cortexm0ds_logic.v(11230)
  and u12666 (n3480, Zsfpw6[19], Cmziu6);  // ../RTL/cortexm0ds_logic.v(11231)
  not u12667 (M1dow6, n3480);  // ../RTL/cortexm0ds_logic.v(11231)
  and u12668 (F1dow6, T1dow6, A2dow6);  // ../RTL/cortexm0ds_logic.v(11232)
  or u12669 (A2dow6, Ft6ow6, S1miu6);  // ../RTL/cortexm0ds_logic.v(11233)
  not u1267 (Bjzhu6, n85);  // ../RTL/cortexm0ds_logic.v(3331)
  and u12670 (S1miu6, H2dow6, O2dow6);  // ../RTL/cortexm0ds_logic.v(11234)
  and u12671 (O2dow6, V2dow6, C3dow6);  // ../RTL/cortexm0ds_logic.v(11235)
  or u12672 (C3dow6, P0cow6, Pzcow6);  // ../RTL/cortexm0ds_logic.v(11236)
  or u12673 (V2dow6, K1cow6, Eccow6);  // ../RTL/cortexm0ds_logic.v(11237)
  and u12674 (H2dow6, J3dow6, Q3dow6);  // ../RTL/cortexm0ds_logic.v(11238)
  or u12675 (Q3dow6, R1cow6, Vacow6);  // ../RTL/cortexm0ds_logic.v(11239)
  or u12676 (J3dow6, Mkziu6, B0cow6);  // ../RTL/cortexm0ds_logic.v(11240)
  and u12677 (n3481, Egziu6, Eafpw6[20]);  // ../RTL/cortexm0ds_logic.v(11241)
  not u12678 (T1dow6, n3481);  // ../RTL/cortexm0ds_logic.v(11241)
  and u12679 (R0dow6, Lccow6, X3dow6);  // ../RTL/cortexm0ds_logic.v(11242)
  and u1268 (Swyhu6, Ijzhu6, Ighpw6[2]);  // ../RTL/cortexm0ds_logic.v(3332)
  and u12680 (n3482, vis_pc_o[19], Jmziu6);  // ../RTL/cortexm0ds_logic.v(11243)
  not u12681 (X3dow6, n3482);  // ../RTL/cortexm0ds_logic.v(11243)
  and u12682 (n3483, E4dow6, L4dow6);  // ../RTL/cortexm0ds_logic.v(11244)
  not u12683 (Umohu6, n3483);  // ../RTL/cortexm0ds_logic.v(11244)
  and u12684 (L4dow6, S4dow6, Z4dow6);  // ../RTL/cortexm0ds_logic.v(11245)
  and u12685 (n3484, Zsfpw6[18], Cmziu6);  // ../RTL/cortexm0ds_logic.v(11246)
  not u12686 (Z4dow6, n3484);  // ../RTL/cortexm0ds_logic.v(11246)
  and u12687 (S4dow6, G5dow6, N5dow6);  // ../RTL/cortexm0ds_logic.v(11247)
  or u12688 (N5dow6, Ft6ow6, R4miu6);  // ../RTL/cortexm0ds_logic.v(11248)
  and u12689 (R4miu6, U5dow6, B6dow6);  // ../RTL/cortexm0ds_logic.v(11249)
  and u1269 (n86, Mdhpw6[3], Pjzhu6);  // ../RTL/cortexm0ds_logic.v(3333)
  and u12690 (B6dow6, I6dow6, P6dow6);  // ../RTL/cortexm0ds_logic.v(11250)
  or u12691 (P6dow6, Mkziu6, Kfcow6);  // ../RTL/cortexm0ds_logic.v(11251)
  or u12692 (I6dow6, Tgcow6, Vacow6);  // ../RTL/cortexm0ds_logic.v(11252)
  and u12693 (U5dow6, W6dow6, D7dow6);  // ../RTL/cortexm0ds_logic.v(11253)
  or u12694 (D7dow6, Ahcow6, Eccow6);  // ../RTL/cortexm0ds_logic.v(11254)
  or u12695 (W6dow6, Yfcow6, Pzcow6);  // ../RTL/cortexm0ds_logic.v(11255)
  and u12696 (n3485, Egziu6, Eafpw6[19]);  // ../RTL/cortexm0ds_logic.v(11256)
  not u12697 (G5dow6, n3485);  // ../RTL/cortexm0ds_logic.v(11256)
  and u12698 (E4dow6, Lccow6, K7dow6);  // ../RTL/cortexm0ds_logic.v(11257)
  and u12699 (n3486, vis_pc_o[18], Jmziu6);  // ../RTL/cortexm0ds_logic.v(11258)
  buf u127 (Vbgpw6[29], Kojpw6);  // ../RTL/cortexm0ds_logic.v(3092)
  not u1270 (Uizhu6, n86);  // ../RTL/cortexm0ds_logic.v(3333)
  not u12700 (K7dow6, n3486);  // ../RTL/cortexm0ds_logic.v(11258)
  and u12701 (n3487, R7dow6, Y7dow6);  // ../RTL/cortexm0ds_logic.v(11259)
  not u12702 (Nmohu6, n3487);  // ../RTL/cortexm0ds_logic.v(11259)
  and u12703 (Y7dow6, F8dow6, M8dow6);  // ../RTL/cortexm0ds_logic.v(11260)
  and u12704 (n3488, Zsfpw6[17], Cmziu6);  // ../RTL/cortexm0ds_logic.v(11261)
  not u12705 (M8dow6, n3488);  // ../RTL/cortexm0ds_logic.v(11261)
  and u12706 (F8dow6, T8dow6, A9dow6);  // ../RTL/cortexm0ds_logic.v(11262)
  or u12707 (A9dow6, Ft6ow6, Q7miu6);  // ../RTL/cortexm0ds_logic.v(11263)
  and u12708 (Q7miu6, H9dow6, O9dow6);  // ../RTL/cortexm0ds_logic.v(11264)
  and u12709 (O9dow6, V9dow6, Cadow6);  // ../RTL/cortexm0ds_logic.v(11265)
  and u1271 (n87, Wjzhu6, Dkzhu6);  // ../RTL/cortexm0ds_logic.v(3334)
  or u12710 (Cadow6, Vacow6, Plcow6);  // ../RTL/cortexm0ds_logic.v(11266)
  or u12711 (V9dow6, Pzcow6, Ukcow6);  // ../RTL/cortexm0ds_logic.v(11267)
  and u12712 (H9dow6, Jadow6, Qadow6);  // ../RTL/cortexm0ds_logic.v(11269)
  or u12713 (Qadow6, Mkziu6, Gkcow6);  // ../RTL/cortexm0ds_logic.v(11270)
  or u12714 (Jadow6, Eccow6, Wlcow6);  // ../RTL/cortexm0ds_logic.v(11272)
  and u12715 (n3489, Egziu6, Eafpw6[18]);  // ../RTL/cortexm0ds_logic.v(11273)
  not u12716 (T8dow6, n3489);  // ../RTL/cortexm0ds_logic.v(11273)
  and u12717 (R7dow6, Lccow6, Xadow6);  // ../RTL/cortexm0ds_logic.v(11274)
  and u12718 (n3490, vis_pc_o[17], Jmziu6);  // ../RTL/cortexm0ds_logic.v(11275)
  not u12719 (Xadow6, n3490);  // ../RTL/cortexm0ds_logic.v(11275)
  not u1272 (Pjzhu6, n87);  // ../RTL/cortexm0ds_logic.v(3334)
  and u12720 (n3491, Ebdow6, Lbdow6);  // ../RTL/cortexm0ds_logic.v(11276)
  not u12721 (Gmohu6, n3491);  // ../RTL/cortexm0ds_logic.v(11276)
  and u12722 (Lbdow6, Sbdow6, Zbdow6);  // ../RTL/cortexm0ds_logic.v(11277)
  and u12723 (n3492, Zsfpw6[16], Cmziu6);  // ../RTL/cortexm0ds_logic.v(11278)
  not u12724 (Zbdow6, n3492);  // ../RTL/cortexm0ds_logic.v(11278)
  and u12725 (Sbdow6, Gcdow6, Ncdow6);  // ../RTL/cortexm0ds_logic.v(11279)
  or u12726 (Ncdow6, Ft6ow6, Pamiu6);  // ../RTL/cortexm0ds_logic.v(11280)
  and u12727 (Pamiu6, Ucdow6, Bddow6);  // ../RTL/cortexm0ds_logic.v(11281)
  and u12728 (Bddow6, Iddow6, Pddow6);  // ../RTL/cortexm0ds_logic.v(11282)
  and u12729 (n3493, Xbcow6, Ew6ow6);  // ../RTL/cortexm0ds_logic.v(11283)
  or u1273 (n88, Kkzhu6, Hgyhu6);  // ../RTL/cortexm0ds_logic.v(3335)
  not u12730 (Pddow6, n3493);  // ../RTL/cortexm0ds_logic.v(11283)
  or u12731 (Iddow6, Xv6ow6, Vacow6);  // ../RTL/cortexm0ds_logic.v(11284)
  and u12732 (Ucdow6, Wddow6, Dedow6);  // ../RTL/cortexm0ds_logic.v(11285)
  or u12733 (Dedow6, Ou6ow6, Eccow6);  // ../RTL/cortexm0ds_logic.v(11286)
  and u12734 (n3494, Cv6ow6, Cbcow6);  // ../RTL/cortexm0ds_logic.v(11287)
  not u12735 (Wddow6, n3494);  // ../RTL/cortexm0ds_logic.v(11287)
  and u12736 (n3495, Egziu6, Eafpw6[17]);  // ../RTL/cortexm0ds_logic.v(11288)
  not u12737 (Gcdow6, n3495);  // ../RTL/cortexm0ds_logic.v(11288)
  and u12738 (Ebdow6, Lccow6, Kedow6);  // ../RTL/cortexm0ds_logic.v(11289)
  and u12739 (n3496, vis_pc_o[16], Jmziu6);  // ../RTL/cortexm0ds_logic.v(11290)
  not u1274 (Dkzhu6, n88);  // ../RTL/cortexm0ds_logic.v(3335)
  not u12740 (Kedow6, n3496);  // ../RTL/cortexm0ds_logic.v(11290)
  and u12741 (n3497, Redow6, Yedow6);  // ../RTL/cortexm0ds_logic.v(11291)
  not u12742 (Zlohu6, n3497);  // ../RTL/cortexm0ds_logic.v(11291)
  and u12743 (Yedow6, Ffdow6, Mfdow6);  // ../RTL/cortexm0ds_logic.v(11292)
  and u12744 (n3498, Zsfpw6[15], Cmziu6);  // ../RTL/cortexm0ds_logic.v(11293)
  not u12745 (Mfdow6, n3498);  // ../RTL/cortexm0ds_logic.v(11293)
  and u12746 (Ffdow6, Tfdow6, Agdow6);  // ../RTL/cortexm0ds_logic.v(11294)
  or u12747 (Agdow6, Ft6ow6, Odmiu6);  // ../RTL/cortexm0ds_logic.v(11295)
  and u12748 (Odmiu6, Hgdow6, Ogdow6);  // ../RTL/cortexm0ds_logic.v(11296)
  and u12749 (Ogdow6, Vgdow6, Chdow6);  // ../RTL/cortexm0ds_logic.v(11297)
  and u1275 (Hgyhu6, Rkzhu6, Zazhu6);  // ../RTL/cortexm0ds_logic.v(3336)
  and u12750 (n3499, Xbcow6, Tdliu6);  // ../RTL/cortexm0ds_logic.v(11298)
  not u12751 (Chdow6, n3499);  // ../RTL/cortexm0ds_logic.v(11298)
  or u12752 (Vgdow6, Rcliu6, Vacow6);  // ../RTL/cortexm0ds_logic.v(11299)
  and u12753 (Hgdow6, Jhdow6, Qhdow6);  // ../RTL/cortexm0ds_logic.v(11300)
  or u12754 (Qhdow6, Veliu6, Eccow6);  // ../RTL/cortexm0ds_logic.v(11301)
  and u12755 (n3500, Jfliu6, Cbcow6);  // ../RTL/cortexm0ds_logic.v(11302)
  not u12756 (Jhdow6, n3500);  // ../RTL/cortexm0ds_logic.v(11302)
  and u12757 (n3501, Egziu6, Eafpw6[16]);  // ../RTL/cortexm0ds_logic.v(11303)
  not u12758 (Tfdow6, n3501);  // ../RTL/cortexm0ds_logic.v(11303)
  and u12759 (Redow6, Lccow6, Xhdow6);  // ../RTL/cortexm0ds_logic.v(11304)
  and u1276 (n89, Tfyhu6, Wryhu6);  // ../RTL/cortexm0ds_logic.v(3337)
  and u12760 (n3502, vis_pc_o[15], Jmziu6);  // ../RTL/cortexm0ds_logic.v(11305)
  not u12761 (Xhdow6, n3502);  // ../RTL/cortexm0ds_logic.v(11305)
  and u12762 (n3503, Eidow6, Lidow6);  // ../RTL/cortexm0ds_logic.v(11306)
  not u12763 (Slohu6, n3503);  // ../RTL/cortexm0ds_logic.v(11306)
  and u12764 (Lidow6, Sidow6, Zidow6);  // ../RTL/cortexm0ds_logic.v(11307)
  and u12765 (n3504, Egziu6, Eafpw6[14]);  // ../RTL/cortexm0ds_logic.v(11308)
  not u12766 (Zidow6, n3504);  // ../RTL/cortexm0ds_logic.v(11308)
  and u12767 (Sidow6, Gjdow6, Sgziu6);  // ../RTL/cortexm0ds_logic.v(11309)
  and u12768 (n3505, Zgziu6, Yimiu6);  // ../RTL/cortexm0ds_logic.v(11310)
  not u12769 (Gjdow6, n3505);  // ../RTL/cortexm0ds_logic.v(11310)
  not u1277 (Kkzhu6, n89);  // ../RTL/cortexm0ds_logic.v(3337)
  and u12770 (n3506, Njdow6, Ujdow6);  // ../RTL/cortexm0ds_logic.v(11311)
  not u12771 (Yimiu6, n3506);  // ../RTL/cortexm0ds_logic.v(11311)
  and u12772 (Ujdow6, Bkdow6, Ikdow6);  // ../RTL/cortexm0ds_logic.v(11312)
  or u12773 (Ikdow6, L5cow6, Pkdow6);  // ../RTL/cortexm0ds_logic.v(11313)
  and u12774 (Bkdow6, Wkdow6, Dldow6);  // ../RTL/cortexm0ds_logic.v(11314)
  or u12775 (Wkdow6, G6cow6, Kldow6);  // ../RTL/cortexm0ds_logic.v(11315)
  and u12776 (Njdow6, Rldow6, Yldow6);  // ../RTL/cortexm0ds_logic.v(11316)
  and u12777 (n3507, X4cow6, Fmdow6);  // ../RTL/cortexm0ds_logic.v(11317)
  not u12778 (Yldow6, n3507);  // ../RTL/cortexm0ds_logic.v(11317)
  and u12779 (n3508, N6cow6, Mmdow6);  // ../RTL/cortexm0ds_logic.v(11318)
  and u1278 (n90, Ykzhu6, Epyhu6);  // ../RTL/cortexm0ds_logic.v(3338)
  not u12780 (Rldow6, n3508);  // ../RTL/cortexm0ds_logic.v(11318)
  and u12781 (Eidow6, Tmdow6, Andow6);  // ../RTL/cortexm0ds_logic.v(11319)
  and u12782 (n3509, Zsfpw6[13], Cmziu6);  // ../RTL/cortexm0ds_logic.v(11320)
  not u12783 (Andow6, n3509);  // ../RTL/cortexm0ds_logic.v(11320)
  and u12784 (n3510, vis_pc_o[13], Jmziu6);  // ../RTL/cortexm0ds_logic.v(11321)
  not u12785 (Tmdow6, n3510);  // ../RTL/cortexm0ds_logic.v(11321)
  and u12786 (n3511, Hndow6, Ondow6);  // ../RTL/cortexm0ds_logic.v(11322)
  not u12787 (Llohu6, n3511);  // ../RTL/cortexm0ds_logic.v(11322)
  and u12788 (Ondow6, Vndow6, Codow6);  // ../RTL/cortexm0ds_logic.v(11323)
  and u12789 (n3512, Egziu6, Eafpw6[13]);  // ../RTL/cortexm0ds_logic.v(11324)
  not u1279 (Wryhu6, n90);  // ../RTL/cortexm0ds_logic.v(3338)
  not u12790 (Codow6, n3512);  // ../RTL/cortexm0ds_logic.v(11324)
  and u12791 (Vndow6, Jodow6, Sgziu6);  // ../RTL/cortexm0ds_logic.v(11325)
  and u12792 (n3513, Zgziu6, Qlmiu6);  // ../RTL/cortexm0ds_logic.v(11326)
  not u12793 (Jodow6, n3513);  // ../RTL/cortexm0ds_logic.v(11326)
  and u12794 (n3514, Qodow6, Xodow6);  // ../RTL/cortexm0ds_logic.v(11327)
  not u12795 (Qlmiu6, n3514);  // ../RTL/cortexm0ds_logic.v(11327)
  and u12796 (Xodow6, Epdow6, Lpdow6);  // ../RTL/cortexm0ds_logic.v(11328)
  or u12797 (Lpdow6, Rjziu6, Spdow6);  // ../RTL/cortexm0ds_logic.v(11329)
  and u12798 (Epdow6, Zpdow6, Dldow6);  // ../RTL/cortexm0ds_logic.v(11330)
  or u12799 (Zpdow6, Tkziu6, Pkdow6);  // ../RTL/cortexm0ds_logic.v(11331)
  buf u128 (Vbgpw6[28], Usipw6);  // ../RTL/cortexm0ds_logic.v(3092)
  or u1280 (n91, Vuyhu6, Deyhu6);  // ../RTL/cortexm0ds_logic.v(3339)
  and u12800 (Qodow6, Gqdow6, Nqdow6);  // ../RTL/cortexm0ds_logic.v(11332)
  or u12801 (Nqdow6, Alziu6, Kldow6);  // ../RTL/cortexm0ds_logic.v(11333)
  or u12802 (Gqdow6, Piziu6, Uqdow6);  // ../RTL/cortexm0ds_logic.v(11334)
  and u12803 (Hndow6, Brdow6, Irdow6);  // ../RTL/cortexm0ds_logic.v(11335)
  and u12804 (n3515, Zsfpw6[12], Cmziu6);  // ../RTL/cortexm0ds_logic.v(11336)
  not u12805 (Irdow6, n3515);  // ../RTL/cortexm0ds_logic.v(11336)
  and u12806 (n3516, vis_pc_o[12], Jmziu6);  // ../RTL/cortexm0ds_logic.v(11337)
  not u12807 (Brdow6, n3516);  // ../RTL/cortexm0ds_logic.v(11337)
  and u12808 (n3517, Prdow6, Wrdow6);  // ../RTL/cortexm0ds_logic.v(11338)
  not u12809 (Elohu6, n3517);  // ../RTL/cortexm0ds_logic.v(11338)
  not u1281 (Ykzhu6, n91);  // ../RTL/cortexm0ds_logic.v(3339)
  and u12810 (Wrdow6, Dsdow6, Ksdow6);  // ../RTL/cortexm0ds_logic.v(11339)
  and u12811 (n3518, Egziu6, Eafpw6[12]);  // ../RTL/cortexm0ds_logic.v(11340)
  not u12812 (Ksdow6, n3518);  // ../RTL/cortexm0ds_logic.v(11340)
  and u12813 (Dsdow6, Rsdow6, Sgziu6);  // ../RTL/cortexm0ds_logic.v(11341)
  and u12814 (n3519, Zgziu6, Iomiu6);  // ../RTL/cortexm0ds_logic.v(11342)
  not u12815 (Rsdow6, n3519);  // ../RTL/cortexm0ds_logic.v(11342)
  and u12816 (n3520, Ysdow6, Ftdow6);  // ../RTL/cortexm0ds_logic.v(11343)
  not u12817 (Iomiu6, n3520);  // ../RTL/cortexm0ds_logic.v(11343)
  and u12818 (Ftdow6, Mtdow6, Ttdow6);  // ../RTL/cortexm0ds_logic.v(11344)
  or u12819 (Ttdow6, K1cow6, Kldow6);  // ../RTL/cortexm0ds_logic.v(11345)
  and u1282 (n92, Rkzhu6, Ighpw6[0]);  // ../RTL/cortexm0ds_logic.v(3340)
  and u12820 (Mtdow6, Audow6, Dldow6);  // ../RTL/cortexm0ds_logic.v(11346)
  or u12821 (Audow6, P0cow6, Spdow6);  // ../RTL/cortexm0ds_logic.v(11347)
  and u12822 (Ysdow6, Hudow6, Oudow6);  // ../RTL/cortexm0ds_logic.v(11348)
  or u12823 (Oudow6, R1cow6, Pkdow6);  // ../RTL/cortexm0ds_logic.v(11349)
  or u12824 (Hudow6, B0cow6, Uqdow6);  // ../RTL/cortexm0ds_logic.v(11350)
  and u12825 (Prdow6, Vudow6, Cvdow6);  // ../RTL/cortexm0ds_logic.v(11351)
  and u12826 (n3521, Zsfpw6[11], Cmziu6);  // ../RTL/cortexm0ds_logic.v(11352)
  not u12827 (Cvdow6, n3521);  // ../RTL/cortexm0ds_logic.v(11352)
  and u12828 (n3522, vis_pc_o[11], Jmziu6);  // ../RTL/cortexm0ds_logic.v(11353)
  not u12829 (Vudow6, n3522);  // ../RTL/cortexm0ds_logic.v(11353)
  not u1283 (Tfyhu6, n92);  // ../RTL/cortexm0ds_logic.v(3340)
  and u12830 (n3523, Jvdow6, Qvdow6);  // ../RTL/cortexm0ds_logic.v(11354)
  not u12831 (Xkohu6, n3523);  // ../RTL/cortexm0ds_logic.v(11354)
  and u12832 (Qvdow6, Xvdow6, Ewdow6);  // ../RTL/cortexm0ds_logic.v(11355)
  and u12833 (n3524, Egziu6, Eafpw6[8]);  // ../RTL/cortexm0ds_logic.v(11356)
  not u12834 (Ewdow6, n3524);  // ../RTL/cortexm0ds_logic.v(11356)
  and u12835 (Xvdow6, Lwdow6, Sgziu6);  // ../RTL/cortexm0ds_logic.v(11357)
  and u12836 (n3525, Zgziu6, E7niu6);  // ../RTL/cortexm0ds_logic.v(11358)
  not u12837 (Lwdow6, n3525);  // ../RTL/cortexm0ds_logic.v(11358)
  and u12838 (n3526, Swdow6, Zwdow6);  // ../RTL/cortexm0ds_logic.v(11359)
  not u12839 (E7niu6, n3526);  // ../RTL/cortexm0ds_logic.v(11359)
  and u1284 (Rkzhu6, Flzhu6, Epyhu6);  // ../RTL/cortexm0ds_logic.v(3341)
  and u12840 (Zwdow6, Gxdow6, Nxdow6);  // ../RTL/cortexm0ds_logic.v(11360)
  or u12841 (Nxdow6, Rcliu6, Pkdow6);  // ../RTL/cortexm0ds_logic.v(11361)
  and u12842 (Rcliu6, Uxdow6, Bydow6);  // ../RTL/cortexm0ds_logic.v(11362)
  or u12843 (Bydow6, Iydow6, W4siu6);  // ../RTL/cortexm0ds_logic.v(11363)
  and u12844 (W4siu6, Pydow6, Wydow6);  // ../RTL/cortexm0ds_logic.v(11364)
  and u12845 (Wydow6, Dzdow6, Kzdow6);  // ../RTL/cortexm0ds_logic.v(11365)
  and u12846 (n3527, Tzfpw6[8], Yvgiu6);  // ../RTL/cortexm0ds_logic.v(11366)
  not u12847 (Kzdow6, n3527);  // ../RTL/cortexm0ds_logic.v(11366)
  and u12848 (Dzdow6, Rzdow6, Yzdow6);  // ../RTL/cortexm0ds_logic.v(11367)
  and u12849 (n3528, F0eow6, Vbgpw6[8]);  // ../RTL/cortexm0ds_logic.v(11368)
  or u1285 (n93, Vuyhu6, Ighpw6[1]);  // ../RTL/cortexm0ds_logic.v(3342)
  not u12850 (Yzdow6, n3528);  // ../RTL/cortexm0ds_logic.v(11368)
  and u12851 (n3529, M0eow6, Odgpw6[8]);  // ../RTL/cortexm0ds_logic.v(11369)
  not u12852 (Rzdow6, n3529);  // ../RTL/cortexm0ds_logic.v(11369)
  and u12853 (Pydow6, T0eow6, A1eow6);  // ../RTL/cortexm0ds_logic.v(11370)
  and u12854 (n3530, Bagpw6[8], M6eiu6);  // ../RTL/cortexm0ds_logic.v(11371)
  not u12855 (A1eow6, n3530);  // ../RTL/cortexm0ds_logic.v(11371)
  and u12856 (n3531, STCALIB[8], H1eow6);  // ../RTL/cortexm0ds_logic.v(11372)
  not u12857 (T0eow6, n3531);  // ../RTL/cortexm0ds_logic.v(11372)
  and u12858 (Uxdow6, O1eow6, V1eow6);  // ../RTL/cortexm0ds_logic.v(11373)
  and u12859 (n3532, Gk3ju6, C2eow6);  // ../RTL/cortexm0ds_logic.v(11374)
  not u1286 (Flzhu6, n93);  // ../RTL/cortexm0ds_logic.v(3342)
  not u12860 (V1eow6, n3532);  // ../RTL/cortexm0ds_logic.v(11374)
  AL_MUX u12861 (
    .i0(Tf4ju6),
    .i1(Cw3ju6),
    .sel(J2eow6),
    .o(Gk3ju6));  // ../RTL/cortexm0ds_logic.v(11375)
  and u12862 (n3533, HRDATA[8], Q2eow6);  // ../RTL/cortexm0ds_logic.v(11376)
  not u12863 (O1eow6, n3533);  // ../RTL/cortexm0ds_logic.v(11376)
  and u12864 (Gxdow6, X2eow6, Dldow6);  // ../RTL/cortexm0ds_logic.v(11377)
  and u12865 (n3534, Tdliu6, Mmdow6);  // ../RTL/cortexm0ds_logic.v(11378)
  not u12866 (X2eow6, n3534);  // ../RTL/cortexm0ds_logic.v(11378)
  and u12867 (n3535, E3eow6, L3eow6);  // ../RTL/cortexm0ds_logic.v(11379)
  not u12868 (Tdliu6, n3535);  // ../RTL/cortexm0ds_logic.v(11379)
  or u12869 (L3eow6, Iydow6, M1xiu6);  // ../RTL/cortexm0ds_logic.v(11380)
  and u1287 (Wjzhu6, Mlzhu6, Tlzhu6);  // ../RTL/cortexm0ds_logic.v(3343)
  and u12870 (M1xiu6, S3eow6, Z3eow6);  // ../RTL/cortexm0ds_logic.v(11381)
  and u12871 (Z3eow6, G4eow6, N4eow6);  // ../RTL/cortexm0ds_logic.v(11382)
  and u12872 (N4eow6, U4eow6, B5eow6);  // ../RTL/cortexm0ds_logic.v(11383)
  and u12873 (n3536, STCALIB[0], H1eow6);  // ../RTL/cortexm0ds_logic.v(11384)
  not u12874 (B5eow6, n3536);  // ../RTL/cortexm0ds_logic.v(11384)
  and u12875 (n3537, ECOREVNUM[0], I5eow6);  // ../RTL/cortexm0ds_logic.v(11385)
  not u12876 (U4eow6, n3537);  // ../RTL/cortexm0ds_logic.v(11385)
  and u12877 (G4eow6, P5eow6, W5eow6);  // ../RTL/cortexm0ds_logic.v(11386)
  and u12878 (n3538, Y5eiu6, Bxghu6);  // ../RTL/cortexm0ds_logic.v(11387)
  not u12879 (W5eow6, n3538);  // ../RTL/cortexm0ds_logic.v(11387)
  and u1288 (n94, M7zhu6, Amzhu6);  // ../RTL/cortexm0ds_logic.v(3344)
  and u12880 (n3539, Yvgiu6, Tzfpw6[0]);  // ../RTL/cortexm0ds_logic.v(11388)
  not u12881 (P5eow6, n3539);  // ../RTL/cortexm0ds_logic.v(11388)
  and u12882 (S3eow6, D6eow6, K6eow6);  // ../RTL/cortexm0ds_logic.v(11389)
  and u12883 (K6eow6, R6eow6, Y6eow6);  // ../RTL/cortexm0ds_logic.v(11390)
  and u12884 (n3540, Bagpw6[0], M6eiu6);  // ../RTL/cortexm0ds_logic.v(11391)
  not u12885 (Y6eow6, n3540);  // ../RTL/cortexm0ds_logic.v(11391)
  and u12886 (n3541, Odgpw6[0], M0eow6);  // ../RTL/cortexm0ds_logic.v(11392)
  not u12887 (R6eow6, n3541);  // ../RTL/cortexm0ds_logic.v(11392)
  and u12888 (D6eow6, F7eow6, M7eow6);  // ../RTL/cortexm0ds_logic.v(11393)
  and u12889 (n3542, T7eow6, vis_ipsr_o[0]);  // ../RTL/cortexm0ds_logic.v(11394)
  not u1289 (Tlzhu6, n94);  // ../RTL/cortexm0ds_logic.v(3344)
  not u12890 (M7eow6, n3542);  // ../RTL/cortexm0ds_logic.v(11394)
  and u12891 (n3543, F0eow6, Vbgpw6[0]);  // ../RTL/cortexm0ds_logic.v(11395)
  not u12892 (F7eow6, n3543);  // ../RTL/cortexm0ds_logic.v(11395)
  and u12893 (E3eow6, A8eow6, H8eow6);  // ../RTL/cortexm0ds_logic.v(11396)
  and u12894 (n3544, C2eow6, Lj3ju6);  // ../RTL/cortexm0ds_logic.v(11397)
  not u12895 (H8eow6, n3544);  // ../RTL/cortexm0ds_logic.v(11397)
  AL_MUX u12896 (
    .i0(O8eow6),
    .i1(Sx3ju6),
    .sel(Hv3ju6),
    .o(Lj3ju6));  // ../RTL/cortexm0ds_logic.v(11398)
  and u12897 (n3545, HRDATA[0], Q2eow6);  // ../RTL/cortexm0ds_logic.v(11399)
  not u12898 (A8eow6, n3545);  // ../RTL/cortexm0ds_logic.v(11399)
  and u12899 (Swdow6, V8eow6, C9eow6);  // ../RTL/cortexm0ds_logic.v(11400)
  buf u129 (G2ohu6, Utqpw6);  // ../RTL/cortexm0ds_logic.v(1938)
  and u1290 (M7zhu6, Hmzhu6, Omzhu6);  // ../RTL/cortexm0ds_logic.v(3345)
  or u12900 (C9eow6, Veliu6, Kldow6);  // ../RTL/cortexm0ds_logic.v(11401)
  and u12901 (Veliu6, J9eow6, Q9eow6);  // ../RTL/cortexm0ds_logic.v(11402)
  or u12902 (Q9eow6, Iydow6, Gntiu6);  // ../RTL/cortexm0ds_logic.v(11403)
  and u12903 (Gntiu6, X9eow6, Eaeow6);  // ../RTL/cortexm0ds_logic.v(11404)
  and u12904 (Eaeow6, Laeow6, Saeow6);  // ../RTL/cortexm0ds_logic.v(11405)
  and u12905 (Saeow6, Zaeow6, Gbeow6);  // ../RTL/cortexm0ds_logic.v(11406)
  and u12906 (n3546, Bagpw6[16], M6eiu6);  // ../RTL/cortexm0ds_logic.v(11407)
  not u12907 (Gbeow6, n3546);  // ../RTL/cortexm0ds_logic.v(11407)
  and u12908 (n3547, Tzfpw6[16], Yvgiu6);  // ../RTL/cortexm0ds_logic.v(11408)
  not u12909 (Zaeow6, n3547);  // ../RTL/cortexm0ds_logic.v(11408)
  or u1291 (n95, Wdyhu6, Vmzhu6);  // ../RTL/cortexm0ds_logic.v(3346)
  and u12910 (Laeow6, Nbeow6, Ubeow6);  // ../RTL/cortexm0ds_logic.v(11409)
  and u12911 (n3548, Krghu6, Y5eiu6);  // ../RTL/cortexm0ds_logic.v(11410)
  not u12912 (Ubeow6, n3548);  // ../RTL/cortexm0ds_logic.v(11410)
  and u12913 (n3549, Odgpw6[16], M0eow6);  // ../RTL/cortexm0ds_logic.v(11411)
  not u12914 (Nbeow6, n3549);  // ../RTL/cortexm0ds_logic.v(11411)
  and u12915 (X9eow6, Bceow6, Iceow6);  // ../RTL/cortexm0ds_logic.v(11412)
  and u12916 (n3550, Pceow6, Wceow6);  // ../RTL/cortexm0ds_logic.v(11413)
  not u12917 (Iceow6, n3550);  // ../RTL/cortexm0ds_logic.v(11413)
  or u12918 (Wceow6, Nzhiu6, Vbgpw6[16]);  // ../RTL/cortexm0ds_logic.v(11414)
  and u12919 (Bceow6, Ddeow6, Kdeow6);  // ../RTL/cortexm0ds_logic.v(11415)
  not u1292 (Hmzhu6, n95);  // ../RTL/cortexm0ds_logic.v(3346)
  and u12920 (n3551, STCALIB[16], H1eow6);  // ../RTL/cortexm0ds_logic.v(11416)
  not u12921 (Kdeow6, n3551);  // ../RTL/cortexm0ds_logic.v(11416)
  or u12922 (Ddeow6, Z4ciu6, Qkgiu6);  // ../RTL/cortexm0ds_logic.v(11417)
  and u12923 (n3552, Rdeow6, Ydeow6);  // ../RTL/cortexm0ds_logic.v(11418)
  not u12924 (Z4ciu6, n3552);  // ../RTL/cortexm0ds_logic.v(11418)
  or u12925 (n3553, Feeow6, Meeow6);  // ../RTL/cortexm0ds_logic.v(11419)
  not u12926 (Rdeow6, n3553);  // ../RTL/cortexm0ds_logic.v(11419)
  and u12927 (J9eow6, Teeow6, Afeow6);  // ../RTL/cortexm0ds_logic.v(11420)
  or u12928 (Afeow6, Uk3ju6, Hfeow6);  // ../RTL/cortexm0ds_logic.v(11421)
  not u12929 (Uk3ju6, Ofeow6);  // ../RTL/cortexm0ds_logic.v(11422)
  and u1293 (Mlzhu6, Cnzhu6, Joyhu6);  // ../RTL/cortexm0ds_logic.v(3347)
  AL_MUX u12930 (
    .i0(Ke4ju6),
    .i1(E44ju6),
    .sel(Hv3ju6),
    .o(Ofeow6));  // ../RTL/cortexm0ds_logic.v(11423)
  and u12931 (n3554, HRDATA[16], Q2eow6);  // ../RTL/cortexm0ds_logic.v(11424)
  not u12932 (Teeow6, n3554);  // ../RTL/cortexm0ds_logic.v(11424)
  and u12933 (n3555, Jfliu6, Fmdow6);  // ../RTL/cortexm0ds_logic.v(11425)
  not u12934 (V8eow6, n3555);  // ../RTL/cortexm0ds_logic.v(11425)
  and u12935 (n3556, Vfeow6, Cgeow6);  // ../RTL/cortexm0ds_logic.v(11426)
  not u12936 (Jfliu6, n3556);  // ../RTL/cortexm0ds_logic.v(11426)
  or u12937 (Cgeow6, Iydow6, P8viu6);  // ../RTL/cortexm0ds_logic.v(11427)
  and u12938 (P8viu6, Jgeow6, Qgeow6);  // ../RTL/cortexm0ds_logic.v(11428)
  and u12939 (Jgeow6, Xgeow6, Eheow6);  // ../RTL/cortexm0ds_logic.v(11429)
  and u1294 (n96, U4zhu6, Jnzhu6);  // ../RTL/cortexm0ds_logic.v(3348)
  and u12940 (n3557, M0eow6, Odgpw6[24]);  // ../RTL/cortexm0ds_logic.v(11430)
  not u12941 (Eheow6, n3557);  // ../RTL/cortexm0ds_logic.v(11430)
  and u12942 (n3558, F0eow6, Vbgpw6[24]);  // ../RTL/cortexm0ds_logic.v(11431)
  not u12943 (Xgeow6, n3558);  // ../RTL/cortexm0ds_logic.v(11431)
  and u12944 (Vfeow6, Lheow6, Sheow6);  // ../RTL/cortexm0ds_logic.v(11432)
  and u12945 (n3559, HRDATA[24], Q2eow6);  // ../RTL/cortexm0ds_logic.v(11433)
  not u12946 (Sheow6, n3559);  // ../RTL/cortexm0ds_logic.v(11433)
  and u12947 (n3560, C2eow6, Eb4ju6);  // ../RTL/cortexm0ds_logic.v(11434)
  not u12948 (Lheow6, n3560);  // ../RTL/cortexm0ds_logic.v(11434)
  and u12949 (n3561, Zheow6, Gieow6);  // ../RTL/cortexm0ds_logic.v(11435)
  not u1295 (Cnzhu6, n96);  // ../RTL/cortexm0ds_logic.v(3348)
  not u12950 (Eb4ju6, n3561);  // ../RTL/cortexm0ds_logic.v(11435)
  and u12951 (n3562, Nieow6, Vh3ju6);  // ../RTL/cortexm0ds_logic.v(11436)
  not u12952 (Gieow6, n3562);  // ../RTL/cortexm0ds_logic.v(11436)
  or u12953 (Zheow6, Nk3ju6, Nieow6);  // ../RTL/cortexm0ds_logic.v(11437)
  or u12954 (n3563, Uieow6, Ii0iu6);  // ../RTL/cortexm0ds_logic.v(11438)
  not u12955 (Nieow6, n3563);  // ../RTL/cortexm0ds_logic.v(11438)
  not u12956 (Nk3ju6, Bjeow6);  // ../RTL/cortexm0ds_logic.v(11439)
  AL_MUX u12957 (
    .i0(V24ju6),
    .i1(Ijeow6),
    .sel(Hv3ju6),
    .o(Bjeow6));  // ../RTL/cortexm0ds_logic.v(11440)
  and u12958 (Jvdow6, Pjeow6, Wjeow6);  // ../RTL/cortexm0ds_logic.v(11441)
  and u12959 (n3564, Zsfpw6[7], Cmziu6);  // ../RTL/cortexm0ds_logic.v(11442)
  and u1296 (n97, Hknhu6, Amzhu6);  // ../RTL/cortexm0ds_logic.v(3349)
  not u12960 (Wjeow6, n3564);  // ../RTL/cortexm0ds_logic.v(11442)
  and u12961 (n3565, vis_pc_o[7], Jmziu6);  // ../RTL/cortexm0ds_logic.v(11443)
  not u12962 (Pjeow6, n3565);  // ../RTL/cortexm0ds_logic.v(11443)
  and u12963 (n3566, Dkeow6, Kkeow6);  // ../RTL/cortexm0ds_logic.v(11444)
  not u12964 (Qkohu6, n3566);  // ../RTL/cortexm0ds_logic.v(11444)
  and u12965 (Kkeow6, Rkeow6, Ykeow6);  // ../RTL/cortexm0ds_logic.v(11445)
  and u12966 (n3567, Egziu6, Eafpw6[6]);  // ../RTL/cortexm0ds_logic.v(11446)
  not u12967 (Ykeow6, n3567);  // ../RTL/cortexm0ds_logic.v(11446)
  and u12968 (Rkeow6, Fleow6, Sgziu6);  // ../RTL/cortexm0ds_logic.v(11447)
  and u12969 (n3568, Zgziu6, Wqkiu6);  // ../RTL/cortexm0ds_logic.v(11448)
  not u1297 (Jnzhu6, n97);  // ../RTL/cortexm0ds_logic.v(3349)
  not u12970 (Fleow6, n3568);  // ../RTL/cortexm0ds_logic.v(11448)
  and u12971 (n3569, Mleow6, Tleow6);  // ../RTL/cortexm0ds_logic.v(11449)
  not u12972 (Wqkiu6, n3569);  // ../RTL/cortexm0ds_logic.v(11449)
  and u12973 (Tleow6, Ameow6, Hmeow6);  // ../RTL/cortexm0ds_logic.v(11450)
  or u12974 (Hmeow6, Cfliu6, G6cow6);  // ../RTL/cortexm0ds_logic.v(11451)
  and u12975 (Ameow6, Omeow6, Mdliu6);  // ../RTL/cortexm0ds_logic.v(11452)
  and u12976 (n3570, Qfliu6, X4cow6);  // ../RTL/cortexm0ds_logic.v(11453)
  not u12977 (Omeow6, n3570);  // ../RTL/cortexm0ds_logic.v(11453)
  and u12978 (Mleow6, Vmeow6, Cneow6);  // ../RTL/cortexm0ds_logic.v(11454)
  or u12979 (Cneow6, Ycliu6, L5cow6);  // ../RTL/cortexm0ds_logic.v(11455)
  and u1298 (n98, Mdhpw6[2], Qnzhu6);  // ../RTL/cortexm0ds_logic.v(3350)
  and u12980 (n3571, Aeliu6, N6cow6);  // ../RTL/cortexm0ds_logic.v(11456)
  not u12981 (Vmeow6, n3571);  // ../RTL/cortexm0ds_logic.v(11456)
  and u12982 (Dkeow6, Jneow6, Qneow6);  // ../RTL/cortexm0ds_logic.v(11457)
  and u12983 (n3572, Zsfpw6[5], Cmziu6);  // ../RTL/cortexm0ds_logic.v(11458)
  not u12984 (Qneow6, n3572);  // ../RTL/cortexm0ds_logic.v(11458)
  and u12985 (n3573, vis_pc_o[5], Jmziu6);  // ../RTL/cortexm0ds_logic.v(11459)
  not u12986 (Jneow6, n3573);  // ../RTL/cortexm0ds_logic.v(11459)
  and u12987 (n3574, Xneow6, Eoeow6);  // ../RTL/cortexm0ds_logic.v(11460)
  not u12988 (Jkohu6, n3574);  // ../RTL/cortexm0ds_logic.v(11460)
  and u12989 (Eoeow6, Loeow6, Soeow6);  // ../RTL/cortexm0ds_logic.v(11461)
  not u1299 (Amzhu6, n98);  // ../RTL/cortexm0ds_logic.v(3350)
  and u12990 (n3575, Egziu6, Eafpw6[5]);  // ../RTL/cortexm0ds_logic.v(11462)
  not u12991 (Soeow6, n3575);  // ../RTL/cortexm0ds_logic.v(11462)
  and u12992 (Loeow6, Zoeow6, Sgziu6);  // ../RTL/cortexm0ds_logic.v(11463)
  or u12993 (Zoeow6, Ft6ow6, Ljbiu6);  // ../RTL/cortexm0ds_logic.v(11464)
  and u12994 (Ljbiu6, Gpeow6, Npeow6);  // ../RTL/cortexm0ds_logic.v(11465)
  and u12995 (Npeow6, Upeow6, Bqeow6);  // ../RTL/cortexm0ds_logic.v(11466)
  or u12996 (Bqeow6, Rjziu6, Iqeow6);  // ../RTL/cortexm0ds_logic.v(11467)
  and u12997 (Rjziu6, Pqeow6, Wqeow6);  // ../RTL/cortexm0ds_logic.v(11468)
  or u12998 (Wqeow6, Iydow6, U6wiu6);  // ../RTL/cortexm0ds_logic.v(11469)
  and u12999 (U6wiu6, Dreow6, Kreow6);  // ../RTL/cortexm0ds_logic.v(11470)
  buf u13 (Qmdhu6, Evhpw6);  // ../RTL/cortexm0ds_logic.v(1769)
  buf u130 (Q7ohu6, Xvqpw6);  // ../RTL/cortexm0ds_logic.v(1939)
  and u1300 (U4zhu6, Xnzhu6, Eozhu6);  // ../RTL/cortexm0ds_logic.v(3352)
  and u13000 (n3576, F0eow6, Vbgpw6[29]);  // ../RTL/cortexm0ds_logic.v(11471)
  not u13001 (Kreow6, n3576);  // ../RTL/cortexm0ds_logic.v(11471)
  and u13002 (Dreow6, Rreow6, Yreow6);  // ../RTL/cortexm0ds_logic.v(11472)
  and u13003 (n3577, Odgpw6[29], M0eow6);  // ../RTL/cortexm0ds_logic.v(11473)
  not u13004 (Rreow6, n3577);  // ../RTL/cortexm0ds_logic.v(11473)
  and u13005 (Pqeow6, Fseow6, Mseow6);  // ../RTL/cortexm0ds_logic.v(11474)
  and u13006 (n3578, C2eow6, Tseow6);  // ../RTL/cortexm0ds_logic.v(11475)
  not u13007 (Mseow6, n3578);  // ../RTL/cortexm0ds_logic.v(11475)
  and u13008 (n3579, T84ju6, Ateow6);  // ../RTL/cortexm0ds_logic.v(11476)
  not u13009 (Tseow6, n3579);  // ../RTL/cortexm0ds_logic.v(11476)
  not u1301 (Pryhu6, U4zhu6);  // ../RTL/cortexm0ds_logic.v(3352)
  or u13010 (Ateow6, Hteow6, Bz3ju6);  // ../RTL/cortexm0ds_logic.v(11477)
  and u13011 (n3580, Oteow6, Vteow6);  // ../RTL/cortexm0ds_logic.v(11478)
  not u13012 (T84ju6, n3580);  // ../RTL/cortexm0ds_logic.v(11478)
  or u13013 (Vteow6, Ex3ju6, J2eow6);  // ../RTL/cortexm0ds_logic.v(11479)
  and u13014 (Oteow6, Cueow6, Hteow6);  // ../RTL/cortexm0ds_logic.v(11480)
  and u13015 (n3581, Jueow6, Queow6);  // ../RTL/cortexm0ds_logic.v(11481)
  not u13016 (Hteow6, n3581);  // ../RTL/cortexm0ds_logic.v(11481)
  and u13017 (Jueow6, Xueow6, Eveow6);  // ../RTL/cortexm0ds_logic.v(11482)
  and u13018 (n3582, Lveow6, Sveow6);  // ../RTL/cortexm0ds_logic.v(11483)
  not u13019 (Eveow6, n3582);  // ../RTL/cortexm0ds_logic.v(11483)
  or u1302 (n99, Vmzhu6, Ighpw6[1]);  // ../RTL/cortexm0ds_logic.v(3353)
  or u13020 (Xueow6, Zveow6, Gweow6);  // ../RTL/cortexm0ds_logic.v(11484)
  and u13021 (n3583, Nweow6, J2eow6);  // ../RTL/cortexm0ds_logic.v(11485)
  not u13022 (Cueow6, n3583);  // ../RTL/cortexm0ds_logic.v(11485)
  and u13023 (n3584, Q2eow6, HRDATA[29]);  // ../RTL/cortexm0ds_logic.v(11486)
  not u13024 (Fseow6, n3584);  // ../RTL/cortexm0ds_logic.v(11486)
  and u13025 (Upeow6, Uweow6, Mdliu6);  // ../RTL/cortexm0ds_logic.v(11487)
  or u13026 (Uweow6, Tkziu6, Ycliu6);  // ../RTL/cortexm0ds_logic.v(11488)
  and u13027 (Tkziu6, Bxeow6, Ixeow6);  // ../RTL/cortexm0ds_logic.v(11489)
  and u13028 (Ixeow6, Pxeow6, Wxeow6);  // ../RTL/cortexm0ds_logic.v(11490)
  and u13029 (n3585, Dyeow6, Ff4ju6);  // ../RTL/cortexm0ds_logic.v(11491)
  not u1303 (Eozhu6, n99);  // ../RTL/cortexm0ds_logic.v(3353)
  not u13030 (Wxeow6, n3585);  // ../RTL/cortexm0ds_logic.v(11491)
  or u13031 (Pxeow6, Iydow6, U2tiu6);  // ../RTL/cortexm0ds_logic.v(11492)
  and u13032 (U2tiu6, Kyeow6, Ryeow6);  // ../RTL/cortexm0ds_logic.v(11493)
  and u13033 (Ryeow6, Yyeow6, Fzeow6);  // ../RTL/cortexm0ds_logic.v(11494)
  and u13034 (n3586, Tzfpw6[13], Yvgiu6);  // ../RTL/cortexm0ds_logic.v(11495)
  not u13035 (Fzeow6, n3586);  // ../RTL/cortexm0ds_logic.v(11495)
  and u13036 (Yyeow6, Mzeow6, Tzeow6);  // ../RTL/cortexm0ds_logic.v(11496)
  and u13037 (n3587, T7eow6, E4ciu6);  // ../RTL/cortexm0ds_logic.v(11497)
  not u13038 (Tzeow6, n3587);  // ../RTL/cortexm0ds_logic.v(11497)
  and u13039 (n3588, A0fow6, H0fow6);  // ../RTL/cortexm0ds_logic.v(11498)
  or u1304 (n100, Zazhu6, Wdyhu6);  // ../RTL/cortexm0ds_logic.v(3354)
  not u13040 (E4ciu6, n3588);  // ../RTL/cortexm0ds_logic.v(11498)
  and u13041 (n3589, O0fow6, V0fow6);  // ../RTL/cortexm0ds_logic.v(11499)
  not u13042 (H0fow6, n3589);  // ../RTL/cortexm0ds_logic.v(11499)
  and u13043 (n3590, C1fow6, J1fow6);  // ../RTL/cortexm0ds_logic.v(11500)
  not u13044 (O0fow6, n3590);  // ../RTL/cortexm0ds_logic.v(11500)
  AL_MUX u13045 (
    .i0(Q1fow6),
    .i1(X1fow6),
    .sel(E2fow6),
    .o(C1fow6));  // ../RTL/cortexm0ds_logic.v(11501)
  and u13046 (X1fow6, L2fow6, S2fow6);  // ../RTL/cortexm0ds_logic.v(11502)
  and u13047 (n3591, Z2fow6, G3fow6);  // ../RTL/cortexm0ds_logic.v(11503)
  not u13048 (S2fow6, n3591);  // ../RTL/cortexm0ds_logic.v(11503)
  AL_MUX u13049 (
    .i0(N3fow6),
    .i1(U3fow6),
    .sel(B4fow6),
    .o(L2fow6));  // ../RTL/cortexm0ds_logic.v(11504)
  not u1305 (Xnzhu6, n100);  // ../RTL/cortexm0ds_logic.v(3354)
  or u13050 (U3fow6, I4fow6, P4fow6);  // ../RTL/cortexm0ds_logic.v(11505)
  AL_MUX u13051 (
    .i0(W4fow6),
    .i1(D5fow6),
    .sel(K5fow6),
    .o(N3fow6));  // ../RTL/cortexm0ds_logic.v(11506)
  and u13052 (Q1fow6, R5fow6, Y5fow6);  // ../RTL/cortexm0ds_logic.v(11507)
  or u13053 (Y5fow6, F6fow6, M6fow6);  // ../RTL/cortexm0ds_logic.v(11508)
  AL_MUX u13054 (
    .i0(T6fow6),
    .i1(A7fow6),
    .sel(H7fow6),
    .o(R5fow6));  // ../RTL/cortexm0ds_logic.v(11509)
  or u13055 (A7fow6, O7fow6, V7fow6);  // ../RTL/cortexm0ds_logic.v(11510)
  or u13056 (n3592, C8fow6, J8fow6);  // ../RTL/cortexm0ds_logic.v(11511)
  not u13057 (T6fow6, n3592);  // ../RTL/cortexm0ds_logic.v(11511)
  or u13058 (n3593, Q8fow6, X8fow6);  // ../RTL/cortexm0ds_logic.v(11512)
  not u13059 (J8fow6, n3593);  // ../RTL/cortexm0ds_logic.v(11512)
  not u1306 (Zazhu6, Ighpw6[0]);  // ../RTL/cortexm0ds_logic.v(3355)
  and u13060 (n3594, Odgpw6[13], M0eow6);  // ../RTL/cortexm0ds_logic.v(11513)
  not u13061 (Mzeow6, n3594);  // ../RTL/cortexm0ds_logic.v(11513)
  and u13062 (Kyeow6, E9fow6, L9fow6);  // ../RTL/cortexm0ds_logic.v(11514)
  and u13063 (n3595, F0eow6, Vbgpw6[13]);  // ../RTL/cortexm0ds_logic.v(11515)
  not u13064 (L9fow6, n3595);  // ../RTL/cortexm0ds_logic.v(11515)
  and u13065 (E9fow6, S9fow6, Z9fow6);  // ../RTL/cortexm0ds_logic.v(11516)
  and u13066 (n3596, STCALIB[13], H1eow6);  // ../RTL/cortexm0ds_logic.v(11517)
  not u13067 (Z9fow6, n3596);  // ../RTL/cortexm0ds_logic.v(11517)
  and u13068 (n3597, Bagpw6[13], M6eiu6);  // ../RTL/cortexm0ds_logic.v(11518)
  not u13069 (S9fow6, n3597);  // ../RTL/cortexm0ds_logic.v(11518)
  and u1307 (n7[0], Gbzhu6, Nbzhu6);  // ../RTL/cortexm0ds_logic.v(3185)
  and u13070 (Bxeow6, Gafow6, Nafow6);  // ../RTL/cortexm0ds_logic.v(11519)
  or u13071 (Nafow6, Uafow6, Uc4ju6);  // ../RTL/cortexm0ds_logic.v(11520)
  and u13072 (n3598, Q2eow6, HRDATA[13]);  // ../RTL/cortexm0ds_logic.v(11521)
  not u13073 (Gafow6, n3598);  // ../RTL/cortexm0ds_logic.v(11521)
  and u13074 (Gpeow6, Bbfow6, Ibfow6);  // ../RTL/cortexm0ds_logic.v(11522)
  or u13075 (Ibfow6, Alziu6, Cfliu6);  // ../RTL/cortexm0ds_logic.v(11523)
  and u13076 (Alziu6, Pbfow6, Wbfow6);  // ../RTL/cortexm0ds_logic.v(11524)
  and u13077 (Wbfow6, Dcfow6, Kcfow6);  // ../RTL/cortexm0ds_logic.v(11525)
  or u13078 (Kcfow6, Rcfow6, J34ju6);  // ../RTL/cortexm0ds_logic.v(11526)
  or u13079 (Dcfow6, Iydow6, Umuiu6);  // ../RTL/cortexm0ds_logic.v(11528)
  buf u1308 (Tnhpw6[0], Qehbx6);  // ../RTL/cortexm0ds_logic.v(2163)
  and u13080 (Umuiu6, Ycfow6, Fdfow6);  // ../RTL/cortexm0ds_logic.v(11529)
  and u13081 (Fdfow6, Mdfow6, Tdfow6);  // ../RTL/cortexm0ds_logic.v(11530)
  and u13082 (n3599, Tzfpw6[21], Yvgiu6);  // ../RTL/cortexm0ds_logic.v(11531)
  not u13083 (Tdfow6, n3599);  // ../RTL/cortexm0ds_logic.v(11531)
  and u13084 (Mdfow6, Aefow6, Hefow6);  // ../RTL/cortexm0ds_logic.v(11532)
  and u13085 (n3600, F0eow6, Vbgpw6[21]);  // ../RTL/cortexm0ds_logic.v(11533)
  not u13086 (Hefow6, n3600);  // ../RTL/cortexm0ds_logic.v(11533)
  and u13087 (n3601, Odgpw6[21], M0eow6);  // ../RTL/cortexm0ds_logic.v(11534)
  not u13088 (Aefow6, n3601);  // ../RTL/cortexm0ds_logic.v(11534)
  and u13089 (Ycfow6, Oefow6, Vefow6);  // ../RTL/cortexm0ds_logic.v(11535)
  and u1309 (n102, Zozhu6, Gpzhu6);  // ../RTL/cortexm0ds_logic.v(3357)
  and u13090 (n3602, Bagpw6[21], M6eiu6);  // ../RTL/cortexm0ds_logic.v(11536)
  not u13091 (Vefow6, n3602);  // ../RTL/cortexm0ds_logic.v(11536)
  and u13092 (n3603, STCALIB[21], H1eow6);  // ../RTL/cortexm0ds_logic.v(11537)
  not u13093 (Oefow6, n3603);  // ../RTL/cortexm0ds_logic.v(11537)
  and u13094 (Pbfow6, Cffow6, Jffow6);  // ../RTL/cortexm0ds_logic.v(11538)
  or u13095 (Jffow6, Uafow6, F14ju6);  // ../RTL/cortexm0ds_logic.v(11539)
  and u13096 (n3604, HRDATA[21], Q2eow6);  // ../RTL/cortexm0ds_logic.v(11540)
  not u13097 (Cffow6, n3604);  // ../RTL/cortexm0ds_logic.v(11540)
  or u13098 (Bbfow6, Piziu6, Qffow6);  // ../RTL/cortexm0ds_logic.v(11541)
  and u13099 (Piziu6, Xffow6, Egfow6);  // ../RTL/cortexm0ds_logic.v(11542)
  buf u131 (Lznhu6, Xxqpw6);  // ../RTL/cortexm0ds_logic.v(1940)
  not u1310 (Sozhu6, n102);  // ../RTL/cortexm0ds_logic.v(3357)
  and u13100 (Egfow6, Lgfow6, Sgfow6);  // ../RTL/cortexm0ds_logic.v(11543)
  and u13101 (n3605, Dyeow6, Hg4ju6);  // ../RTL/cortexm0ds_logic.v(11544)
  not u13102 (Sgfow6, n3605);  // ../RTL/cortexm0ds_logic.v(11544)
  or u13103 (Lgfow6, Iydow6, Eariu6);  // ../RTL/cortexm0ds_logic.v(11545)
  and u13104 (Eariu6, Zgfow6, Ghfow6);  // ../RTL/cortexm0ds_logic.v(11546)
  and u13105 (Ghfow6, Nhfow6, Uhfow6);  // ../RTL/cortexm0ds_logic.v(11547)
  and u13106 (n3606, Tzfpw6[5], Yvgiu6);  // ../RTL/cortexm0ds_logic.v(11548)
  not u13107 (Uhfow6, n3606);  // ../RTL/cortexm0ds_logic.v(11548)
  and u13108 (Nhfow6, Bifow6, Iifow6);  // ../RTL/cortexm0ds_logic.v(11549)
  and u13109 (n3607, Bagpw6[5], M6eiu6);  // ../RTL/cortexm0ds_logic.v(11550)
  and u1311 (n103, Npzhu6, Upzhu6);  // ../RTL/cortexm0ds_logic.v(3358)
  not u13110 (Iifow6, n3607);  // ../RTL/cortexm0ds_logic.v(11550)
  and u13111 (n3608, Odgpw6[5], M0eow6);  // ../RTL/cortexm0ds_logic.v(11551)
  not u13112 (Bifow6, n3608);  // ../RTL/cortexm0ds_logic.v(11551)
  and u13113 (Zgfow6, Pifow6, Wifow6);  // ../RTL/cortexm0ds_logic.v(11552)
  and u13114 (n3609, F0eow6, Vbgpw6[5]);  // ../RTL/cortexm0ds_logic.v(11553)
  not u13115 (Wifow6, n3609);  // ../RTL/cortexm0ds_logic.v(11553)
  and u13116 (Pifow6, Djfow6, Kjfow6);  // ../RTL/cortexm0ds_logic.v(11554)
  and u13117 (n3610, STCALIB[5], H1eow6);  // ../RTL/cortexm0ds_logic.v(11555)
  not u13118 (Kjfow6, n3610);  // ../RTL/cortexm0ds_logic.v(11555)
  or u13119 (Djfow6, Qkgiu6, Vhbiu6);  // ../RTL/cortexm0ds_logic.v(11556)
  not u1312 (Zozhu6, n103);  // ../RTL/cortexm0ds_logic.v(3358)
  and u13120 (Xffow6, Rjfow6, Yjfow6);  // ../RTL/cortexm0ds_logic.v(11557)
  or u13121 (Yjfow6, Uafow6, Mu3ju6);  // ../RTL/cortexm0ds_logic.v(11558)
  and u13122 (n3611, HRDATA[5], Q2eow6);  // ../RTL/cortexm0ds_logic.v(11559)
  not u13123 (Rjfow6, n3611);  // ../RTL/cortexm0ds_logic.v(11559)
  and u13124 (Xneow6, Fkfow6, Mkfow6);  // ../RTL/cortexm0ds_logic.v(11560)
  and u13125 (n3612, Zsfpw6[4], Cmziu6);  // ../RTL/cortexm0ds_logic.v(11561)
  not u13126 (Mkfow6, n3612);  // ../RTL/cortexm0ds_logic.v(11561)
  and u13127 (n3613, vis_pc_o[4], Jmziu6);  // ../RTL/cortexm0ds_logic.v(11562)
  not u13128 (Fkfow6, n3613);  // ../RTL/cortexm0ds_logic.v(11562)
  and u13129 (n3614, Tkfow6, Alfow6);  // ../RTL/cortexm0ds_logic.v(11563)
  and u1313 (n104, Bqzhu6, Iqzhu6);  // ../RTL/cortexm0ds_logic.v(3359)
  not u13130 (Ckohu6, n3614);  // ../RTL/cortexm0ds_logic.v(11563)
  and u13131 (Alfow6, Hlfow6, Olfow6);  // ../RTL/cortexm0ds_logic.v(11564)
  and u13132 (n3615, Egziu6, Eafpw6[4]);  // ../RTL/cortexm0ds_logic.v(11565)
  not u13133 (Olfow6, n3615);  // ../RTL/cortexm0ds_logic.v(11565)
  and u13134 (Hlfow6, Vlfow6, Sgziu6);  // ../RTL/cortexm0ds_logic.v(11566)
  or u13135 (Vlfow6, Ft6ow6, Y4fiu6);  // ../RTL/cortexm0ds_logic.v(11567)
  and u13136 (Y4fiu6, Cmfow6, Jmfow6);  // ../RTL/cortexm0ds_logic.v(11568)
  and u13137 (Jmfow6, Qmfow6, Xmfow6);  // ../RTL/cortexm0ds_logic.v(11569)
  or u13138 (Xmfow6, K1cow6, Cfliu6);  // ../RTL/cortexm0ds_logic.v(11570)
  and u13139 (K1cow6, Enfow6, Lnfow6);  // ../RTL/cortexm0ds_logic.v(11571)
  not u1314 (Upzhu6, n104);  // ../RTL/cortexm0ds_logic.v(3359)
  and u13140 (Lnfow6, Snfow6, Znfow6);  // ../RTL/cortexm0ds_logic.v(11572)
  and u13141 (n3616, Dyeow6, V24ju6);  // ../RTL/cortexm0ds_logic.v(11573)
  not u13142 (Znfow6, n3616);  // ../RTL/cortexm0ds_logic.v(11573)
  and u13143 (n3617, Gofow6, Nofow6);  // ../RTL/cortexm0ds_logic.v(11574)
  not u13144 (V24ju6, n3617);  // ../RTL/cortexm0ds_logic.v(11574)
  and u13145 (Nofow6, Uofow6, Bpfow6);  // ../RTL/cortexm0ds_logic.v(11575)
  or u13146 (Bpfow6, Ipfow6, A70iu6);  // ../RTL/cortexm0ds_logic.v(11576)
  or u13147 (Uofow6, Ppfow6, V70iu6);  // ../RTL/cortexm0ds_logic.v(11577)
  and u13148 (Gofow6, Wpfow6, Dqfow6);  // ../RTL/cortexm0ds_logic.v(11578)
  or u13149 (Dqfow6, Kqfow6, O70iu6);  // ../RTL/cortexm0ds_logic.v(11579)
  or u1315 (V9xiu6, Pqzhu6, Wqzhu6);  // ../RTL/cortexm0ds_logic.v(3360)
  or u13150 (Wpfow6, Rqfow6, H70iu6);  // ../RTL/cortexm0ds_logic.v(11580)
  or u13151 (Snfow6, Iydow6, Bguiu6);  // ../RTL/cortexm0ds_logic.v(11581)
  and u13152 (Bguiu6, Yqfow6, Frfow6);  // ../RTL/cortexm0ds_logic.v(11582)
  and u13153 (Frfow6, Mrfow6, Trfow6);  // ../RTL/cortexm0ds_logic.v(11583)
  and u13154 (n3618, Tzfpw6[20], Yvgiu6);  // ../RTL/cortexm0ds_logic.v(11584)
  not u13155 (Trfow6, n3618);  // ../RTL/cortexm0ds_logic.v(11584)
  and u13156 (Mrfow6, Asfow6, Hsfow6);  // ../RTL/cortexm0ds_logic.v(11585)
  and u13157 (n3619, F0eow6, Vbgpw6[20]);  // ../RTL/cortexm0ds_logic.v(11586)
  not u13158 (Hsfow6, n3619);  // ../RTL/cortexm0ds_logic.v(11586)
  and u13159 (n3620, Odgpw6[20], M0eow6);  // ../RTL/cortexm0ds_logic.v(11587)
  not u1316 (Bqzhu6, V9xiu6);  // ../RTL/cortexm0ds_logic.v(3360)
  not u13160 (Asfow6, n3620);  // ../RTL/cortexm0ds_logic.v(11587)
  and u13161 (Yqfow6, Osfow6, Vsfow6);  // ../RTL/cortexm0ds_logic.v(11588)
  and u13162 (n3621, Bagpw6[20], M6eiu6);  // ../RTL/cortexm0ds_logic.v(11589)
  not u13163 (Vsfow6, n3621);  // ../RTL/cortexm0ds_logic.v(11589)
  and u13164 (n3622, STCALIB[20], H1eow6);  // ../RTL/cortexm0ds_logic.v(11590)
  not u13165 (Osfow6, n3622);  // ../RTL/cortexm0ds_logic.v(11590)
  and u13166 (Enfow6, Ctfow6, Jtfow6);  // ../RTL/cortexm0ds_logic.v(11591)
  and u13167 (n3623, Qtfow6, E44ju6);  // ../RTL/cortexm0ds_logic.v(11592)
  not u13168 (Jtfow6, n3623);  // ../RTL/cortexm0ds_logic.v(11592)
  and u13169 (n3624, Xtfow6, Eufow6);  // ../RTL/cortexm0ds_logic.v(11593)
  and u1317 (n105, Drzhu6, Krzhu6);  // ../RTL/cortexm0ds_logic.v(3361)
  not u13170 (E44ju6, n3624);  // ../RTL/cortexm0ds_logic.v(11593)
  and u13171 (Eufow6, Lufow6, Sufow6);  // ../RTL/cortexm0ds_logic.v(11594)
  or u13172 (Sufow6, Ipfow6, C80iu6);  // ../RTL/cortexm0ds_logic.v(11595)
  or u13173 (Lufow6, Rqfow6, J80iu6);  // ../RTL/cortexm0ds_logic.v(11596)
  and u13174 (Xtfow6, Zufow6, Gvfow6);  // ../RTL/cortexm0ds_logic.v(11597)
  or u13175 (Gvfow6, Ppfow6, X80iu6);  // ../RTL/cortexm0ds_logic.v(11598)
  or u13176 (Zufow6, Kqfow6, Q80iu6);  // ../RTL/cortexm0ds_logic.v(11599)
  and u13177 (n3625, HRDATA[20], Q2eow6);  // ../RTL/cortexm0ds_logic.v(11600)
  not u13178 (Ctfow6, n3625);  // ../RTL/cortexm0ds_logic.v(11600)
  and u13179 (Qmfow6, Nvfow6, Mdliu6);  // ../RTL/cortexm0ds_logic.v(11601)
  not u1318 (Lozhu6, n105);  // ../RTL/cortexm0ds_logic.v(3361)
  or u13180 (Nvfow6, P0cow6, Iqeow6);  // ../RTL/cortexm0ds_logic.v(11602)
  and u13181 (P0cow6, Uvfow6, Bwfow6);  // ../RTL/cortexm0ds_logic.v(11603)
  or u13182 (Bwfow6, Iydow6, I0wiu6);  // ../RTL/cortexm0ds_logic.v(11604)
  and u13183 (I0wiu6, Iwfow6, Pwfow6);  // ../RTL/cortexm0ds_logic.v(11605)
  and u13184 (n3626, Pceow6, Wwfow6);  // ../RTL/cortexm0ds_logic.v(11606)
  not u13185 (Pwfow6, n3626);  // ../RTL/cortexm0ds_logic.v(11606)
  or u13186 (Wwfow6, Nzhiu6, Vbgpw6[28]);  // ../RTL/cortexm0ds_logic.v(11607)
  and u13187 (Iwfow6, Dxfow6, Kxfow6);  // ../RTL/cortexm0ds_logic.v(11608)
  or u13188 (Kxfow6, Jh5iu6, Qkgiu6);  // ../RTL/cortexm0ds_logic.v(11609)
  not u13189 (Jh5iu6, Ikghu6);  // ../RTL/cortexm0ds_logic.v(11610)
  buf u1319 (Vbgpw6[25], Pv0bx6);  // ../RTL/cortexm0ds_logic.v(3092)
  and u13190 (n3627, Odgpw6[28], M0eow6);  // ../RTL/cortexm0ds_logic.v(11611)
  not u13191 (Dxfow6, n3627);  // ../RTL/cortexm0ds_logic.v(11611)
  and u13192 (Uvfow6, Rxfow6, Yxfow6);  // ../RTL/cortexm0ds_logic.v(11612)
  and u13193 (n3628, C2eow6, Xa4ju6);  // ../RTL/cortexm0ds_logic.v(11613)
  not u13194 (Yxfow6, n3628);  // ../RTL/cortexm0ds_logic.v(11613)
  AL_MUX u13195 (
    .i0(Fyfow6),
    .i1(Vh3ju6),
    .sel(Myfow6),
    .o(Xa4ju6));  // ../RTL/cortexm0ds_logic.v(11614)
  and u13196 (Myfow6, Tyfow6, Cyfpw6[3]);  // ../RTL/cortexm0ds_logic.v(11615)
  and u13197 (Tyfow6, Azfow6, Hzfow6);  // ../RTL/cortexm0ds_logic.v(11616)
  AL_MUX u13198 (
    .i0(Ijeow6),
    .i1(O8eow6),
    .sel(Hv3ju6),
    .o(Fyfow6));  // ../RTL/cortexm0ds_logic.v(11617)
  and u13199 (n3629, Ozfow6, Vzfow6);  // ../RTL/cortexm0ds_logic.v(11618)
  buf u132 (vis_r6_o[0], Kloax6);  // ../RTL/cortexm0ds_logic.v(2523)
  buf u1320 (Vbgpw6[26], X5upw6);  // ../RTL/cortexm0ds_logic.v(3092)
  not u13200 (O8eow6, n3629);  // ../RTL/cortexm0ds_logic.v(11618)
  and u13201 (Vzfow6, C0gow6, J0gow6);  // ../RTL/cortexm0ds_logic.v(11619)
  or u13202 (J0gow6, Rqfow6, F60iu6);  // ../RTL/cortexm0ds_logic.v(11620)
  or u13203 (C0gow6, Ipfow6, K50iu6);  // ../RTL/cortexm0ds_logic.v(11621)
  and u13204 (Ozfow6, Q0gow6, X0gow6);  // ../RTL/cortexm0ds_logic.v(11622)
  or u13205 (X0gow6, Ppfow6, Dc0iu6);  // ../RTL/cortexm0ds_logic.v(11623)
  or u13206 (Q0gow6, Kqfow6, E90iu6);  // ../RTL/cortexm0ds_logic.v(11624)
  and u13207 (n3630, E1gow6, L1gow6);  // ../RTL/cortexm0ds_logic.v(11625)
  not u13208 (Ijeow6, n3630);  // ../RTL/cortexm0ds_logic.v(11625)
  and u13209 (L1gow6, S1gow6, Z1gow6);  // ../RTL/cortexm0ds_logic.v(11626)
  and u1321 (n106, Krzhu6, Fszhu6);  // ../RTL/cortexm0ds_logic.v(3363)
  or u13210 (Z1gow6, Ipfow6, R50iu6);  // ../RTL/cortexm0ds_logic.v(11627)
  or u13211 (S1gow6, Ppfow6, T60iu6);  // ../RTL/cortexm0ds_logic.v(11628)
  and u13212 (E1gow6, G2gow6, N2gow6);  // ../RTL/cortexm0ds_logic.v(11629)
  or u13213 (N2gow6, Kqfow6, M60iu6);  // ../RTL/cortexm0ds_logic.v(11630)
  or u13214 (G2gow6, Rqfow6, Y50iu6);  // ../RTL/cortexm0ds_logic.v(11631)
  and u13215 (n3631, HRDATA[28], Q2eow6);  // ../RTL/cortexm0ds_logic.v(11632)
  not u13216 (Rxfow6, n3631);  // ../RTL/cortexm0ds_logic.v(11632)
  and u13217 (Cmfow6, U2gow6, B3gow6);  // ../RTL/cortexm0ds_logic.v(11633)
  or u13218 (B3gow6, R1cow6, Ycliu6);  // ../RTL/cortexm0ds_logic.v(11634)
  and u13219 (R1cow6, I3gow6, P3gow6);  // ../RTL/cortexm0ds_logic.v(11635)
  not u1322 (Yrzhu6, n106);  // ../RTL/cortexm0ds_logic.v(3363)
  and u13220 (P3gow6, W3gow6, D4gow6);  // ../RTL/cortexm0ds_logic.v(11636)
  and u13221 (n3632, Dyeow6, Ke4ju6);  // ../RTL/cortexm0ds_logic.v(11637)
  not u13222 (D4gow6, n3632);  // ../RTL/cortexm0ds_logic.v(11637)
  and u13223 (n3633, K4gow6, R4gow6);  // ../RTL/cortexm0ds_logic.v(11638)
  not u13224 (Ke4ju6, n3633);  // ../RTL/cortexm0ds_logic.v(11638)
  and u13225 (R4gow6, Y4gow6, F5gow6);  // ../RTL/cortexm0ds_logic.v(11639)
  or u13226 (F5gow6, Ipfow6, L90iu6);  // ../RTL/cortexm0ds_logic.v(11640)
  or u13227 (Y4gow6, Rqfow6, S90iu6);  // ../RTL/cortexm0ds_logic.v(11641)
  and u13228 (K4gow6, M5gow6, T5gow6);  // ../RTL/cortexm0ds_logic.v(11642)
  or u13229 (T5gow6, Ppfow6, Ga0iu6);  // ../RTL/cortexm0ds_logic.v(11643)
  or u1323 (n107, Mszhu6, Tszhu6);  // ../RTL/cortexm0ds_logic.v(3364)
  or u13230 (M5gow6, Kqfow6, Z90iu6);  // ../RTL/cortexm0ds_logic.v(11644)
  or u13231 (W3gow6, Iydow6, Nvsiu6);  // ../RTL/cortexm0ds_logic.v(11645)
  and u13232 (Nvsiu6, A6gow6, H6gow6);  // ../RTL/cortexm0ds_logic.v(11646)
  and u13233 (H6gow6, O6gow6, V6gow6);  // ../RTL/cortexm0ds_logic.v(11647)
  and u13234 (n3634, Bagpw6[12], M6eiu6);  // ../RTL/cortexm0ds_logic.v(11648)
  not u13235 (V6gow6, n3634);  // ../RTL/cortexm0ds_logic.v(11648)
  and u13236 (O6gow6, C7gow6, J7gow6);  // ../RTL/cortexm0ds_logic.v(11649)
  or u13237 (J7gow6, Kmbiu6, Qkgiu6);  // ../RTL/cortexm0ds_logic.v(11650)
  and u13238 (n3635, Q7gow6, Te6iu6);  // ../RTL/cortexm0ds_logic.v(11651)
  not u13239 (Kmbiu6, n3635);  // ../RTL/cortexm0ds_logic.v(11651)
  not u1324 (Rrzhu6, n107);  // ../RTL/cortexm0ds_logic.v(3364)
  and u13240 (n3636, X7gow6, E8gow6);  // ../RTL/cortexm0ds_logic.v(11652)
  not u13241 (Q7gow6, n3636);  // ../RTL/cortexm0ds_logic.v(11652)
  and u13242 (n3637, L8gow6, S8gow6);  // ../RTL/cortexm0ds_logic.v(11653)
  not u13243 (E8gow6, n3637);  // ../RTL/cortexm0ds_logic.v(11653)
  or u13244 (S8gow6, Z8gow6, Feeow6);  // ../RTL/cortexm0ds_logic.v(11654)
  AL_MUX u13245 (
    .i0(G9gow6),
    .i1(N9gow6),
    .sel(Meeow6),
    .o(Z8gow6));  // ../RTL/cortexm0ds_logic.v(11655)
  AL_MUX u13246 (
    .i0(U9gow6),
    .i1(Bagow6),
    .sel(H7fow6),
    .o(N9gow6));  // ../RTL/cortexm0ds_logic.v(11656)
  AL_MUX u13247 (
    .i0(Iagow6),
    .i1(Pagow6),
    .sel(O7fow6),
    .o(Bagow6));  // ../RTL/cortexm0ds_logic.v(11657)
  AL_MUX u13248 (
    .i0(Wagow6),
    .i1(Dbgow6),
    .sel(M6fow6),
    .o(Pagow6));  // ../RTL/cortexm0ds_logic.v(11658)
  AL_MUX u13249 (
    .i0(Kbgow6),
    .i1(Rbgow6),
    .sel(V7fow6),
    .o(Iagow6));  // ../RTL/cortexm0ds_logic.v(11659)
  and u1325 (Mszhu6, Atzhu6, Iqzhu6);  // ../RTL/cortexm0ds_logic.v(3365)
  and u13250 (n3638, Ybgow6, Fcgow6);  // ../RTL/cortexm0ds_logic.v(11660)
  not u13251 (U9gow6, n3638);  // ../RTL/cortexm0ds_logic.v(11660)
  and u13252 (n3639, C8fow6, Mcgow6);  // ../RTL/cortexm0ds_logic.v(11661)
  not u13253 (Fcgow6, n3639);  // ../RTL/cortexm0ds_logic.v(11661)
  AL_MUX u13254 (
    .i0(Tcgow6),
    .i1(Adgow6),
    .sel(Hdgow6),
    .o(Ybgow6));  // ../RTL/cortexm0ds_logic.v(11662)
  AL_MUX u13255 (
    .i0(Odgow6),
    .i1(Vdgow6),
    .sel(Cegow6),
    .o(Adgow6));  // ../RTL/cortexm0ds_logic.v(11663)
  or u13256 (Tcgow6, Jegow6, Qegow6);  // ../RTL/cortexm0ds_logic.v(11664)
  not u13257 (G9gow6, Xegow6);  // ../RTL/cortexm0ds_logic.v(11665)
  AL_MUX u13258 (
    .i0(Lfgow6),
    .i1(Efgow6),
    .sel(B4fow6),
    .o(Xegow6));  // ../RTL/cortexm0ds_logic.v(11666)
  AL_MUX u13259 (
    .i0(Zfgow6),
    .i1(Gggow6),
    .sel(Nggow6),
    .o(Lfgow6));  // ../RTL/cortexm0ds_logic.v(11667)
  or u1326 (n108, Sqhpw6[0], Sqhpw6[1]);  // ../RTL/cortexm0ds_logic.v(3366)
  AL_MUX u13260 (
    .i0(Bhgow6),
    .i1(Uggow6),
    .sel(W4fow6),
    .o(Gggow6));  // ../RTL/cortexm0ds_logic.v(11668)
  AL_MUX u13261 (
    .i0(Phgow6),
    .i1(Whgow6),
    .sel(Digow6),
    .o(Zfgow6));  // ../RTL/cortexm0ds_logic.v(11669)
  AL_MUX u13262 (
    .i0(Kigow6),
    .i1(Rigow6),
    .sel(Yigow6),
    .o(Efgow6));  // ../RTL/cortexm0ds_logic.v(11670)
  AL_MUX u13263 (
    .i0(Fjgow6),
    .i1(Mjgow6),
    .sel(Tjgow6),
    .o(Rigow6));  // ../RTL/cortexm0ds_logic.v(11671)
  AL_MUX u13264 (
    .i0(Akgow6),
    .i1(Hkgow6),
    .sel(G3fow6),
    .o(Kigow6));  // ../RTL/cortexm0ds_logic.v(11672)
  and u13265 (L8gow6, Okgow6, V0fow6);  // ../RTL/cortexm0ds_logic.v(11673)
  and u13266 (n3640, Tzfpw6[12], Yvgiu6);  // ../RTL/cortexm0ds_logic.v(11674)
  not u13267 (C7gow6, n3640);  // ../RTL/cortexm0ds_logic.v(11674)
  and u13268 (A6gow6, Vkgow6, Clgow6);  // ../RTL/cortexm0ds_logic.v(11675)
  and u13269 (n3641, F0eow6, Vbgpw6[12]);  // ../RTL/cortexm0ds_logic.v(11676)
  not u1327 (Atzhu6, n108);  // ../RTL/cortexm0ds_logic.v(3366)
  not u13270 (Clgow6, n3641);  // ../RTL/cortexm0ds_logic.v(11676)
  and u13271 (Vkgow6, Jlgow6, Qlgow6);  // ../RTL/cortexm0ds_logic.v(11677)
  and u13272 (n3642, STCALIB[12], H1eow6);  // ../RTL/cortexm0ds_logic.v(11678)
  not u13273 (Qlgow6, n3642);  // ../RTL/cortexm0ds_logic.v(11678)
  and u13274 (n3643, Odgpw6[12], M0eow6);  // ../RTL/cortexm0ds_logic.v(11679)
  not u13275 (Jlgow6, n3643);  // ../RTL/cortexm0ds_logic.v(11679)
  and u13276 (I3gow6, Xlgow6, Emgow6);  // ../RTL/cortexm0ds_logic.v(11680)
  and u13277 (n3644, Qtfow6, Tf4ju6);  // ../RTL/cortexm0ds_logic.v(11681)
  not u13278 (Emgow6, n3644);  // ../RTL/cortexm0ds_logic.v(11681)
  and u13279 (n3645, Lmgow6, Smgow6);  // ../RTL/cortexm0ds_logic.v(11682)
  and u1328 (n101[0], Rrzhu6, Yrzhu6);  // ../RTL/cortexm0ds_logic.v(3356)
  not u13280 (Tf4ju6, n3645);  // ../RTL/cortexm0ds_logic.v(11682)
  and u13281 (Smgow6, Zmgow6, Gngow6);  // ../RTL/cortexm0ds_logic.v(11683)
  or u13282 (Gngow6, Ipfow6, Na0iu6);  // ../RTL/cortexm0ds_logic.v(11684)
  or u13283 (Zmgow6, Rqfow6, Ua0iu6);  // ../RTL/cortexm0ds_logic.v(11685)
  and u13284 (Lmgow6, Nngow6, Ungow6);  // ../RTL/cortexm0ds_logic.v(11686)
  or u13285 (Ungow6, Ppfow6, Ib0iu6);  // ../RTL/cortexm0ds_logic.v(11687)
  or u13286 (Nngow6, Kqfow6, Bb0iu6);  // ../RTL/cortexm0ds_logic.v(11688)
  and u13287 (n3646, HRDATA[12], Q2eow6);  // ../RTL/cortexm0ds_logic.v(11689)
  not u13288 (Xlgow6, n3646);  // ../RTL/cortexm0ds_logic.v(11689)
  or u13289 (U2gow6, B0cow6, Qffow6);  // ../RTL/cortexm0ds_logic.v(11690)
  buf u1329 (K7hpw6[20], Fldbx6);  // ../RTL/cortexm0ds_logic.v(2366)
  and u13290 (B0cow6, Bogow6, Iogow6);  // ../RTL/cortexm0ds_logic.v(11691)
  and u13291 (Iogow6, Pogow6, Wogow6);  // ../RTL/cortexm0ds_logic.v(11692)
  and u13292 (n3647, Dyeow6, Cw3ju6);  // ../RTL/cortexm0ds_logic.v(11693)
  not u13293 (Wogow6, n3647);  // ../RTL/cortexm0ds_logic.v(11693)
  and u13294 (n3648, Dpgow6, Kpgow6);  // ../RTL/cortexm0ds_logic.v(11694)
  not u13295 (Cw3ju6, n3648);  // ../RTL/cortexm0ds_logic.v(11694)
  and u13296 (Kpgow6, Rpgow6, Ypgow6);  // ../RTL/cortexm0ds_logic.v(11695)
  or u13297 (Ypgow6, Ppfow6, B40iu6);  // ../RTL/cortexm0ds_logic.v(11696)
  or u13298 (Rpgow6, Ipfow6, Pb0iu6);  // ../RTL/cortexm0ds_logic.v(11697)
  and u13299 (Dpgow6, Fqgow6, Mqgow6);  // ../RTL/cortexm0ds_logic.v(11698)
  buf u133 (vis_r8_o[1], Pqrax6);  // ../RTL/cortexm0ds_logic.v(2579)
  buf u1330 (K7hpw6[21], M4ebx6);  // ../RTL/cortexm0ds_logic.v(2366)
  or u13300 (Mqgow6, Rqfow6, Wb0iu6);  // ../RTL/cortexm0ds_logic.v(11699)
  or u13301 (Fqgow6, Kqfow6, U30iu6);  // ../RTL/cortexm0ds_logic.v(11700)
  or u13302 (Pogow6, Iydow6, Yzqiu6);  // ../RTL/cortexm0ds_logic.v(11701)
  and u13303 (Yzqiu6, Tqgow6, Argow6);  // ../RTL/cortexm0ds_logic.v(11702)
  and u13304 (Argow6, Hrgow6, Orgow6);  // ../RTL/cortexm0ds_logic.v(11703)
  and u13305 (Orgow6, Vrgow6, Csgow6);  // ../RTL/cortexm0ds_logic.v(11704)
  and u13306 (n3649, Odgpw6[4], M0eow6);  // ../RTL/cortexm0ds_logic.v(11705)
  not u13307 (Csgow6, n3649);  // ../RTL/cortexm0ds_logic.v(11705)
  and u13308 (n3650, STCALIB[4], H1eow6);  // ../RTL/cortexm0ds_logic.v(11706)
  not u13309 (Vrgow6, n3650);  // ../RTL/cortexm0ds_logic.v(11706)
  buf u1331 (K7hpw6[22], Tjfbx6);  // ../RTL/cortexm0ds_logic.v(2366)
  and u13310 (Hrgow6, Jsgow6, Qsgow6);  // ../RTL/cortexm0ds_logic.v(11707)
  and u13311 (n3651, T7eow6, vis_ipsr_o[4]);  // ../RTL/cortexm0ds_logic.v(11708)
  not u13312 (Qsgow6, n3651);  // ../RTL/cortexm0ds_logic.v(11708)
  and u13313 (n3652, F0eow6, Vbgpw6[4]);  // ../RTL/cortexm0ds_logic.v(11709)
  not u13314 (Jsgow6, n3652);  // ../RTL/cortexm0ds_logic.v(11709)
  and u13315 (Tqgow6, Xsgow6, Etgow6);  // ../RTL/cortexm0ds_logic.v(11710)
  and u13316 (n3653, Fpgiu6, Gfghu6);  // ../RTL/cortexm0ds_logic.v(11711)
  not u13317 (Etgow6, n3653);  // ../RTL/cortexm0ds_logic.v(11711)
  and u13318 (Xsgow6, Ltgow6, Stgow6);  // ../RTL/cortexm0ds_logic.v(11712)
  and u13319 (n3654, Bagpw6[4], M6eiu6);  // ../RTL/cortexm0ds_logic.v(11713)
  buf u1332 (K7hpw6[23], Zvgbx6);  // ../RTL/cortexm0ds_logic.v(2366)
  not u13320 (Stgow6, n3654);  // ../RTL/cortexm0ds_logic.v(11713)
  and u13321 (n3655, Tzfpw6[4], Yvgiu6);  // ../RTL/cortexm0ds_logic.v(11714)
  not u13322 (Ltgow6, n3655);  // ../RTL/cortexm0ds_logic.v(11714)
  and u13323 (Bogow6, Ztgow6, Gugow6);  // ../RTL/cortexm0ds_logic.v(11715)
  and u13324 (n3656, Qtfow6, Sx3ju6);  // ../RTL/cortexm0ds_logic.v(11716)
  not u13325 (Gugow6, n3656);  // ../RTL/cortexm0ds_logic.v(11716)
  and u13326 (n3657, Nugow6, Uugow6);  // ../RTL/cortexm0ds_logic.v(11717)
  not u13327 (Sx3ju6, n3657);  // ../RTL/cortexm0ds_logic.v(11717)
  and u13328 (Uugow6, Bvgow6, Ivgow6);  // ../RTL/cortexm0ds_logic.v(11718)
  or u13329 (Ivgow6, Ipfow6, I40iu6);  // ../RTL/cortexm0ds_logic.v(11719)
  buf u1333 (K7hpw6[24], D99ax6);  // ../RTL/cortexm0ds_logic.v(2366)
  or u13330 (Bvgow6, Kqfow6, W40iu6);  // ../RTL/cortexm0ds_logic.v(11720)
  and u13331 (Nugow6, Pvgow6, Wvgow6);  // ../RTL/cortexm0ds_logic.v(11721)
  or u13332 (Wvgow6, Ppfow6, D50iu6);  // ../RTL/cortexm0ds_logic.v(11722)
  or u13333 (Pvgow6, Rqfow6, P40iu6);  // ../RTL/cortexm0ds_logic.v(11723)
  and u13334 (n3658, HRDATA[4], Q2eow6);  // ../RTL/cortexm0ds_logic.v(11724)
  not u13335 (Ztgow6, n3658);  // ../RTL/cortexm0ds_logic.v(11724)
  and u13336 (Tkfow6, Dwgow6, Kwgow6);  // ../RTL/cortexm0ds_logic.v(11725)
  and u13337 (n3659, Zsfpw6[3], Cmziu6);  // ../RTL/cortexm0ds_logic.v(11726)
  not u13338 (Kwgow6, n3659);  // ../RTL/cortexm0ds_logic.v(11726)
  and u13339 (n3660, vis_pc_o[3], Jmziu6);  // ../RTL/cortexm0ds_logic.v(11727)
  buf u1334 (K7hpw6[25], G79ax6);  // ../RTL/cortexm0ds_logic.v(2366)
  not u13340 (Dwgow6, n3660);  // ../RTL/cortexm0ds_logic.v(11727)
  and u13341 (n3661, Rwgow6, Ywgow6);  // ../RTL/cortexm0ds_logic.v(11728)
  not u13342 (Vjohu6, n3661);  // ../RTL/cortexm0ds_logic.v(11728)
  and u13343 (Ywgow6, Fxgow6, Mxgow6);  // ../RTL/cortexm0ds_logic.v(11729)
  and u13344 (n3662, Egziu6, Eafpw6[3]);  // ../RTL/cortexm0ds_logic.v(11730)
  not u13345 (Mxgow6, n3662);  // ../RTL/cortexm0ds_logic.v(11730)
  and u13346 (Fxgow6, Txgow6, Sgziu6);  // ../RTL/cortexm0ds_logic.v(11731)
  or u13347 (Txgow6, Ft6ow6, Kifiu6);  // ../RTL/cortexm0ds_logic.v(11732)
  and u13348 (Kifiu6, Aygow6, Hygow6);  // ../RTL/cortexm0ds_logic.v(11733)
  and u13349 (Hygow6, Oygow6, Vygow6);  // ../RTL/cortexm0ds_logic.v(11734)
  buf u1335 (K7hpw6[26], Facbx6);  // ../RTL/cortexm0ds_logic.v(2366)
  or u13350 (Vygow6, Cfliu6, Ahcow6);  // ../RTL/cortexm0ds_logic.v(11735)
  and u13351 (Oygow6, Czgow6, Mdliu6);  // ../RTL/cortexm0ds_logic.v(11736)
  or u13352 (Czgow6, Iqeow6, Yfcow6);  // ../RTL/cortexm0ds_logic.v(11737)
  and u13353 (Aygow6, Jzgow6, Qzgow6);  // ../RTL/cortexm0ds_logic.v(11738)
  or u13354 (Qzgow6, Ycliu6, Tgcow6);  // ../RTL/cortexm0ds_logic.v(11739)
  or u13355 (Jzgow6, Qffow6, Kfcow6);  // ../RTL/cortexm0ds_logic.v(11740)
  and u13356 (Rwgow6, Xzgow6, E0how6);  // ../RTL/cortexm0ds_logic.v(11741)
  and u13357 (n3663, Zsfpw6[2], Cmziu6);  // ../RTL/cortexm0ds_logic.v(11742)
  not u13358 (E0how6, n3663);  // ../RTL/cortexm0ds_logic.v(11742)
  and u13359 (n3664, vis_pc_o[2], Jmziu6);  // ../RTL/cortexm0ds_logic.v(11743)
  and u1336 (n109, Htzhu6, Otzhu6);  // ../RTL/cortexm0ds_logic.v(3375)
  not u13360 (Xzgow6, n3664);  // ../RTL/cortexm0ds_logic.v(11743)
  and u13361 (n3665, L0how6, S0how6);  // ../RTL/cortexm0ds_logic.v(11744)
  not u13362 (Ojohu6, n3665);  // ../RTL/cortexm0ds_logic.v(11744)
  and u13363 (S0how6, Z0how6, G1how6);  // ../RTL/cortexm0ds_logic.v(11745)
  and u13364 (n3666, Egziu6, Eafpw6[2]);  // ../RTL/cortexm0ds_logic.v(11746)
  not u13365 (G1how6, n3666);  // ../RTL/cortexm0ds_logic.v(11746)
  and u13366 (Z0how6, N1how6, Sgziu6);  // ../RTL/cortexm0ds_logic.v(11747)
  or u13367 (N1how6, Ft6ow6, Ogciu6);  // ../RTL/cortexm0ds_logic.v(11748)
  and u13368 (Ogciu6, U1how6, B2how6);  // ../RTL/cortexm0ds_logic.v(11749)
  and u13369 (B2how6, I2how6, P2how6);  // ../RTL/cortexm0ds_logic.v(11750)
  not u1337 (R0ghu6, n109);  // ../RTL/cortexm0ds_logic.v(3375)
  or u13370 (P2how6, Cfliu6, Wlcow6);  // ../RTL/cortexm0ds_logic.v(11751)
  and u13371 (Cfliu6, W2how6, D3how6);  // ../RTL/cortexm0ds_logic.v(11752)
  or u13372 (D3how6, K3how6, R3how6);  // ../RTL/cortexm0ds_logic.v(11753)
  and u13373 (W2how6, Y3how6, F4how6);  // ../RTL/cortexm0ds_logic.v(11754)
  and u13374 (n3667, M4how6, T4how6);  // ../RTL/cortexm0ds_logic.v(11755)
  not u13375 (Y3how6, n3667);  // ../RTL/cortexm0ds_logic.v(11755)
  or u13376 (n3668, Iwfpw6[0], Y7ghu6);  // ../RTL/cortexm0ds_logic.v(11756)
  not u13377 (M4how6, n3668);  // ../RTL/cortexm0ds_logic.v(11756)
  and u13378 (I2how6, A5how6, Mdliu6);  // ../RTL/cortexm0ds_logic.v(11757)
  and u13379 (n3669, H5how6, O5how6);  // ../RTL/cortexm0ds_logic.v(11758)
  and u1338 (n110, Vtzhu6, Cuzhu6);  // ../RTL/cortexm0ds_logic.v(3376)
  not u13380 (Mdliu6, n3669);  // ../RTL/cortexm0ds_logic.v(11758)
  and u13381 (n3670, V5how6, C6how6);  // ../RTL/cortexm0ds_logic.v(11759)
  not u13382 (O5how6, n3670);  // ../RTL/cortexm0ds_logic.v(11759)
  and u13383 (n3671, J6how6, Q6how6);  // ../RTL/cortexm0ds_logic.v(11760)
  not u13384 (V5how6, n3671);  // ../RTL/cortexm0ds_logic.v(11760)
  and u13385 (Q6how6, Ny3ju6, Tucow6);  // ../RTL/cortexm0ds_logic.v(11761)
  and u13386 (J6how6, Z44ju6, X6how6);  // ../RTL/cortexm0ds_logic.v(11762)
  or u13387 (Z44ju6, R3how6, E7how6);  // ../RTL/cortexm0ds_logic.v(11763)
  and u13388 (E7how6, Avcow6, L7how6);  // ../RTL/cortexm0ds_logic.v(11764)
  or u13389 (A5how6, Iqeow6, Ukcow6);  // ../RTL/cortexm0ds_logic.v(11765)
  not u1339 (Otzhu6, n110);  // ../RTL/cortexm0ds_logic.v(3376)
  and u13390 (Iqeow6, S7how6, Z7how6);  // ../RTL/cortexm0ds_logic.v(11767)
  not u13391 (Qfliu6, Iqeow6);  // ../RTL/cortexm0ds_logic.v(11767)
  and u13392 (n3672, G8how6, Iwfpw6[1]);  // ../RTL/cortexm0ds_logic.v(11768)
  not u13393 (Z7how6, n3672);  // ../RTL/cortexm0ds_logic.v(11768)
  and u13394 (S7how6, N8how6, Dtcow6);  // ../RTL/cortexm0ds_logic.v(11769)
  or u13395 (N8how6, X6how6, Ktcow6);  // ../RTL/cortexm0ds_logic.v(11770)
  and u13396 (U1how6, U8how6, B9how6);  // ../RTL/cortexm0ds_logic.v(11771)
  or u13397 (B9how6, Ycliu6, Plcow6);  // ../RTL/cortexm0ds_logic.v(11772)
  and u13398 (Ycliu6, I9how6, P9how6);  // ../RTL/cortexm0ds_logic.v(11773)
  and u13399 (P9how6, W9how6, Dahow6);  // ../RTL/cortexm0ds_logic.v(11774)
  buf u134 (vis_r8_o[29], Kmjpw6);  // ../RTL/cortexm0ds_logic.v(2579)
  or u1340 (Htzhu6, Juzhu6, Quzhu6);  // ../RTL/cortexm0ds_logic.v(3377)
  and u13400 (I9how6, Kahow6, Rahow6);  // ../RTL/cortexm0ds_logic.v(11775)
  and u13401 (n3673, G8how6, Yahow6);  // ../RTL/cortexm0ds_logic.v(11776)
  not u13402 (Kahow6, n3673);  // ../RTL/cortexm0ds_logic.v(11776)
  and u13403 (G8how6, Fbhow6, Mbhow6);  // ../RTL/cortexm0ds_logic.v(11777)
  or u13404 (n3674, Cyfpw6[1], Y7ghu6);  // ../RTL/cortexm0ds_logic.v(11778)
  not u13405 (Mbhow6, n3674);  // ../RTL/cortexm0ds_logic.v(11778)
  or u13406 (n3675, Tbhow6, Tucow6);  // ../RTL/cortexm0ds_logic.v(11779)
  not u13407 (Fbhow6, n3675);  // ../RTL/cortexm0ds_logic.v(11779)
  not u13408 (Tbhow6, Iwfpw6[0]);  // ../RTL/cortexm0ds_logic.v(11780)
  or u13409 (U8how6, Qffow6, Gkcow6);  // ../RTL/cortexm0ds_logic.v(11781)
  buf u1341 (vis_apsr_o[1], Qijpw6);  // ../RTL/cortexm0ds_logic.v(1880)
  and u13410 (Qffow6, Eccow6, Achow6);  // ../RTL/cortexm0ds_logic.v(11783)
  not u13411 (Aeliu6, Qffow6);  // ../RTL/cortexm0ds_logic.v(11783)
  and u13412 (n3676, Ktcow6, Hchow6);  // ../RTL/cortexm0ds_logic.v(11784)
  not u13413 (Achow6, n3676);  // ../RTL/cortexm0ds_logic.v(11784)
  and u13414 (n3677, Ochow6, Vchow6);  // ../RTL/cortexm0ds_logic.v(11785)
  not u13415 (Hchow6, n3677);  // ../RTL/cortexm0ds_logic.v(11785)
  and u13416 (Vchow6, Cdhow6, Eu0iu6);  // ../RTL/cortexm0ds_logic.v(11786)
  not u13417 (Eu0iu6, Jdhow6);  // ../RTL/cortexm0ds_logic.v(11787)
  and u13418 (n3678, Qdhow6, Xdhow6);  // ../RTL/cortexm0ds_logic.v(11788)
  not u13419 (Cdhow6, n3678);  // ../RTL/cortexm0ds_logic.v(11788)
  buf u1342 (vis_r6_o[21], E7pax6);  // ../RTL/cortexm0ds_logic.v(2523)
  and u13420 (n3679, Cyfpw6[1], Eehow6);  // ../RTL/cortexm0ds_logic.v(11789)
  not u13421 (Xdhow6, n3679);  // ../RTL/cortexm0ds_logic.v(11789)
  or u13422 (Eehow6, Cyfpw6[0], Cyfpw6[3]);  // ../RTL/cortexm0ds_logic.v(11790)
  or u13423 (Phnow6, Iwfpw6[0], Iwfpw6[1]);  // ../RTL/cortexm0ds_logic.v(11791)
  not u13424 (Qdhow6, Phnow6);  // ../RTL/cortexm0ds_logic.v(11791)
  and u13425 (Ochow6, Cyfpw6[5], Lehow6);  // ../RTL/cortexm0ds_logic.v(11792)
  or u13426 (Lehow6, Nlaiu6, Tfjiu6);  // ../RTL/cortexm0ds_logic.v(11793)
  and u13427 (L0how6, Sehow6, Zehow6);  // ../RTL/cortexm0ds_logic.v(11794)
  and u13428 (n3680, Zsfpw6[1], Cmziu6);  // ../RTL/cortexm0ds_logic.v(11795)
  not u13429 (Zehow6, n3680);  // ../RTL/cortexm0ds_logic.v(11795)
  buf u1343 (vis_apsr_o[2], Bfjpw6);  // ../RTL/cortexm0ds_logic.v(1880)
  or u13430 (Sehow6, Quzhu6, Ar8iu6);  // ../RTL/cortexm0ds_logic.v(11796)
  not u13431 (Quzhu6, vis_pc_o[1]);  // ../RTL/cortexm0ds_logic.v(11797)
  and u13432 (n3681, Gfhow6, Nfhow6);  // ../RTL/cortexm0ds_logic.v(11798)
  not u13433 (Hjohu6, n3681);  // ../RTL/cortexm0ds_logic.v(11798)
  and u13434 (n3682, Ufhow6, Ophiu6);  // ../RTL/cortexm0ds_logic.v(11799)
  not u13435 (Nfhow6, n3682);  // ../RTL/cortexm0ds_logic.v(11799)
  and u13436 (n3683, Juzhu6, Bghow6);  // ../RTL/cortexm0ds_logic.v(11800)
  not u13437 (Ufhow6, n3683);  // ../RTL/cortexm0ds_logic.v(11800)
  or u13438 (Bghow6, N6piu6, Eh6iu6);  // ../RTL/cortexm0ds_logic.v(11801)
  and u13439 (n3684, Sufpw6[1], Eh6iu6);  // ../RTL/cortexm0ds_logic.v(11802)
  buf u1344 (vis_r6_o[22], T7fbx6);  // ../RTL/cortexm0ds_logic.v(2523)
  not u13440 (Gfhow6, n3684);  // ../RTL/cortexm0ds_logic.v(11802)
  not u13441 (Ajohu6, Ighow6);  // ../RTL/cortexm0ds_logic.v(11803)
  AL_MUX u13442 (
    .i0(Sijiu6),
    .i1(X5phu6),
    .sel(F2biu6),
    .o(Ighow6));  // ../RTL/cortexm0ds_logic.v(11804)
  or u13443 (n3685, Eh6iu6, K9aiu6);  // ../RTL/cortexm0ds_logic.v(11805)
  not u13444 (F2biu6, n3685);  // ../RTL/cortexm0ds_logic.v(11805)
  and u13445 (n3686, Ivfhu6, Pghow6);  // ../RTL/cortexm0ds_logic.v(11806)
  not u13446 (X5phu6, n3686);  // ../RTL/cortexm0ds_logic.v(11806)
  and u13447 (n3687, Wghow6, Dhhow6);  // ../RTL/cortexm0ds_logic.v(11807)
  not u13448 (Pghow6, n3687);  // ../RTL/cortexm0ds_logic.v(11807)
  and u13449 (Dhhow6, Khhow6, Rhhow6);  // ../RTL/cortexm0ds_logic.v(11808)
  buf u1345 (vis_apsr_o[3], Arnpw6);  // ../RTL/cortexm0ds_logic.v(1880)
  or u13450 (n3688, Ppfpw6[8], Ppfpw6[9]);  // ../RTL/cortexm0ds_logic.v(11809)
  not u13451 (Rhhow6, n3688);  // ../RTL/cortexm0ds_logic.v(11809)
  or u13452 (n3689, Ppfpw6[6], Ppfpw6[7]);  // ../RTL/cortexm0ds_logic.v(11810)
  not u13453 (Khhow6, n3689);  // ../RTL/cortexm0ds_logic.v(11810)
  and u13454 (Wghow6, Yhhow6, Fihow6);  // ../RTL/cortexm0ds_logic.v(11811)
  or u13455 (n3690, Ppfpw6[12], Ppfpw6[13]);  // ../RTL/cortexm0ds_logic.v(11812)
  not u13456 (Fihow6, n3690);  // ../RTL/cortexm0ds_logic.v(11812)
  or u13457 (n3691, Ppfpw6[10], Ppfpw6[11]);  // ../RTL/cortexm0ds_logic.v(11813)
  not u13458 (Yhhow6, n3691);  // ../RTL/cortexm0ds_logic.v(11813)
  AL_MUX u13459 (
    .i0(Mihow6),
    .i1(T6ehu6),
    .sel(Eh6iu6),
    .o(Tiohu6));  // ../RTL/cortexm0ds_logic.v(11814)
  buf u1346 (vis_r6_o[23], Kfoax6);  // ../RTL/cortexm0ds_logic.v(2523)
  and u13460 (n3692, Tihow6, Ajhow6);  // ../RTL/cortexm0ds_logic.v(11815)
  not u13461 (Mihow6, n3692);  // ../RTL/cortexm0ds_logic.v(11815)
  and u13462 (n3693, H4oiu6, Hjhow6);  // ../RTL/cortexm0ds_logic.v(11816)
  not u13463 (Ajhow6, n3693);  // ../RTL/cortexm0ds_logic.v(11816)
  or u13464 (n3694, Xkaow6, R75iu6);  // ../RTL/cortexm0ds_logic.v(11817)
  not u13465 (Hjhow6, n3694);  // ../RTL/cortexm0ds_logic.v(11817)
  or u13466 (n3695, K9bow6, G7oiu6);  // ../RTL/cortexm0ds_logic.v(11818)
  not u13467 (H4oiu6, n3695);  // ../RTL/cortexm0ds_logic.v(11818)
  and u13468 (n3696, Ojhow6, Vjhow6);  // ../RTL/cortexm0ds_logic.v(11819)
  not u13469 (Tihow6, n3696);  // ../RTL/cortexm0ds_logic.v(11819)
  buf u1347 (Dhgpw6[1], Xnbax6);  // ../RTL/cortexm0ds_logic.v(2280)
  or u13470 (n3697, P1bow6, Y2oiu6);  // ../RTL/cortexm0ds_logic.v(11820)
  not u13471 (Ojhow6, n3697);  // ../RTL/cortexm0ds_logic.v(11820)
  or u13472 (Miohu6, Ckhow6, Jkhow6);  // ../RTL/cortexm0ds_logic.v(11821)
  or u13473 (n3698, Qkhow6, Dk7ow6);  // ../RTL/cortexm0ds_logic.v(11822)
  not u13474 (Jkhow6, n3698);  // ../RTL/cortexm0ds_logic.v(11822)
  not u13475 (Qkhow6, Xkhow6);  // ../RTL/cortexm0ds_logic.v(11823)
  AL_MUX u13476 (
    .i0(Elhow6),
    .i1(S8fpw6[7]),
    .sel(Rk7ow6),
    .o(Ckhow6));  // ../RTL/cortexm0ds_logic.v(11824)
  and u13477 (n3699, Llhow6, Slhow6);  // ../RTL/cortexm0ds_logic.v(11825)
  not u13478 (Elhow6, n3699);  // ../RTL/cortexm0ds_logic.v(11825)
  and u13479 (n3700, D7fpw6[7], Zlhow6);  // ../RTL/cortexm0ds_logic.v(11826)
  buf u1348 (vis_r6_o[24], Fvoax6);  // ../RTL/cortexm0ds_logic.v(2523)
  not u13480 (Slhow6, n3700);  // ../RTL/cortexm0ds_logic.v(11826)
  or u13481 (Llhow6, Ad8iu6, Cn7ow6);  // ../RTL/cortexm0ds_logic.v(11827)
  AL_MUX u13482 (
    .i0(W7cow6),
    .i1(Dxfhu6),
    .sel(Eh6iu6),
    .o(Fiohu6));  // ../RTL/cortexm0ds_logic.v(11828)
  AL_MUX u13483 (
    .i0(Wz4iu6),
    .i1(Hrfpw6[16]),
    .sel(Qqhiu6),
    .o(Yhohu6));  // ../RTL/cortexm0ds_logic.v(11829)
  and u13484 (n3701, Gmhow6, Nmhow6);  // ../RTL/cortexm0ds_logic.v(11830)
  not u13485 (Rhohu6, n3701);  // ../RTL/cortexm0ds_logic.v(11830)
  and u13486 (n3702, Umhow6, HRDATA[16]);  // ../RTL/cortexm0ds_logic.v(11831)
  not u13487 (Nmhow6, n3702);  // ../RTL/cortexm0ds_logic.v(11831)
  and u13488 (n3703, Hrfpw6[0], Qqhiu6);  // ../RTL/cortexm0ds_logic.v(11832)
  not u13489 (Gmhow6, n3703);  // ../RTL/cortexm0ds_logic.v(11832)
  buf u1349 (Dhgpw6[2], Rkbax6);  // ../RTL/cortexm0ds_logic.v(2280)
  and u13490 (n3704, Bnhow6, Inhow6);  // ../RTL/cortexm0ds_logic.v(11833)
  not u13491 (Khohu6, n3704);  // ../RTL/cortexm0ds_logic.v(11833)
  and u13492 (n3705, Umhow6, HRDATA[31]);  // ../RTL/cortexm0ds_logic.v(11834)
  not u13493 (Inhow6, n3705);  // ../RTL/cortexm0ds_logic.v(11834)
  and u13494 (n3706, Hrfpw6[15], Qqhiu6);  // ../RTL/cortexm0ds_logic.v(11835)
  not u13495 (Bnhow6, n3706);  // ../RTL/cortexm0ds_logic.v(11835)
  and u13496 (n3707, Pnhow6, Wnhow6);  // ../RTL/cortexm0ds_logic.v(11836)
  not u13497 (Dhohu6, n3707);  // ../RTL/cortexm0ds_logic.v(11836)
  and u13498 (n3708, Umhow6, HRDATA[29]);  // ../RTL/cortexm0ds_logic.v(11837)
  not u13499 (Wnhow6, n3708);  // ../RTL/cortexm0ds_logic.v(11837)
  buf u135 (Uthpw6[20], Cydbx6);  // ../RTL/cortexm0ds_logic.v(1882)
  buf u1350 (vis_r6_o[25], E5pax6);  // ../RTL/cortexm0ds_logic.v(2523)
  and u13500 (n3709, Hrfpw6[13], Qqhiu6);  // ../RTL/cortexm0ds_logic.v(11838)
  not u13501 (Pnhow6, n3709);  // ../RTL/cortexm0ds_logic.v(11838)
  and u13502 (n3710, Dohow6, Kohow6);  // ../RTL/cortexm0ds_logic.v(11839)
  not u13503 (Wgohu6, n3710);  // ../RTL/cortexm0ds_logic.v(11839)
  and u13504 (n3711, Umhow6, HRDATA[28]);  // ../RTL/cortexm0ds_logic.v(11840)
  not u13505 (Kohow6, n3711);  // ../RTL/cortexm0ds_logic.v(11840)
  and u13506 (n3712, Hrfpw6[12], Qqhiu6);  // ../RTL/cortexm0ds_logic.v(11841)
  not u13507 (Dohow6, n3712);  // ../RTL/cortexm0ds_logic.v(11841)
  and u13508 (n3713, Rohow6, Yohow6);  // ../RTL/cortexm0ds_logic.v(11842)
  not u13509 (Pgohu6, n3713);  // ../RTL/cortexm0ds_logic.v(11842)
  buf u1351 (Dhgpw6[3], Thiax6);  // ../RTL/cortexm0ds_logic.v(2280)
  and u13510 (n3714, Umhow6, HRDATA[27]);  // ../RTL/cortexm0ds_logic.v(11843)
  not u13511 (Yohow6, n3714);  // ../RTL/cortexm0ds_logic.v(11843)
  and u13512 (n3715, Hrfpw6[11], Qqhiu6);  // ../RTL/cortexm0ds_logic.v(11844)
  not u13513 (Rohow6, n3715);  // ../RTL/cortexm0ds_logic.v(11844)
  and u13514 (n3716, Fphow6, Mphow6);  // ../RTL/cortexm0ds_logic.v(11845)
  not u13515 (Igohu6, n3716);  // ../RTL/cortexm0ds_logic.v(11845)
  and u13516 (n3717, Umhow6, HRDATA[26]);  // ../RTL/cortexm0ds_logic.v(11846)
  not u13517 (Mphow6, n3717);  // ../RTL/cortexm0ds_logic.v(11846)
  and u13518 (n3718, Hrfpw6[10], Qqhiu6);  // ../RTL/cortexm0ds_logic.v(11847)
  not u13519 (Fphow6, n3718);  // ../RTL/cortexm0ds_logic.v(11847)
  buf u1352 (vis_r6_o[26], Fxoax6);  // ../RTL/cortexm0ds_logic.v(2523)
  and u13520 (n3719, Tphow6, Aqhow6);  // ../RTL/cortexm0ds_logic.v(11848)
  not u13521 (Bgohu6, n3719);  // ../RTL/cortexm0ds_logic.v(11848)
  and u13522 (n3720, Umhow6, HRDATA[25]);  // ../RTL/cortexm0ds_logic.v(11849)
  not u13523 (Aqhow6, n3720);  // ../RTL/cortexm0ds_logic.v(11849)
  and u13524 (n3721, Hrfpw6[9], Qqhiu6);  // ../RTL/cortexm0ds_logic.v(11850)
  not u13525 (Tphow6, n3721);  // ../RTL/cortexm0ds_logic.v(11850)
  and u13526 (n3722, Hqhow6, Oqhow6);  // ../RTL/cortexm0ds_logic.v(11851)
  not u13527 (Ufohu6, n3722);  // ../RTL/cortexm0ds_logic.v(11851)
  and u13528 (n3723, Umhow6, HRDATA[24]);  // ../RTL/cortexm0ds_logic.v(11852)
  not u13529 (Oqhow6, n3723);  // ../RTL/cortexm0ds_logic.v(11852)
  buf u1353 (Dhgpw6[4], Hmbax6);  // ../RTL/cortexm0ds_logic.v(2280)
  and u13530 (n3724, Hrfpw6[8], Qqhiu6);  // ../RTL/cortexm0ds_logic.v(11853)
  not u13531 (Hqhow6, n3724);  // ../RTL/cortexm0ds_logic.v(11853)
  and u13532 (n3725, Vqhow6, Crhow6);  // ../RTL/cortexm0ds_logic.v(11854)
  not u13533 (Nfohu6, n3725);  // ../RTL/cortexm0ds_logic.v(11854)
  and u13534 (n3726, Umhow6, HRDATA[23]);  // ../RTL/cortexm0ds_logic.v(11855)
  not u13535 (Crhow6, n3726);  // ../RTL/cortexm0ds_logic.v(11855)
  and u13536 (n3727, Hrfpw6[7], Qqhiu6);  // ../RTL/cortexm0ds_logic.v(11856)
  not u13537 (Vqhow6, n3727);  // ../RTL/cortexm0ds_logic.v(11856)
  AL_MUX u13538 (
    .i0(Jrhow6),
    .i1(H2fpw6[3]),
    .sel(G81ju6),
    .o(Gfohu6));  // ../RTL/cortexm0ds_logic.v(11857)
  and u13539 (n3728, HREADY, Qrhow6);  // ../RTL/cortexm0ds_logic.v(11858)
  buf u1354 (vis_r6_o[27], Fzoax6);  // ../RTL/cortexm0ds_logic.v(2523)
  not u13540 (G81ju6, n3728);  // ../RTL/cortexm0ds_logic.v(11858)
  and u13541 (n3729, Xrhow6, Eshow6);  // ../RTL/cortexm0ds_logic.v(11859)
  not u13542 (Qrhow6, n3729);  // ../RTL/cortexm0ds_logic.v(11859)
  and u13543 (Eshow6, Lshow6, Sshow6);  // ../RTL/cortexm0ds_logic.v(11860)
  and u13544 (Sshow6, Zshow6, Gthow6);  // ../RTL/cortexm0ds_logic.v(11861)
  and u13545 (n3730, Nthow6, Lraiu6);  // ../RTL/cortexm0ds_logic.v(11862)
  not u13546 (Gthow6, n3730);  // ../RTL/cortexm0ds_logic.v(11862)
  and u13547 (Nthow6, Uu9ow6, Uthow6);  // ../RTL/cortexm0ds_logic.v(11863)
  and u13548 (n3731, D7fpw6[15], Buhow6);  // ../RTL/cortexm0ds_logic.v(11864)
  not u13549 (Uthow6, n3731);  // ../RTL/cortexm0ds_logic.v(11864)
  buf u1355 (Ppfpw6[0], Xdspw6);  // ../RTL/cortexm0ds_logic.v(2461)
  and u13550 (n3732, Iuhow6, Bkjiu6);  // ../RTL/cortexm0ds_logic.v(11865)
  not u13551 (Buhow6, n3732);  // ../RTL/cortexm0ds_logic.v(11865)
  or u13552 (Iuhow6, Rg2ju6, D7fpw6[3]);  // ../RTL/cortexm0ds_logic.v(11866)
  not u13553 (Uu9ow6, X5aiu6);  // ../RTL/cortexm0ds_logic.v(11867)
  or u13554 (X5aiu6, Puhow6, Ttciu6);  // ../RTL/cortexm0ds_logic.v(11868)
  not u13555 (Ttciu6, T0hhu6);  // ../RTL/cortexm0ds_logic.v(11869)
  or u13556 (Puhow6, E45iu6, Ii0iu6);  // ../RTL/cortexm0ds_logic.v(11870)
  not u13557 (E45iu6, N20ju6);  // ../RTL/cortexm0ds_logic.v(11871)
  and u13558 (n3733, Wuhow6, Vviiu6);  // ../RTL/cortexm0ds_logic.v(11872)
  not u13559 (Zshow6, n3733);  // ../RTL/cortexm0ds_logic.v(11872)
  not u1356 (Mifpw6[0], n112[0]);  // ../RTL/cortexm0ds_logic.v(3417)
  or u13560 (n3734, D7fpw6[10], D7fpw6[8]);  // ../RTL/cortexm0ds_logic.v(11873)
  not u13561 (Wuhow6, n3734);  // ../RTL/cortexm0ds_logic.v(11873)
  and u13562 (Lshow6, Dvhow6, Kvhow6);  // ../RTL/cortexm0ds_logic.v(11874)
  and u13563 (n3735, Y31ju6, Rvhow6);  // ../RTL/cortexm0ds_logic.v(11875)
  not u13564 (Kvhow6, n3735);  // ../RTL/cortexm0ds_logic.v(11875)
  and u13565 (n3736, Yvhow6, Fwhow6);  // ../RTL/cortexm0ds_logic.v(11876)
  not u13566 (Rvhow6, n3736);  // ../RTL/cortexm0ds_logic.v(11876)
  and u13567 (Fwhow6, Mwhow6, Twhow6);  // ../RTL/cortexm0ds_logic.v(11877)
  and u13568 (n3737, Axhow6, Ftjiu6);  // ../RTL/cortexm0ds_logic.v(11878)
  not u13569 (Twhow6, n3737);  // ../RTL/cortexm0ds_logic.v(11878)
  buf u1357 (Iahpw6[10], Gw6bx6);  // ../RTL/cortexm0ds_logic.v(1883)
  and u13570 (n3738, N38ow6, Hxhow6);  // ../RTL/cortexm0ds_logic.v(11879)
  not u13571 (Axhow6, n3738);  // ../RTL/cortexm0ds_logic.v(11879)
  and u13572 (n3739, C0ehu6, An6ow6);  // ../RTL/cortexm0ds_logic.v(11880)
  not u13573 (Hxhow6, n3739);  // ../RTL/cortexm0ds_logic.v(11880)
  or u13574 (An6ow6, D7fpw6[11], D7fpw6[7]);  // ../RTL/cortexm0ds_logic.v(11881)
  or u13575 (n3740, Oxhow6, Evyiu6);  // ../RTL/cortexm0ds_logic.v(11882)
  not u13576 (Mwhow6, n3740);  // ../RTL/cortexm0ds_logic.v(11882)
  and u13577 (Oxhow6, Quyiu6, Ejiiu6);  // ../RTL/cortexm0ds_logic.v(11883)
  and u13578 (Ejiiu6, C0ehu6, D7fpw6[12]);  // ../RTL/cortexm0ds_logic.v(11884)
  or u13579 (n3741, X1ziu6, D7fpw6[11]);  // ../RTL/cortexm0ds_logic.v(11885)
  buf u1358 (Cjhpw6[3], J0gax6);  // ../RTL/cortexm0ds_logic.v(2365)
  not u13580 (Quyiu6, n3741);  // ../RTL/cortexm0ds_logic.v(11885)
  and u13581 (Yvhow6, Vxhow6, Cyhow6);  // ../RTL/cortexm0ds_logic.v(11886)
  or u13582 (Cyhow6, S80ju6, D7fpw6[8]);  // ../RTL/cortexm0ds_logic.v(11887)
  not u13583 (S80ju6, P0piu6);  // ../RTL/cortexm0ds_logic.v(11888)
  or u13584 (Vxhow6, Yb9ow6, Qxoiu6);  // ../RTL/cortexm0ds_logic.v(11889)
  and u13585 (n3742, P0piu6, W0piu6);  // ../RTL/cortexm0ds_logic.v(11891)
  not u13586 (Dvhow6, n3742);  // ../RTL/cortexm0ds_logic.v(11891)
  and u13587 (Xrhow6, Jyhow6, M1jiu6);  // ../RTL/cortexm0ds_logic.v(11892)
  and u13588 (M1jiu6, Qyhow6, Xyhow6);  // ../RTL/cortexm0ds_logic.v(11893)
  or u13589 (n3743, Ezhow6, Wkjiu6);  // ../RTL/cortexm0ds_logic.v(11894)
  buf u1359 (L1gpw6[1], Gz6ax6);  // ../RTL/cortexm0ds_logic.v(2191)
  not u13590 (Xyhow6, n3743);  // ../RTL/cortexm0ds_logic.v(11894)
  and u13591 (Wkjiu6, Lzhow6, Y31ju6);  // ../RTL/cortexm0ds_logic.v(11895)
  and u13592 (Qyhow6, Szhow6, Zzhow6);  // ../RTL/cortexm0ds_logic.v(11896)
  and u13593 (n3744, Hviiu6, G0iow6);  // ../RTL/cortexm0ds_logic.v(11897)
  not u13594 (Zzhow6, n3744);  // ../RTL/cortexm0ds_logic.v(11897)
  and u13595 (n3745, O7ziu6, Zt9ow6);  // ../RTL/cortexm0ds_logic.v(11898)
  not u13596 (G0iow6, n3745);  // ../RTL/cortexm0ds_logic.v(11898)
  or u13597 (Zt9ow6, Od0ju6, L01ju6);  // ../RTL/cortexm0ds_logic.v(11899)
  not u13598 (Od0ju6, Sdbow6);  // ../RTL/cortexm0ds_logic.v(11900)
  and u13599 (Sdbow6, Jwiiu6, Ndiiu6);  // ../RTL/cortexm0ds_logic.v(11901)
  buf u136 (E1hpw6[8], Vlaax6);  // ../RTL/cortexm0ds_logic.v(2367)
  buf u1360 (vis_r6_o[28], Rlibx6);  // ../RTL/cortexm0ds_logic.v(2523)
  not u13600 (Ndiiu6, D7fpw6[8]);  // ../RTL/cortexm0ds_logic.v(11902)
  and u13601 (Jwiiu6, D7fpw6[9], I6jiu6);  // ../RTL/cortexm0ds_logic.v(11903)
  not u13602 (O7ziu6, Db0ju6);  // ../RTL/cortexm0ds_logic.v(11904)
  and u13603 (n3746, Wliiu6, W0piu6);  // ../RTL/cortexm0ds_logic.v(11905)
  not u13604 (Szhow6, n3746);  // ../RTL/cortexm0ds_logic.v(11905)
  and u13605 (Jyhow6, Onjiu6, N0iow6);  // ../RTL/cortexm0ds_logic.v(11906)
  or u13606 (N0iow6, Jojiu6, Cyfpw6[7]);  // ../RTL/cortexm0ds_logic.v(11907)
  or u13607 (Onjiu6, Yn2ju6, Kq0iu6);  // ../RTL/cortexm0ds_logic.v(11908)
  and u13608 (n3747, Ir6ow6, U0iow6);  // ../RTL/cortexm0ds_logic.v(11909)
  not u13609 (Jrhow6, n3747);  // ../RTL/cortexm0ds_logic.v(11909)
  buf u1361 (Iahpw6[11], Wq8ax6);  // ../RTL/cortexm0ds_logic.v(1883)
  and u13610 (n3748, D7fpw6[7], B1iow6);  // ../RTL/cortexm0ds_logic.v(11910)
  not u13611 (U0iow6, n3748);  // ../RTL/cortexm0ds_logic.v(11910)
  and u13612 (n3749, Uvziu6, I1iow6);  // ../RTL/cortexm0ds_logic.v(11911)
  not u13613 (B1iow6, n3749);  // ../RTL/cortexm0ds_logic.v(11911)
  and u13614 (n3750, Srbow6, D7fpw6[10]);  // ../RTL/cortexm0ds_logic.v(11912)
  not u13615 (I1iow6, n3750);  // ../RTL/cortexm0ds_logic.v(11912)
  and u13616 (Ir6ow6, P1iow6, W1iow6);  // ../RTL/cortexm0ds_logic.v(11913)
  and u13617 (W1iow6, D2iow6, K2iow6);  // ../RTL/cortexm0ds_logic.v(11914)
  and u13618 (n3751, Y7ghu6, R2iow6);  // ../RTL/cortexm0ds_logic.v(11915)
  not u13619 (K2iow6, n3751);  // ../RTL/cortexm0ds_logic.v(11915)
  buf u1362 (vis_r6_o[1], F3pax6);  // ../RTL/cortexm0ds_logic.v(2523)
  or u13620 (R2iow6, Ii0iu6, D7fpw6[3]);  // ../RTL/cortexm0ds_logic.v(11916)
  and u13621 (D2iow6, Y2iow6, Faaiu6);  // ../RTL/cortexm0ds_logic.v(11917)
  and u13622 (n3752, Aujiu6, F3iow6);  // ../RTL/cortexm0ds_logic.v(11918)
  not u13623 (Y2iow6, n3752);  // ../RTL/cortexm0ds_logic.v(11918)
  or u13624 (F3iow6, Tniiu6, Gaziu6);  // ../RTL/cortexm0ds_logic.v(11919)
  and u13625 (P1iow6, Mb1ju6, M3iow6);  // ../RTL/cortexm0ds_logic.v(11920)
  buf u13626 (Ocfhu6, Ozkbx6[9]);  // ../RTL/cortexm0ds_logic.v(3176)
  not u13627 (M3iow6, Ka1ju6);  // ../RTL/cortexm0ds_logic.v(11921)
  and u13628 (Mb1ju6, T3iow6, A4iow6);  // ../RTL/cortexm0ds_logic.v(11922)
  or u13629 (A4iow6, Bkjiu6, Uvziu6);  // ../RTL/cortexm0ds_logic.v(11923)
  buf u1363 (Iahpw6[12], Oh8ax6);  // ../RTL/cortexm0ds_logic.v(1883)
  and u13630 (n3753, R9aiu6, D7fpw6[3]);  // ../RTL/cortexm0ds_logic.v(11924)
  not u13631 (Bkjiu6, n3753);  // ../RTL/cortexm0ds_logic.v(11924)
  or u13632 (n3754, H4iow6, Hs8ow6);  // ../RTL/cortexm0ds_logic.v(11925)
  not u13633 (T3iow6, n3754);  // ../RTL/cortexm0ds_logic.v(11925)
  and u13634 (Hs8ow6, O4iow6, Aujiu6);  // ../RTL/cortexm0ds_logic.v(11926)
  or u13635 (n3755, X1ziu6, Jcaiu6);  // ../RTL/cortexm0ds_logic.v(11927)
  not u13636 (O4iow6, n3755);  // ../RTL/cortexm0ds_logic.v(11927)
  and u13637 (H4iow6, Srbow6, V4iow6);  // ../RTL/cortexm0ds_logic.v(11928)
  or u13638 (V4iow6, D7fpw6[11], Q6aow6);  // ../RTL/cortexm0ds_logic.v(11929)
  and u13639 (Srbow6, C5iow6, J5iow6);  // ../RTL/cortexm0ds_logic.v(11930)
  buf u1364 (vis_r6_o[2], Mboax6);  // ../RTL/cortexm0ds_logic.v(2523)
  or u13640 (n3756, Jcaiu6, D7fpw6[12]);  // ../RTL/cortexm0ds_logic.v(11931)
  not u13641 (C5iow6, n3756);  // ../RTL/cortexm0ds_logic.v(11931)
  and u13642 (n3757, Q5iow6, X5iow6);  // ../RTL/cortexm0ds_logic.v(11932)
  not u13643 (Zeohu6, n3757);  // ../RTL/cortexm0ds_logic.v(11932)
  and u13644 (n3758, Umhow6, HRDATA[22]);  // ../RTL/cortexm0ds_logic.v(11933)
  not u13645 (X5iow6, n3758);  // ../RTL/cortexm0ds_logic.v(11933)
  and u13646 (n3759, Hrfpw6[6], Qqhiu6);  // ../RTL/cortexm0ds_logic.v(11934)
  not u13647 (Q5iow6, n3759);  // ../RTL/cortexm0ds_logic.v(11934)
  and u13648 (n3760, E6iow6, L6iow6);  // ../RTL/cortexm0ds_logic.v(11935)
  not u13649 (Seohu6, n3760);  // ../RTL/cortexm0ds_logic.v(11935)
  buf u1365 (Iahpw6[13], Xf8ax6);  // ../RTL/cortexm0ds_logic.v(1883)
  and u13650 (n3761, Umhow6, HRDATA[21]);  // ../RTL/cortexm0ds_logic.v(11936)
  not u13651 (L6iow6, n3761);  // ../RTL/cortexm0ds_logic.v(11936)
  and u13652 (n3762, Hrfpw6[5], Qqhiu6);  // ../RTL/cortexm0ds_logic.v(11937)
  not u13653 (E6iow6, n3762);  // ../RTL/cortexm0ds_logic.v(11937)
  or u13654 (Leohu6, S6iow6, Z6iow6);  // ../RTL/cortexm0ds_logic.v(11938)
  or u13655 (n3763, G7iow6, Dk7ow6);  // ../RTL/cortexm0ds_logic.v(11939)
  not u13656 (Z6iow6, n3763);  // ../RTL/cortexm0ds_logic.v(11939)
  and u13657 (Dk7ow6, N7iow6, S3kiu6);  // ../RTL/cortexm0ds_logic.v(11940)
  and u13658 (S3kiu6, U7iow6, B8iow6);  // ../RTL/cortexm0ds_logic.v(11941)
  and u13659 (n3764, Toaiu6, It2ju6);  // ../RTL/cortexm0ds_logic.v(11942)
  buf u1366 (vis_r6_o[3], Jnoax6);  // ../RTL/cortexm0ds_logic.v(2523)
  not u13660 (B8iow6, n3764);  // ../RTL/cortexm0ds_logic.v(11942)
  buf u13661 (Cefhu6, Ozkbx6[8]);  // ../RTL/cortexm0ds_logic.v(3176)
  and u13662 (N7iow6, I8iow6, Et0ju6);  // ../RTL/cortexm0ds_logic.v(11944)
  and u13663 (n3765, L45iu6, Llaow6);  // ../RTL/cortexm0ds_logic.v(11945)
  not u13664 (I8iow6, n3765);  // ../RTL/cortexm0ds_logic.v(11945)
  AL_MUX u13665 (
    .i0(P8iow6),
    .i1(S8fpw6[6]),
    .sel(Rk7ow6),
    .o(S6iow6));  // ../RTL/cortexm0ds_logic.v(11946)
  and u13666 (n3766, HREADY, W8iow6);  // ../RTL/cortexm0ds_logic.v(11947)
  not u13667 (Rk7ow6, n3766);  // ../RTL/cortexm0ds_logic.v(11947)
  and u13668 (n3767, D9iow6, K9iow6);  // ../RTL/cortexm0ds_logic.v(11948)
  not u13669 (W8iow6, n3767);  // ../RTL/cortexm0ds_logic.v(11948)
  buf u1367 (Iahpw6[14], E97ax6);  // ../RTL/cortexm0ds_logic.v(1883)
  and u13670 (K9iow6, R9iow6, Y9iow6);  // ../RTL/cortexm0ds_logic.v(11949)
  and u13671 (Y9iow6, Faiow6, Maiow6);  // ../RTL/cortexm0ds_logic.v(11950)
  and u13672 (n3768, Taiow6, N2ghu6);  // ../RTL/cortexm0ds_logic.v(11951)
  not u13673 (Maiow6, n3768);  // ../RTL/cortexm0ds_logic.v(11951)
  or u13674 (n3769, D9oiu6, Kq0iu6);  // ../RTL/cortexm0ds_logic.v(11952)
  not u13675 (Taiow6, n3769);  // ../RTL/cortexm0ds_logic.v(11952)
  not u13676 (D9oiu6, Whfiu6);  // ../RTL/cortexm0ds_logic.v(11953)
  and u13677 (n3770, Abiow6, Ae0iu6);  // ../RTL/cortexm0ds_logic.v(11954)
  not u13678 (Faiow6, n3770);  // ../RTL/cortexm0ds_logic.v(11954)
  and u13679 (Abiow6, Pthiu6, Mr0iu6);  // ../RTL/cortexm0ds_logic.v(11955)
  buf u1368 (vis_r6_o[4], Ldoax6);  // ../RTL/cortexm0ds_logic.v(2523)
  and u13680 (R9iow6, Hbiow6, Obiow6);  // ../RTL/cortexm0ds_logic.v(11956)
  and u13681 (n3771, Vbiow6, Xzmiu6);  // ../RTL/cortexm0ds_logic.v(11957)
  not u13682 (Obiow6, n3771);  // ../RTL/cortexm0ds_logic.v(11957)
  and u13683 (n3772, Hviiu6, Gaziu6);  // ../RTL/cortexm0ds_logic.v(11958)
  not u13684 (Hbiow6, n3772);  // ../RTL/cortexm0ds_logic.v(11958)
  and u13685 (D9iow6, Cciow6, T1jiu6);  // ../RTL/cortexm0ds_logic.v(11959)
  and u13686 (T1jiu6, Jciow6, Qciow6);  // ../RTL/cortexm0ds_logic.v(11960)
  and u13687 (n3773, Us2ju6, Yljiu6);  // ../RTL/cortexm0ds_logic.v(11961)
  not u13688 (Qciow6, n3773);  // ../RTL/cortexm0ds_logic.v(11961)
  and u13689 (Jciow6, Xciow6, Ediow6);  // ../RTL/cortexm0ds_logic.v(11962)
  buf u1369 (Iahpw6[15], Hlwpw6);  // ../RTL/cortexm0ds_logic.v(1883)
  and u13690 (n3774, Ldiow6, S6aiu6);  // ../RTL/cortexm0ds_logic.v(11963)
  not u13691 (Ediow6, n3774);  // ../RTL/cortexm0ds_logic.v(11963)
  buf u13692 (Qffhu6, Ozkbx6[7]);  // ../RTL/cortexm0ds_logic.v(3176)
  not u13693 (Ldiow6, Eehow6);  // ../RTL/cortexm0ds_logic.v(11964)
  and u13694 (n3775, Zzniu6, Qu7ow6);  // ../RTL/cortexm0ds_logic.v(11965)
  not u13695 (Xciow6, n3775);  // ../RTL/cortexm0ds_logic.v(11965)
  or u13696 (n3776, R2aiu6, Mjfiu6);  // ../RTL/cortexm0ds_logic.v(11966)
  not u13697 (Zzniu6, n3776);  // ../RTL/cortexm0ds_logic.v(11966)
  and u13698 (Cciow6, Epjiu6, Sdiow6);  // ../RTL/cortexm0ds_logic.v(11967)
  or u13699 (Sdiow6, Wmaiu6, Nloiu6);  // ../RTL/cortexm0ds_logic.v(11968)
  buf u137 (E1hpw6[7], Rnaax6);  // ../RTL/cortexm0ds_logic.v(2367)
  buf u1370 (vis_r6_o[5], Ipoax6);  // ../RTL/cortexm0ds_logic.v(2523)
  and u13700 (Epjiu6, Zdiow6, Geiow6);  // ../RTL/cortexm0ds_logic.v(11969)
  and u13701 (Geiow6, Neiow6, Ueiow6);  // ../RTL/cortexm0ds_logic.v(11970)
  and u13702 (Ueiow6, Bfiow6, Ifiow6);  // ../RTL/cortexm0ds_logic.v(11971)
  and u13703 (n3777, Lzhow6, Raaow6);  // ../RTL/cortexm0ds_logic.v(11972)
  not u13704 (Ifiow6, n3777);  // ../RTL/cortexm0ds_logic.v(11972)
  and u13705 (Raaow6, Uyiiu6, Uriiu6);  // ../RTL/cortexm0ds_logic.v(11973)
  and u13706 (Lzhow6, Nbkiu6, X1ziu6);  // ../RTL/cortexm0ds_logic.v(11974)
  and u13707 (Bfiow6, E2ziu6, Oe8ow6);  // ../RTL/cortexm0ds_logic.v(11975)
  and u13708 (n3778, Pfiow6, Jjhiu6);  // ../RTL/cortexm0ds_logic.v(11976)
  not u13709 (E2ziu6, n3778);  // ../RTL/cortexm0ds_logic.v(11976)
  buf u1371 (Iahpw6[16], Ufbbx6);  // ../RTL/cortexm0ds_logic.v(1883)
  and u13710 (Neiow6, Wfiow6, Dgiow6);  // ../RTL/cortexm0ds_logic.v(11977)
  and u13711 (n3779, Vviiu6, Kgiow6);  // ../RTL/cortexm0ds_logic.v(11978)
  not u13712 (Dgiow6, n3779);  // ../RTL/cortexm0ds_logic.v(11978)
  and u13713 (n3780, X1ziu6, Rgiow6);  // ../RTL/cortexm0ds_logic.v(11979)
  not u13714 (Kgiow6, n3780);  // ../RTL/cortexm0ds_logic.v(11979)
  or u13715 (Rgiow6, D7fpw6[8], D7fpw6[9]);  // ../RTL/cortexm0ds_logic.v(11980)
  and u13716 (Vviiu6, Uyiiu6, J9kiu6);  // ../RTL/cortexm0ds_logic.v(11981)
  and u13717 (n3781, Hviiu6, Db0ju6);  // ../RTL/cortexm0ds_logic.v(11982)
  not u13718 (Wfiow6, n3781);  // ../RTL/cortexm0ds_logic.v(11982)
  and u13719 (Db0ju6, D7fpw6[10], Tniiu6);  // ../RTL/cortexm0ds_logic.v(11983)
  buf u1372 (vis_r6_o[6], Hroax6);  // ../RTL/cortexm0ds_logic.v(2523)
  and u13720 (Hviiu6, Ygiow6, J9kiu6);  // ../RTL/cortexm0ds_logic.v(11984)
  or u13721 (n3782, Lraiu6, D7fpw6[14]);  // ../RTL/cortexm0ds_logic.v(11985)
  not u13722 (Ygiow6, n3782);  // ../RTL/cortexm0ds_logic.v(11985)
  and u13723 (Zdiow6, Fhiow6, Mhiow6);  // ../RTL/cortexm0ds_logic.v(11986)
  and u13724 (Mhiow6, Thiow6, Aiiow6);  // ../RTL/cortexm0ds_logic.v(11987)
  and u13725 (n3783, Y31ju6, Hiiow6);  // ../RTL/cortexm0ds_logic.v(11988)
  not u13726 (Aiiow6, n3783);  // ../RTL/cortexm0ds_logic.v(11988)
  and u13727 (n3784, Oiiow6, Viiow6);  // ../RTL/cortexm0ds_logic.v(11989)
  not u13728 (Hiiow6, n3784);  // ../RTL/cortexm0ds_logic.v(11989)
  or u13729 (Viiow6, N38ow6, D7fpw6[15]);  // ../RTL/cortexm0ds_logic.v(11990)
  buf u1373 (Iahpw6[17], Puwpw6);  // ../RTL/cortexm0ds_logic.v(1883)
  or u13730 (n3785, Cjiow6, J1ziu6);  // ../RTL/cortexm0ds_logic.v(11991)
  not u13731 (Oiiow6, n3785);  // ../RTL/cortexm0ds_logic.v(11991)
  and u13732 (Cjiow6, Jjiow6, P0piu6);  // ../RTL/cortexm0ds_logic.v(11992)
  or u13733 (n3786, Qjiow6, O95iu6);  // ../RTL/cortexm0ds_logic.v(11993)
  not u13734 (Jjiow6, n3786);  // ../RTL/cortexm0ds_logic.v(11993)
  or u13735 (Thiow6, O4aiu6, D7fpw6[3]);  // ../RTL/cortexm0ds_logic.v(11994)
  and u13736 (Fhiow6, D0jiu6, Veziu6);  // ../RTL/cortexm0ds_logic.v(11995)
  and u13737 (Veziu6, B1aiu6, Xjiow6);  // ../RTL/cortexm0ds_logic.v(11996)
  and u13738 (n3787, Y0jiu6, Tfjiu6);  // ../RTL/cortexm0ds_logic.v(11997)
  not u13739 (Xjiow6, n3787);  // ../RTL/cortexm0ds_logic.v(11997)
  buf u1374 (vis_r6_o[7], Gtoax6);  // ../RTL/cortexm0ds_logic.v(2523)
  not u13740 (B1aiu6, Ezhow6);  // ../RTL/cortexm0ds_logic.v(11998)
  and u13741 (Ezhow6, O4oiu6, Taaiu6);  // ../RTL/cortexm0ds_logic.v(11999)
  and u13742 (D0jiu6, Ekiow6, Lkiow6);  // ../RTL/cortexm0ds_logic.v(12000)
  and u13743 (Lkiow6, Skiow6, Zkiow6);  // ../RTL/cortexm0ds_logic.v(12001)
  and u13744 (n3788, Gliow6, Nliow6);  // ../RTL/cortexm0ds_logic.v(12002)
  not u13745 (Zkiow6, n3788);  // ../RTL/cortexm0ds_logic.v(12002)
  or u13746 (n3789, Qxoiu6, D7fpw6[13]);  // ../RTL/cortexm0ds_logic.v(12003)
  not u13747 (Nliow6, n3789);  // ../RTL/cortexm0ds_logic.v(12003)
  and u13748 (Gliow6, J9kiu6, Q5aiu6);  // ../RTL/cortexm0ds_logic.v(12004)
  and u13749 (n3790, De6ow6, F9aju6);  // ../RTL/cortexm0ds_logic.v(12005)
  buf u1375 (Iahpw6[18], Ldvpw6);  // ../RTL/cortexm0ds_logic.v(1883)
  not u13750 (Skiow6, n3790);  // ../RTL/cortexm0ds_logic.v(12005)
  and u13751 (Ekiow6, Uliow6, Bmiow6);  // ../RTL/cortexm0ds_logic.v(12006)
  and u13752 (n3791, Evyiu6, W0piu6);  // ../RTL/cortexm0ds_logic.v(12007)
  not u13753 (Bmiow6, n3791);  // ../RTL/cortexm0ds_logic.v(12007)
  or u13754 (n3792, Ftjiu6, Lraiu6);  // ../RTL/cortexm0ds_logic.v(12008)
  not u13755 (W0piu6, n3792);  // ../RTL/cortexm0ds_logic.v(12008)
  and u13756 (Evyiu6, Mtjiu6, X1ziu6);  // ../RTL/cortexm0ds_logic.v(12009)
  or u13757 (Uliow6, O4aiu6, Cyfpw6[0]);  // ../RTL/cortexm0ds_logic.v(12010)
  and u13758 (n3793, Nu9ow6, K9aiu6);  // ../RTL/cortexm0ds_logic.v(12011)
  not u13759 (O4aiu6, n3793);  // ../RTL/cortexm0ds_logic.v(12011)
  buf u1376 (vis_r6_o[8], Dtpax6);  // ../RTL/cortexm0ds_logic.v(2523)
  and u13760 (Nu9ow6, Imiow6, Pmiow6);  // ../RTL/cortexm0ds_logic.v(12012)
  or u13761 (n3794, D7fpw6[14], Cyfpw6[3]);  // ../RTL/cortexm0ds_logic.v(12013)
  not u13762 (Pmiow6, n3794);  // ../RTL/cortexm0ds_logic.v(12013)
  and u13763 (Imiow6, Ya1ju6, Hzziu6);  // ../RTL/cortexm0ds_logic.v(12014)
  and u13764 (n3795, Wmiow6, Dniow6);  // ../RTL/cortexm0ds_logic.v(12015)
  not u13765 (P8iow6, n3795);  // ../RTL/cortexm0ds_logic.v(12015)
  or u13766 (Dniow6, Ad8iu6, Hm7ow6);  // ../RTL/cortexm0ds_logic.v(12016)
  or u13767 (n3796, Zlhow6, Th2ju6);  // ../RTL/cortexm0ds_logic.v(12017)
  not u13768 (Hm7ow6, n3796);  // ../RTL/cortexm0ds_logic.v(12017)
  and u13769 (n3797, Kniow6, Rniow6);  // ../RTL/cortexm0ds_logic.v(12018)
  buf u1377 (Iahpw6[19], Jfdbx6);  // ../RTL/cortexm0ds_logic.v(1883)
  not u13770 (Zlhow6, n3797);  // ../RTL/cortexm0ds_logic.v(12018)
  and u13771 (Rniow6, Yniow6, Foiow6);  // ../RTL/cortexm0ds_logic.v(12019)
  buf u13772 (Dhfhu6, Ozkbx6[6]);  // ../RTL/cortexm0ds_logic.v(3176)
  and u13773 (Yniow6, Moiow6, S4jiu6);  // ../RTL/cortexm0ds_logic.v(12021)
  and u13774 (n3798, Toiow6, Ia8iu6);  // ../RTL/cortexm0ds_logic.v(12022)
  not u13775 (S4jiu6, n3798);  // ../RTL/cortexm0ds_logic.v(12022)
  or u13776 (n3799, C27ow6, Ftjiu6);  // ../RTL/cortexm0ds_logic.v(12023)
  not u13777 (Toiow6, n3799);  // ../RTL/cortexm0ds_logic.v(12023)
  not u13778 (C27ow6, Wliiu6);  // ../RTL/cortexm0ds_logic.v(12024)
  and u13779 (n3800, J1ziu6, Ia8iu6);  // ../RTL/cortexm0ds_logic.v(12025)
  buf u1378 (vis_r6_o[9], Erpax6);  // ../RTL/cortexm0ds_logic.v(2523)
  not u13780 (Moiow6, n3800);  // ../RTL/cortexm0ds_logic.v(12025)
  and u13781 (J1ziu6, Wliiu6, D7fpw6[11]);  // ../RTL/cortexm0ds_logic.v(12026)
  and u13782 (Wliiu6, Mtjiu6, Gaziu6);  // ../RTL/cortexm0ds_logic.v(12027)
  not u13783 (Gaziu6, D7fpw6[13]);  // ../RTL/cortexm0ds_logic.v(12028)
  and u13784 (Kniow6, Ubkiu6, Apiow6);  // ../RTL/cortexm0ds_logic.v(12029)
  or u13785 (Apiow6, E4jiu6, Ae0iu6);  // ../RTL/cortexm0ds_logic.v(12030)
  and u13786 (Ubkiu6, Ymiiu6, Hpiow6);  // ../RTL/cortexm0ds_logic.v(12031)
  or u13787 (Hpiow6, Hujiu6, Aujiu6);  // ../RTL/cortexm0ds_logic.v(12032)
  not u13788 (Hujiu6, Th2ju6);  // ../RTL/cortexm0ds_logic.v(12033)
  and u13789 (Th2ju6, Xiiiu6, Kxziu6);  // ../RTL/cortexm0ds_logic.v(12034)
  buf u1379 (Iahpw6[20], Sddbx6);  // ../RTL/cortexm0ds_logic.v(1883)
  or u13790 (Ymiiu6, Xl0ju6, Qpaju6);  // ../RTL/cortexm0ds_logic.v(12035)
  not u13791 (Xl0ju6, R7jiu6);  // ../RTL/cortexm0ds_logic.v(12037)
  or u13792 (Wmiow6, Dzjiu6, Cn7ow6);  // ../RTL/cortexm0ds_logic.v(12038)
  and u13793 (Cn7ow6, Opiow6, Oaiiu6);  // ../RTL/cortexm0ds_logic.v(12039)
  and u13794 (Ry7ow6, Vpiow6, J9kiu6);  // ../RTL/cortexm0ds_logic.v(12040)
  not u13795 (Oaiiu6, Ry7ow6);  // ../RTL/cortexm0ds_logic.v(12040)
  or u13796 (n3801, Co6ow6, Ae0iu6);  // ../RTL/cortexm0ds_logic.v(12041)
  not u13797 (Vpiow6, n3801);  // ../RTL/cortexm0ds_logic.v(12041)
  and u13798 (n3802, Ia8iu6, Ozziu6);  // ../RTL/cortexm0ds_logic.v(12042)
  not u13799 (Opiow6, n3802);  // ../RTL/cortexm0ds_logic.v(12042)
  buf u138 (vis_r1_o[9], Ir1qw6);  // ../RTL/cortexm0ds_logic.v(1876)
  buf u1380 (vis_r6_o[10], Eppax6);  // ../RTL/cortexm0ds_logic.v(2523)
  and u13800 (n3803, Cqiow6, Jqiow6);  // ../RTL/cortexm0ds_logic.v(12043)
  not u13801 (Eeohu6, n3803);  // ../RTL/cortexm0ds_logic.v(12043)
  and u13802 (n3804, Umhow6, HRDATA[20]);  // ../RTL/cortexm0ds_logic.v(12044)
  not u13803 (Jqiow6, n3804);  // ../RTL/cortexm0ds_logic.v(12044)
  and u13804 (n3805, Hrfpw6[4], Qqhiu6);  // ../RTL/cortexm0ds_logic.v(12045)
  not u13805 (Cqiow6, n3805);  // ../RTL/cortexm0ds_logic.v(12045)
  AL_MUX u13806 (
    .i0(Qqiow6),
    .i1(Sufpw6[0]),
    .sel(Eh6iu6),
    .o(Xdohu6));  // ../RTL/cortexm0ds_logic.v(12046)
  and u13807 (Qqiow6, Xqiow6, Ophiu6);  // ../RTL/cortexm0ds_logic.v(12047)
  or u13808 (Xqiow6, N6piu6, Sufpw6[1]);  // ../RTL/cortexm0ds_logic.v(12048)
  AL_MUX u13809 (
    .i0(Fnpiu6),
    .i1(L3ehu6),
    .sel(Eh6iu6),
    .o(Qdohu6));  // ../RTL/cortexm0ds_logic.v(12049)
  buf u1381 (Cjhpw6[1], Nrqpw6);  // ../RTL/cortexm0ds_logic.v(2365)
  not u13810 (Fnpiu6, Ejpiu6);  // ../RTL/cortexm0ds_logic.v(12050)
  and u13811 (n3806, Eriow6, Lriow6);  // ../RTL/cortexm0ds_logic.v(12051)
  not u13812 (Jdohu6, n3806);  // ../RTL/cortexm0ds_logic.v(12051)
  and u13813 (Lriow6, Sriow6, Zriow6);  // ../RTL/cortexm0ds_logic.v(12052)
  and u13814 (n3807, Egziu6, Eafpw6[11]);  // ../RTL/cortexm0ds_logic.v(12053)
  not u13815 (Zriow6, n3807);  // ../RTL/cortexm0ds_logic.v(12053)
  and u13816 (Sriow6, Gsiow6, Sgziu6);  // ../RTL/cortexm0ds_logic.v(12054)
  and u13817 (n3808, Zgziu6, Uumiu6);  // ../RTL/cortexm0ds_logic.v(12055)
  not u13818 (Gsiow6, n3808);  // ../RTL/cortexm0ds_logic.v(12055)
  and u13819 (n3809, Nsiow6, Usiow6);  // ../RTL/cortexm0ds_logic.v(12056)
  buf u1382 (vis_r6_o[29], F1pax6);  // ../RTL/cortexm0ds_logic.v(2523)
  not u13820 (Uumiu6, n3809);  // ../RTL/cortexm0ds_logic.v(12056)
  and u13821 (Usiow6, Btiow6, Itiow6);  // ../RTL/cortexm0ds_logic.v(12057)
  or u13822 (Itiow6, Tgcow6, Pkdow6);  // ../RTL/cortexm0ds_logic.v(12058)
  and u13823 (Tgcow6, Ptiow6, Wtiow6);  // ../RTL/cortexm0ds_logic.v(12059)
  and u13824 (Wtiow6, Duiow6, Kuiow6);  // ../RTL/cortexm0ds_logic.v(12060)
  and u13825 (n3810, Dyeow6, Re4ju6);  // ../RTL/cortexm0ds_logic.v(12061)
  not u13826 (Kuiow6, n3810);  // ../RTL/cortexm0ds_logic.v(12061)
  or u13827 (Duiow6, Iydow6, Uosiu6);  // ../RTL/cortexm0ds_logic.v(12062)
  and u13828 (Uosiu6, Ruiow6, Yuiow6);  // ../RTL/cortexm0ds_logic.v(12063)
  and u13829 (Yuiow6, Fviow6, Mviow6);  // ../RTL/cortexm0ds_logic.v(12064)
  buf u1383 (Iahpw6[21], Bcdbx6);  // ../RTL/cortexm0ds_logic.v(1883)
  and u13830 (n3811, Tzfpw6[11], Yvgiu6);  // ../RTL/cortexm0ds_logic.v(12065)
  not u13831 (Mviow6, n3811);  // ../RTL/cortexm0ds_logic.v(12065)
  and u13832 (Fviow6, Tviow6, Awiow6);  // ../RTL/cortexm0ds_logic.v(12066)
  and u13833 (n3812, F0eow6, Vbgpw6[11]);  // ../RTL/cortexm0ds_logic.v(12067)
  not u13834 (Awiow6, n3812);  // ../RTL/cortexm0ds_logic.v(12067)
  and u13835 (n3813, Odgpw6[11], M0eow6);  // ../RTL/cortexm0ds_logic.v(12068)
  not u13836 (Tviow6, n3813);  // ../RTL/cortexm0ds_logic.v(12068)
  and u13837 (Ruiow6, Hwiow6, Owiow6);  // ../RTL/cortexm0ds_logic.v(12069)
  and u13838 (n3814, Bagpw6[11], M6eiu6);  // ../RTL/cortexm0ds_logic.v(12070)
  not u13839 (Owiow6, n3814);  // ../RTL/cortexm0ds_logic.v(12070)
  buf u1384 (vis_r6_o[11], Cm7bx6);  // ../RTL/cortexm0ds_logic.v(2523)
  and u13840 (n3815, STCALIB[11], H1eow6);  // ../RTL/cortexm0ds_logic.v(12071)
  not u13841 (Hwiow6, n3815);  // ../RTL/cortexm0ds_logic.v(12071)
  and u13842 (Ptiow6, Vwiow6, Cxiow6);  // ../RTL/cortexm0ds_logic.v(12072)
  and u13843 (n3816, Qtfow6, Ag4ju6);  // ../RTL/cortexm0ds_logic.v(12073)
  not u13844 (Cxiow6, n3816);  // ../RTL/cortexm0ds_logic.v(12073)
  and u13845 (n3817, HRDATA[11], Q2eow6);  // ../RTL/cortexm0ds_logic.v(12074)
  not u13846 (Vwiow6, n3817);  // ../RTL/cortexm0ds_logic.v(12074)
  and u13847 (Btiow6, Jxiow6, Dldow6);  // ../RTL/cortexm0ds_logic.v(12075)
  or u13848 (Jxiow6, Kfcow6, Uqdow6);  // ../RTL/cortexm0ds_logic.v(12076)
  and u13849 (Kfcow6, Qxiow6, Xxiow6);  // ../RTL/cortexm0ds_logic.v(12077)
  buf u1385 (Iahpw6[22], Kadbx6);  // ../RTL/cortexm0ds_logic.v(1883)
  and u13850 (Xxiow6, Eyiow6, Lyiow6);  // ../RTL/cortexm0ds_logic.v(12078)
  and u13851 (n3818, Dyeow6, Jw3ju6);  // ../RTL/cortexm0ds_logic.v(12079)
  not u13852 (Lyiow6, n3818);  // ../RTL/cortexm0ds_logic.v(12079)
  or u13853 (Eyiow6, Iydow6, Tmqiu6);  // ../RTL/cortexm0ds_logic.v(12080)
  and u13854 (Tmqiu6, Syiow6, Zyiow6);  // ../RTL/cortexm0ds_logic.v(12081)
  and u13855 (Zyiow6, Gziow6, Nziow6);  // ../RTL/cortexm0ds_logic.v(12082)
  and u13856 (Nziow6, Uziow6, B0jow6);  // ../RTL/cortexm0ds_logic.v(12083)
  and u13857 (n3819, STCALIB[3], H1eow6);  // ../RTL/cortexm0ds_logic.v(12084)
  not u13858 (Uziow6, n3819);  // ../RTL/cortexm0ds_logic.v(12084)
  and u13859 (Gziow6, I0jow6, P0jow6);  // ../RTL/cortexm0ds_logic.v(12085)
  buf u1386 (vis_r6_o[12], Enpax6);  // ../RTL/cortexm0ds_logic.v(2523)
  and u13860 (n3820, Odgpw6[3], M0eow6);  // ../RTL/cortexm0ds_logic.v(12086)
  not u13861 (P0jow6, n3820);  // ../RTL/cortexm0ds_logic.v(12086)
  and u13862 (n3821, Tzfpw6[3], Yvgiu6);  // ../RTL/cortexm0ds_logic.v(12087)
  not u13863 (I0jow6, n3821);  // ../RTL/cortexm0ds_logic.v(12087)
  and u13864 (Syiow6, W0jow6, D1jow6);  // ../RTL/cortexm0ds_logic.v(12088)
  and u13865 (D1jow6, K1jow6, R1jow6);  // ../RTL/cortexm0ds_logic.v(12089)
  and u13866 (n3822, Bagpw6[3], M6eiu6);  // ../RTL/cortexm0ds_logic.v(12090)
  not u13867 (R1jow6, n3822);  // ../RTL/cortexm0ds_logic.v(12090)
  and u13868 (n3823, F0eow6, Vbgpw6[3]);  // ../RTL/cortexm0ds_logic.v(12091)
  not u13869 (K1jow6, n3823);  // ../RTL/cortexm0ds_logic.v(12091)
  buf u1387 (Iahpw6[23], Stkpw6);  // ../RTL/cortexm0ds_logic.v(1883)
  and u13870 (W0jow6, Y1jow6, F2jow6);  // ../RTL/cortexm0ds_logic.v(12092)
  or u13871 (F2jow6, Qkgiu6, Ngfiu6);  // ../RTL/cortexm0ds_logic.v(12093)
  and u13872 (n3824, ECOREVNUM[3], I5eow6);  // ../RTL/cortexm0ds_logic.v(12094)
  not u13873 (Y1jow6, n3824);  // ../RTL/cortexm0ds_logic.v(12094)
  and u13874 (Qxiow6, M2jow6, T2jow6);  // ../RTL/cortexm0ds_logic.v(12095)
  and u13875 (n3825, Qtfow6, Lx3ju6);  // ../RTL/cortexm0ds_logic.v(12096)
  not u13876 (T2jow6, n3825);  // ../RTL/cortexm0ds_logic.v(12096)
  and u13877 (n3826, HRDATA[3], Q2eow6);  // ../RTL/cortexm0ds_logic.v(12097)
  not u13878 (M2jow6, n3826);  // ../RTL/cortexm0ds_logic.v(12097)
  and u13879 (Nsiow6, A3jow6, H3jow6);  // ../RTL/cortexm0ds_logic.v(12098)
  buf u1388 (vis_r6_o[13], Elpax6);  // ../RTL/cortexm0ds_logic.v(2523)
  or u13880 (H3jow6, Ahcow6, Kldow6);  // ../RTL/cortexm0ds_logic.v(12099)
  and u13881 (Ahcow6, O3jow6, V3jow6);  // ../RTL/cortexm0ds_logic.v(12100)
  and u13882 (V3jow6, C4jow6, J4jow6);  // ../RTL/cortexm0ds_logic.v(12101)
  or u13883 (J4jow6, Rcfow6, C34ju6);  // ../RTL/cortexm0ds_logic.v(12102)
  or u13884 (C4jow6, Iydow6, U8uiu6);  // ../RTL/cortexm0ds_logic.v(12103)
  and u13885 (U8uiu6, Q4jow6, X4jow6);  // ../RTL/cortexm0ds_logic.v(12104)
  and u13886 (X4jow6, E5jow6, L5jow6);  // ../RTL/cortexm0ds_logic.v(12105)
  and u13887 (n3827, STCALIB[19], H1eow6);  // ../RTL/cortexm0ds_logic.v(12106)
  not u13888 (L5jow6, n3827);  // ../RTL/cortexm0ds_logic.v(12106)
  and u13889 (E5jow6, S5jow6, Z5jow6);  // ../RTL/cortexm0ds_logic.v(12107)
  buf u1389 (Iahpw6[24], Kn2qw6);  // ../RTL/cortexm0ds_logic.v(1883)
  and u13890 (n3828, Tzfpw6[19], Yvgiu6);  // ../RTL/cortexm0ds_logic.v(12108)
  not u13891 (Z5jow6, n3828);  // ../RTL/cortexm0ds_logic.v(12108)
  and u13892 (n3829, Bagpw6[19], M6eiu6);  // ../RTL/cortexm0ds_logic.v(12109)
  not u13893 (S5jow6, n3829);  // ../RTL/cortexm0ds_logic.v(12109)
  or u13894 (n3830, G6jow6, I5eow6);  // ../RTL/cortexm0ds_logic.v(12110)
  not u13895 (Q4jow6, n3830);  // ../RTL/cortexm0ds_logic.v(12110)
  and u13896 (n3831, N6jow6, U6jow6);  // ../RTL/cortexm0ds_logic.v(12111)
  not u13897 (G6jow6, n3831);  // ../RTL/cortexm0ds_logic.v(12111)
  and u13898 (n3832, Odgpw6[19], M0eow6);  // ../RTL/cortexm0ds_logic.v(12112)
  not u13899 (U6jow6, n3832);  // ../RTL/cortexm0ds_logic.v(12112)
  buf u139 (vis_r12_o[12], Eutax6);  // ../RTL/cortexm0ds_logic.v(2599)
  buf u1390 (vis_r6_o[14], Ejpax6);  // ../RTL/cortexm0ds_logic.v(2523)
  and u13900 (n3833, F0eow6, Vbgpw6[19]);  // ../RTL/cortexm0ds_logic.v(12113)
  not u13901 (N6jow6, n3833);  // ../RTL/cortexm0ds_logic.v(12113)
  and u13902 (O3jow6, B7jow6, I7jow6);  // ../RTL/cortexm0ds_logic.v(12114)
  and u13903 (n3834, Qtfow6, L44ju6);  // ../RTL/cortexm0ds_logic.v(12115)
  not u13904 (I7jow6, n3834);  // ../RTL/cortexm0ds_logic.v(12115)
  and u13905 (n3835, HRDATA[19], Q2eow6);  // ../RTL/cortexm0ds_logic.v(12116)
  not u13906 (B7jow6, n3835);  // ../RTL/cortexm0ds_logic.v(12116)
  or u13907 (A3jow6, Yfcow6, Spdow6);  // ../RTL/cortexm0ds_logic.v(12117)
  and u13908 (Yfcow6, P7jow6, W7jow6);  // ../RTL/cortexm0ds_logic.v(12118)
  or u13909 (W7jow6, Iydow6, Wtviu6);  // ../RTL/cortexm0ds_logic.v(12119)
  buf u1391 (Iahpw6[25], J4cbx6);  // ../RTL/cortexm0ds_logic.v(1883)
  and u13910 (Wtviu6, D8jow6, K8jow6);  // ../RTL/cortexm0ds_logic.v(12120)
  and u13911 (n3836, F0eow6, Vbgpw6[27]);  // ../RTL/cortexm0ds_logic.v(12121)
  not u13912 (K8jow6, n3836);  // ../RTL/cortexm0ds_logic.v(12121)
  and u13913 (D8jow6, R8jow6, Yreow6);  // ../RTL/cortexm0ds_logic.v(12122)
  and u13914 (n3837, Odgpw6[27], M0eow6);  // ../RTL/cortexm0ds_logic.v(12123)
  not u13915 (R8jow6, n3837);  // ../RTL/cortexm0ds_logic.v(12123)
  and u13916 (P7jow6, Y8jow6, F9jow6);  // ../RTL/cortexm0ds_logic.v(12124)
  and u13917 (n3838, C2eow6, M9jow6);  // ../RTL/cortexm0ds_logic.v(12125)
  not u13918 (F9jow6, n3838);  // ../RTL/cortexm0ds_logic.v(12125)
  and u13919 (n3839, O94ju6, T9jow6);  // ../RTL/cortexm0ds_logic.v(12126)
  buf u1392 (vis_r6_o[15], Zb8bx6);  // ../RTL/cortexm0ds_logic.v(2523)
  not u13920 (M9jow6, n3839);  // ../RTL/cortexm0ds_logic.v(12126)
  or u13921 (T9jow6, Aajow6, Bz3ju6);  // ../RTL/cortexm0ds_logic.v(12127)
  and u13922 (n3840, Hajow6, Oajow6);  // ../RTL/cortexm0ds_logic.v(12128)
  not u13923 (O94ju6, n3840);  // ../RTL/cortexm0ds_logic.v(12128)
  or u13924 (Oajow6, Vajow6, J2eow6);  // ../RTL/cortexm0ds_logic.v(12129)
  and u13925 (Hajow6, Cbjow6, Aajow6);  // ../RTL/cortexm0ds_logic.v(12130)
  and u13926 (n3841, Jbjow6, Qbjow6);  // ../RTL/cortexm0ds_logic.v(12131)
  not u13927 (Aajow6, n3841);  // ../RTL/cortexm0ds_logic.v(12131)
  and u13928 (n3842, Xbjow6, Ecjow6);  // ../RTL/cortexm0ds_logic.v(12132)
  not u13929 (Cbjow6, n3842);  // ../RTL/cortexm0ds_logic.v(12132)
  buf u1393 (Iahpw6[26], S2cbx6);  // ../RTL/cortexm0ds_logic.v(1883)
  and u13930 (Xbjow6, J2eow6, Lcjow6);  // ../RTL/cortexm0ds_logic.v(12133)
  and u13931 (n3843, HRDATA[27], Q2eow6);  // ../RTL/cortexm0ds_logic.v(12134)
  not u13932 (Y8jow6, n3843);  // ../RTL/cortexm0ds_logic.v(12134)
  and u13933 (Eriow6, Scjow6, Zcjow6);  // ../RTL/cortexm0ds_logic.v(12135)
  and u13934 (n3844, Zsfpw6[10], Cmziu6);  // ../RTL/cortexm0ds_logic.v(12136)
  not u13935 (Zcjow6, n3844);  // ../RTL/cortexm0ds_logic.v(12136)
  and u13936 (n3845, vis_pc_o[10], Jmziu6);  // ../RTL/cortexm0ds_logic.v(12137)
  not u13937 (Scjow6, n3845);  // ../RTL/cortexm0ds_logic.v(12137)
  and u13938 (n3846, Gdjow6, Ndjow6);  // ../RTL/cortexm0ds_logic.v(12138)
  not u13939 (Cdohu6, n3846);  // ../RTL/cortexm0ds_logic.v(12138)
  buf u1394 (vis_r6_o[16], Ehpax6);  // ../RTL/cortexm0ds_logic.v(2523)
  and u13940 (Ndjow6, Udjow6, Bejow6);  // ../RTL/cortexm0ds_logic.v(12139)
  and u13941 (n3847, Egziu6, Eafpw6[9]);  // ../RTL/cortexm0ds_logic.v(12140)
  not u13942 (Bejow6, n3847);  // ../RTL/cortexm0ds_logic.v(12140)
  and u13943 (Udjow6, Iejow6, Sgziu6);  // ../RTL/cortexm0ds_logic.v(12141)
  and u13944 (n3848, Zgziu6, S0niu6);  // ../RTL/cortexm0ds_logic.v(12142)
  not u13945 (Iejow6, n3848);  // ../RTL/cortexm0ds_logic.v(12142)
  and u13946 (n3849, Pejow6, Wejow6);  // ../RTL/cortexm0ds_logic.v(12143)
  not u13947 (S0niu6, n3849);  // ../RTL/cortexm0ds_logic.v(12143)
  and u13948 (Wejow6, Dfjow6, Kfjow6);  // ../RTL/cortexm0ds_logic.v(12144)
  and u13949 (n3850, Mmdow6, Ew6ow6);  // ../RTL/cortexm0ds_logic.v(12145)
  buf u1395 (Iahpw6[27], Nfqpw6);  // ../RTL/cortexm0ds_logic.v(1883)
  not u13950 (Kfjow6, n3850);  // ../RTL/cortexm0ds_logic.v(12145)
  and u13951 (n3851, Rfjow6, Yfjow6);  // ../RTL/cortexm0ds_logic.v(12146)
  not u13952 (Ew6ow6, n3851);  // ../RTL/cortexm0ds_logic.v(12146)
  and u13953 (Yfjow6, Fgjow6, Mgjow6);  // ../RTL/cortexm0ds_logic.v(12147)
  or u13954 (Mgjow6, Rcfow6, Mu3ju6);  // ../RTL/cortexm0ds_logic.v(12148)
  and u13955 (Mu3ju6, Tgjow6, Ahjow6);  // ../RTL/cortexm0ds_logic.v(12149)
  and u13956 (Ahjow6, Hhjow6, Ohjow6);  // ../RTL/cortexm0ds_logic.v(12150)
  or u13957 (Ohjow6, Rqfow6, I40iu6);  // ../RTL/cortexm0ds_logic.v(12151)
  or u13958 (Hhjow6, Ipfow6, B40iu6);  // ../RTL/cortexm0ds_logic.v(12152)
  and u13959 (Tgjow6, Vhjow6, Cijow6);  // ../RTL/cortexm0ds_logic.v(12153)
  buf u1396 (vis_r6_o[17], Efpax6);  // ../RTL/cortexm0ds_logic.v(2523)
  or u13960 (Cijow6, Ppfow6, W40iu6);  // ../RTL/cortexm0ds_logic.v(12154)
  or u13961 (Vhjow6, Kqfow6, P40iu6);  // ../RTL/cortexm0ds_logic.v(12155)
  or u13962 (Fgjow6, Iydow6, Ovpiu6);  // ../RTL/cortexm0ds_logic.v(12156)
  and u13963 (Ovpiu6, Jijow6, Qijow6);  // ../RTL/cortexm0ds_logic.v(12157)
  and u13964 (Qijow6, Xijow6, Ejjow6);  // ../RTL/cortexm0ds_logic.v(12158)
  and u13965 (Ejjow6, Ljjow6, Sjjow6);  // ../RTL/cortexm0ds_logic.v(12159)
  and u13966 (n3852, Odgpw6[1], M0eow6);  // ../RTL/cortexm0ds_logic.v(12160)
  not u13967 (Sjjow6, n3852);  // ../RTL/cortexm0ds_logic.v(12160)
  and u13968 (Ljjow6, Zjjow6, Gkjow6);  // ../RTL/cortexm0ds_logic.v(12161)
  and u13969 (n3853, Fpgiu6, Qqdhu6);  // ../RTL/cortexm0ds_logic.v(12162)
  buf u1397 (Iahpw6[28], Wt3qw6);  // ../RTL/cortexm0ds_logic.v(1883)
  not u13970 (Gkjow6, n3853);  // ../RTL/cortexm0ds_logic.v(12162)
  and u13971 (n3854, Tzfpw6[1], Yvgiu6);  // ../RTL/cortexm0ds_logic.v(12163)
  not u13972 (Zjjow6, n3854);  // ../RTL/cortexm0ds_logic.v(12163)
  and u13973 (Xijow6, Nkjow6, Ukjow6);  // ../RTL/cortexm0ds_logic.v(12164)
  and u13974 (n3855, ECOREVNUM[1], I5eow6);  // ../RTL/cortexm0ds_logic.v(12165)
  not u13975 (Ukjow6, n3855);  // ../RTL/cortexm0ds_logic.v(12165)
  and u13976 (n3856, Y5eiu6, Dvghu6);  // ../RTL/cortexm0ds_logic.v(12166)
  not u13977 (Nkjow6, n3856);  // ../RTL/cortexm0ds_logic.v(12166)
  and u13978 (Jijow6, Bljow6, Iljow6);  // ../RTL/cortexm0ds_logic.v(12167)
  and u13979 (Iljow6, Pljow6, Wljow6);  // ../RTL/cortexm0ds_logic.v(12168)
  buf u1398 (vis_r6_o[18], Edpax6);  // ../RTL/cortexm0ds_logic.v(2523)
  and u13980 (n3857, F0eow6, Vbgpw6[1]);  // ../RTL/cortexm0ds_logic.v(12169)
  not u13981 (Wljow6, n3857);  // ../RTL/cortexm0ds_logic.v(12169)
  and u13982 (n3858, Bagpw6[1], M6eiu6);  // ../RTL/cortexm0ds_logic.v(12170)
  not u13983 (Pljow6, n3858);  // ../RTL/cortexm0ds_logic.v(12170)
  and u13984 (Bljow6, Dmjow6, Kmjow6);  // ../RTL/cortexm0ds_logic.v(12171)
  and u13985 (n3859, STCALIB[1], H1eow6);  // ../RTL/cortexm0ds_logic.v(12172)
  not u13986 (Kmjow6, n3859);  // ../RTL/cortexm0ds_logic.v(12172)
  or u13987 (Dmjow6, Qkgiu6, Siciu6);  // ../RTL/cortexm0ds_logic.v(12173)
  and u13988 (Rfjow6, Rmjow6, Ymjow6);  // ../RTL/cortexm0ds_logic.v(12174)
  and u13989 (n3860, Qtfow6, Ex3ju6);  // ../RTL/cortexm0ds_logic.v(12175)
  buf u1399 (Iahpw6[29], C72qw6);  // ../RTL/cortexm0ds_logic.v(1883)
  not u13990 (Ymjow6, n3860);  // ../RTL/cortexm0ds_logic.v(12175)
  and u13991 (n3861, Fnjow6, Mnjow6);  // ../RTL/cortexm0ds_logic.v(12176)
  not u13992 (Ex3ju6, n3861);  // ../RTL/cortexm0ds_logic.v(12176)
  and u13993 (Mnjow6, Tnjow6, Aojow6);  // ../RTL/cortexm0ds_logic.v(12177)
  or u13994 (Aojow6, Kqfow6, F60iu6);  // ../RTL/cortexm0ds_logic.v(12178)
  or u13995 (Tnjow6, Ipfow6, D50iu6);  // ../RTL/cortexm0ds_logic.v(12179)
  and u13996 (Fnjow6, Hojow6, Oojow6);  // ../RTL/cortexm0ds_logic.v(12180)
  or u13997 (Oojow6, Rqfow6, K50iu6);  // ../RTL/cortexm0ds_logic.v(12181)
  or u13998 (Hojow6, Ppfow6, E90iu6);  // ../RTL/cortexm0ds_logic.v(12182)
  and u13999 (n3862, HRDATA[1], Q2eow6);  // ../RTL/cortexm0ds_logic.v(12183)
  buf u14 (Pndhu6, Hwhpw6);  // ../RTL/cortexm0ds_logic.v(1770)
  buf u140 (S1ehu6, Hgrpw6);  // ../RTL/cortexm0ds_logic.v(1949)
  buf u1400 (vis_r6_o[19], Ebpax6);  // ../RTL/cortexm0ds_logic.v(2523)
  not u14000 (Rmjow6, n3862);  // ../RTL/cortexm0ds_logic.v(12183)
  and u14001 (Dfjow6, Vojow6, Dldow6);  // ../RTL/cortexm0ds_logic.v(12184)
  or u14002 (Vojow6, Pkdow6, Xv6ow6);  // ../RTL/cortexm0ds_logic.v(12185)
  and u14003 (Xv6ow6, Cpjow6, Jpjow6);  // ../RTL/cortexm0ds_logic.v(12186)
  and u14004 (Jpjow6, Qpjow6, Xpjow6);  // ../RTL/cortexm0ds_logic.v(12187)
  or u14005 (Xpjow6, Rcfow6, Uc4ju6);  // ../RTL/cortexm0ds_logic.v(12188)
  and u14006 (Uc4ju6, Eqjow6, Lqjow6);  // ../RTL/cortexm0ds_logic.v(12189)
  and u14007 (Lqjow6, Sqjow6, Zqjow6);  // ../RTL/cortexm0ds_logic.v(12190)
  or u14008 (Zqjow6, Ipfow6, Ga0iu6);  // ../RTL/cortexm0ds_logic.v(12191)
  or u14009 (Sqjow6, Ppfow6, Bb0iu6);  // ../RTL/cortexm0ds_logic.v(12192)
  buf u1401 (Iahpw6[30], Zwnpw6);  // ../RTL/cortexm0ds_logic.v(1883)
  and u14010 (Eqjow6, Grjow6, Nrjow6);  // ../RTL/cortexm0ds_logic.v(12193)
  or u14011 (Nrjow6, Kqfow6, Ua0iu6);  // ../RTL/cortexm0ds_logic.v(12194)
  or u14012 (Grjow6, Rqfow6, Na0iu6);  // ../RTL/cortexm0ds_logic.v(12195)
  or u14013 (Qpjow6, Iydow6, Ibsiu6);  // ../RTL/cortexm0ds_logic.v(12196)
  and u14014 (Ibsiu6, Urjow6, Bsjow6);  // ../RTL/cortexm0ds_logic.v(12197)
  and u14015 (Bsjow6, Isjow6, Psjow6);  // ../RTL/cortexm0ds_logic.v(12198)
  and u14016 (Psjow6, Wsjow6, B0jow6);  // ../RTL/cortexm0ds_logic.v(12199)
  and u14017 (n3863, Rzciu6, Dtjow6);  // ../RTL/cortexm0ds_logic.v(12200)
  not u14018 (B0jow6, n3863);  // ../RTL/cortexm0ds_logic.v(12200)
  and u14019 (n3864, Bagpw6[9], M6eiu6);  // ../RTL/cortexm0ds_logic.v(12201)
  buf u1402 (vis_r6_o[20], E9pax6);  // ../RTL/cortexm0ds_logic.v(2523)
  not u14020 (Wsjow6, n3864);  // ../RTL/cortexm0ds_logic.v(12201)
  and u14021 (Isjow6, Ktjow6, Rtjow6);  // ../RTL/cortexm0ds_logic.v(12202)
  and u14022 (n3865, Tzfpw6[9], Yvgiu6);  // ../RTL/cortexm0ds_logic.v(12203)
  not u14023 (Rtjow6, n3865);  // ../RTL/cortexm0ds_logic.v(12203)
  and u14024 (n3866, F0eow6, Vbgpw6[9]);  // ../RTL/cortexm0ds_logic.v(12204)
  not u14025 (Ktjow6, n3866);  // ../RTL/cortexm0ds_logic.v(12204)
  and u14026 (Urjow6, Ytjow6, Qgeow6);  // ../RTL/cortexm0ds_logic.v(12205)
  and u14027 (Ytjow6, Fujow6, Mujow6);  // ../RTL/cortexm0ds_logic.v(12206)
  and u14028 (n3867, STCALIB[9], H1eow6);  // ../RTL/cortexm0ds_logic.v(12207)
  not u14029 (Mujow6, n3867);  // ../RTL/cortexm0ds_logic.v(12207)
  buf u1403 (Cjhpw6[2], Nmfax6);  // ../RTL/cortexm0ds_logic.v(2365)
  and u14030 (n3868, M0eow6, Odgpw6[9]);  // ../RTL/cortexm0ds_logic.v(12208)
  not u14031 (Fujow6, n3868);  // ../RTL/cortexm0ds_logic.v(12208)
  and u14032 (Cpjow6, Tujow6, Avjow6);  // ../RTL/cortexm0ds_logic.v(12209)
  and u14033 (n3869, Qtfow6, Hg4ju6);  // ../RTL/cortexm0ds_logic.v(12210)
  not u14034 (Avjow6, n3869);  // ../RTL/cortexm0ds_logic.v(12210)
  and u14035 (n3870, Hvjow6, Ovjow6);  // ../RTL/cortexm0ds_logic.v(12211)
  not u14036 (Hg4ju6, n3870);  // ../RTL/cortexm0ds_logic.v(12211)
  and u14037 (Ovjow6, Vvjow6, Cwjow6);  // ../RTL/cortexm0ds_logic.v(12212)
  or u14038 (Cwjow6, Rqfow6, Pb0iu6);  // ../RTL/cortexm0ds_logic.v(12213)
  or u14039 (Vvjow6, Ppfow6, U30iu6);  // ../RTL/cortexm0ds_logic.v(12214)
  buf u1404 (vis_r6_o[30], Khoax6);  // ../RTL/cortexm0ds_logic.v(2523)
  and u14040 (Hvjow6, Jwjow6, Qwjow6);  // ../RTL/cortexm0ds_logic.v(12215)
  or u14041 (Qwjow6, Kqfow6, Wb0iu6);  // ../RTL/cortexm0ds_logic.v(12216)
  or u14042 (Jwjow6, Ipfow6, Ib0iu6);  // ../RTL/cortexm0ds_logic.v(12217)
  and u14043 (n3871, HRDATA[9], Q2eow6);  // ../RTL/cortexm0ds_logic.v(12218)
  not u14044 (Tujow6, n3871);  // ../RTL/cortexm0ds_logic.v(12218)
  and u14045 (Pejow6, Xwjow6, Exjow6);  // ../RTL/cortexm0ds_logic.v(12219)
  and u14046 (n3872, Fmdow6, Cv6ow6);  // ../RTL/cortexm0ds_logic.v(12220)
  not u14047 (Exjow6, n3872);  // ../RTL/cortexm0ds_logic.v(12220)
  and u14048 (n3873, Lxjow6, Sxjow6);  // ../RTL/cortexm0ds_logic.v(12221)
  not u14049 (Cv6ow6, n3873);  // ../RTL/cortexm0ds_logic.v(12221)
  buf u1405 (vis_pc_o[10], Mw5bx6);  // ../RTL/cortexm0ds_logic.v(2011)
  or u14050 (Sxjow6, Iydow6, Wfviu6);  // ../RTL/cortexm0ds_logic.v(12222)
  and u14051 (Wfviu6, Zxjow6, Gyjow6);  // ../RTL/cortexm0ds_logic.v(12223)
  and u14052 (n3874, F0eow6, Vbgpw6[25]);  // ../RTL/cortexm0ds_logic.v(12224)
  not u14053 (Gyjow6, n3874);  // ../RTL/cortexm0ds_logic.v(12224)
  and u14054 (Zxjow6, Nyjow6, Yreow6);  // ../RTL/cortexm0ds_logic.v(12225)
  and u14055 (n3875, M0eow6, Odgpw6[25]);  // ../RTL/cortexm0ds_logic.v(12226)
  not u14056 (Nyjow6, n3875);  // ../RTL/cortexm0ds_logic.v(12226)
  and u14057 (Lxjow6, Uyjow6, Bzjow6);  // ../RTL/cortexm0ds_logic.v(12227)
  and u14058 (n3876, C2eow6, Izjow6);  // ../RTL/cortexm0ds_logic.v(12228)
  not u14059 (Bzjow6, n3876);  // ../RTL/cortexm0ds_logic.v(12228)
  buf u1406 (S8fpw6[11], Rkkax6);  // ../RTL/cortexm0ds_logic.v(2451)
  and u14060 (n3877, Pzjow6, Wzjow6);  // ../RTL/cortexm0ds_logic.v(12229)
  not u14061 (Izjow6, n3877);  // ../RTL/cortexm0ds_logic.v(12229)
  or u14062 (Wzjow6, D0kow6, Bz3ju6);  // ../RTL/cortexm0ds_logic.v(12230)
  and u14063 (n3878, M84ju6, K0kow6);  // ../RTL/cortexm0ds_logic.v(12231)
  not u14064 (Pzjow6, n3878);  // ../RTL/cortexm0ds_logic.v(12231)
  or u14065 (K0kow6, V94ju6, Hv3ju6);  // ../RTL/cortexm0ds_logic.v(12232)
  and u14066 (J34ju6, R0kow6, Y0kow6);  // ../RTL/cortexm0ds_logic.v(12233)
  not u14067 (V94ju6, J34ju6);  // ../RTL/cortexm0ds_logic.v(12233)
  and u14068 (Y0kow6, F1kow6, M1kow6);  // ../RTL/cortexm0ds_logic.v(12234)
  or u14069 (M1kow6, Ipfow6, T60iu6);  // ../RTL/cortexm0ds_logic.v(12235)
  buf u1407 (vis_pc_o[11], Knhax6);  // ../RTL/cortexm0ds_logic.v(2011)
  or u14070 (F1kow6, Ppfow6, O70iu6);  // ../RTL/cortexm0ds_logic.v(12236)
  and u14071 (R0kow6, T1kow6, A2kow6);  // ../RTL/cortexm0ds_logic.v(12237)
  or u14072 (A2kow6, Kqfow6, H70iu6);  // ../RTL/cortexm0ds_logic.v(12238)
  or u14073 (T1kow6, Rqfow6, A70iu6);  // ../RTL/cortexm0ds_logic.v(12239)
  and u14074 (M84ju6, H2kow6, D0kow6);  // ../RTL/cortexm0ds_logic.v(12240)
  and u14075 (n3879, O2kow6, Jbjow6);  // ../RTL/cortexm0ds_logic.v(12241)
  not u14076 (D0kow6, n3879);  // ../RTL/cortexm0ds_logic.v(12241)
  AL_MUX u14077 (
    .i0(Qbjow6),
    .i1(V2kow6),
    .sel(Sveow6),
    .o(O2kow6));  // ../RTL/cortexm0ds_logic.v(12242)
  or u14078 (Sveow6, C3kow6, Gweow6);  // ../RTL/cortexm0ds_logic.v(12243)
  and u14079 (n3880, Nweow6, Hv3ju6);  // ../RTL/cortexm0ds_logic.v(12244)
  buf u1408 (Iahpw6[1], Li7ax6);  // ../RTL/cortexm0ds_logic.v(1883)
  not u14080 (H2kow6, n3880);  // ../RTL/cortexm0ds_logic.v(12244)
  and u14081 (Nweow6, J3kow6, Q3kow6);  // ../RTL/cortexm0ds_logic.v(12245)
  and u14082 (Q3kow6, X3kow6, E4kow6);  // ../RTL/cortexm0ds_logic.v(12246)
  or u14083 (E4kow6, Ipfow6, Dc0iu6);  // ../RTL/cortexm0ds_logic.v(12247)
  or u14084 (X3kow6, Rqfow6, R50iu6);  // ../RTL/cortexm0ds_logic.v(12248)
  and u14085 (J3kow6, L4kow6, S4kow6);  // ../RTL/cortexm0ds_logic.v(12249)
  or u14086 (S4kow6, Ppfow6, M60iu6);  // ../RTL/cortexm0ds_logic.v(12250)
  or u14087 (L4kow6, Kqfow6, Y50iu6);  // ../RTL/cortexm0ds_logic.v(12251)
  and u14088 (n3881, HRDATA[25], Q2eow6);  // ../RTL/cortexm0ds_logic.v(12252)
  not u14089 (Uyjow6, n3881);  // ../RTL/cortexm0ds_logic.v(12252)
  buf u1409 (vis_pc_o[12], Nlhax6);  // ../RTL/cortexm0ds_logic.v(2011)
  or u14090 (Xwjow6, Kldow6, Ou6ow6);  // ../RTL/cortexm0ds_logic.v(12253)
  and u14091 (Ou6ow6, Z4kow6, G5kow6);  // ../RTL/cortexm0ds_logic.v(12254)
  and u14092 (G5kow6, N5kow6, U5kow6);  // ../RTL/cortexm0ds_logic.v(12255)
  or u14093 (U5kow6, Rcfow6, F14ju6);  // ../RTL/cortexm0ds_logic.v(12256)
  and u14094 (F14ju6, B6kow6, I6kow6);  // ../RTL/cortexm0ds_logic.v(12257)
  and u14095 (I6kow6, P6kow6, W6kow6);  // ../RTL/cortexm0ds_logic.v(12258)
  or u14096 (W6kow6, Ipfow6, V70iu6);  // ../RTL/cortexm0ds_logic.v(12259)
  or u14097 (P6kow6, Rqfow6, C80iu6);  // ../RTL/cortexm0ds_logic.v(12260)
  and u14098 (B6kow6, D7kow6, K7kow6);  // ../RTL/cortexm0ds_logic.v(12261)
  or u14099 (K7kow6, Ppfow6, Q80iu6);  // ../RTL/cortexm0ds_logic.v(12262)
  buf u141 (H4ghu6, Hirpw6);  // ../RTL/cortexm0ds_logic.v(1950)
  buf u1410 (Iahpw6[2], Bx2qw6);  // ../RTL/cortexm0ds_logic.v(1883)
  or u14100 (D7kow6, Kqfow6, J80iu6);  // ../RTL/cortexm0ds_logic.v(12263)
  or u14101 (N5kow6, Iydow6, Nutiu6);  // ../RTL/cortexm0ds_logic.v(12264)
  and u14102 (Nutiu6, R7kow6, Y7kow6);  // ../RTL/cortexm0ds_logic.v(12265)
  and u14103 (Y7kow6, F8kow6, M8kow6);  // ../RTL/cortexm0ds_logic.v(12266)
  and u14104 (n3882, Tzfpw6[17], Yvgiu6);  // ../RTL/cortexm0ds_logic.v(12267)
  not u14105 (M8kow6, n3882);  // ../RTL/cortexm0ds_logic.v(12267)
  and u14106 (F8kow6, T8kow6, A9kow6);  // ../RTL/cortexm0ds_logic.v(12268)
  or u14107 (A9kow6, W6ciu6, Qkgiu6);  // ../RTL/cortexm0ds_logic.v(12269)
  and u14108 (n3883, H9kow6, Ydeow6);  // ../RTL/cortexm0ds_logic.v(12270)
  not u14109 (W6ciu6, n3883);  // ../RTL/cortexm0ds_logic.v(12270)
  buf u1411 (vis_pc_o[13], Qjhax6);  // ../RTL/cortexm0ds_logic.v(2011)
  or u14110 (n3884, Feeow6, E2fow6);  // ../RTL/cortexm0ds_logic.v(12271)
  not u14111 (H9kow6, n3884);  // ../RTL/cortexm0ds_logic.v(12271)
  and u14112 (n3885, Odgpw6[17], M0eow6);  // ../RTL/cortexm0ds_logic.v(12272)
  not u14113 (T8kow6, n3885);  // ../RTL/cortexm0ds_logic.v(12272)
  and u14114 (R7kow6, O9kow6, V9kow6);  // ../RTL/cortexm0ds_logic.v(12273)
  and u14115 (n3886, F0eow6, Vbgpw6[17]);  // ../RTL/cortexm0ds_logic.v(12274)
  not u14116 (V9kow6, n3886);  // ../RTL/cortexm0ds_logic.v(12274)
  and u14117 (O9kow6, Cakow6, Jakow6);  // ../RTL/cortexm0ds_logic.v(12275)
  and u14118 (n3887, STCALIB[17], H1eow6);  // ../RTL/cortexm0ds_logic.v(12276)
  not u14119 (Jakow6, n3887);  // ../RTL/cortexm0ds_logic.v(12276)
  buf u1412 (Iahpw6[3], Z73qw6);  // ../RTL/cortexm0ds_logic.v(1883)
  and u14120 (n3888, Bagpw6[17], M6eiu6);  // ../RTL/cortexm0ds_logic.v(12277)
  not u14121 (Cakow6, n3888);  // ../RTL/cortexm0ds_logic.v(12277)
  and u14122 (Z4kow6, Qakow6, Xakow6);  // ../RTL/cortexm0ds_logic.v(12278)
  and u14123 (n3889, Qtfow6, Ff4ju6);  // ../RTL/cortexm0ds_logic.v(12279)
  not u14124 (Xakow6, n3889);  // ../RTL/cortexm0ds_logic.v(12279)
  and u14125 (n3890, Ebkow6, Lbkow6);  // ../RTL/cortexm0ds_logic.v(12280)
  not u14126 (Ff4ju6, n3890);  // ../RTL/cortexm0ds_logic.v(12280)
  and u14127 (Lbkow6, Sbkow6, Zbkow6);  // ../RTL/cortexm0ds_logic.v(12281)
  or u14128 (Zbkow6, Ipfow6, X80iu6);  // ../RTL/cortexm0ds_logic.v(12282)
  or u14129 (Sbkow6, Rqfow6, L90iu6);  // ../RTL/cortexm0ds_logic.v(12283)
  buf u1413 (vis_pc_o[14], Cq7bx6);  // ../RTL/cortexm0ds_logic.v(2011)
  and u14130 (Ebkow6, Gckow6, Nckow6);  // ../RTL/cortexm0ds_logic.v(12284)
  or u14131 (Nckow6, Ppfow6, Z90iu6);  // ../RTL/cortexm0ds_logic.v(12285)
  or u14132 (Gckow6, Kqfow6, S90iu6);  // ../RTL/cortexm0ds_logic.v(12286)
  and u14133 (n3891, HRDATA[17], Q2eow6);  // ../RTL/cortexm0ds_logic.v(12287)
  not u14134 (Qakow6, n3891);  // ../RTL/cortexm0ds_logic.v(12287)
  and u14135 (Gdjow6, Uckow6, Bdkow6);  // ../RTL/cortexm0ds_logic.v(12288)
  and u14136 (n3892, Zsfpw6[8], Cmziu6);  // ../RTL/cortexm0ds_logic.v(12289)
  not u14137 (Bdkow6, n3892);  // ../RTL/cortexm0ds_logic.v(12289)
  and u14138 (n3893, vis_pc_o[8], Jmziu6);  // ../RTL/cortexm0ds_logic.v(12290)
  not u14139 (Uckow6, n3893);  // ../RTL/cortexm0ds_logic.v(12290)
  buf u1414 (Iahpw6[4], D2opw6);  // ../RTL/cortexm0ds_logic.v(1883)
  and u14140 (n3894, Idkow6, Pdkow6);  // ../RTL/cortexm0ds_logic.v(12291)
  not u14141 (Vcohu6, n3894);  // ../RTL/cortexm0ds_logic.v(12291)
  and u14142 (Pdkow6, Wdkow6, Dekow6);  // ../RTL/cortexm0ds_logic.v(12292)
  and u14143 (n3895, Egziu6, Eafpw6[15]);  // ../RTL/cortexm0ds_logic.v(12293)
  not u14144 (Dekow6, n3895);  // ../RTL/cortexm0ds_logic.v(12293)
  and u14145 (Wdkow6, Kekow6, Sgziu6);  // ../RTL/cortexm0ds_logic.v(12294)
  or u14146 (Kekow6, Ft6ow6, Ggmiu6);  // ../RTL/cortexm0ds_logic.v(12295)
  and u14147 (Ggmiu6, Rekow6, Yekow6);  // ../RTL/cortexm0ds_logic.v(12296)
  and u14148 (Yekow6, Ffkow6, Mfkow6);  // ../RTL/cortexm0ds_logic.v(12297)
  or u14149 (Mfkow6, H78ow6, Kldow6);  // ../RTL/cortexm0ds_logic.v(12298)
  buf u1415 (vis_pc_o[15], Thhax6);  // ../RTL/cortexm0ds_logic.v(2011)
  and u14150 (Ffkow6, Tfkow6, Dldow6);  // ../RTL/cortexm0ds_logic.v(12299)
  and u14151 (n3896, Mmdow6, X88ow6);  // ../RTL/cortexm0ds_logic.v(12300)
  not u14152 (Tfkow6, n3896);  // ../RTL/cortexm0ds_logic.v(12300)
  and u14153 (Rekow6, Agkow6, Hgkow6);  // ../RTL/cortexm0ds_logic.v(12301)
  and u14154 (n3897, V78ow6, Fmdow6);  // ../RTL/cortexm0ds_logic.v(12302)
  not u14155 (Hgkow6, n3897);  // ../RTL/cortexm0ds_logic.v(12302)
  or u14156 (Agkow6, Q88ow6, Pkdow6);  // ../RTL/cortexm0ds_logic.v(12303)
  and u14157 (Idkow6, Ogkow6, Vgkow6);  // ../RTL/cortexm0ds_logic.v(12304)
  and u14158 (n3898, Zsfpw6[14], Cmziu6);  // ../RTL/cortexm0ds_logic.v(12305)
  not u14159 (Vgkow6, n3898);  // ../RTL/cortexm0ds_logic.v(12305)
  buf u1416 (Iahpw6[5], Zgfax6);  // ../RTL/cortexm0ds_logic.v(1883)
  and u14160 (n3899, vis_pc_o[14], Jmziu6);  // ../RTL/cortexm0ds_logic.v(12306)
  not u14161 (Ogkow6, n3899);  // ../RTL/cortexm0ds_logic.v(12306)
  and u14162 (n3900, Chkow6, Jhkow6);  // ../RTL/cortexm0ds_logic.v(12307)
  not u14163 (Ocohu6, n3900);  // ../RTL/cortexm0ds_logic.v(12307)
  and u14164 (Jhkow6, Qhkow6, Xhkow6);  // ../RTL/cortexm0ds_logic.v(12308)
  and u14165 (n3901, Zsfpw6[21], Cmziu6);  // ../RTL/cortexm0ds_logic.v(12309)
  not u14166 (Xhkow6, n3901);  // ../RTL/cortexm0ds_logic.v(12309)
  and u14167 (Qhkow6, Eikow6, Likow6);  // ../RTL/cortexm0ds_logic.v(12310)
  or u14168 (Likow6, Ft6ow6, Nvliu6);  // ../RTL/cortexm0ds_logic.v(12311)
  and u14169 (Nvliu6, Sikow6, Zikow6);  // ../RTL/cortexm0ds_logic.v(12312)
  buf u1417 (vis_pc_o[16], Wfhax6);  // ../RTL/cortexm0ds_logic.v(2011)
  and u14170 (Zikow6, Gjkow6, Njkow6);  // ../RTL/cortexm0ds_logic.v(12313)
  or u14171 (Njkow6, G6cow6, Eccow6);  // ../RTL/cortexm0ds_logic.v(12314)
  and u14172 (G6cow6, Ujkow6, Bkkow6);  // ../RTL/cortexm0ds_logic.v(12315)
  and u14173 (Bkkow6, Ikkow6, Pkkow6);  // ../RTL/cortexm0ds_logic.v(12316)
  or u14174 (Pkkow6, Rcfow6, Wkkow6);  // ../RTL/cortexm0ds_logic.v(12317)
  or u14175 (Ikkow6, Iydow6, Ntuiu6);  // ../RTL/cortexm0ds_logic.v(12319)
  and u14176 (Ntuiu6, Dlkow6, Klkow6);  // ../RTL/cortexm0ds_logic.v(12320)
  and u14177 (Klkow6, Rlkow6, Ylkow6);  // ../RTL/cortexm0ds_logic.v(12321)
  and u14178 (Ylkow6, Fmkow6, Mmkow6);  // ../RTL/cortexm0ds_logic.v(12322)
  and u14179 (Mmkow6, Tmkow6, Ankow6);  // ../RTL/cortexm0ds_logic.v(12323)
  buf u1418 (Iahpw6[6], Yzlpw6);  // ../RTL/cortexm0ds_logic.v(1883)
  and u14180 (n3902, Odgpw6[22], M0eow6);  // ../RTL/cortexm0ds_logic.v(12324)
  not u14181 (Ankow6, n3902);  // ../RTL/cortexm0ds_logic.v(12324)
  and u14182 (n3903, STCALIB[22], H1eow6);  // ../RTL/cortexm0ds_logic.v(12325)
  not u14183 (Tmkow6, n3903);  // ../RTL/cortexm0ds_logic.v(12325)
  and u14184 (Fmkow6, Hnkow6, Onkow6);  // ../RTL/cortexm0ds_logic.v(12326)
  and u14185 (n3904, Tzdiu6, R4gpw6[4]);  // ../RTL/cortexm0ds_logic.v(12327)
  not u14186 (Onkow6, n3904);  // ../RTL/cortexm0ds_logic.v(12327)
  and u14187 (n3905, I3fiu6, R4gpw6[12]);  // ../RTL/cortexm0ds_logic.v(12328)
  not u14188 (Hnkow6, n3905);  // ../RTL/cortexm0ds_logic.v(12328)
  and u14189 (Rlkow6, Vnkow6, Cokow6);  // ../RTL/cortexm0ds_logic.v(12329)
  or u1419 (n111[0], Xuzhu6, N30iu6);  // ../RTL/cortexm0ds_logic.v(3385)
  and u14190 (Cokow6, Jokow6, Qokow6);  // ../RTL/cortexm0ds_logic.v(12330)
  and u14191 (n3906, Tzfpw6[22], Yvgiu6);  // ../RTL/cortexm0ds_logic.v(12331)
  not u14192 (Qokow6, n3906);  // ../RTL/cortexm0ds_logic.v(12331)
  and u14193 (n3907, Hqgiu6, L1gpw6[0]);  // ../RTL/cortexm0ds_logic.v(12332)
  not u14194 (Jokow6, n3907);  // ../RTL/cortexm0ds_logic.v(12332)
  and u14195 (Vnkow6, Xokow6, Epkow6);  // ../RTL/cortexm0ds_logic.v(12333)
  and u14196 (n3908, S1fiu6, R4gpw6[36]);  // ../RTL/cortexm0ds_logic.v(12334)
  not u14197 (Epkow6, n3908);  // ../RTL/cortexm0ds_logic.v(12334)
  and u14198 (n3909, G2fiu6, R4gpw6[28]);  // ../RTL/cortexm0ds_logic.v(12335)
  not u14199 (Xokow6, n3909);  // ../RTL/cortexm0ds_logic.v(12335)
  buf u142 (vis_r2_o[10], U8rax6);  // ../RTL/cortexm0ds_logic.v(2551)
  buf u1420 (Fkfpw6[0], I1lpw6);  // ../RTL/cortexm0ds_logic.v(1881)
  and u14200 (Dlkow6, Lpkow6, Spkow6);  // ../RTL/cortexm0ds_logic.v(12336)
  and u14201 (Spkow6, Zpkow6, Gqkow6);  // ../RTL/cortexm0ds_logic.v(12337)
  and u14202 (Gqkow6, Nqkow6, Uqkow6);  // ../RTL/cortexm0ds_logic.v(12338)
  and u14203 (n3910, C0fiu6, R4gpw6[60]);  // ../RTL/cortexm0ds_logic.v(12339)
  not u14204 (Uqkow6, n3910);  // ../RTL/cortexm0ds_logic.v(12339)
  and u14205 (n3911, F0eow6, Vbgpw6[22]);  // ../RTL/cortexm0ds_logic.v(12340)
  not u14206 (Nqkow6, n3911);  // ../RTL/cortexm0ds_logic.v(12340)
  and u14207 (Zpkow6, Brkow6, Irkow6);  // ../RTL/cortexm0ds_logic.v(12341)
  and u14208 (n3912, Bagpw6[22], M6eiu6);  // ../RTL/cortexm0ds_logic.v(12342)
  not u14209 (Irkow6, n3912);  // ../RTL/cortexm0ds_logic.v(12342)
  buf u1421 (vis_psp_o[18], X4jpw6);  // ../RTL/cortexm0ds_logic.v(2085)
  and u14210 (n3913, E1fiu6, R4gpw6[44]);  // ../RTL/cortexm0ds_logic.v(12343)
  not u14211 (Brkow6, n3913);  // ../RTL/cortexm0ds_logic.v(12343)
  and u14212 (Lpkow6, Prkow6, Wrkow6);  // ../RTL/cortexm0ds_logic.v(12344)
  and u14213 (n3914, T7eow6, Dskow6);  // ../RTL/cortexm0ds_logic.v(12345)
  not u14214 (Wrkow6, n3914);  // ../RTL/cortexm0ds_logic.v(12345)
  and u14215 (n3915, Kskow6, Rskow6);  // ../RTL/cortexm0ds_logic.v(12346)
  not u14216 (Dskow6, n3915);  // ../RTL/cortexm0ds_logic.v(12346)
  and u14217 (Rskow6, Yskow6, Ftkow6);  // ../RTL/cortexm0ds_logic.v(12347)
  and u14218 (Ftkow6, Mtkow6, Ttkow6);  // ../RTL/cortexm0ds_logic.v(12348)
  and u14219 (Ttkow6, Aukow6, Hukow6);  // ../RTL/cortexm0ds_logic.v(12349)
  buf u1422 (vis_pc_o[20], I8hax6);  // ../RTL/cortexm0ds_logic.v(2011)
  or u14220 (n3916, Odgpw6[8], Odgpw6[9]);  // ../RTL/cortexm0ds_logic.v(12350)
  not u14221 (Hukow6, n3916);  // ../RTL/cortexm0ds_logic.v(12350)
  or u14222 (n3917, Odgpw6[6], Odgpw6[7]);  // ../RTL/cortexm0ds_logic.v(12351)
  not u14223 (Aukow6, n3917);  // ../RTL/cortexm0ds_logic.v(12351)
  and u14224 (Mtkow6, Oukow6, Vukow6);  // ../RTL/cortexm0ds_logic.v(12352)
  or u14225 (n3918, Odgpw6[4], Odgpw6[5]);  // ../RTL/cortexm0ds_logic.v(12353)
  not u14226 (Vukow6, n3918);  // ../RTL/cortexm0ds_logic.v(12353)
  or u14227 (n3919, Odgpw6[31], Odgpw6[3]);  // ../RTL/cortexm0ds_logic.v(12354)
  not u14228 (Oukow6, n3919);  // ../RTL/cortexm0ds_logic.v(12354)
  and u14229 (Yskow6, Cvkow6, Jvkow6);  // ../RTL/cortexm0ds_logic.v(12355)
  buf u1423 (vis_pc_o[17], Zdhax6);  // ../RTL/cortexm0ds_logic.v(2011)
  and u14230 (Jvkow6, Qvkow6, Xvkow6);  // ../RTL/cortexm0ds_logic.v(12356)
  or u14231 (n3920, Odgpw6[2], Odgpw6[30]);  // ../RTL/cortexm0ds_logic.v(12357)
  not u14232 (Xvkow6, n3920);  // ../RTL/cortexm0ds_logic.v(12357)
  or u14233 (n3921, Odgpw6[28], Odgpw6[29]);  // ../RTL/cortexm0ds_logic.v(12358)
  not u14234 (Qvkow6, n3921);  // ../RTL/cortexm0ds_logic.v(12358)
  and u14235 (Cvkow6, Ewkow6, Lwkow6);  // ../RTL/cortexm0ds_logic.v(12359)
  or u14236 (n3922, Odgpw6[26], Odgpw6[27]);  // ../RTL/cortexm0ds_logic.v(12360)
  not u14237 (Lwkow6, n3922);  // ../RTL/cortexm0ds_logic.v(12360)
  or u14238 (n3923, Odgpw6[24], Odgpw6[25]);  // ../RTL/cortexm0ds_logic.v(12361)
  not u14239 (Ewkow6, n3923);  // ../RTL/cortexm0ds_logic.v(12361)
  buf u1424 (Iahpw6[7], Qa1qw6);  // ../RTL/cortexm0ds_logic.v(1883)
  and u14240 (Kskow6, Swkow6, Zwkow6);  // ../RTL/cortexm0ds_logic.v(12362)
  and u14241 (Zwkow6, Gxkow6, Nxkow6);  // ../RTL/cortexm0ds_logic.v(12363)
  and u14242 (Nxkow6, Uxkow6, Bykow6);  // ../RTL/cortexm0ds_logic.v(12364)
  or u14243 (n3924, Odgpw6[22], Odgpw6[23]);  // ../RTL/cortexm0ds_logic.v(12365)
  not u14244 (Bykow6, n3924);  // ../RTL/cortexm0ds_logic.v(12365)
  or u14245 (n3925, Odgpw6[20], Odgpw6[21]);  // ../RTL/cortexm0ds_logic.v(12366)
  not u14246 (Uxkow6, n3925);  // ../RTL/cortexm0ds_logic.v(12366)
  and u14247 (Gxkow6, Iykow6, Pykow6);  // ../RTL/cortexm0ds_logic.v(12367)
  or u14248 (n3926, Odgpw6[19], Odgpw6[1]);  // ../RTL/cortexm0ds_logic.v(12368)
  not u14249 (Pykow6, n3926);  // ../RTL/cortexm0ds_logic.v(12368)
  buf u1425 (vis_psp_o[19], Rfkpw6);  // ../RTL/cortexm0ds_logic.v(2085)
  or u14250 (n3927, Odgpw6[17], Odgpw6[18]);  // ../RTL/cortexm0ds_logic.v(12369)
  not u14251 (Iykow6, n3927);  // ../RTL/cortexm0ds_logic.v(12369)
  and u14252 (Swkow6, Wykow6, Dzkow6);  // ../RTL/cortexm0ds_logic.v(12370)
  and u14253 (Dzkow6, Kzkow6, Rzkow6);  // ../RTL/cortexm0ds_logic.v(12371)
  or u14254 (n3928, Odgpw6[15], Odgpw6[16]);  // ../RTL/cortexm0ds_logic.v(12372)
  not u14255 (Rzkow6, n3928);  // ../RTL/cortexm0ds_logic.v(12372)
  or u14256 (n3929, Odgpw6[13], Odgpw6[14]);  // ../RTL/cortexm0ds_logic.v(12373)
  not u14257 (Kzkow6, n3929);  // ../RTL/cortexm0ds_logic.v(12373)
  and u14258 (Wykow6, Yzkow6, F0low6);  // ../RTL/cortexm0ds_logic.v(12374)
  or u14259 (n3930, Odgpw6[11], Odgpw6[12]);  // ../RTL/cortexm0ds_logic.v(12375)
  buf u1426 (vis_pc_o[21], Nxabx6);  // ../RTL/cortexm0ds_logic.v(2011)
  not u14260 (F0low6, n3930);  // ../RTL/cortexm0ds_logic.v(12375)
  or u14261 (n3931, Odgpw6[0], Odgpw6[10]);  // ../RTL/cortexm0ds_logic.v(12376)
  not u14262 (Yzkow6, n3931);  // ../RTL/cortexm0ds_logic.v(12376)
  and u14263 (Prkow6, M0low6, T0low6);  // ../RTL/cortexm0ds_logic.v(12377)
  and u14264 (n3932, Q0fiu6, R4gpw6[52]);  // ../RTL/cortexm0ds_logic.v(12378)
  not u14265 (T0low6, n3932);  // ../RTL/cortexm0ds_logic.v(12378)
  and u14266 (n3933, U2fiu6, R4gpw6[20]);  // ../RTL/cortexm0ds_logic.v(12379)
  not u14267 (M0low6, n3933);  // ../RTL/cortexm0ds_logic.v(12379)
  and u14268 (Ujkow6, A1low6, H1low6);  // ../RTL/cortexm0ds_logic.v(12380)
  or u14269 (H1low6, Uafow6, R04ju6);  // ../RTL/cortexm0ds_logic.v(12381)
  buf u1427 (vis_psp_o[20], Thfbx6);  // ../RTL/cortexm0ds_logic.v(2085)
  and u14270 (n3934, HRDATA[22], Q2eow6);  // ../RTL/cortexm0ds_logic.v(12382)
  not u14271 (A1low6, n3934);  // ../RTL/cortexm0ds_logic.v(12382)
  or u14272 (Gjkow6, L5cow6, Vacow6);  // ../RTL/cortexm0ds_logic.v(12383)
  and u14273 (Vacow6, O1low6, Dtcow6);  // ../RTL/cortexm0ds_logic.v(12384)
  and u14274 (L5cow6, V1low6, C2low6);  // ../RTL/cortexm0ds_logic.v(12385)
  and u14275 (C2low6, J2low6, Q2low6);  // ../RTL/cortexm0ds_logic.v(12386)
  and u14276 (n3935, Dyeow6, Ye4ju6);  // ../RTL/cortexm0ds_logic.v(12387)
  not u14277 (Q2low6, n3935);  // ../RTL/cortexm0ds_logic.v(12387)
  or u14278 (J2low6, Iydow6, N9tiu6);  // ../RTL/cortexm0ds_logic.v(12388)
  and u14279 (N9tiu6, X2low6, E3low6);  // ../RTL/cortexm0ds_logic.v(12389)
  buf u1428 (vis_pc_o[22], C37ax6);  // ../RTL/cortexm0ds_logic.v(2011)
  and u14280 (E3low6, L3low6, S3low6);  // ../RTL/cortexm0ds_logic.v(12390)
  and u14281 (S3low6, Z3low6, G4low6);  // ../RTL/cortexm0ds_logic.v(12391)
  and u14282 (G4low6, N4low6, U4low6);  // ../RTL/cortexm0ds_logic.v(12392)
  and u14283 (n3936, Tzdiu6, R4gpw6[2]);  // ../RTL/cortexm0ds_logic.v(12393)
  not u14284 (U4low6, n3936);  // ../RTL/cortexm0ds_logic.v(12393)
  and u14285 (n3937, S1fiu6, R4gpw6[34]);  // ../RTL/cortexm0ds_logic.v(12394)
  not u14286 (N4low6, n3937);  // ../RTL/cortexm0ds_logic.v(12394)
  and u14287 (Z3low6, B5low6, I5low6);  // ../RTL/cortexm0ds_logic.v(12395)
  and u14288 (n3938, STCALIB[14], H1eow6);  // ../RTL/cortexm0ds_logic.v(12396)
  not u14289 (I5low6, n3938);  // ../RTL/cortexm0ds_logic.v(12396)
  buf u1429 (vis_psp_o[21], Gr6ax6);  // ../RTL/cortexm0ds_logic.v(2085)
  and u14290 (n3939, F0eow6, Vbgpw6[14]);  // ../RTL/cortexm0ds_logic.v(12397)
  not u14291 (B5low6, n3939);  // ../RTL/cortexm0ds_logic.v(12397)
  and u14292 (L3low6, P5low6, W5low6);  // ../RTL/cortexm0ds_logic.v(12398)
  and u14293 (W5low6, D6low6, K6low6);  // ../RTL/cortexm0ds_logic.v(12399)
  and u14294 (n3940, U2fiu6, R4gpw6[18]);  // ../RTL/cortexm0ds_logic.v(12400)
  not u14295 (K6low6, n3940);  // ../RTL/cortexm0ds_logic.v(12400)
  and u14296 (n3941, I3fiu6, R4gpw6[10]);  // ../RTL/cortexm0ds_logic.v(12401)
  not u14297 (D6low6, n3941);  // ../RTL/cortexm0ds_logic.v(12401)
  and u14298 (P5low6, R6low6, Y6low6);  // ../RTL/cortexm0ds_logic.v(12402)
  or u14299 (Y6low6, U5ciu6, Qkgiu6);  // ../RTL/cortexm0ds_logic.v(12403)
  buf u143 (Trgpw6[17], Hpbbx6);  // ../RTL/cortexm0ds_logic.v(2376)
  buf u1430 (vis_pc_o[23], L6hax6);  // ../RTL/cortexm0ds_logic.v(2011)
  and u14300 (n3942, Ydeow6, F7low6);  // ../RTL/cortexm0ds_logic.v(12404)
  not u14301 (U5ciu6, n3942);  // ../RTL/cortexm0ds_logic.v(12404)
  and u14302 (n3943, Okgow6, M7low6);  // ../RTL/cortexm0ds_logic.v(12405)
  not u14303 (F7low6, n3943);  // ../RTL/cortexm0ds_logic.v(12405)
  and u14304 (n3944, T7low6, A8low6);  // ../RTL/cortexm0ds_logic.v(12406)
  not u14305 (M7low6, n3944);  // ../RTL/cortexm0ds_logic.v(12406)
  and u14306 (n3945, H8low6, O8low6);  // ../RTL/cortexm0ds_logic.v(12407)
  not u14307 (T7low6, n3945);  // ../RTL/cortexm0ds_logic.v(12407)
  AL_MUX u14308 (
    .i0(V8low6),
    .i1(C9low6),
    .sel(E2fow6),
    .o(H8low6));  // ../RTL/cortexm0ds_logic.v(12408)
  or u14309 (n3946, Z2fow6, J9low6);  // ../RTL/cortexm0ds_logic.v(12409)
  buf u1431 (vis_psp_o[22], Z8zpw6);  // ../RTL/cortexm0ds_logic.v(2085)
  not u14310 (C9low6, n3946);  // ../RTL/cortexm0ds_logic.v(12409)
  or u14311 (n3947, B4fow6, Nggow6);  // ../RTL/cortexm0ds_logic.v(12410)
  not u14312 (J9low6, n3947);  // ../RTL/cortexm0ds_logic.v(12410)
  and u14313 (V8low6, F6fow6, Q9low6);  // ../RTL/cortexm0ds_logic.v(12411)
  or u14314 (Q9low6, H7fow6, Hdgow6);  // ../RTL/cortexm0ds_logic.v(12412)
  and u14315 (n3948, Q0fiu6, R4gpw6[50]);  // ../RTL/cortexm0ds_logic.v(12413)
  not u14316 (R6low6, n3948);  // ../RTL/cortexm0ds_logic.v(12413)
  and u14317 (X2low6, X9low6, Ealow6);  // ../RTL/cortexm0ds_logic.v(12414)
  and u14318 (Ealow6, Lalow6, Salow6);  // ../RTL/cortexm0ds_logic.v(12415)
  and u14319 (Salow6, Zalow6, Gblow6);  // ../RTL/cortexm0ds_logic.v(12416)
  buf u1432 (vis_pc_o[24], O4hax6);  // ../RTL/cortexm0ds_logic.v(2011)
  and u14320 (n3949, Tzfpw6[14], Yvgiu6);  // ../RTL/cortexm0ds_logic.v(12417)
  not u14321 (Gblow6, n3949);  // ../RTL/cortexm0ds_logic.v(12417)
  and u14322 (n3950, Odgpw6[14], M0eow6);  // ../RTL/cortexm0ds_logic.v(12418)
  not u14323 (Zalow6, n3950);  // ../RTL/cortexm0ds_logic.v(12418)
  and u14324 (Lalow6, Nblow6, Ublow6);  // ../RTL/cortexm0ds_logic.v(12419)
  and u14325 (n3951, C0fiu6, R4gpw6[58]);  // ../RTL/cortexm0ds_logic.v(12420)
  not u14326 (Ublow6, n3951);  // ../RTL/cortexm0ds_logic.v(12420)
  and u14327 (n3952, E1fiu6, R4gpw6[42]);  // ../RTL/cortexm0ds_logic.v(12421)
  not u14328 (Nblow6, n3952);  // ../RTL/cortexm0ds_logic.v(12421)
  and u14329 (X9low6, Bclow6, Qgeow6);  // ../RTL/cortexm0ds_logic.v(12422)
  buf u1433 (vis_psp_o[23], Zbtpw6);  // ../RTL/cortexm0ds_logic.v(2085)
  and u14330 (Bclow6, Iclow6, Pclow6);  // ../RTL/cortexm0ds_logic.v(12423)
  and u14331 (n3953, Bagpw6[14], M6eiu6);  // ../RTL/cortexm0ds_logic.v(12424)
  not u14332 (Pclow6, n3953);  // ../RTL/cortexm0ds_logic.v(12424)
  and u14333 (n3954, G2fiu6, R4gpw6[26]);  // ../RTL/cortexm0ds_logic.v(12425)
  not u14334 (Iclow6, n3954);  // ../RTL/cortexm0ds_logic.v(12425)
  and u14335 (V1low6, Wclow6, Ddlow6);  // ../RTL/cortexm0ds_logic.v(12426)
  or u14336 (Ddlow6, Uafow6, Id4ju6);  // ../RTL/cortexm0ds_logic.v(12427)
  and u14337 (n3955, HRDATA[14], Q2eow6);  // ../RTL/cortexm0ds_logic.v(12428)
  not u14338 (Wclow6, n3955);  // ../RTL/cortexm0ds_logic.v(12428)
  and u14339 (Sikow6, Kdlow6, Rdlow6);  // ../RTL/cortexm0ds_logic.v(12429)
  buf u1434 (vis_pc_o[25], R2hax6);  // ../RTL/cortexm0ds_logic.v(2011)
  and u14340 (n3956, X4cow6, Cbcow6);  // ../RTL/cortexm0ds_logic.v(12430)
  not u14341 (Rdlow6, n3956);  // ../RTL/cortexm0ds_logic.v(12430)
  and u14342 (Pzcow6, Ydlow6, W9how6);  // ../RTL/cortexm0ds_logic.v(12431)
  not u14343 (Cbcow6, Pzcow6);  // ../RTL/cortexm0ds_logic.v(12431)
  and u14344 (n3957, Felow6, Melow6);  // ../RTL/cortexm0ds_logic.v(12432)
  not u14345 (X4cow6, n3957);  // ../RTL/cortexm0ds_logic.v(12432)
  or u14346 (Melow6, Iydow6, Bewiu6);  // ../RTL/cortexm0ds_logic.v(12433)
  and u14347 (Bewiu6, Telow6, Aflow6);  // ../RTL/cortexm0ds_logic.v(12434)
  and u14348 (Aflow6, Hflow6, Oflow6);  // ../RTL/cortexm0ds_logic.v(12435)
  and u14349 (Oflow6, Vflow6, Cglow6);  // ../RTL/cortexm0ds_logic.v(12436)
  buf u1435 (vis_psp_o[24], Zazpw6);  // ../RTL/cortexm0ds_logic.v(2085)
  and u14350 (Cglow6, Jglow6, Qglow6);  // ../RTL/cortexm0ds_logic.v(12437)
  and u14351 (n3958, Odgpw6[30], M0eow6);  // ../RTL/cortexm0ds_logic.v(12438)
  not u14352 (Qglow6, n3958);  // ../RTL/cortexm0ds_logic.v(12438)
  or u14353 (Jglow6, Tpgiu6, Xglow6);  // ../RTL/cortexm0ds_logic.v(12439)
  and u14354 (Vflow6, Ehlow6, Lhlow6);  // ../RTL/cortexm0ds_logic.v(12440)
  and u14355 (n3959, E1fiu6, R4gpw6[46]);  // ../RTL/cortexm0ds_logic.v(12441)
  not u14356 (Lhlow6, n3959);  // ../RTL/cortexm0ds_logic.v(12441)
  and u14357 (n3960, Tzdiu6, R4gpw6[6]);  // ../RTL/cortexm0ds_logic.v(12442)
  not u14358 (Ehlow6, n3960);  // ../RTL/cortexm0ds_logic.v(12442)
  and u14359 (Hflow6, Shlow6, Zhlow6);  // ../RTL/cortexm0ds_logic.v(12443)
  buf u1436 (vis_pc_o[26], U0hax6);  // ../RTL/cortexm0ds_logic.v(2011)
  and u14360 (n3961, U2fiu6, R4gpw6[22]);  // ../RTL/cortexm0ds_logic.v(12444)
  not u14361 (Zhlow6, n3961);  // ../RTL/cortexm0ds_logic.v(12444)
  and u14362 (Shlow6, Gilow6, Nilow6);  // ../RTL/cortexm0ds_logic.v(12445)
  and u14363 (n3962, STCALIB[24], H1eow6);  // ../RTL/cortexm0ds_logic.v(12446)
  not u14364 (Nilow6, n3962);  // ../RTL/cortexm0ds_logic.v(12446)
  and u14365 (n3963, G2fiu6, R4gpw6[30]);  // ../RTL/cortexm0ds_logic.v(12447)
  not u14366 (Gilow6, n3963);  // ../RTL/cortexm0ds_logic.v(12447)
  and u14367 (Telow6, Uilow6, Bjlow6);  // ../RTL/cortexm0ds_logic.v(12448)
  and u14368 (Bjlow6, Ijlow6, Pjlow6);  // ../RTL/cortexm0ds_logic.v(12449)
  and u14369 (Pjlow6, Wjlow6, Dklow6);  // ../RTL/cortexm0ds_logic.v(12450)
  buf u1437 (vis_psp_o[25], Zczpw6);  // ../RTL/cortexm0ds_logic.v(2085)
  and u14370 (n3964, Hqgiu6, H8gpw6[0]);  // ../RTL/cortexm0ds_logic.v(12451)
  not u14371 (Dklow6, n3964);  // ../RTL/cortexm0ds_logic.v(12451)
  and u14372 (n3965, I3fiu6, R4gpw6[14]);  // ../RTL/cortexm0ds_logic.v(12452)
  not u14373 (Wjlow6, n3965);  // ../RTL/cortexm0ds_logic.v(12452)
  and u14374 (Ijlow6, Kklow6, Rklow6);  // ../RTL/cortexm0ds_logic.v(12453)
  and u14375 (n3966, C0fiu6, R4gpw6[62]);  // ../RTL/cortexm0ds_logic.v(12454)
  not u14376 (Rklow6, n3966);  // ../RTL/cortexm0ds_logic.v(12454)
  and u14377 (n3967, S1fiu6, R4gpw6[38]);  // ../RTL/cortexm0ds_logic.v(12455)
  not u14378 (Kklow6, n3967);  // ../RTL/cortexm0ds_logic.v(12455)
  and u14379 (Uilow6, Yklow6, Qgeow6);  // ../RTL/cortexm0ds_logic.v(12456)
  buf u1438 (vis_pc_o[27], D12qw6);  // ../RTL/cortexm0ds_logic.v(2011)
  and u14380 (Yklow6, Fllow6, Mllow6);  // ../RTL/cortexm0ds_logic.v(12457)
  and u14381 (n3968, Q0fiu6, R4gpw6[54]);  // ../RTL/cortexm0ds_logic.v(12458)
  not u14382 (Mllow6, n3968);  // ../RTL/cortexm0ds_logic.v(12458)
  and u14383 (n3969, Pceow6, Tllow6);  // ../RTL/cortexm0ds_logic.v(12459)
  not u14384 (Fllow6, n3969);  // ../RTL/cortexm0ds_logic.v(12459)
  or u14385 (Tllow6, Nzhiu6, Vbgpw6[30]);  // ../RTL/cortexm0ds_logic.v(12460)
  and u14386 (Felow6, Amlow6, Hmlow6);  // ../RTL/cortexm0ds_logic.v(12461)
  and u14387 (n3970, C2eow6, Omlow6);  // ../RTL/cortexm0ds_logic.v(12462)
  not u14388 (Hmlow6, n3970);  // ../RTL/cortexm0ds_logic.v(12462)
  and u14389 (n3971, Vmlow6, A94ju6);  // ../RTL/cortexm0ds_logic.v(12463)
  buf u1439 (vis_psp_o[26], Rtibx6);  // ../RTL/cortexm0ds_logic.v(2085)
  not u14390 (Omlow6, n3971);  // ../RTL/cortexm0ds_logic.v(12463)
  and u14391 (n3972, Cnlow6, Jnlow6);  // ../RTL/cortexm0ds_logic.v(12464)
  not u14392 (A94ju6, n3972);  // ../RTL/cortexm0ds_logic.v(12464)
  and u14393 (n3973, Qnlow6, Queow6);  // ../RTL/cortexm0ds_logic.v(12465)
  not u14394 (Jnlow6, n3973);  // ../RTL/cortexm0ds_logic.v(12465)
  and u14395 (Qnlow6, Xnlow6, Zveow6);  // ../RTL/cortexm0ds_logic.v(12466)
  or u14396 (Xnlow6, Azfow6, Kqfow6);  // ../RTL/cortexm0ds_logic.v(12467)
  AL_MUX u14397 (
    .i0(Zx3ju6),
    .i1(Eolow6),
    .sel(J2eow6),
    .o(Cnlow6));  // ../RTL/cortexm0ds_logic.v(12468)
  and u14398 (n3974, Lolow6, Vh3ju6);  // ../RTL/cortexm0ds_logic.v(12469)
  not u14399 (Vmlow6, n3974);  // ../RTL/cortexm0ds_logic.v(12469)
  buf u144 (Jshpw6[9], Yf1qw6);  // ../RTL/cortexm0ds_logic.v(2372)
  buf u1440 (vis_pc_o[28], Lqjpw6);  // ../RTL/cortexm0ds_logic.v(2011)
  and u14400 (Lolow6, Queow6, Zveow6);  // ../RTL/cortexm0ds_logic.v(12470)
  or u14401 (Zveow6, Solow6, C3kow6);  // ../RTL/cortexm0ds_logic.v(12471)
  and u14402 (n3975, HRDATA[30], Q2eow6);  // ../RTL/cortexm0ds_logic.v(12472)
  not u14403 (Amlow6, n3975);  // ../RTL/cortexm0ds_logic.v(12472)
  and u14404 (n3976, Xbcow6, N6cow6);  // ../RTL/cortexm0ds_logic.v(12473)
  not u14405 (Kdlow6, n3976);  // ../RTL/cortexm0ds_logic.v(12473)
  and u14406 (n3977, Zolow6, Gplow6);  // ../RTL/cortexm0ds_logic.v(12474)
  not u14407 (N6cow6, n3977);  // ../RTL/cortexm0ds_logic.v(12474)
  and u14408 (Gplow6, Nplow6, Uplow6);  // ../RTL/cortexm0ds_logic.v(12475)
  and u14409 (n3978, Dyeow6, Og4ju6);  // ../RTL/cortexm0ds_logic.v(12476)
  buf u1441 (vis_psp_o[27], Zezpw6);  // ../RTL/cortexm0ds_logic.v(2085)
  not u14410 (Uplow6, n3978);  // ../RTL/cortexm0ds_logic.v(12476)
  or u14411 (Nplow6, Iydow6, Kkriu6);  // ../RTL/cortexm0ds_logic.v(12477)
  and u14412 (Kkriu6, Bqlow6, Iqlow6);  // ../RTL/cortexm0ds_logic.v(12478)
  and u14413 (Iqlow6, Pqlow6, Wqlow6);  // ../RTL/cortexm0ds_logic.v(12479)
  and u14414 (Wqlow6, Drlow6, Krlow6);  // ../RTL/cortexm0ds_logic.v(12480)
  and u14415 (Krlow6, Rrlow6, Yrlow6);  // ../RTL/cortexm0ds_logic.v(12481)
  and u14416 (n3979, Odgpw6[6], M0eow6);  // ../RTL/cortexm0ds_logic.v(12482)
  not u14417 (Yrlow6, n3979);  // ../RTL/cortexm0ds_logic.v(12482)
  and u14418 (n3980, Q0fiu6, R4gpw6[48]);  // ../RTL/cortexm0ds_logic.v(12483)
  not u14419 (Rrlow6, n3980);  // ../RTL/cortexm0ds_logic.v(12483)
  buf u1442 (vis_pc_o[29], A32qw6);  // ../RTL/cortexm0ds_logic.v(2011)
  and u14420 (Drlow6, Fslow6, Mslow6);  // ../RTL/cortexm0ds_logic.v(12484)
  and u14421 (n3981, Bagpw6[6], M6eiu6);  // ../RTL/cortexm0ds_logic.v(12485)
  not u14422 (Mslow6, n3981);  // ../RTL/cortexm0ds_logic.v(12485)
  and u14423 (n3982, C0fiu6, R4gpw6[56]);  // ../RTL/cortexm0ds_logic.v(12486)
  not u14424 (Fslow6, n3982);  // ../RTL/cortexm0ds_logic.v(12486)
  and u14425 (Pqlow6, Tslow6, Atlow6);  // ../RTL/cortexm0ds_logic.v(12487)
  and u14426 (n3983, E1fiu6, R4gpw6[40]);  // ../RTL/cortexm0ds_logic.v(12488)
  not u14427 (Atlow6, n3983);  // ../RTL/cortexm0ds_logic.v(12488)
  and u14428 (Tslow6, Htlow6, Otlow6);  // ../RTL/cortexm0ds_logic.v(12489)
  and u14429 (n3984, Tzfpw6[6], Yvgiu6);  // ../RTL/cortexm0ds_logic.v(12490)
  buf u1443 (vis_psp_o[28], Exypw6);  // ../RTL/cortexm0ds_logic.v(2085)
  not u14430 (Otlow6, n3984);  // ../RTL/cortexm0ds_logic.v(12490)
  and u14431 (n3985, STCALIB[6], H1eow6);  // ../RTL/cortexm0ds_logic.v(12491)
  not u14432 (Htlow6, n3985);  // ../RTL/cortexm0ds_logic.v(12491)
  and u14433 (Bqlow6, Vtlow6, Culow6);  // ../RTL/cortexm0ds_logic.v(12492)
  and u14434 (Culow6, Julow6, Qulow6);  // ../RTL/cortexm0ds_logic.v(12493)
  and u14435 (n3986, F0eow6, Vbgpw6[6]);  // ../RTL/cortexm0ds_logic.v(12494)
  not u14436 (Qulow6, n3986);  // ../RTL/cortexm0ds_logic.v(12494)
  and u14437 (Julow6, Xulow6, Evlow6);  // ../RTL/cortexm0ds_logic.v(12495)
  and u14438 (n3987, S1fiu6, R4gpw6[32]);  // ../RTL/cortexm0ds_logic.v(12496)
  not u14439 (Evlow6, n3987);  // ../RTL/cortexm0ds_logic.v(12496)
  buf u1444 (vis_pc_o[30], Awupw6);  // ../RTL/cortexm0ds_logic.v(2011)
  and u14440 (n3988, G2fiu6, R4gpw6[24]);  // ../RTL/cortexm0ds_logic.v(12497)
  not u14441 (Xulow6, n3988);  // ../RTL/cortexm0ds_logic.v(12497)
  and u14442 (Vtlow6, Lvlow6, Svlow6);  // ../RTL/cortexm0ds_logic.v(12498)
  and u14443 (n3989, U2fiu6, R4gpw6[16]);  // ../RTL/cortexm0ds_logic.v(12499)
  not u14444 (Svlow6, n3989);  // ../RTL/cortexm0ds_logic.v(12499)
  and u14445 (Lvlow6, Zvlow6, Gwlow6);  // ../RTL/cortexm0ds_logic.v(12500)
  and u14446 (n3990, I3fiu6, R4gpw6[8]);  // ../RTL/cortexm0ds_logic.v(12501)
  not u14447 (Gwlow6, n3990);  // ../RTL/cortexm0ds_logic.v(12501)
  and u14448 (n3991, Tzdiu6, R4gpw6[0]);  // ../RTL/cortexm0ds_logic.v(12502)
  not u14449 (Zvlow6, n3991);  // ../RTL/cortexm0ds_logic.v(12502)
  buf u1445 (vis_pc_o[18], Cchax6);  // ../RTL/cortexm0ds_logic.v(2011)
  and u14450 (Zolow6, Nwlow6, Uwlow6);  // ../RTL/cortexm0ds_logic.v(12503)
  or u14451 (Uwlow6, Uafow6, Yt3ju6);  // ../RTL/cortexm0ds_logic.v(12504)
  and u14452 (n3992, HRDATA[6], Q2eow6);  // ../RTL/cortexm0ds_logic.v(12506)
  not u14453 (Nwlow6, n3992);  // ../RTL/cortexm0ds_logic.v(12506)
  or u14454 (Mkziu6, K3how6, Df3ju6);  // ../RTL/cortexm0ds_logic.v(12507)
  not u14455 (Xbcow6, Mkziu6);  // ../RTL/cortexm0ds_logic.v(12507)
  and u14456 (n3993, Egziu6, Eafpw6[22]);  // ../RTL/cortexm0ds_logic.v(12508)
  not u14457 (Eikow6, n3993);  // ../RTL/cortexm0ds_logic.v(12508)
  and u14458 (Chkow6, Lccow6, Bxlow6);  // ../RTL/cortexm0ds_logic.v(12509)
  and u14459 (n3994, vis_pc_o[21], Jmziu6);  // ../RTL/cortexm0ds_logic.v(12510)
  buf u1446 (Iahpw6[8], Qj1qw6);  // ../RTL/cortexm0ds_logic.v(1883)
  not u14460 (Bxlow6, n3994);  // ../RTL/cortexm0ds_logic.v(12510)
  and u14461 (Lccow6, Sgziu6, Ixlow6);  // ../RTL/cortexm0ds_logic.v(12511)
  or u14462 (Ixlow6, Svkiu6, Ft6ow6);  // ../RTL/cortexm0ds_logic.v(12512)
  and u14463 (n3995, Pxlow6, Ytcow6);  // ../RTL/cortexm0ds_logic.v(12514)
  not u14464 (Svkiu6, n3995);  // ../RTL/cortexm0ds_logic.v(12514)
  and u14465 (Ytcow6, Wxlow6, H5how6);  // ../RTL/cortexm0ds_logic.v(12515)
  AL_MUX u14466 (
    .i0(Dylow6),
    .i1(Oh3ju6),
    .sel(Tucow6),
    .o(Wxlow6));  // ../RTL/cortexm0ds_logic.v(12516)
  and u14467 (Oh3ju6, Kylow6, Kf3ju6);  // ../RTL/cortexm0ds_logic.v(12517)
  or u14468 (Kylow6, L7how6, Df3ju6);  // ../RTL/cortexm0ds_logic.v(12518)
  and u14469 (n3996, Rylow6, Yylow6);  // ../RTL/cortexm0ds_logic.v(12519)
  buf u1447 (vis_psp_o[29], Evypw6);  // ../RTL/cortexm0ds_logic.v(2085)
  not u14470 (Dylow6, n3996);  // ../RTL/cortexm0ds_logic.v(12519)
  and u14471 (n3997, Fzlow6, C0ehu6);  // ../RTL/cortexm0ds_logic.v(12520)
  not u14472 (Yylow6, n3997);  // ../RTL/cortexm0ds_logic.v(12520)
  and u14473 (Fzlow6, Pthiu6, Cyfpw6[5]);  // ../RTL/cortexm0ds_logic.v(12521)
  and u14474 (Rylow6, C6how6, Mzlow6);  // ../RTL/cortexm0ds_logic.v(12522)
  and u14475 (Pxlow6, Ydlow6, Tzlow6);  // ../RTL/cortexm0ds_logic.v(12523)
  or u14476 (Ydlow6, Avcow6, Ktcow6);  // ../RTL/cortexm0ds_logic.v(12524)
  and u14477 (n3998, A0mow6, H0mow6);  // ../RTL/cortexm0ds_logic.v(12525)
  not u14478 (Hcohu6, n3998);  // ../RTL/cortexm0ds_logic.v(12525)
  and u14479 (H0mow6, O0mow6, V0mow6);  // ../RTL/cortexm0ds_logic.v(12526)
  buf u1448 (S8fpw6[1], R9mpw6);  // ../RTL/cortexm0ds_logic.v(2451)
  and u14480 (n3999, Egziu6, Eafpw6[10]);  // ../RTL/cortexm0ds_logic.v(12527)
  not u14481 (V0mow6, n3999);  // ../RTL/cortexm0ds_logic.v(12527)
  and u14482 (Egziu6, Ar8iu6, Et8iu6);  // ../RTL/cortexm0ds_logic.v(12528)
  and u14483 (O0mow6, C1mow6, Sgziu6);  // ../RTL/cortexm0ds_logic.v(12529)
  and u14484 (n4000, Ar8iu6, J1mow6);  // ../RTL/cortexm0ds_logic.v(12530)
  not u14485 (Sgziu6, n4000);  // ../RTL/cortexm0ds_logic.v(12530)
  and u14486 (n4001, Q1mow6, X1mow6);  // ../RTL/cortexm0ds_logic.v(12531)
  not u14487 (J1mow6, n4001);  // ../RTL/cortexm0ds_logic.v(12531)
  and u14488 (n4002, Jydhu6, Zmfiu6);  // ../RTL/cortexm0ds_logic.v(12532)
  not u14489 (X1mow6, n4002);  // ../RTL/cortexm0ds_logic.v(12532)
  buf u1449 (vis_pc_o[1], Nyhax6);  // ../RTL/cortexm0ds_logic.v(2011)
  and u14490 (Q1mow6, E2mow6, Dp8iu6);  // ../RTL/cortexm0ds_logic.v(12534)
  and u14491 (n4003, Qwdhu6, M2biu6);  // ../RTL/cortexm0ds_logic.v(12535)
  not u14492 (E2mow6, n4003);  // ../RTL/cortexm0ds_logic.v(12535)
  and u14493 (n4004, Zgziu6, Oymiu6);  // ../RTL/cortexm0ds_logic.v(12537)
  not u14494 (C1mow6, n4004);  // ../RTL/cortexm0ds_logic.v(12537)
  and u14495 (n4005, L2mow6, S2mow6);  // ../RTL/cortexm0ds_logic.v(12538)
  not u14496 (Oymiu6, n4005);  // ../RTL/cortexm0ds_logic.v(12538)
  and u14497 (S2mow6, Z2mow6, G3mow6);  // ../RTL/cortexm0ds_logic.v(12539)
  or u14498 (G3mow6, Plcow6, Pkdow6);  // ../RTL/cortexm0ds_logic.v(12540)
  and u14499 (Pkdow6, Eccow6, N3mow6);  // ../RTL/cortexm0ds_logic.v(12541)
  buf u145 (K7hpw6[19], Ab9ax6);  // ../RTL/cortexm0ds_logic.v(2366)
  buf u1450 (S8fpw6[2], Rskax6);  // ../RTL/cortexm0ds_logic.v(2451)
  and u14500 (n4006, Ktcow6, U3mow6);  // ../RTL/cortexm0ds_logic.v(12542)
  not u14501 (N3mow6, n4006);  // ../RTL/cortexm0ds_logic.v(12542)
  and u14502 (n4007, B4mow6, I4mow6);  // ../RTL/cortexm0ds_logic.v(12543)
  not u14503 (U3mow6, n4007);  // ../RTL/cortexm0ds_logic.v(12543)
  and u14504 (n4008, P4mow6, Yahow6);  // ../RTL/cortexm0ds_logic.v(12544)
  not u14505 (I4mow6, n4008);  // ../RTL/cortexm0ds_logic.v(12544)
  or u14506 (P4mow6, E6oiu6, W4mow6);  // ../RTL/cortexm0ds_logic.v(12545)
  and u14507 (W4mow6, F9aju6, Nlaiu6);  // ../RTL/cortexm0ds_logic.v(12546)
  and u14508 (E6oiu6, Cyfpw6[3], Tr0iu6);  // ../RTL/cortexm0ds_logic.v(12547)
  or u14509 (n4009, Jdhow6, K2aiu6);  // ../RTL/cortexm0ds_logic.v(12548)
  buf u1451 (vis_pc_o[2], Rwhax6);  // ../RTL/cortexm0ds_logic.v(2011)
  not u14510 (B4mow6, n4009);  // ../RTL/cortexm0ds_logic.v(12548)
  and u14511 (Jdhow6, T23ju6, Cyfpw6[3]);  // ../RTL/cortexm0ds_logic.v(12549)
  or u14512 (n4010, Tfjiu6, Tr0iu6);  // ../RTL/cortexm0ds_logic.v(12550)
  not u14513 (T23ju6, n4010);  // ../RTL/cortexm0ds_logic.v(12550)
  and u14514 (Eccow6, Tzlow6, D5mow6);  // ../RTL/cortexm0ds_logic.v(12551)
  not u14515 (D5mow6, Ovcow6);  // ../RTL/cortexm0ds_logic.v(12552)
  and u14516 (Ovcow6, Ktcow6, K5mow6);  // ../RTL/cortexm0ds_logic.v(12553)
  and u14517 (n4011, C0ehu6, R5mow6);  // ../RTL/cortexm0ds_logic.v(12554)
  not u14518 (K5mow6, n4011);  // ../RTL/cortexm0ds_logic.v(12554)
  and u14519 (n4012, G7oiu6, Y5mow6);  // ../RTL/cortexm0ds_logic.v(12555)
  buf u1452 (S8fpw6[3], U1kpw6);  // ../RTL/cortexm0ds_logic.v(2451)
  not u14520 (R5mow6, n4012);  // ../RTL/cortexm0ds_logic.v(12555)
  or u14521 (Y5mow6, Y2oiu6, Tr0iu6);  // ../RTL/cortexm0ds_logic.v(12556)
  and u14522 (Plcow6, F6mow6, M6mow6);  // ../RTL/cortexm0ds_logic.v(12557)
  and u14523 (M6mow6, T6mow6, A7mow6);  // ../RTL/cortexm0ds_logic.v(12558)
  or u14524 (A7mow6, Rcfow6, Id4ju6);  // ../RTL/cortexm0ds_logic.v(12559)
  and u14525 (Id4ju6, H7mow6, O7mow6);  // ../RTL/cortexm0ds_logic.v(12560)
  and u14526 (O7mow6, V7mow6, C8mow6);  // ../RTL/cortexm0ds_logic.v(12561)
  or u14527 (C8mow6, Ipfow6, Z90iu6);  // ../RTL/cortexm0ds_logic.v(12562)
  or u14528 (V7mow6, Kqfow6, Na0iu6);  // ../RTL/cortexm0ds_logic.v(12563)
  and u14529 (H7mow6, J8mow6, Q8mow6);  // ../RTL/cortexm0ds_logic.v(12564)
  buf u1453 (vis_pc_o[3], Vuhax6);  // ../RTL/cortexm0ds_logic.v(2011)
  or u14530 (Q8mow6, Rqfow6, Ga0iu6);  // ../RTL/cortexm0ds_logic.v(12565)
  or u14531 (J8mow6, Ppfow6, Ua0iu6);  // ../RTL/cortexm0ds_logic.v(12566)
  or u14532 (T6mow6, Iydow6, Bisiu6);  // ../RTL/cortexm0ds_logic.v(12567)
  and u14533 (Bisiu6, X8mow6, E9mow6);  // ../RTL/cortexm0ds_logic.v(12568)
  and u14534 (E9mow6, L9mow6, S9mow6);  // ../RTL/cortexm0ds_logic.v(12569)
  and u14535 (n4013, Tzfpw6[10], Yvgiu6);  // ../RTL/cortexm0ds_logic.v(12570)
  not u14536 (S9mow6, n4013);  // ../RTL/cortexm0ds_logic.v(12570)
  and u14537 (L9mow6, Z9mow6, Gamow6);  // ../RTL/cortexm0ds_logic.v(12571)
  and u14538 (n4014, F0eow6, Vbgpw6[10]);  // ../RTL/cortexm0ds_logic.v(12572)
  not u14539 (Gamow6, n4014);  // ../RTL/cortexm0ds_logic.v(12572)
  buf u1454 (S8fpw6[4], Ubypw6);  // ../RTL/cortexm0ds_logic.v(2451)
  and u14540 (n4015, Odgpw6[10], M0eow6);  // ../RTL/cortexm0ds_logic.v(12573)
  not u14541 (Z9mow6, n4015);  // ../RTL/cortexm0ds_logic.v(12573)
  and u14542 (X8mow6, Namow6, Uamow6);  // ../RTL/cortexm0ds_logic.v(12574)
  and u14543 (n4016, Bagpw6[10], M6eiu6);  // ../RTL/cortexm0ds_logic.v(12575)
  not u14544 (Uamow6, n4016);  // ../RTL/cortexm0ds_logic.v(12575)
  and u14545 (n4017, STCALIB[10], H1eow6);  // ../RTL/cortexm0ds_logic.v(12576)
  not u14546 (Namow6, n4017);  // ../RTL/cortexm0ds_logic.v(12576)
  and u14547 (F6mow6, Bbmow6, Ibmow6);  // ../RTL/cortexm0ds_logic.v(12577)
  and u14548 (n4018, Qtfow6, Og4ju6);  // ../RTL/cortexm0ds_logic.v(12578)
  not u14549 (Ibmow6, n4018);  // ../RTL/cortexm0ds_logic.v(12578)
  buf u1455 (vis_pc_o[4], Zshax6);  // ../RTL/cortexm0ds_logic.v(2011)
  and u14550 (n4019, Pbmow6, Wbmow6);  // ../RTL/cortexm0ds_logic.v(12579)
  not u14551 (Og4ju6, n4019);  // ../RTL/cortexm0ds_logic.v(12579)
  and u14552 (Wbmow6, Dcmow6, Kcmow6);  // ../RTL/cortexm0ds_logic.v(12580)
  or u14553 (Kcmow6, Kqfow6, Pb0iu6);  // ../RTL/cortexm0ds_logic.v(12581)
  or u14554 (Dcmow6, Ppfow6, Wb0iu6);  // ../RTL/cortexm0ds_logic.v(12582)
  and u14555 (Pbmow6, Rcmow6, Ycmow6);  // ../RTL/cortexm0ds_logic.v(12583)
  or u14556 (Ycmow6, Ipfow6, Bb0iu6);  // ../RTL/cortexm0ds_logic.v(12584)
  or u14557 (Rcmow6, Rqfow6, Ib0iu6);  // ../RTL/cortexm0ds_logic.v(12585)
  and u14558 (n4020, HRDATA[10], Q2eow6);  // ../RTL/cortexm0ds_logic.v(12586)
  not u14559 (Bbmow6, n4020);  // ../RTL/cortexm0ds_logic.v(12586)
  buf u1456 (S8fpw6[5], Fkrpw6);  // ../RTL/cortexm0ds_logic.v(2451)
  and u14560 (Z2mow6, Fdmow6, Dldow6);  // ../RTL/cortexm0ds_logic.v(12587)
  and u14561 (n4021, H5how6, Mdmow6);  // ../RTL/cortexm0ds_logic.v(12588)
  not u14562 (Dldow6, n4021);  // ../RTL/cortexm0ds_logic.v(12588)
  and u14563 (n4022, Tdmow6, C6how6);  // ../RTL/cortexm0ds_logic.v(12589)
  not u14564 (Mdmow6, n4022);  // ../RTL/cortexm0ds_logic.v(12589)
  and u14565 (n4023, Aemow6, V3xhu6);  // ../RTL/cortexm0ds_logic.v(12590)
  not u14566 (C6how6, n4023);  // ../RTL/cortexm0ds_logic.v(12590)
  and u14567 (Aemow6, Hemow6, Ktcow6);  // ../RTL/cortexm0ds_logic.v(12591)
  and u14568 (n4024, Oemow6, Vemow6);  // ../RTL/cortexm0ds_logic.v(12592)
  not u14569 (Tdmow6, n4024);  // ../RTL/cortexm0ds_logic.v(12592)
  buf u1457 (vis_pc_o[5], Drhax6);  // ../RTL/cortexm0ds_logic.v(2011)
  and u14570 (Vemow6, Cfmow6, Dahow6);  // ../RTL/cortexm0ds_logic.v(12593)
  and u14571 (Cfmow6, Tzlow6, K3how6);  // ../RTL/cortexm0ds_logic.v(12594)
  or u14572 (Tzlow6, Ny3ju6, Ktcow6);  // ../RTL/cortexm0ds_logic.v(12595)
  or u14573 (Ny3ju6, Fg3ju6, R3how6);  // ../RTL/cortexm0ds_logic.v(12596)
  and u14574 (n4025, Jfmow6, Ej3ju6);  // ../RTL/cortexm0ds_logic.v(12597)
  not u14575 (Fg3ju6, n4025);  // ../RTL/cortexm0ds_logic.v(12597)
  and u14576 (Oemow6, Qfmow6, O1low6);  // ../RTL/cortexm0ds_logic.v(12598)
  and u14577 (n4026, Xfmow6, Ktcow6);  // ../RTL/cortexm0ds_logic.v(12599)
  not u14578 (Qfmow6, n4026);  // ../RTL/cortexm0ds_logic.v(12599)
  and u14579 (Xfmow6, Egmow6, Lgmow6);  // ../RTL/cortexm0ds_logic.v(12600)
  buf u1458 (S8fpw6[6], Umkax6);  // ../RTL/cortexm0ds_logic.v(2451)
  and u14580 (n4027, Sgmow6, C0ehu6);  // ../RTL/cortexm0ds_logic.v(12601)
  not u14581 (Lgmow6, n4027);  // ../RTL/cortexm0ds_logic.v(12601)
  or u14582 (n4028, Mjfiu6, Cyfpw6[0]);  // ../RTL/cortexm0ds_logic.v(12602)
  not u14583 (Sgmow6, n4028);  // ../RTL/cortexm0ds_logic.v(12602)
  or u14584 (Egmow6, Rn2ju6, Tfjiu6);  // ../RTL/cortexm0ds_logic.v(12603)
  and u14585 (n4029, Zgmow6, Ghmow6);  // ../RTL/cortexm0ds_logic.v(12604)
  not u14586 (H5how6, n4029);  // ../RTL/cortexm0ds_logic.v(12604)
  and u14587 (Ghmow6, Nhmow6, Uhmow6);  // ../RTL/cortexm0ds_logic.v(12605)
  or u14588 (Uhmow6, Bimow6, Q88ow6);  // ../RTL/cortexm0ds_logic.v(12606)
  and u14589 (Q88ow6, Iimow6, Pimow6);  // ../RTL/cortexm0ds_logic.v(12607)
  buf u1459 (vis_pc_o[6], Equpw6);  // ../RTL/cortexm0ds_logic.v(2011)
  or u14590 (Pimow6, Iydow6, Ggtiu6);  // ../RTL/cortexm0ds_logic.v(12608)
  and u14591 (Ggtiu6, Wimow6, Djmow6);  // ../RTL/cortexm0ds_logic.v(12609)
  and u14592 (Djmow6, Kjmow6, Rjmow6);  // ../RTL/cortexm0ds_logic.v(12610)
  and u14593 (Rjmow6, Yjmow6, Fkmow6);  // ../RTL/cortexm0ds_logic.v(12611)
  and u14594 (Fkmow6, Mkmow6, Tkmow6);  // ../RTL/cortexm0ds_logic.v(12612)
  and u14595 (n4030, E1fiu6, R4gpw6[43]);  // ../RTL/cortexm0ds_logic.v(12613)
  not u14596 (Tkmow6, n4030);  // ../RTL/cortexm0ds_logic.v(12613)
  and u14597 (n4031, Q0fiu6, R4gpw6[51]);  // ../RTL/cortexm0ds_logic.v(12614)
  not u14598 (Mkmow6, n4031);  // ../RTL/cortexm0ds_logic.v(12614)
  and u14599 (Yjmow6, Almow6, Hlmow6);  // ../RTL/cortexm0ds_logic.v(12615)
  buf u146 (vis_r2_o[30], A1qax6);  // ../RTL/cortexm0ds_logic.v(2551)
  buf u1460 (S8fpw6[7], V6jax6);  // ../RTL/cortexm0ds_logic.v(2451)
  and u14600 (n4032, Tzdiu6, R4gpw6[3]);  // ../RTL/cortexm0ds_logic.v(12616)
  not u14601 (Hlmow6, n4032);  // ../RTL/cortexm0ds_logic.v(12616)
  and u14602 (n4033, STCALIB[15], H1eow6);  // ../RTL/cortexm0ds_logic.v(12617)
  not u14603 (Almow6, n4033);  // ../RTL/cortexm0ds_logic.v(12617)
  and u14604 (Kjmow6, Olmow6, Vlmow6);  // ../RTL/cortexm0ds_logic.v(12618)
  and u14605 (Vlmow6, Cmmow6, Jmmow6);  // ../RTL/cortexm0ds_logic.v(12619)
  or u14606 (Jmmow6, P6ciu6, Qkgiu6);  // ../RTL/cortexm0ds_logic.v(12620)
  and u14607 (n4034, Ydeow6, Qmmow6);  // ../RTL/cortexm0ds_logic.v(12621)
  not u14608 (P6ciu6, n4034);  // ../RTL/cortexm0ds_logic.v(12621)
  and u14609 (n4035, Xmmow6, J1fow6);  // ../RTL/cortexm0ds_logic.v(12622)
  buf u1461 (vis_pc_o[7], Hphax6);  // ../RTL/cortexm0ds_logic.v(2011)
  not u14610 (Qmmow6, n4035);  // ../RTL/cortexm0ds_logic.v(12622)
  and u14611 (J1fow6, O8low6, A8low6);  // ../RTL/cortexm0ds_logic.v(12624)
  not u14612 (Feeow6, J1fow6);  // ../RTL/cortexm0ds_logic.v(12624)
  AL_MUX u14613 (
    .i0(B4fow6),
    .i1(H7fow6),
    .sel(Meeow6),
    .o(Xmmow6));  // ../RTL/cortexm0ds_logic.v(12625)
  and u14614 (Ydeow6, A0fow6, V0fow6);  // ../RTL/cortexm0ds_logic.v(12626)
  or u14615 (n4036, Righu6, Ahghu6);  // ../RTL/cortexm0ds_logic.v(12627)
  not u14616 (A0fow6, n4036);  // ../RTL/cortexm0ds_logic.v(12627)
  and u14617 (n4037, I3fiu6, R4gpw6[11]);  // ../RTL/cortexm0ds_logic.v(12628)
  not u14618 (Cmmow6, n4037);  // ../RTL/cortexm0ds_logic.v(12628)
  and u14619 (Olmow6, Enmow6, Lnmow6);  // ../RTL/cortexm0ds_logic.v(12629)
  buf u1462 (S8fpw6[8], Iekax6);  // ../RTL/cortexm0ds_logic.v(2451)
  and u14620 (n4038, G2fiu6, R4gpw6[27]);  // ../RTL/cortexm0ds_logic.v(12630)
  not u14621 (Lnmow6, n4038);  // ../RTL/cortexm0ds_logic.v(12630)
  and u14622 (n4039, U2fiu6, R4gpw6[19]);  // ../RTL/cortexm0ds_logic.v(12631)
  not u14623 (Enmow6, n4039);  // ../RTL/cortexm0ds_logic.v(12631)
  and u14624 (Wimow6, Snmow6, Znmow6);  // ../RTL/cortexm0ds_logic.v(12632)
  and u14625 (Znmow6, Gomow6, Nomow6);  // ../RTL/cortexm0ds_logic.v(12633)
  and u14626 (Nomow6, Uomow6, Bpmow6);  // ../RTL/cortexm0ds_logic.v(12634)
  and u14627 (n4040, Odgpw6[15], M0eow6);  // ../RTL/cortexm0ds_logic.v(12635)
  not u14628 (Bpmow6, n4040);  // ../RTL/cortexm0ds_logic.v(12635)
  and u14629 (n4041, Tzfpw6[15], Yvgiu6);  // ../RTL/cortexm0ds_logic.v(12636)
  buf u1463 (vis_pc_o[8], J06bx6);  // ../RTL/cortexm0ds_logic.v(2011)
  not u14630 (Uomow6, n4041);  // ../RTL/cortexm0ds_logic.v(12636)
  and u14631 (Gomow6, Ipmow6, Ppmow6);  // ../RTL/cortexm0ds_logic.v(12637)
  and u14632 (n4042, F0eow6, Vbgpw6[15]);  // ../RTL/cortexm0ds_logic.v(12638)
  not u14633 (Ppmow6, n4042);  // ../RTL/cortexm0ds_logic.v(12638)
  and u14634 (n4043, Bagpw6[15], M6eiu6);  // ../RTL/cortexm0ds_logic.v(12639)
  not u14635 (Ipmow6, n4043);  // ../RTL/cortexm0ds_logic.v(12639)
  and u14636 (Snmow6, Wpmow6, Dqmow6);  // ../RTL/cortexm0ds_logic.v(12640)
  and u14637 (Dqmow6, Kqmow6, Rqmow6);  // ../RTL/cortexm0ds_logic.v(12641)
  and u14638 (n4044, C0fiu6, R4gpw6[59]);  // ../RTL/cortexm0ds_logic.v(12642)
  not u14639 (Rqmow6, n4044);  // ../RTL/cortexm0ds_logic.v(12642)
  buf u1464 (S8fpw6[9], Lgkax6);  // ../RTL/cortexm0ds_logic.v(2451)
  and u14640 (n4045, Zlghu6, Xrgiu6);  // ../RTL/cortexm0ds_logic.v(12643)
  not u14641 (Kqmow6, n4045);  // ../RTL/cortexm0ds_logic.v(12643)
  and u14642 (Xrgiu6, Yqmow6, Ynhiu6);  // ../RTL/cortexm0ds_logic.v(12644)
  and u14643 (Yqmow6, K5eiu6, Jfgpw6[4]);  // ../RTL/cortexm0ds_logic.v(12645)
  and u14644 (Wpmow6, Qgeow6, Frmow6);  // ../RTL/cortexm0ds_logic.v(12646)
  and u14645 (n4046, S1fiu6, R4gpw6[35]);  // ../RTL/cortexm0ds_logic.v(12647)
  not u14646 (Frmow6, n4046);  // ../RTL/cortexm0ds_logic.v(12647)
  and u14647 (Iimow6, Mrmow6, Trmow6);  // ../RTL/cortexm0ds_logic.v(12648)
  or u14648 (Trmow6, We3ju6, Hfeow6);  // ../RTL/cortexm0ds_logic.v(12649)
  not u14649 (We3ju6, Y83ju6);  // ../RTL/cortexm0ds_logic.v(12650)
  buf u1465 (vis_pc_o[9], P7bbx6);  // ../RTL/cortexm0ds_logic.v(2011)
  AL_MUX u14650 (
    .i0(Re4ju6),
    .i1(L44ju6),
    .sel(Hv3ju6),
    .o(Y83ju6));  // ../RTL/cortexm0ds_logic.v(12651)
  and u14651 (n4047, Asmow6, Hsmow6);  // ../RTL/cortexm0ds_logic.v(12652)
  not u14652 (L44ju6, n4047);  // ../RTL/cortexm0ds_logic.v(12652)
  and u14653 (Hsmow6, Osmow6, Vsmow6);  // ../RTL/cortexm0ds_logic.v(12653)
  or u14654 (Vsmow6, Ipfow6, J80iu6);  // ../RTL/cortexm0ds_logic.v(12654)
  or u14655 (Osmow6, Rqfow6, Q80iu6);  // ../RTL/cortexm0ds_logic.v(12655)
  and u14656 (Asmow6, Ctmow6, Jtmow6);  // ../RTL/cortexm0ds_logic.v(12656)
  or u14657 (Jtmow6, Ppfow6, L90iu6);  // ../RTL/cortexm0ds_logic.v(12657)
  or u14658 (Ctmow6, Kqfow6, X80iu6);  // ../RTL/cortexm0ds_logic.v(12658)
  and u14659 (n4048, Qtmow6, Xtmow6);  // ../RTL/cortexm0ds_logic.v(12659)
  buf u1466 (S8fpw6[10], Oikax6);  // ../RTL/cortexm0ds_logic.v(2451)
  not u14660 (Re4ju6, n4048);  // ../RTL/cortexm0ds_logic.v(12659)
  and u14661 (Xtmow6, Eumow6, Lumow6);  // ../RTL/cortexm0ds_logic.v(12660)
  or u14662 (Lumow6, Ipfow6, S90iu6);  // ../RTL/cortexm0ds_logic.v(12661)
  or u14663 (Eumow6, Rqfow6, Z90iu6);  // ../RTL/cortexm0ds_logic.v(12662)
  and u14664 (Qtmow6, Sumow6, Zumow6);  // ../RTL/cortexm0ds_logic.v(12663)
  or u14665 (Zumow6, Ppfow6, Na0iu6);  // ../RTL/cortexm0ds_logic.v(12664)
  or u14666 (Sumow6, Kqfow6, Ga0iu6);  // ../RTL/cortexm0ds_logic.v(12665)
  and u14667 (n4049, Q2eow6, HRDATA[15]);  // ../RTL/cortexm0ds_logic.v(12666)
  not u14668 (Mrmow6, n4049);  // ../RTL/cortexm0ds_logic.v(12666)
  and u14669 (Bimow6, Gvmow6, Nvmow6);  // ../RTL/cortexm0ds_logic.v(12667)
  buf u1467 (vis_pc_o[19], Fahax6);  // ../RTL/cortexm0ds_logic.v(2011)
  and u14670 (n4050, S2ziu6, Cyfpw6[3]);  // ../RTL/cortexm0ds_logic.v(12668)
  not u14671 (Nvmow6, n4050);  // ../RTL/cortexm0ds_logic.v(12668)
  or u14672 (n4051, Tfjiu6, Hs0iu6);  // ../RTL/cortexm0ds_logic.v(12669)
  not u14673 (S2ziu6, n4051);  // ../RTL/cortexm0ds_logic.v(12669)
  and u14674 (n4052, Uvmow6, Yahow6);  // ../RTL/cortexm0ds_logic.v(12670)
  not u14675 (Gvmow6, n4052);  // ../RTL/cortexm0ds_logic.v(12670)
  and u14676 (Nhmow6, Bwmow6, Bz3ju6);  // ../RTL/cortexm0ds_logic.v(12671)
  and u14677 (n4053, Iwmow6, X88ow6);  // ../RTL/cortexm0ds_logic.v(12672)
  not u14678 (Bwmow6, n4053);  // ../RTL/cortexm0ds_logic.v(12672)
  and u14679 (n4054, Pwmow6, Wwmow6);  // ../RTL/cortexm0ds_logic.v(12673)
  buf u1468 (Iahpw6[9], L0ypw6);  // ../RTL/cortexm0ds_logic.v(1883)
  not u14680 (X88ow6, n4054);  // ../RTL/cortexm0ds_logic.v(12673)
  or u14681 (Wwmow6, Iydow6, Pxriu6);  // ../RTL/cortexm0ds_logic.v(12674)
  and u14682 (Pxriu6, Dxmow6, Kxmow6);  // ../RTL/cortexm0ds_logic.v(12675)
  and u14683 (Kxmow6, Rxmow6, Yxmow6);  // ../RTL/cortexm0ds_logic.v(12676)
  and u14684 (Yxmow6, Fymow6, Mymow6);  // ../RTL/cortexm0ds_logic.v(12677)
  and u14685 (Mymow6, Tymow6, Azmow6);  // ../RTL/cortexm0ds_logic.v(12678)
  and u14686 (n4055, Odgpw6[7], M0eow6);  // ../RTL/cortexm0ds_logic.v(12679)
  not u14687 (Azmow6, n4055);  // ../RTL/cortexm0ds_logic.v(12679)
  and u14688 (n4056, Q0fiu6, R4gpw6[49]);  // ../RTL/cortexm0ds_logic.v(12680)
  not u14689 (Tymow6, n4056);  // ../RTL/cortexm0ds_logic.v(12680)
  and u1469 (Xuzhu6, Kc0iu6, Rc0iu6);  // ../RTL/cortexm0ds_logic.v(3442)
  and u14690 (Fymow6, Hzmow6, Ozmow6);  // ../RTL/cortexm0ds_logic.v(12681)
  and u14691 (n4057, Bagpw6[7], M6eiu6);  // ../RTL/cortexm0ds_logic.v(12682)
  not u14692 (Ozmow6, n4057);  // ../RTL/cortexm0ds_logic.v(12682)
  and u14693 (n4058, C0fiu6, R4gpw6[57]);  // ../RTL/cortexm0ds_logic.v(12683)
  not u14694 (Hzmow6, n4058);  // ../RTL/cortexm0ds_logic.v(12683)
  and u14695 (Rxmow6, Vzmow6, C0now6);  // ../RTL/cortexm0ds_logic.v(12684)
  and u14696 (n4059, E1fiu6, R4gpw6[41]);  // ../RTL/cortexm0ds_logic.v(12685)
  not u14697 (C0now6, n4059);  // ../RTL/cortexm0ds_logic.v(12685)
  and u14698 (Vzmow6, J0now6, Q0now6);  // ../RTL/cortexm0ds_logic.v(12686)
  and u14699 (n4060, Tzfpw6[7], Yvgiu6);  // ../RTL/cortexm0ds_logic.v(12687)
  buf u147 (vis_r1_o[2], Untpw6);  // ../RTL/cortexm0ds_logic.v(1876)
  and u1470 (n113, Yc0iu6, Fd0iu6);  // ../RTL/cortexm0ds_logic.v(3443)
  not u14700 (Q0now6, n4060);  // ../RTL/cortexm0ds_logic.v(12687)
  and u14701 (n4061, STCALIB[7], H1eow6);  // ../RTL/cortexm0ds_logic.v(12688)
  not u14702 (J0now6, n4061);  // ../RTL/cortexm0ds_logic.v(12688)
  and u14703 (Dxmow6, X0now6, E1now6);  // ../RTL/cortexm0ds_logic.v(12689)
  and u14704 (E1now6, L1now6, S1now6);  // ../RTL/cortexm0ds_logic.v(12690)
  and u14705 (n4062, F0eow6, Vbgpw6[7]);  // ../RTL/cortexm0ds_logic.v(12691)
  not u14706 (S1now6, n4062);  // ../RTL/cortexm0ds_logic.v(12691)
  and u14707 (L1now6, Z1now6, G2now6);  // ../RTL/cortexm0ds_logic.v(12692)
  and u14708 (n4063, S1fiu6, R4gpw6[33]);  // ../RTL/cortexm0ds_logic.v(12693)
  not u14709 (G2now6, n4063);  // ../RTL/cortexm0ds_logic.v(12693)
  not u1471 (Rc0iu6, n113);  // ../RTL/cortexm0ds_logic.v(3443)
  and u14710 (n4064, G2fiu6, R4gpw6[25]);  // ../RTL/cortexm0ds_logic.v(12694)
  not u14711 (Z1now6, n4064);  // ../RTL/cortexm0ds_logic.v(12694)
  and u14712 (X0now6, N2now6, U2now6);  // ../RTL/cortexm0ds_logic.v(12695)
  and u14713 (n4065, U2fiu6, R4gpw6[17]);  // ../RTL/cortexm0ds_logic.v(12696)
  not u14714 (U2now6, n4065);  // ../RTL/cortexm0ds_logic.v(12696)
  and u14715 (N2now6, B3now6, I3now6);  // ../RTL/cortexm0ds_logic.v(12697)
  and u14716 (n4066, I3fiu6, R4gpw6[9]);  // ../RTL/cortexm0ds_logic.v(12698)
  not u14717 (I3now6, n4066);  // ../RTL/cortexm0ds_logic.v(12698)
  and u14718 (n4067, Tzdiu6, R4gpw6[1]);  // ../RTL/cortexm0ds_logic.v(12699)
  not u14719 (B3now6, n4067);  // ../RTL/cortexm0ds_logic.v(12699)
  and u1472 (Yc0iu6, C0ehu6, Md0iu6);  // ../RTL/cortexm0ds_logic.v(3444)
  and u14720 (Pwmow6, P3now6, W3now6);  // ../RTL/cortexm0ds_logic.v(12700)
  and u14721 (n4068, C2eow6, Jb3ju6);  // ../RTL/cortexm0ds_logic.v(12701)
  not u14722 (W3now6, n4068);  // ../RTL/cortexm0ds_logic.v(12701)
  AL_MUX u14723 (
    .i0(Jw3ju6),
    .i1(Ag4ju6),
    .sel(Hv3ju6),
    .o(Jb3ju6));  // ../RTL/cortexm0ds_logic.v(12702)
  and u14724 (n4069, D4now6, K4now6);  // ../RTL/cortexm0ds_logic.v(12703)
  not u14725 (Ag4ju6, n4069);  // ../RTL/cortexm0ds_logic.v(12703)
  and u14726 (K4now6, R4now6, Y4now6);  // ../RTL/cortexm0ds_logic.v(12704)
  or u14727 (Y4now6, Ppfow6, Pb0iu6);  // ../RTL/cortexm0ds_logic.v(12705)
  and u14728 (Pb0iu6, F5now6, M5now6);  // ../RTL/cortexm0ds_logic.v(12706)
  and u14729 (M5now6, T5now6, A6now6);  // ../RTL/cortexm0ds_logic.v(12707)
  or u1473 (Kc0iu6, Td0iu6, Ae0iu6);  // ../RTL/cortexm0ds_logic.v(3445)
  and u14730 (A6now6, H6now6, O6now6);  // ../RTL/cortexm0ds_logic.v(12708)
  and u14731 (n4070, V6now6, vis_r2_o[11]);  // ../RTL/cortexm0ds_logic.v(12709)
  not u14732 (O6now6, n4070);  // ../RTL/cortexm0ds_logic.v(12709)
  and u14733 (n4071, C7now6, vis_r6_o[11]);  // ../RTL/cortexm0ds_logic.v(12710)
  not u14734 (H6now6, n4071);  // ../RTL/cortexm0ds_logic.v(12710)
  and u14735 (T5now6, J7now6, Q7now6);  // ../RTL/cortexm0ds_logic.v(12711)
  and u14736 (n4072, X7now6, vis_r5_o[11]);  // ../RTL/cortexm0ds_logic.v(12712)
  not u14737 (Q7now6, n4072);  // ../RTL/cortexm0ds_logic.v(12712)
  and u14738 (n4073, E8now6, vis_r4_o[11]);  // ../RTL/cortexm0ds_logic.v(12713)
  not u14739 (J7now6, n4073);  // ../RTL/cortexm0ds_logic.v(12713)
  buf u1474 (Bagpw6[4], Imhbx6);  // ../RTL/cortexm0ds_logic.v(2680)
  and u14740 (F5now6, L8now6, S8now6);  // ../RTL/cortexm0ds_logic.v(12714)
  and u14741 (S8now6, Z8now6, G9now6);  // ../RTL/cortexm0ds_logic.v(12715)
  and u14742 (n4074, N9now6, vis_r1_o[11]);  // ../RTL/cortexm0ds_logic.v(12716)
  not u14743 (G9now6, n4074);  // ../RTL/cortexm0ds_logic.v(12716)
  and u14744 (n4075, U9now6, vis_r0_o[11]);  // ../RTL/cortexm0ds_logic.v(12717)
  not u14745 (Z8now6, n4075);  // ../RTL/cortexm0ds_logic.v(12717)
  and u14746 (L8now6, Banow6, Ianow6);  // ../RTL/cortexm0ds_logic.v(12718)
  and u14747 (n4076, Panow6, vis_r3_o[11]);  // ../RTL/cortexm0ds_logic.v(12719)
  not u14748 (Ianow6, n4076);  // ../RTL/cortexm0ds_logic.v(12719)
  and u14749 (n4077, Wanow6, vis_r7_o[11]);  // ../RTL/cortexm0ds_logic.v(12720)
  buf u1475 (vis_r10_o[17], Wfmax6);  // ../RTL/cortexm0ds_logic.v(2469)
  not u14750 (Banow6, n4077);  // ../RTL/cortexm0ds_logic.v(12720)
  or u14751 (R4now6, Ipfow6, Ua0iu6);  // ../RTL/cortexm0ds_logic.v(12721)
  and u14752 (D4now6, Dbnow6, Kbnow6);  // ../RTL/cortexm0ds_logic.v(12722)
  or u14753 (Kbnow6, Rqfow6, Bb0iu6);  // ../RTL/cortexm0ds_logic.v(12723)
  or u14754 (Dbnow6, Kqfow6, Ib0iu6);  // ../RTL/cortexm0ds_logic.v(12724)
  and u14755 (n4078, Rbnow6, Ybnow6);  // ../RTL/cortexm0ds_logic.v(12725)
  not u14756 (Jw3ju6, n4078);  // ../RTL/cortexm0ds_logic.v(12725)
  and u14757 (Ybnow6, Fcnow6, Mcnow6);  // ../RTL/cortexm0ds_logic.v(12726)
  or u14758 (Mcnow6, Ppfow6, I40iu6);  // ../RTL/cortexm0ds_logic.v(12727)
  or u14759 (Fcnow6, Kqfow6, B40iu6);  // ../RTL/cortexm0ds_logic.v(12728)
  and u1476 (Vnfpw6[7], Ppfpw6[13], Ivfhu6);  // ../RTL/cortexm0ds_logic.v(3367)
  and u14760 (Rbnow6, Tcnow6, Adnow6);  // ../RTL/cortexm0ds_logic.v(12729)
  or u14761 (Adnow6, Ipfow6, Wb0iu6);  // ../RTL/cortexm0ds_logic.v(12730)
  and u14762 (Wb0iu6, Hdnow6, Odnow6);  // ../RTL/cortexm0ds_logic.v(12731)
  and u14763 (Odnow6, Vdnow6, Cenow6);  // ../RTL/cortexm0ds_logic.v(12732)
  and u14764 (Cenow6, Jenow6, Qenow6);  // ../RTL/cortexm0ds_logic.v(12733)
  and u14765 (n4079, V6now6, vis_r2_o[10]);  // ../RTL/cortexm0ds_logic.v(12734)
  not u14766 (Qenow6, n4079);  // ../RTL/cortexm0ds_logic.v(12734)
  and u14767 (n4080, C7now6, vis_r6_o[10]);  // ../RTL/cortexm0ds_logic.v(12735)
  not u14768 (Jenow6, n4080);  // ../RTL/cortexm0ds_logic.v(12735)
  and u14769 (Vdnow6, Xenow6, Efnow6);  // ../RTL/cortexm0ds_logic.v(12736)
  buf u1477 (vis_r10_o[18], Wdmax6);  // ../RTL/cortexm0ds_logic.v(2469)
  and u14770 (n4081, X7now6, vis_r5_o[10]);  // ../RTL/cortexm0ds_logic.v(12737)
  not u14771 (Efnow6, n4081);  // ../RTL/cortexm0ds_logic.v(12737)
  and u14772 (n4082, E8now6, vis_r4_o[10]);  // ../RTL/cortexm0ds_logic.v(12738)
  not u14773 (Xenow6, n4082);  // ../RTL/cortexm0ds_logic.v(12738)
  and u14774 (Hdnow6, Lfnow6, Sfnow6);  // ../RTL/cortexm0ds_logic.v(12739)
  and u14775 (Sfnow6, Zfnow6, Ggnow6);  // ../RTL/cortexm0ds_logic.v(12740)
  and u14776 (n4083, N9now6, vis_r1_o[10]);  // ../RTL/cortexm0ds_logic.v(12741)
  not u14777 (Ggnow6, n4083);  // ../RTL/cortexm0ds_logic.v(12741)
  and u14778 (n4084, U9now6, vis_r0_o[10]);  // ../RTL/cortexm0ds_logic.v(12742)
  not u14779 (Zfnow6, n4084);  // ../RTL/cortexm0ds_logic.v(12742)
  buf u1478 (vis_ipsr_o[1], Pcrpw6);  // ../RTL/cortexm0ds_logic.v(1815)
  and u14780 (Lfnow6, Ngnow6, Ugnow6);  // ../RTL/cortexm0ds_logic.v(12743)
  and u14781 (n4085, Panow6, vis_r3_o[10]);  // ../RTL/cortexm0ds_logic.v(12744)
  not u14782 (Ugnow6, n4085);  // ../RTL/cortexm0ds_logic.v(12744)
  and u14783 (n4086, Wanow6, vis_r7_o[10]);  // ../RTL/cortexm0ds_logic.v(12745)
  not u14784 (Ngnow6, n4086);  // ../RTL/cortexm0ds_logic.v(12745)
  or u14785 (Tcnow6, Rqfow6, U30iu6);  // ../RTL/cortexm0ds_logic.v(12746)
  and u14786 (n4087, HRDATA[7], Q2eow6);  // ../RTL/cortexm0ds_logic.v(12747)
  not u14787 (P3now6, n4087);  // ../RTL/cortexm0ds_logic.v(12747)
  and u14788 (n4088, Rn2ju6, Bhnow6);  // ../RTL/cortexm0ds_logic.v(12748)
  not u14789 (Iwmow6, n4088);  // ../RTL/cortexm0ds_logic.v(12748)
  buf u1479 (Bagpw6[5], X5opw6);  // ../RTL/cortexm0ds_logic.v(2680)
  and u14790 (n4089, Ihnow6, Tfjiu6);  // ../RTL/cortexm0ds_logic.v(12749)
  not u14791 (Bhnow6, n4089);  // ../RTL/cortexm0ds_logic.v(12749)
  and u14792 (n4090, Tr0iu6, Phnow6);  // ../RTL/cortexm0ds_logic.v(12750)
  not u14793 (Ihnow6, n4090);  // ../RTL/cortexm0ds_logic.v(12750)
  buf u14794 (Qifhu6, Ozkbx6[5]);  // ../RTL/cortexm0ds_logic.v(3176)
  not u14795 (Rn2ju6, A3aju6);  // ../RTL/cortexm0ds_logic.v(12752)
  and u14796 (Zgmow6, Whnow6, Dinow6);  // ../RTL/cortexm0ds_logic.v(12753)
  and u14797 (n4091, Iwfpw6[1], Kinow6);  // ../RTL/cortexm0ds_logic.v(12754)
  not u14798 (Dinow6, n4091);  // ../RTL/cortexm0ds_logic.v(12754)
  and u14799 (n4092, Rinow6, Yinow6);  // ../RTL/cortexm0ds_logic.v(12755)
  buf u148 (Uthpw6[4], V53qw6);  // ../RTL/cortexm0ds_logic.v(1882)
  buf u1480 (vis_r10_o[19], Wbmax6);  // ../RTL/cortexm0ds_logic.v(2469)
  not u14800 (Kinow6, n4092);  // ../RTL/cortexm0ds_logic.v(12755)
  and u14801 (n4093, Fjnow6, Qyniu6);  // ../RTL/cortexm0ds_logic.v(12756)
  not u14802 (Yinow6, n4093);  // ../RTL/cortexm0ds_logic.v(12756)
  or u14803 (n4094, H78ow6, Iwfpw6[0]);  // ../RTL/cortexm0ds_logic.v(12757)
  not u14804 (Fjnow6, n4094);  // ../RTL/cortexm0ds_logic.v(12757)
  and u14805 (H78ow6, Mjnow6, Tjnow6);  // ../RTL/cortexm0ds_logic.v(12758)
  or u14806 (Tjnow6, Iydow6, N0viu6);  // ../RTL/cortexm0ds_logic.v(12759)
  and u14807 (N0viu6, Aknow6, Hknow6);  // ../RTL/cortexm0ds_logic.v(12760)
  and u14808 (Hknow6, Oknow6, Vknow6);  // ../RTL/cortexm0ds_logic.v(12761)
  and u14809 (Vknow6, Clnow6, Jlnow6);  // ../RTL/cortexm0ds_logic.v(12762)
  buf u1481 (vis_ipsr_o[2], Aniax6);  // ../RTL/cortexm0ds_logic.v(1815)
  and u14810 (Jlnow6, Qlnow6, Xlnow6);  // ../RTL/cortexm0ds_logic.v(12763)
  and u14811 (n4095, Odgpw6[23], M0eow6);  // ../RTL/cortexm0ds_logic.v(12764)
  not u14812 (Xlnow6, n4095);  // ../RTL/cortexm0ds_logic.v(12764)
  and u14813 (n4096, Q0fiu6, R4gpw6[53]);  // ../RTL/cortexm0ds_logic.v(12765)
  not u14814 (Qlnow6, n4096);  // ../RTL/cortexm0ds_logic.v(12765)
  and u14815 (Clnow6, Emnow6, Lmnow6);  // ../RTL/cortexm0ds_logic.v(12766)
  and u14816 (n4097, Tzdiu6, R4gpw6[5]);  // ../RTL/cortexm0ds_logic.v(12767)
  not u14817 (Lmnow6, n4097);  // ../RTL/cortexm0ds_logic.v(12767)
  and u14818 (n4098, I3fiu6, R4gpw6[13]);  // ../RTL/cortexm0ds_logic.v(12768)
  not u14819 (Emnow6, n4098);  // ../RTL/cortexm0ds_logic.v(12768)
  buf u1482 (vis_r10_o[20], W9max6);  // ../RTL/cortexm0ds_logic.v(2469)
  and u14820 (Oknow6, Smnow6, Zmnow6);  // ../RTL/cortexm0ds_logic.v(12769)
  and u14821 (Zmnow6, Gnnow6, Nnnow6);  // ../RTL/cortexm0ds_logic.v(12770)
  and u14822 (n4099, Hqgiu6, L1gpw6[1]);  // ../RTL/cortexm0ds_logic.v(12771)
  not u14823 (Nnnow6, n4099);  // ../RTL/cortexm0ds_logic.v(12771)
  and u14824 (n4100, STCALIB[23], H1eow6);  // ../RTL/cortexm0ds_logic.v(12772)
  not u14825 (Gnnow6, n4100);  // ../RTL/cortexm0ds_logic.v(12772)
  and u14826 (Smnow6, Unnow6, Bonow6);  // ../RTL/cortexm0ds_logic.v(12773)
  and u14827 (n4101, G2fiu6, R4gpw6[29]);  // ../RTL/cortexm0ds_logic.v(12774)
  not u14828 (Bonow6, n4101);  // ../RTL/cortexm0ds_logic.v(12774)
  and u14829 (n4102, U2fiu6, R4gpw6[21]);  // ../RTL/cortexm0ds_logic.v(12775)
  buf u1483 (vis_ipsr_o[3], Qhmpw6);  // ../RTL/cortexm0ds_logic.v(1815)
  not u14830 (Unnow6, n4102);  // ../RTL/cortexm0ds_logic.v(12775)
  and u14831 (Aknow6, Ionow6, Ponow6);  // ../RTL/cortexm0ds_logic.v(12776)
  and u14832 (Ponow6, Wonow6, Dpnow6);  // ../RTL/cortexm0ds_logic.v(12777)
  and u14833 (Dpnow6, Kpnow6, Rpnow6);  // ../RTL/cortexm0ds_logic.v(12778)
  and u14834 (n4103, Tzfpw6[23], Yvgiu6);  // ../RTL/cortexm0ds_logic.v(12779)
  not u14835 (Rpnow6, n4103);  // ../RTL/cortexm0ds_logic.v(12779)
  or u14836 (Kpnow6, Qkgiu6, U6piu6);  // ../RTL/cortexm0ds_logic.v(12780)
  and u14837 (Wonow6, Ypnow6, Fqnow6);  // ../RTL/cortexm0ds_logic.v(12781)
  and u14838 (n4104, Bagpw6[23], M6eiu6);  // ../RTL/cortexm0ds_logic.v(12782)
  not u14839 (Fqnow6, n4104);  // ../RTL/cortexm0ds_logic.v(12782)
  buf u1484 (vis_r10_o[21], W7max6);  // ../RTL/cortexm0ds_logic.v(2469)
  and u14840 (n4105, E1fiu6, R4gpw6[45]);  // ../RTL/cortexm0ds_logic.v(12783)
  not u14841 (Ypnow6, n4105);  // ../RTL/cortexm0ds_logic.v(12783)
  and u14842 (Ionow6, Mqnow6, Tqnow6);  // ../RTL/cortexm0ds_logic.v(12784)
  and u14843 (n4106, S1fiu6, R4gpw6[37]);  // ../RTL/cortexm0ds_logic.v(12785)
  not u14844 (Tqnow6, n4106);  // ../RTL/cortexm0ds_logic.v(12785)
  and u14845 (Mqnow6, Arnow6, Hrnow6);  // ../RTL/cortexm0ds_logic.v(12786)
  and u14846 (n4107, C0fiu6, R4gpw6[61]);  // ../RTL/cortexm0ds_logic.v(12787)
  not u14847 (Hrnow6, n4107);  // ../RTL/cortexm0ds_logic.v(12787)
  and u14848 (n4108, F0eow6, Vbgpw6[23]);  // ../RTL/cortexm0ds_logic.v(12788)
  not u14849 (Arnow6, n4108);  // ../RTL/cortexm0ds_logic.v(12788)
  buf u1485 (vis_ipsr_o[4], Ijiax6);  // ../RTL/cortexm0ds_logic.v(1815)
  and u14850 (Mjnow6, Ornow6, Vrnow6);  // ../RTL/cortexm0ds_logic.v(12789)
  or u14851 (Vrnow6, Hfeow6, Ha3ju6);  // ../RTL/cortexm0ds_logic.v(12790)
  AL_MUX u14852 (
    .i0(C34ju6),
    .i1(Csnow6),
    .sel(Hv3ju6),
    .o(Ha3ju6));  // ../RTL/cortexm0ds_logic.v(12791)
  and u14853 (Csnow6, Ecjow6, Lcjow6);  // ../RTL/cortexm0ds_logic.v(12792)
  and u14854 (Lcjow6, Jsnow6, Qsnow6);  // ../RTL/cortexm0ds_logic.v(12793)
  or u14855 (Qsnow6, Ipfow6, Y50iu6);  // ../RTL/cortexm0ds_logic.v(12794)
  or u14856 (Jsnow6, Rqfow6, M60iu6);  // ../RTL/cortexm0ds_logic.v(12795)
  and u14857 (Ecjow6, Xsnow6, Etnow6);  // ../RTL/cortexm0ds_logic.v(12796)
  or u14858 (Etnow6, Ppfow6, A70iu6);  // ../RTL/cortexm0ds_logic.v(12797)
  and u14859 (n4109, C3kow6, Ltnow6);  // ../RTL/cortexm0ds_logic.v(12798)
  or u1486 (n112[0], Xuzhu6, Dc0iu6);  // ../RTL/cortexm0ds_logic.v(3417)
  not u14860 (Xsnow6, n4109);  // ../RTL/cortexm0ds_logic.v(12798)
  and u14861 (C34ju6, Stnow6, Ztnow6);  // ../RTL/cortexm0ds_logic.v(12799)
  and u14862 (Ztnow6, Gunow6, Nunow6);  // ../RTL/cortexm0ds_logic.v(12800)
  or u14863 (Nunow6, Ipfow6, H70iu6);  // ../RTL/cortexm0ds_logic.v(12801)
  or u14864 (Gunow6, Rqfow6, O70iu6);  // ../RTL/cortexm0ds_logic.v(12802)
  and u14865 (Stnow6, Uunow6, Bvnow6);  // ../RTL/cortexm0ds_logic.v(12803)
  or u14866 (Bvnow6, Ppfow6, C80iu6);  // ../RTL/cortexm0ds_logic.v(12804)
  or u14867 (Uunow6, Kqfow6, V70iu6);  // ../RTL/cortexm0ds_logic.v(12805)
  and u14868 (n4110, HRDATA[23], Q2eow6);  // ../RTL/cortexm0ds_logic.v(12806)
  not u14869 (Ornow6, n4110);  // ../RTL/cortexm0ds_logic.v(12806)
  not u1487 (Tgfpw6[0], n111[0]);  // ../RTL/cortexm0ds_logic.v(3385)
  and u14870 (n4111, Uvmow6, V78ow6);  // ../RTL/cortexm0ds_logic.v(12807)
  not u14871 (Rinow6, n4111);  // ../RTL/cortexm0ds_logic.v(12807)
  and u14872 (n4112, Ivnow6, Pvnow6);  // ../RTL/cortexm0ds_logic.v(12808)
  not u14873 (V78ow6, n4112);  // ../RTL/cortexm0ds_logic.v(12808)
  or u14874 (Pvnow6, Iydow6, Rw1iu6);  // ../RTL/cortexm0ds_logic.v(12809)
  and u14875 (Rw1iu6, Wvnow6, Dwnow6);  // ../RTL/cortexm0ds_logic.v(12810)
  and u14876 (Dwnow6, Kwnow6, Rwnow6);  // ../RTL/cortexm0ds_logic.v(12811)
  and u14877 (Rwnow6, Ywnow6, Fxnow6);  // ../RTL/cortexm0ds_logic.v(12812)
  and u14878 (Fxnow6, Mxnow6, Txnow6);  // ../RTL/cortexm0ds_logic.v(12813)
  or u14879 (Txnow6, Te6iu6, Qkgiu6);  // ../RTL/cortexm0ds_logic.v(12814)
  buf u1488 (Bagpw6[6], Ox9bx6);  // ../RTL/cortexm0ds_logic.v(2680)
  and u14880 (n4113, Hqgiu6, H8gpw6[1]);  // ../RTL/cortexm0ds_logic.v(12815)
  not u14881 (Mxnow6, n4113);  // ../RTL/cortexm0ds_logic.v(12815)
  and u14882 (Hqgiu6, Aynow6, Ynhiu6);  // ../RTL/cortexm0ds_logic.v(12816)
  and u14883 (Aynow6, K5eiu6, U89iu6);  // ../RTL/cortexm0ds_logic.v(12817)
  and u14884 (Ywnow6, Hynow6, Oynow6);  // ../RTL/cortexm0ds_logic.v(12818)
  and u14885 (n4114, STCALIB[25], H1eow6);  // ../RTL/cortexm0ds_logic.v(12819)
  not u14886 (Oynow6, n4114);  // ../RTL/cortexm0ds_logic.v(12819)
  and u14887 (n4115, C0fiu6, R4gpw6[63]);  // ../RTL/cortexm0ds_logic.v(12820)
  not u14888 (Hynow6, n4115);  // ../RTL/cortexm0ds_logic.v(12820)
  and u14889 (C0fiu6, Vynow6, Cznow6);  // ../RTL/cortexm0ds_logic.v(12821)
  and u1489 (Zg0iu6, Nh0iu6, Oe0iu6);  // ../RTL/cortexm0ds_logic.v(3455)
  and u14890 (Kwnow6, Jznow6, Qznow6);  // ../RTL/cortexm0ds_logic.v(12822)
  and u14891 (n4116, S1fiu6, R4gpw6[39]);  // ../RTL/cortexm0ds_logic.v(12823)
  not u14892 (Qznow6, n4116);  // ../RTL/cortexm0ds_logic.v(12823)
  and u14893 (S1fiu6, Xznow6, Vynow6);  // ../RTL/cortexm0ds_logic.v(12824)
  and u14894 (Jznow6, E0oow6, L0oow6);  // ../RTL/cortexm0ds_logic.v(12825)
  and u14895 (n4117, Tzdiu6, R4gpw6[7]);  // ../RTL/cortexm0ds_logic.v(12826)
  not u14896 (L0oow6, n4117);  // ../RTL/cortexm0ds_logic.v(12826)
  and u14897 (Tzdiu6, Xznow6, Pjyiu6);  // ../RTL/cortexm0ds_logic.v(12827)
  and u14898 (n4118, Q0fiu6, R4gpw6[55]);  // ../RTL/cortexm0ds_logic.v(12828)
  not u14899 (E0oow6, n4118);  // ../RTL/cortexm0ds_logic.v(12828)
  buf u149 (Jshpw6[28], Vqgax6);  // ../RTL/cortexm0ds_logic.v(2372)
  and u1490 (n115, Uh0iu6, H6ghu6);  // ../RTL/cortexm0ds_logic.v(3456)
  and u14900 (Q0fiu6, S0oow6, Vynow6);  // ../RTL/cortexm0ds_logic.v(12829)
  and u14901 (Wvnow6, Z0oow6, G1oow6);  // ../RTL/cortexm0ds_logic.v(12830)
  and u14902 (G1oow6, N1oow6, U1oow6);  // ../RTL/cortexm0ds_logic.v(12831)
  and u14903 (U1oow6, B2oow6, I2oow6);  // ../RTL/cortexm0ds_logic.v(12832)
  and u14904 (n4119, Pceow6, P2oow6);  // ../RTL/cortexm0ds_logic.v(12833)
  not u14905 (I2oow6, n4119);  // ../RTL/cortexm0ds_logic.v(12833)
  or u14906 (P2oow6, Nzhiu6, Vbgpw6[31]);  // ../RTL/cortexm0ds_logic.v(12834)
  and u14907 (n4120, G2fiu6, R4gpw6[31]);  // ../RTL/cortexm0ds_logic.v(12835)
  not u14908 (B2oow6, n4120);  // ../RTL/cortexm0ds_logic.v(12835)
  and u14909 (G2fiu6, Pjyiu6, Cznow6);  // ../RTL/cortexm0ds_logic.v(12836)
  not u1491 (Nh0iu6, n115);  // ../RTL/cortexm0ds_logic.v(3456)
  and u14910 (N1oow6, W2oow6, D3oow6);  // ../RTL/cortexm0ds_logic.v(12837)
  and u14911 (n4121, U2fiu6, R4gpw6[23]);  // ../RTL/cortexm0ds_logic.v(12838)
  not u14912 (D3oow6, n4121);  // ../RTL/cortexm0ds_logic.v(12838)
  and u14913 (U2fiu6, S0oow6, Pjyiu6);  // ../RTL/cortexm0ds_logic.v(12839)
  and u14914 (S0oow6, K3oow6, Jfgpw6[3]);  // ../RTL/cortexm0ds_logic.v(12840)
  or u14915 (n4122, Jfgpw6[2], Jfgpw6[4]);  // ../RTL/cortexm0ds_logic.v(12841)
  not u14916 (K3oow6, n4122);  // ../RTL/cortexm0ds_logic.v(12841)
  and u14917 (n4123, E1fiu6, R4gpw6[47]);  // ../RTL/cortexm0ds_logic.v(12842)
  not u14918 (W2oow6, n4123);  // ../RTL/cortexm0ds_logic.v(12842)
  and u14919 (E1fiu6, Vynow6, Dtjow6);  // ../RTL/cortexm0ds_logic.v(12843)
  and u1492 (Uh0iu6, Bi0iu6, Ii0iu6);  // ../RTL/cortexm0ds_logic.v(3457)
  and u14920 (Z0oow6, R3oow6, Y3oow6);  // ../RTL/cortexm0ds_logic.v(12844)
  or u14921 (Y3oow6, Tpgiu6, F4oow6);  // ../RTL/cortexm0ds_logic.v(12845)
  and u14922 (n4124, Rzciu6, Cznow6);  // ../RTL/cortexm0ds_logic.v(12846)
  not u14923 (Tpgiu6, n4124);  // ../RTL/cortexm0ds_logic.v(12846)
  and u14924 (R3oow6, M4oow6, T4oow6);  // ../RTL/cortexm0ds_logic.v(12847)
  and u14925 (n4125, I3fiu6, R4gpw6[15]);  // ../RTL/cortexm0ds_logic.v(12848)
  not u14926 (T4oow6, n4125);  // ../RTL/cortexm0ds_logic.v(12848)
  and u14927 (I3fiu6, Pjyiu6, Dtjow6);  // ../RTL/cortexm0ds_logic.v(12849)
  and u14928 (n4126, Odgpw6[31], M0eow6);  // ../RTL/cortexm0ds_logic.v(12850)
  not u14929 (M4oow6, n4126);  // ../RTL/cortexm0ds_logic.v(12850)
  buf u1493 (vis_r6_o[31], Kjoax6);  // ../RTL/cortexm0ds_logic.v(2523)
  and u14930 (Ivnow6, A5oow6, H5oow6);  // ../RTL/cortexm0ds_logic.v(12851)
  or u14931 (H5oow6, Hfeow6, Mg3ju6);  // ../RTL/cortexm0ds_logic.v(12852)
  not u14932 (Mg3ju6, O5oow6);  // ../RTL/cortexm0ds_logic.v(12853)
  AL_MUX u14933 (
    .i0(Qb3ju6),
    .i1(Vh3ju6),
    .sel(V5oow6),
    .o(O5oow6));  // ../RTL/cortexm0ds_logic.v(12854)
  and u14934 (V5oow6, Queow6, Solow6);  // ../RTL/cortexm0ds_logic.v(12855)
  and u14935 (n4127, V2kow6, Ppfow6);  // ../RTL/cortexm0ds_logic.v(12856)
  not u14936 (Solow6, n4127);  // ../RTL/cortexm0ds_logic.v(12856)
  and u14937 (Queow6, C6oow6, Cyfpw6[3]);  // ../RTL/cortexm0ds_logic.v(12857)
  and u14938 (C6oow6, J6oow6, Hzfow6);  // ../RTL/cortexm0ds_logic.v(12858)
  or u14939 (J6oow6, Azfow6, Ppfow6);  // ../RTL/cortexm0ds_logic.v(12859)
  buf u1494 (vis_r10_o[23], Cglax6);  // ../RTL/cortexm0ds_logic.v(2469)
  AL_MUX u14940 (
    .i0(Vajow6),
    .i1(Lx3ju6),
    .sel(Hv3ju6),
    .o(Qb3ju6));  // ../RTL/cortexm0ds_logic.v(12861)
  and u14941 (n4128, Q6oow6, X6oow6);  // ../RTL/cortexm0ds_logic.v(12862)
  not u14942 (Lx3ju6, n4128);  // ../RTL/cortexm0ds_logic.v(12862)
  and u14943 (X6oow6, E7oow6, L7oow6);  // ../RTL/cortexm0ds_logic.v(12863)
  or u14944 (L7oow6, Rqfow6, W40iu6);  // ../RTL/cortexm0ds_logic.v(12864)
  or u14945 (E7oow6, Kqfow6, D50iu6);  // ../RTL/cortexm0ds_logic.v(12865)
  and u14946 (Q6oow6, S7oow6, Z7oow6);  // ../RTL/cortexm0ds_logic.v(12866)
  or u14947 (Z7oow6, Ppfow6, K50iu6);  // ../RTL/cortexm0ds_logic.v(12867)
  or u14948 (S7oow6, Ipfow6, P40iu6);  // ../RTL/cortexm0ds_logic.v(12868)
  and u14949 (n4129, G8oow6, N8oow6);  // ../RTL/cortexm0ds_logic.v(12869)
  buf u1495 (vis_r10_o[1], X3max6);  // ../RTL/cortexm0ds_logic.v(2469)
  not u14950 (Vajow6, n4129);  // ../RTL/cortexm0ds_logic.v(12869)
  and u14951 (N8oow6, U8oow6, B9oow6);  // ../RTL/cortexm0ds_logic.v(12870)
  or u14952 (B9oow6, Ipfow6, F60iu6);  // ../RTL/cortexm0ds_logic.v(12871)
  or u14953 (U8oow6, Rqfow6, E90iu6);  // ../RTL/cortexm0ds_logic.v(12872)
  and u14954 (G8oow6, I9oow6, P9oow6);  // ../RTL/cortexm0ds_logic.v(12873)
  or u14955 (P9oow6, Ppfow6, R50iu6);  // ../RTL/cortexm0ds_logic.v(12874)
  or u14956 (I9oow6, Kqfow6, Dc0iu6);  // ../RTL/cortexm0ds_logic.v(12875)
  and u14957 (n4130, Q2eow6, HRDATA[31]);  // ../RTL/cortexm0ds_logic.v(12876)
  not u14958 (A5oow6, n4130);  // ../RTL/cortexm0ds_logic.v(12876)
  and u14959 (n4131, W9oow6, Daoow6);  // ../RTL/cortexm0ds_logic.v(12877)
  buf u1496 (vis_r10_o[24], Xvlax6);  // ../RTL/cortexm0ds_logic.v(2469)
  not u14960 (Uvmow6, n4131);  // ../RTL/cortexm0ds_logic.v(12877)
  or u14961 (Daoow6, X5oiu6, Cyfpw6[0]);  // ../RTL/cortexm0ds_logic.v(12878)
  and u14962 (n4132, Iwfpw6[0], Qyniu6);  // ../RTL/cortexm0ds_logic.v(12879)
  not u14963 (W9oow6, n4132);  // ../RTL/cortexm0ds_logic.v(12879)
  and u14964 (n4133, V3xhu6, Hemow6);  // ../RTL/cortexm0ds_logic.v(12880)
  not u14965 (Whnow6, n4133);  // ../RTL/cortexm0ds_logic.v(12880)
  or u14966 (Fdmow6, Gkcow6, Uqdow6);  // ../RTL/cortexm0ds_logic.v(12881)
  and u14967 (Uqdow6, Hlziu6, Rahow6);  // ../RTL/cortexm0ds_logic.v(12883)
  not u14968 (Mmdow6, Uqdow6);  // ../RTL/cortexm0ds_logic.v(12883)
  and u14969 (n4134, Kaoow6, Ktcow6);  // ../RTL/cortexm0ds_logic.v(12884)
  buf u1497 (Bagpw6[1], Wnxax6);  // ../RTL/cortexm0ds_logic.v(2680)
  not u14970 (Rahow6, n4134);  // ../RTL/cortexm0ds_logic.v(12884)
  and u14971 (Kaoow6, Fd0iu6, Pthiu6);  // ../RTL/cortexm0ds_logic.v(12885)
  and u14972 (Hlziu6, O1low6, W9how6);  // ../RTL/cortexm0ds_logic.v(12886)
  and u14973 (n4135, Ktcow6, Vxniu6);  // ../RTL/cortexm0ds_logic.v(12887)
  not u14974 (W9how6, n4135);  // ../RTL/cortexm0ds_logic.v(12887)
  or u14975 (O1low6, Kf3ju6, Ktcow6);  // ../RTL/cortexm0ds_logic.v(12888)
  or u14976 (Kf3ju6, X6how6, Df3ju6);  // ../RTL/cortexm0ds_logic.v(12889)
  and u14977 (n4136, Raoow6, Oa3ju6);  // ../RTL/cortexm0ds_logic.v(12890)
  not u14978 (X6how6, n4136);  // ../RTL/cortexm0ds_logic.v(12890)
  and u14979 (Raoow6, F93ju6, U54ju6);  // ../RTL/cortexm0ds_logic.v(12891)
  buf u1498 (Bagpw6[2], Vlxax6);  // ../RTL/cortexm0ds_logic.v(2680)
  and u14980 (Gkcow6, Yaoow6, Fboow6);  // ../RTL/cortexm0ds_logic.v(12892)
  and u14981 (Fboow6, Mboow6, Tboow6);  // ../RTL/cortexm0ds_logic.v(12893)
  or u14982 (Tboow6, Rcfow6, Yt3ju6);  // ../RTL/cortexm0ds_logic.v(12894)
  and u14983 (Yt3ju6, Acoow6, Hcoow6);  // ../RTL/cortexm0ds_logic.v(12895)
  and u14984 (Hcoow6, Ocoow6, Vcoow6);  // ../RTL/cortexm0ds_logic.v(12896)
  or u14985 (Vcoow6, Kqfow6, I40iu6);  // ../RTL/cortexm0ds_logic.v(12897)
  and u14986 (I40iu6, Cdoow6, Jdoow6);  // ../RTL/cortexm0ds_logic.v(12898)
  and u14987 (Jdoow6, Qdoow6, Xdoow6);  // ../RTL/cortexm0ds_logic.v(12899)
  and u14988 (Xdoow6, Eeoow6, Leoow6);  // ../RTL/cortexm0ds_logic.v(12900)
  and u14989 (n4137, V6now6, vis_r2_o[7]);  // ../RTL/cortexm0ds_logic.v(12901)
  buf u1499 (Bagpw6[3], Oyhbx6);  // ../RTL/cortexm0ds_logic.v(2680)
  not u14990 (Leoow6, n4137);  // ../RTL/cortexm0ds_logic.v(12901)
  and u14991 (n4138, C7now6, vis_r6_o[7]);  // ../RTL/cortexm0ds_logic.v(12902)
  not u14992 (Eeoow6, n4138);  // ../RTL/cortexm0ds_logic.v(12902)
  and u14993 (Qdoow6, Seoow6, Zeoow6);  // ../RTL/cortexm0ds_logic.v(12903)
  and u14994 (n4139, X7now6, vis_r5_o[7]);  // ../RTL/cortexm0ds_logic.v(12904)
  not u14995 (Zeoow6, n4139);  // ../RTL/cortexm0ds_logic.v(12904)
  and u14996 (n4140, E8now6, vis_r4_o[7]);  // ../RTL/cortexm0ds_logic.v(12905)
  not u14997 (Seoow6, n4140);  // ../RTL/cortexm0ds_logic.v(12905)
  and u14998 (Cdoow6, Gfoow6, Nfoow6);  // ../RTL/cortexm0ds_logic.v(12906)
  and u14999 (Nfoow6, Ufoow6, Bgoow6);  // ../RTL/cortexm0ds_logic.v(12907)
  buf u15 (Oodhu6, Kxhpw6);  // ../RTL/cortexm0ds_logic.v(1771)
  buf u150 (vis_r0_o[30], Gvmpw6);  // ../RTL/cortexm0ds_logic.v(1875)
  buf u1500 (vis_r10_o[2], Eclax6);  // ../RTL/cortexm0ds_logic.v(2469)
  and u15000 (n4141, N9now6, vis_r1_o[7]);  // ../RTL/cortexm0ds_logic.v(12908)
  not u15001 (Bgoow6, n4141);  // ../RTL/cortexm0ds_logic.v(12908)
  and u15002 (n4142, U9now6, vis_r0_o[7]);  // ../RTL/cortexm0ds_logic.v(12909)
  not u15003 (Ufoow6, n4142);  // ../RTL/cortexm0ds_logic.v(12909)
  and u15004 (Gfoow6, Igoow6, Pgoow6);  // ../RTL/cortexm0ds_logic.v(12910)
  and u15005 (n4143, Panow6, vis_r3_o[7]);  // ../RTL/cortexm0ds_logic.v(12911)
  not u15006 (Pgoow6, n4143);  // ../RTL/cortexm0ds_logic.v(12911)
  and u15007 (n4144, Wanow6, vis_r7_o[7]);  // ../RTL/cortexm0ds_logic.v(12912)
  not u15008 (Igoow6, n4144);  // ../RTL/cortexm0ds_logic.v(12912)
  or u15009 (Ocoow6, Rqfow6, B40iu6);  // ../RTL/cortexm0ds_logic.v(12913)
  buf u1501 (vis_r10_o[25], W5max6);  // ../RTL/cortexm0ds_logic.v(2469)
  and u15010 (B40iu6, Wgoow6, Dhoow6);  // ../RTL/cortexm0ds_logic.v(12914)
  and u15011 (Dhoow6, Khoow6, Rhoow6);  // ../RTL/cortexm0ds_logic.v(12915)
  and u15012 (Rhoow6, Yhoow6, Fioow6);  // ../RTL/cortexm0ds_logic.v(12916)
  and u15013 (n4145, V6now6, vis_r2_o[8]);  // ../RTL/cortexm0ds_logic.v(12917)
  not u15014 (Fioow6, n4145);  // ../RTL/cortexm0ds_logic.v(12917)
  and u15015 (n4146, C7now6, vis_r6_o[8]);  // ../RTL/cortexm0ds_logic.v(12918)
  not u15016 (Yhoow6, n4146);  // ../RTL/cortexm0ds_logic.v(12918)
  and u15017 (Khoow6, Mioow6, Tioow6);  // ../RTL/cortexm0ds_logic.v(12919)
  and u15018 (n4147, X7now6, vis_r5_o[8]);  // ../RTL/cortexm0ds_logic.v(12920)
  not u15019 (Tioow6, n4147);  // ../RTL/cortexm0ds_logic.v(12920)
  buf u1502 (vis_r10_o[3], Bolax6);  // ../RTL/cortexm0ds_logic.v(2469)
  and u15020 (n4148, E8now6, vis_r4_o[8]);  // ../RTL/cortexm0ds_logic.v(12921)
  not u15021 (Mioow6, n4148);  // ../RTL/cortexm0ds_logic.v(12921)
  and u15022 (Wgoow6, Ajoow6, Hjoow6);  // ../RTL/cortexm0ds_logic.v(12922)
  and u15023 (Hjoow6, Ojoow6, Vjoow6);  // ../RTL/cortexm0ds_logic.v(12923)
  and u15024 (n4149, N9now6, vis_r1_o[8]);  // ../RTL/cortexm0ds_logic.v(12924)
  not u15025 (Vjoow6, n4149);  // ../RTL/cortexm0ds_logic.v(12924)
  and u15026 (n4150, U9now6, vis_r0_o[8]);  // ../RTL/cortexm0ds_logic.v(12925)
  not u15027 (Ojoow6, n4150);  // ../RTL/cortexm0ds_logic.v(12925)
  and u15028 (Ajoow6, Ckoow6, Jkoow6);  // ../RTL/cortexm0ds_logic.v(12926)
  and u15029 (n4151, Panow6, vis_r3_o[8]);  // ../RTL/cortexm0ds_logic.v(12927)
  buf u1503 (vis_r10_o[26], Xxlax6);  // ../RTL/cortexm0ds_logic.v(2469)
  not u15030 (Jkoow6, n4151);  // ../RTL/cortexm0ds_logic.v(12927)
  and u15031 (n4152, Wanow6, vis_r7_o[8]);  // ../RTL/cortexm0ds_logic.v(12928)
  not u15032 (Ckoow6, n4152);  // ../RTL/cortexm0ds_logic.v(12928)
  and u15033 (Acoow6, Qkoow6, Xkoow6);  // ../RTL/cortexm0ds_logic.v(12929)
  or u15034 (Xkoow6, Ipfow6, U30iu6);  // ../RTL/cortexm0ds_logic.v(12930)
  or u15035 (Qkoow6, Ppfow6, P40iu6);  // ../RTL/cortexm0ds_logic.v(12931)
  or u15036 (Mboow6, Iydow6, Jaqiu6);  // ../RTL/cortexm0ds_logic.v(12932)
  and u15037 (Jaqiu6, Eloow6, Lloow6);  // ../RTL/cortexm0ds_logic.v(12933)
  and u15038 (Lloow6, Sloow6, Zloow6);  // ../RTL/cortexm0ds_logic.v(12934)
  and u15039 (Zloow6, Gmoow6, Nmoow6);  // ../RTL/cortexm0ds_logic.v(12935)
  buf u1504 (vis_r10_o[4], Delax6);  // ../RTL/cortexm0ds_logic.v(2469)
  and u15040 (n4153, Odgpw6[2], M0eow6);  // ../RTL/cortexm0ds_logic.v(12936)
  not u15041 (Nmoow6, n4153);  // ../RTL/cortexm0ds_logic.v(12936)
  and u15042 (Gmoow6, Umoow6, Bnoow6);  // ../RTL/cortexm0ds_logic.v(12937)
  and u15043 (n4154, Ndghu6, Fpgiu6);  // ../RTL/cortexm0ds_logic.v(12938)
  not u15044 (Bnoow6, n4154);  // ../RTL/cortexm0ds_logic.v(12938)
  and u15045 (Fpgiu6, Rzciu6, Xznow6);  // ../RTL/cortexm0ds_logic.v(12939)
  and u15046 (n4155, STCALIB[2], H1eow6);  // ../RTL/cortexm0ds_logic.v(12940)
  not u15047 (Umoow6, n4155);  // ../RTL/cortexm0ds_logic.v(12940)
  and u15048 (Sloow6, Inoow6, Pnoow6);  // ../RTL/cortexm0ds_logic.v(12941)
  and u15049 (n4156, ECOREVNUM[2], I5eow6);  // ../RTL/cortexm0ds_logic.v(12942)
  buf u1505 (vis_r10_o[27], Xzlax6);  // ../RTL/cortexm0ds_logic.v(2469)
  not u15050 (Pnoow6, n4156);  // ../RTL/cortexm0ds_logic.v(12942)
  and u15051 (n4157, Y5eiu6, Wnoow6);  // ../RTL/cortexm0ds_logic.v(12943)
  not u15052 (Inoow6, n4157);  // ../RTL/cortexm0ds_logic.v(12943)
  or u15053 (Wnoow6, STCALIB[25], Ftghu6);  // ../RTL/cortexm0ds_logic.v(12944)
  and u15054 (Y5eiu6, Vynow6, Wjyiu6);  // ../RTL/cortexm0ds_logic.v(12945)
  and u15055 (Eloow6, Dooow6, Kooow6);  // ../RTL/cortexm0ds_logic.v(12946)
  and u15056 (Kooow6, Rooow6, Yooow6);  // ../RTL/cortexm0ds_logic.v(12947)
  and u15057 (n4158, F0eow6, Vbgpw6[2]);  // ../RTL/cortexm0ds_logic.v(12948)
  not u15058 (Yooow6, n4158);  // ../RTL/cortexm0ds_logic.v(12948)
  and u15059 (n4159, Bagpw6[2], M6eiu6);  // ../RTL/cortexm0ds_logic.v(12949)
  buf u1506 (vis_r10_o[5], Aqlax6);  // ../RTL/cortexm0ds_logic.v(2469)
  not u15060 (Rooow6, n4159);  // ../RTL/cortexm0ds_logic.v(12949)
  and u15061 (Dooow6, Fpoow6, Mpoow6);  // ../RTL/cortexm0ds_logic.v(12950)
  and u15062 (n4160, Tzfpw6[2], Yvgiu6);  // ../RTL/cortexm0ds_logic.v(12951)
  not u15063 (Mpoow6, n4160);  // ../RTL/cortexm0ds_logic.v(12951)
  or u15064 (Fpoow6, Qkgiu6, Tfciu6);  // ../RTL/cortexm0ds_logic.v(12952)
  and u15065 (Yaoow6, Tpoow6, Aqoow6);  // ../RTL/cortexm0ds_logic.v(12953)
  and u15066 (n4161, Qtfow6, Zx3ju6);  // ../RTL/cortexm0ds_logic.v(12954)
  not u15067 (Aqoow6, n4161);  // ../RTL/cortexm0ds_logic.v(12954)
  and u15068 (n4162, Hqoow6, Oqoow6);  // ../RTL/cortexm0ds_logic.v(12955)
  not u15069 (Zx3ju6, n4162);  // ../RTL/cortexm0ds_logic.v(12955)
  buf u1507 (vis_r10_o[28], Rfibx6);  // ../RTL/cortexm0ds_logic.v(2469)
  and u15070 (Oqoow6, Vqoow6, Croow6);  // ../RTL/cortexm0ds_logic.v(12956)
  or u15071 (Croow6, Ipfow6, W40iu6);  // ../RTL/cortexm0ds_logic.v(12957)
  and u15072 (W40iu6, Jroow6, Qroow6);  // ../RTL/cortexm0ds_logic.v(12958)
  and u15073 (Qroow6, Xroow6, Esoow6);  // ../RTL/cortexm0ds_logic.v(12959)
  and u15074 (Esoow6, Lsoow6, Ssoow6);  // ../RTL/cortexm0ds_logic.v(12960)
  and u15075 (n4163, V6now6, vis_r2_o[5]);  // ../RTL/cortexm0ds_logic.v(12961)
  not u15076 (Ssoow6, n4163);  // ../RTL/cortexm0ds_logic.v(12961)
  and u15077 (n4164, C7now6, vis_r6_o[5]);  // ../RTL/cortexm0ds_logic.v(12962)
  not u15078 (Lsoow6, n4164);  // ../RTL/cortexm0ds_logic.v(12962)
  and u15079 (Xroow6, Zsoow6, Gtoow6);  // ../RTL/cortexm0ds_logic.v(12963)
  buf u1508 (vis_r10_o[6], Zrlax6);  // ../RTL/cortexm0ds_logic.v(2469)
  and u15080 (n4165, X7now6, vis_r5_o[5]);  // ../RTL/cortexm0ds_logic.v(12964)
  not u15081 (Gtoow6, n4165);  // ../RTL/cortexm0ds_logic.v(12964)
  and u15082 (n4166, E8now6, vis_r4_o[5]);  // ../RTL/cortexm0ds_logic.v(12965)
  not u15083 (Zsoow6, n4166);  // ../RTL/cortexm0ds_logic.v(12965)
  and u15084 (Jroow6, Ntoow6, Utoow6);  // ../RTL/cortexm0ds_logic.v(12966)
  and u15085 (Utoow6, Buoow6, Iuoow6);  // ../RTL/cortexm0ds_logic.v(12967)
  and u15086 (n4167, N9now6, vis_r1_o[5]);  // ../RTL/cortexm0ds_logic.v(12968)
  not u15087 (Iuoow6, n4167);  // ../RTL/cortexm0ds_logic.v(12968)
  and u15088 (n4168, U9now6, vis_r0_o[5]);  // ../RTL/cortexm0ds_logic.v(12969)
  not u15089 (Buoow6, n4168);  // ../RTL/cortexm0ds_logic.v(12969)
  buf u1509 (vis_r10_o[29], X1max6);  // ../RTL/cortexm0ds_logic.v(2469)
  and u15090 (Ntoow6, Puoow6, Wuoow6);  // ../RTL/cortexm0ds_logic.v(12970)
  and u15091 (n4169, Panow6, vis_r3_o[5]);  // ../RTL/cortexm0ds_logic.v(12971)
  not u15092 (Wuoow6, n4169);  // ../RTL/cortexm0ds_logic.v(12971)
  and u15093 (n4170, Wanow6, vis_r7_o[5]);  // ../RTL/cortexm0ds_logic.v(12972)
  not u15094 (Puoow6, n4170);  // ../RTL/cortexm0ds_logic.v(12972)
  or u15095 (Vqoow6, Kqfow6, K50iu6);  // ../RTL/cortexm0ds_logic.v(12973)
  and u15096 (K50iu6, Dvoow6, Kvoow6);  // ../RTL/cortexm0ds_logic.v(12974)
  and u15097 (Kvoow6, Rvoow6, Yvoow6);  // ../RTL/cortexm0ds_logic.v(12975)
  and u15098 (Yvoow6, Fwoow6, Mwoow6);  // ../RTL/cortexm0ds_logic.v(12976)
  and u15099 (n4171, V6now6, vis_r2_o[3]);  // ../RTL/cortexm0ds_logic.v(12977)
  buf u151 (Gqgpw6[27], W0dbx6);  // ../RTL/cortexm0ds_logic.v(2377)
  buf u1510 (vis_r10_o[22], Tzebx6);  // ../RTL/cortexm0ds_logic.v(2469)
  not u15100 (Mwoow6, n4171);  // ../RTL/cortexm0ds_logic.v(12977)
  and u15101 (n4172, C7now6, vis_r6_o[3]);  // ../RTL/cortexm0ds_logic.v(12978)
  not u15102 (Fwoow6, n4172);  // ../RTL/cortexm0ds_logic.v(12978)
  and u15103 (Rvoow6, Twoow6, Axoow6);  // ../RTL/cortexm0ds_logic.v(12979)
  and u15104 (n4173, X7now6, vis_r5_o[3]);  // ../RTL/cortexm0ds_logic.v(12980)
  not u15105 (Axoow6, n4173);  // ../RTL/cortexm0ds_logic.v(12980)
  and u15106 (n4174, E8now6, vis_r4_o[3]);  // ../RTL/cortexm0ds_logic.v(12981)
  not u15107 (Twoow6, n4174);  // ../RTL/cortexm0ds_logic.v(12981)
  and u15108 (Dvoow6, Hxoow6, Oxoow6);  // ../RTL/cortexm0ds_logic.v(12982)
  and u15109 (Oxoow6, Vxoow6, Cyoow6);  // ../RTL/cortexm0ds_logic.v(12983)
  buf u1511 (vis_ipsr_o[5], Vbkpw6);  // ../RTL/cortexm0ds_logic.v(1815)
  and u15110 (n4175, N9now6, vis_r1_o[3]);  // ../RTL/cortexm0ds_logic.v(12984)
  not u15111 (Cyoow6, n4175);  // ../RTL/cortexm0ds_logic.v(12984)
  and u15112 (n4176, U9now6, vis_r0_o[3]);  // ../RTL/cortexm0ds_logic.v(12985)
  not u15113 (Vxoow6, n4176);  // ../RTL/cortexm0ds_logic.v(12985)
  and u15114 (Hxoow6, Jyoow6, Qyoow6);  // ../RTL/cortexm0ds_logic.v(12986)
  and u15115 (n4177, Panow6, vis_r3_o[3]);  // ../RTL/cortexm0ds_logic.v(12987)
  not u15116 (Qyoow6, n4177);  // ../RTL/cortexm0ds_logic.v(12987)
  and u15117 (n4178, Wanow6, vis_r7_o[3]);  // ../RTL/cortexm0ds_logic.v(12988)
  not u15118 (Jyoow6, n4178);  // ../RTL/cortexm0ds_logic.v(12988)
  and u15119 (Hqoow6, Xyoow6, Ezoow6);  // ../RTL/cortexm0ds_logic.v(12989)
  buf u1512 (vis_r10_o[7], Ytlax6);  // ../RTL/cortexm0ds_logic.v(2469)
  or u15120 (Ezoow6, Ppfow6, F60iu6);  // ../RTL/cortexm0ds_logic.v(12990)
  and u15121 (F60iu6, Lzoow6, Szoow6);  // ../RTL/cortexm0ds_logic.v(12991)
  and u15122 (Szoow6, Zzoow6, G0pow6);  // ../RTL/cortexm0ds_logic.v(12992)
  and u15123 (G0pow6, N0pow6, U0pow6);  // ../RTL/cortexm0ds_logic.v(12993)
  and u15124 (n4179, V6now6, vis_r2_o[2]);  // ../RTL/cortexm0ds_logic.v(12994)
  not u15125 (U0pow6, n4179);  // ../RTL/cortexm0ds_logic.v(12994)
  and u15126 (n4180, C7now6, vis_r6_o[2]);  // ../RTL/cortexm0ds_logic.v(12995)
  not u15127 (N0pow6, n4180);  // ../RTL/cortexm0ds_logic.v(12995)
  and u15128 (Zzoow6, B1pow6, I1pow6);  // ../RTL/cortexm0ds_logic.v(12996)
  and u15129 (n4181, X7now6, vis_r5_o[2]);  // ../RTL/cortexm0ds_logic.v(12997)
  buf u1513 (vis_r10_o[30], Cilax6);  // ../RTL/cortexm0ds_logic.v(2469)
  not u15130 (I1pow6, n4181);  // ../RTL/cortexm0ds_logic.v(12997)
  and u15131 (n4182, E8now6, vis_r4_o[2]);  // ../RTL/cortexm0ds_logic.v(12998)
  not u15132 (B1pow6, n4182);  // ../RTL/cortexm0ds_logic.v(12998)
  and u15133 (Lzoow6, P1pow6, W1pow6);  // ../RTL/cortexm0ds_logic.v(12999)
  and u15134 (W1pow6, D2pow6, K2pow6);  // ../RTL/cortexm0ds_logic.v(13000)
  and u15135 (n4183, N9now6, vis_r1_o[2]);  // ../RTL/cortexm0ds_logic.v(13001)
  not u15136 (K2pow6, n4183);  // ../RTL/cortexm0ds_logic.v(13001)
  and u15137 (n4184, U9now6, vis_r0_o[2]);  // ../RTL/cortexm0ds_logic.v(13002)
  not u15138 (D2pow6, n4184);  // ../RTL/cortexm0ds_logic.v(13002)
  and u15139 (P1pow6, R2pow6, Y2pow6);  // ../RTL/cortexm0ds_logic.v(13003)
  buf u1514 (vis_r10_o[8], Vtmax6);  // ../RTL/cortexm0ds_logic.v(2469)
  and u15140 (n4185, Panow6, vis_r3_o[2]);  // ../RTL/cortexm0ds_logic.v(13004)
  not u15141 (Y2pow6, n4185);  // ../RTL/cortexm0ds_logic.v(13004)
  and u15142 (n4186, Wanow6, vis_r7_o[2]);  // ../RTL/cortexm0ds_logic.v(13005)
  not u15143 (R2pow6, n4186);  // ../RTL/cortexm0ds_logic.v(13005)
  or u15144 (Xyoow6, Rqfow6, D50iu6);  // ../RTL/cortexm0ds_logic.v(13006)
  and u15145 (D50iu6, F3pow6, M3pow6);  // ../RTL/cortexm0ds_logic.v(13007)
  and u15146 (M3pow6, T3pow6, A4pow6);  // ../RTL/cortexm0ds_logic.v(13008)
  and u15147 (A4pow6, H4pow6, O4pow6);  // ../RTL/cortexm0ds_logic.v(13009)
  and u15148 (n4187, V6now6, vis_r2_o[4]);  // ../RTL/cortexm0ds_logic.v(13010)
  not u15149 (O4pow6, n4187);  // ../RTL/cortexm0ds_logic.v(13010)
  buf u1515 (vis_r10_o[31], Cklax6);  // ../RTL/cortexm0ds_logic.v(2469)
  and u15150 (n4188, C7now6, vis_r6_o[4]);  // ../RTL/cortexm0ds_logic.v(13011)
  not u15151 (H4pow6, n4188);  // ../RTL/cortexm0ds_logic.v(13011)
  and u15152 (T3pow6, V4pow6, C5pow6);  // ../RTL/cortexm0ds_logic.v(13012)
  and u15153 (n4189, X7now6, vis_r5_o[4]);  // ../RTL/cortexm0ds_logic.v(13013)
  not u15154 (C5pow6, n4189);  // ../RTL/cortexm0ds_logic.v(13013)
  and u15155 (n4190, E8now6, vis_r4_o[4]);  // ../RTL/cortexm0ds_logic.v(13014)
  not u15156 (V4pow6, n4190);  // ../RTL/cortexm0ds_logic.v(13014)
  and u15157 (F3pow6, J5pow6, Q5pow6);  // ../RTL/cortexm0ds_logic.v(13015)
  and u15158 (Q5pow6, X5pow6, E6pow6);  // ../RTL/cortexm0ds_logic.v(13016)
  and u15159 (n4191, N9now6, vis_r1_o[4]);  // ../RTL/cortexm0ds_logic.v(13017)
  buf u1516 (vis_r10_o[9], Wrmax6);  // ../RTL/cortexm0ds_logic.v(2469)
  not u15160 (E6pow6, n4191);  // ../RTL/cortexm0ds_logic.v(13017)
  and u15161 (n4192, U9now6, vis_r0_o[4]);  // ../RTL/cortexm0ds_logic.v(13018)
  not u15162 (X5pow6, n4192);  // ../RTL/cortexm0ds_logic.v(13018)
  and u15163 (J5pow6, L6pow6, S6pow6);  // ../RTL/cortexm0ds_logic.v(13019)
  and u15164 (n4193, Panow6, vis_r3_o[4]);  // ../RTL/cortexm0ds_logic.v(13020)
  not u15165 (S6pow6, n4193);  // ../RTL/cortexm0ds_logic.v(13020)
  and u15166 (n4194, Wanow6, vis_r7_o[4]);  // ../RTL/cortexm0ds_logic.v(13021)
  not u15167 (L6pow6, n4194);  // ../RTL/cortexm0ds_logic.v(13021)
  and u15168 (n4195, HRDATA[2], Q2eow6);  // ../RTL/cortexm0ds_logic.v(13022)
  not u15169 (Tpoow6, n4195);  // ../RTL/cortexm0ds_logic.v(13022)
  buf u1517 (Zbhpw6[28], Ehqpw6);  // ../RTL/cortexm0ds_logic.v(2147)
  and u15170 (L2mow6, Z6pow6, G7pow6);  // ../RTL/cortexm0ds_logic.v(13023)
  or u15171 (G7pow6, Wlcow6, Kldow6);  // ../RTL/cortexm0ds_logic.v(13024)
  and u15172 (Kldow6, Dtcow6, Dahow6);  // ../RTL/cortexm0ds_logic.v(13025)
  or u15173 (Dahow6, Ch4ju6, Ktcow6);  // ../RTL/cortexm0ds_logic.v(13026)
  or u15174 (Ch4ju6, Avcow6, R3how6);  // ../RTL/cortexm0ds_logic.v(13027)
  or u15175 (n4196, Mr0iu6, N7pow6);  // ../RTL/cortexm0ds_logic.v(13028)
  not u15176 (R3how6, n4196);  // ../RTL/cortexm0ds_logic.v(13028)
  and u15177 (n4197, Jfmow6, F93ju6);  // ../RTL/cortexm0ds_logic.v(13029)
  not u15178 (Avcow6, n4197);  // ../RTL/cortexm0ds_logic.v(13029)
  and u15179 (Jfmow6, M93ju6, U54ju6);  // ../RTL/cortexm0ds_logic.v(13030)
  buf u1518 (vis_r10_o[10], Wpmax6);  // ../RTL/cortexm0ds_logic.v(2469)
  not u15180 (M93ju6, Oa3ju6);  // ../RTL/cortexm0ds_logic.v(13031)
  or u15181 (Dtcow6, Tucow6, Qxaiu6);  // ../RTL/cortexm0ds_logic.v(13032)
  and u15182 (Wlcow6, U7pow6, B8pow6);  // ../RTL/cortexm0ds_logic.v(13033)
  and u15183 (B8pow6, I8pow6, P8pow6);  // ../RTL/cortexm0ds_logic.v(13034)
  or u15184 (P8pow6, Rcfow6, R04ju6);  // ../RTL/cortexm0ds_logic.v(13035)
  and u15185 (R04ju6, W8pow6, D9pow6);  // ../RTL/cortexm0ds_logic.v(13036)
  and u15186 (D9pow6, K9pow6, R9pow6);  // ../RTL/cortexm0ds_logic.v(13037)
  or u15187 (R9pow6, Ipfow6, O70iu6);  // ../RTL/cortexm0ds_logic.v(13038)
  or u15188 (K9pow6, Rqfow6, V70iu6);  // ../RTL/cortexm0ds_logic.v(13039)
  and u15189 (W8pow6, Y9pow6, Fapow6);  // ../RTL/cortexm0ds_logic.v(13040)
  buf u1519 (Zbhpw6[30], T82qw6);  // ../RTL/cortexm0ds_logic.v(2147)
  or u15190 (Fapow6, Ppfow6, J80iu6);  // ../RTL/cortexm0ds_logic.v(13041)
  or u15191 (Y9pow6, Kqfow6, C80iu6);  // ../RTL/cortexm0ds_logic.v(13042)
  or u15192 (Rcfow6, Hfeow6, J2eow6);  // ../RTL/cortexm0ds_logic.v(13044)
  not u15193 (Dyeow6, Rcfow6);  // ../RTL/cortexm0ds_logic.v(13044)
  or u15194 (I8pow6, Iydow6, U1uiu6);  // ../RTL/cortexm0ds_logic.v(13045)
  and u15195 (U1uiu6, Mapow6, Tapow6);  // ../RTL/cortexm0ds_logic.v(13046)
  and u15196 (Tapow6, Abpow6, Hbpow6);  // ../RTL/cortexm0ds_logic.v(13047)
  and u15197 (n4198, Pceow6, Obpow6);  // ../RTL/cortexm0ds_logic.v(13048)
  not u15198 (Hbpow6, n4198);  // ../RTL/cortexm0ds_logic.v(13048)
  or u15199 (Obpow6, Nzhiu6, Vbgpw6[18]);  // ../RTL/cortexm0ds_logic.v(13049)
  buf u152 (vis_r0_o[29], E3npw6);  // ../RTL/cortexm0ds_logic.v(1875)
  buf u1520 (vis_r10_o[11], Ce7bx6);  // ../RTL/cortexm0ds_logic.v(2469)
  or u15200 (Pceow6, Nzhiu6, F0eow6);  // ../RTL/cortexm0ds_logic.v(13050)
  and u15201 (Abpow6, Vbpow6, Ccpow6);  // ../RTL/cortexm0ds_logic.v(13051)
  and u15202 (n4199, Tzfpw6[18], Yvgiu6);  // ../RTL/cortexm0ds_logic.v(13052)
  not u15203 (Ccpow6, n4199);  // ../RTL/cortexm0ds_logic.v(13052)
  and u15204 (Yvgiu6, Jcpow6, Vynow6);  // ../RTL/cortexm0ds_logic.v(13053)
  and u15205 (Jcpow6, Ynhiu6, U89iu6);  // ../RTL/cortexm0ds_logic.v(13054)
  and u15206 (n4200, Odgpw6[18], M0eow6);  // ../RTL/cortexm0ds_logic.v(13055)
  not u15207 (Vbpow6, n4200);  // ../RTL/cortexm0ds_logic.v(13055)
  and u15208 (Mapow6, Qcpow6, Qgeow6);  // ../RTL/cortexm0ds_logic.v(13056)
  and u15209 (Qgeow6, Xcpow6, Edpow6);  // ../RTL/cortexm0ds_logic.v(13058)
  and u1521 (Vnfpw6[1], Ppfpw6[7], Ivfhu6);  // ../RTL/cortexm0ds_logic.v(3367)
  not u15210 (I5eow6, Qgeow6);  // ../RTL/cortexm0ds_logic.v(13058)
  and u15211 (n4201, Ldpow6, Cpwiu6);  // ../RTL/cortexm0ds_logic.v(13059)
  not u15212 (Edpow6, n4201);  // ../RTL/cortexm0ds_logic.v(13059)
  and u15213 (Cpwiu6, Sdpow6, X8hpw6[5]);  // ../RTL/cortexm0ds_logic.v(13060)
  or u15214 (n4202, X8hpw6[0], X8hpw6[6]);  // ../RTL/cortexm0ds_logic.v(13061)
  not u15215 (Sdpow6, n4202);  // ../RTL/cortexm0ds_logic.v(13061)
  and u15216 (Ldpow6, Ilwiu6, Q4wiu6);  // ../RTL/cortexm0ds_logic.v(13062)
  or u15217 (n4203, X8hpw6[1], X8hpw6[4]);  // ../RTL/cortexm0ds_logic.v(13063)
  not u15218 (Q4wiu6, n4203);  // ../RTL/cortexm0ds_logic.v(13063)
  and u15219 (Ilwiu6, X8hpw6[2], Vm6iu6);  // ../RTL/cortexm0ds_logic.v(13064)
  buf u1522 (vis_r10_o[12], Wnmax6);  // ../RTL/cortexm0ds_logic.v(2469)
  not u15220 (Vm6iu6, X8hpw6[3]);  // ../RTL/cortexm0ds_logic.v(13065)
  and u15221 (n4204, Xznow6, K5eiu6);  // ../RTL/cortexm0ds_logic.v(13066)
  not u15222 (Xcpow6, n4204);  // ../RTL/cortexm0ds_logic.v(13066)
  and u15223 (Xznow6, Zdpow6, Jfgpw6[2]);  // ../RTL/cortexm0ds_logic.v(13067)
  and u15224 (Qcpow6, Gepow6, Nepow6);  // ../RTL/cortexm0ds_logic.v(13068)
  and u15225 (n4205, Bagpw6[18], M6eiu6);  // ../RTL/cortexm0ds_logic.v(13069)
  not u15226 (Nepow6, n4205);  // ../RTL/cortexm0ds_logic.v(13069)
  and u15227 (M6eiu6, Vynow6, D5eiu6);  // ../RTL/cortexm0ds_logic.v(13070)
  and u15228 (n4206, STCALIB[18], H1eow6);  // ../RTL/cortexm0ds_logic.v(13071)
  not u15229 (Gepow6, n4206);  // ../RTL/cortexm0ds_logic.v(13071)
  and u1523 (Vnfpw6[2], Ppfpw6[8], Ivfhu6);  // ../RTL/cortexm0ds_logic.v(3367)
  and u15230 (H1eow6, Uepow6, Vynow6);  // ../RTL/cortexm0ds_logic.v(13072)
  or u15231 (n4207, Uh7iu6, Jfgpw6[1]);  // ../RTL/cortexm0ds_logic.v(13073)
  not u15232 (Vynow6, n4207);  // ../RTL/cortexm0ds_logic.v(13073)
  and u15233 (Uepow6, Ynhiu6, Jfgpw6[4]);  // ../RTL/cortexm0ds_logic.v(13074)
  and u15234 (Ynhiu6, Jfgpw6[3], Jfgpw6[2]);  // ../RTL/cortexm0ds_logic.v(13075)
  and u15235 (U7pow6, Bfpow6, Ifpow6);  // ../RTL/cortexm0ds_logic.v(13076)
  and u15236 (n4208, Qtfow6, Ye4ju6);  // ../RTL/cortexm0ds_logic.v(13077)
  not u15237 (Ifpow6, n4208);  // ../RTL/cortexm0ds_logic.v(13077)
  and u15238 (n4209, Pfpow6, Wfpow6);  // ../RTL/cortexm0ds_logic.v(13078)
  not u15239 (Ye4ju6, n4209);  // ../RTL/cortexm0ds_logic.v(13078)
  buf u1524 (vis_r10_o[13], Wlmax6);  // ../RTL/cortexm0ds_logic.v(2469)
  and u15240 (Wfpow6, Dgpow6, Kgpow6);  // ../RTL/cortexm0ds_logic.v(13079)
  or u15241 (Kgpow6, Ipfow6, Q80iu6);  // ../RTL/cortexm0ds_logic.v(13080)
  or u15242 (Dgpow6, Ppfow6, S90iu6);  // ../RTL/cortexm0ds_logic.v(13081)
  and u15243 (Pfpow6, Rgpow6, Ygpow6);  // ../RTL/cortexm0ds_logic.v(13082)
  or u15244 (Ygpow6, Kqfow6, L90iu6);  // ../RTL/cortexm0ds_logic.v(13083)
  or u15245 (Rgpow6, Rqfow6, X80iu6);  // ../RTL/cortexm0ds_logic.v(13084)
  or u15246 (Uafow6, Hfeow6, Hv3ju6);  // ../RTL/cortexm0ds_logic.v(13085)
  not u15247 (Qtfow6, Uafow6);  // ../RTL/cortexm0ds_logic.v(13085)
  not u15248 (Hfeow6, C2eow6);  // ../RTL/cortexm0ds_logic.v(13086)
  and u15249 (n4210, HRDATA[18], Q2eow6);  // ../RTL/cortexm0ds_logic.v(13087)
  and u1525 (Vnfpw6[3], Ppfpw6[9], Ivfhu6);  // ../RTL/cortexm0ds_logic.v(3367)
  not u15250 (Bfpow6, n4210);  // ../RTL/cortexm0ds_logic.v(13087)
  or u15251 (Z6pow6, Ukcow6, Spdow6);  // ../RTL/cortexm0ds_logic.v(13088)
  and u15252 (Spdow6, Fhpow6, Mhpow6);  // ../RTL/cortexm0ds_logic.v(13090)
  not u15253 (Fmdow6, Spdow6);  // ../RTL/cortexm0ds_logic.v(13090)
  and u15254 (n4211, T4how6, Cyfpw6[3]);  // ../RTL/cortexm0ds_logic.v(13091)
  not u15255 (Mhpow6, n4211);  // ../RTL/cortexm0ds_logic.v(13091)
  and u15256 (T4how6, Thpow6, Iwfpw6[1]);  // ../RTL/cortexm0ds_logic.v(13092)
  or u15257 (n4212, Tucow6, Cyfpw6[1]);  // ../RTL/cortexm0ds_logic.v(13093)
  not u15258 (Thpow6, n4212);  // ../RTL/cortexm0ds_logic.v(13093)
  and u15259 (Fhpow6, F4how6, K3how6);  // ../RTL/cortexm0ds_logic.v(13094)
  buf u1526 (vis_r10_o[14], Wjmax6);  // ../RTL/cortexm0ds_logic.v(2469)
  or u15260 (K3how6, L7how6, Ktcow6);  // ../RTL/cortexm0ds_logic.v(13095)
  not u15261 (L7how6, Pe3ju6);  // ../RTL/cortexm0ds_logic.v(13097)
  and u15262 (Pe3ju6, Aipow6, Oa3ju6);  // ../RTL/cortexm0ds_logic.v(13098)
  and u15263 (Aipow6, Ej3ju6, U54ju6);  // ../RTL/cortexm0ds_logic.v(13099)
  or u15264 (U54ju6, Ii0iu6, Z53ju6);  // ../RTL/cortexm0ds_logic.v(13100)
  and u15265 (Z53ju6, Hipow6, Oipow6);  // ../RTL/cortexm0ds_logic.v(13102)
  not u15266 (Q43ju6, Z53ju6);  // ../RTL/cortexm0ds_logic.v(13102)
  and u15267 (n4213, Vipow6, Cjpow6);  // ../RTL/cortexm0ds_logic.v(13103)
  not u15268 (Oipow6, n4213);  // ../RTL/cortexm0ds_logic.v(13103)
  and u15269 (Cjpow6, Jjpow6, Qjpow6);  // ../RTL/cortexm0ds_logic.v(13104)
  and u1527 (Vnfpw6[4], Ppfpw6[10], Ivfhu6);  // ../RTL/cortexm0ds_logic.v(3367)
  or u15270 (n4214, S8fpw6[4], H4ghu6);  // ../RTL/cortexm0ds_logic.v(13105)
  not u15271 (Qjpow6, n4214);  // ../RTL/cortexm0ds_logic.v(13105)
  or u15272 (n4215, S8fpw6[2], S8fpw6[3]);  // ../RTL/cortexm0ds_logic.v(13106)
  not u15273 (Jjpow6, n4215);  // ../RTL/cortexm0ds_logic.v(13106)
  and u15274 (Vipow6, Xjpow6, Pugiu6);  // ../RTL/cortexm0ds_logic.v(13107)
  or u15275 (n4216, S8fpw6[0], S8fpw6[1]);  // ../RTL/cortexm0ds_logic.v(13108)
  not u15276 (Xjpow6, n4216);  // ../RTL/cortexm0ds_logic.v(13108)
  and u15277 (Hipow6, Ekpow6, Zc3ju6);  // ../RTL/cortexm0ds_logic.v(13109)
  and u15278 (n4217, Pfoiu6, Lkpow6);  // ../RTL/cortexm0ds_logic.v(13110)
  not u15279 (Zc3ju6, n4217);  // ../RTL/cortexm0ds_logic.v(13110)
  buf u1528 (vis_r10_o[15], Z38bx6);  // ../RTL/cortexm0ds_logic.v(2469)
  and u15280 (n4218, Zvzhu6, Svzhu6);  // ../RTL/cortexm0ds_logic.v(13111)
  not u15281 (Lkpow6, n4218);  // ../RTL/cortexm0ds_logic.v(13111)
  or u15282 (Ekpow6, Yn2ju6, Gwzhu6);  // ../RTL/cortexm0ds_logic.v(13112)
  and u15283 (n4219, Skpow6, Zkpow6);  // ../RTL/cortexm0ds_logic.v(13113)
  not u15284 (F4how6, n4219);  // ../RTL/cortexm0ds_logic.v(13113)
  or u15285 (n4220, Wmaiu6, Tr0iu6);  // ../RTL/cortexm0ds_logic.v(13114)
  not u15286 (Zkpow6, n4220);  // ../RTL/cortexm0ds_logic.v(13114)
  not u15287 (Wmaiu6, Glpow6);  // ../RTL/cortexm0ds_logic.v(13115)
  or u15288 (n4221, Yahow6, Tucow6);  // ../RTL/cortexm0ds_logic.v(13116)
  not u15289 (Skpow6, n4221);  // ../RTL/cortexm0ds_logic.v(13116)
  and u1529 (Vnfpw6[5], Ppfpw6[11], Ivfhu6);  // ../RTL/cortexm0ds_logic.v(3367)
  and u15290 (Ktcow6, Qcoiu6, Nlpow6);  // ../RTL/cortexm0ds_logic.v(13117)
  not u15291 (Tucow6, Ktcow6);  // ../RTL/cortexm0ds_logic.v(13117)
  and u15292 (n4222, Ulpow6, Xkaow6);  // ../RTL/cortexm0ds_logic.v(13118)
  not u15293 (Nlpow6, n4222);  // ../RTL/cortexm0ds_logic.v(13118)
  or u15294 (n4223, Imaiu6, Y7ghu6);  // ../RTL/cortexm0ds_logic.v(13119)
  not u15295 (Ulpow6, n4223);  // ../RTL/cortexm0ds_logic.v(13119)
  not u15296 (Qcoiu6, Bmpow6);  // ../RTL/cortexm0ds_logic.v(13120)
  not u15297 (Yahow6, Iwfpw6[1]);  // ../RTL/cortexm0ds_logic.v(13121)
  and u15298 (Ukcow6, Impow6, Pmpow6);  // ../RTL/cortexm0ds_logic.v(13122)
  or u15299 (Pmpow6, Iydow6, Wmviu6);  // ../RTL/cortexm0ds_logic.v(13123)
  buf u153 (vis_r12_o[18], Ektax6);  // ../RTL/cortexm0ds_logic.v(2599)
  buf u1530 (vis_r10_o[16], Whmax6);  // ../RTL/cortexm0ds_logic.v(2469)
  and u15300 (Wmviu6, Wmpow6, Dnpow6);  // ../RTL/cortexm0ds_logic.v(13124)
  and u15301 (n4224, Odgpw6[26], M0eow6);  // ../RTL/cortexm0ds_logic.v(13125)
  not u15302 (Dnpow6, n4224);  // ../RTL/cortexm0ds_logic.v(13125)
  and u15303 (M0eow6, Pjyiu6, Knpow6);  // ../RTL/cortexm0ds_logic.v(13126)
  and u15304 (Pjyiu6, Jfgpw6[0], Jfgpw6[1]);  // ../RTL/cortexm0ds_logic.v(13127)
  and u15305 (Wmpow6, Rnpow6, Ynpow6);  // ../RTL/cortexm0ds_logic.v(13128)
  and u15306 (n4225, F0eow6, Vbgpw6[26]);  // ../RTL/cortexm0ds_logic.v(13129)
  not u15307 (Ynpow6, n4225);  // ../RTL/cortexm0ds_logic.v(13129)
  and u15308 (F0eow6, K5eiu6, Knpow6);  // ../RTL/cortexm0ds_logic.v(13130)
  or u15309 (Knpow6, Wjyiu6, D5eiu6);  // ../RTL/cortexm0ds_logic.v(13131)
  and u1531 (Vnfpw6[6], Ppfpw6[12], Ivfhu6);  // ../RTL/cortexm0ds_logic.v(3367)
  and u15310 (D5eiu6, Fopow6, Jfgpw6[4]);  // ../RTL/cortexm0ds_logic.v(13132)
  or u15311 (n4226, Jfgpw6[2], Jfgpw6[3]);  // ../RTL/cortexm0ds_logic.v(13133)
  not u15312 (Fopow6, n4226);  // ../RTL/cortexm0ds_logic.v(13133)
  and u15313 (n4227, Yyghu6, T7eow6);  // ../RTL/cortexm0ds_logic.v(13134)
  not u15314 (Rnpow6, n4227);  // ../RTL/cortexm0ds_logic.v(13134)
  and u15315 (T7eow6, K5eiu6, Dtjow6);  // ../RTL/cortexm0ds_logic.v(13136)
  not u15316 (Qkgiu6, T7eow6);  // ../RTL/cortexm0ds_logic.v(13136)
  and u15317 (Dtjow6, Mopow6, Jfgpw6[4]);  // ../RTL/cortexm0ds_logic.v(13137)
  or u15318 (n4228, Ka9iu6, Jfgpw6[3]);  // ../RTL/cortexm0ds_logic.v(13138)
  not u15319 (Mopow6, n4228);  // ../RTL/cortexm0ds_logic.v(13138)
  buf u1532 (Bagpw6[7], Thxax6);  // ../RTL/cortexm0ds_logic.v(2680)
  and u15320 (n4229, Hemow6, Topow6);  // ../RTL/cortexm0ds_logic.v(13139)
  not u15321 (Iydow6, n4229);  // ../RTL/cortexm0ds_logic.v(13139)
  and u15322 (Ytwiu6, Rzciu6, Wjyiu6);  // ../RTL/cortexm0ds_logic.v(13140)
  not u15323 (Topow6, Ytwiu6);  // ../RTL/cortexm0ds_logic.v(13140)
  and u15324 (Impow6, Appow6, Hppow6);  // ../RTL/cortexm0ds_logic.v(13141)
  and u15325 (n4230, C2eow6, Oppow6);  // ../RTL/cortexm0ds_logic.v(13142)
  not u15326 (Hppow6, n4230);  // ../RTL/cortexm0ds_logic.v(13142)
  and u15327 (n4231, Vppow6, Cqpow6);  // ../RTL/cortexm0ds_logic.v(13143)
  not u15328 (Oppow6, n4231);  // ../RTL/cortexm0ds_logic.v(13143)
  or u15329 (Cqpow6, Jqpow6, Bz3ju6);  // ../RTL/cortexm0ds_logic.v(13144)
  and u1533 (Dqfhu6, H6ghu6, No0iu6);  // ../RTL/cortexm0ds_logic.v(3481)
  and u15330 (Vh3ju6, Qqpow6, E5ehu6);  // ../RTL/cortexm0ds_logic.v(13145)
  not u15331 (Bz3ju6, Vh3ju6);  // ../RTL/cortexm0ds_logic.v(13145)
  or u15332 (n4232, Xqpow6, R50iu6);  // ../RTL/cortexm0ds_logic.v(13146)
  not u15333 (Qqpow6, n4232);  // ../RTL/cortexm0ds_logic.v(13146)
  or u15334 (n4233, F3aiu6, Pt2ju6);  // ../RTL/cortexm0ds_logic.v(13147)
  not u15335 (Xqpow6, n4233);  // ../RTL/cortexm0ds_logic.v(13147)
  and u15336 (n4234, F84ju6, Erpow6);  // ../RTL/cortexm0ds_logic.v(13148)
  not u15337 (Vppow6, n4234);  // ../RTL/cortexm0ds_logic.v(13148)
  or u15338 (Erpow6, O24ju6, Hv3ju6);  // ../RTL/cortexm0ds_logic.v(13149)
  and u15339 (Wkkow6, Lrpow6, Srpow6);  // ../RTL/cortexm0ds_logic.v(13150)
  and u1534 (n116, Uo0iu6, Bp0iu6);  // ../RTL/cortexm0ds_logic.v(3482)
  not u15340 (O24ju6, Wkkow6);  // ../RTL/cortexm0ds_logic.v(13150)
  and u15341 (Srpow6, Zrpow6, Gspow6);  // ../RTL/cortexm0ds_logic.v(13151)
  or u15342 (Gspow6, Ipfow6, M60iu6);  // ../RTL/cortexm0ds_logic.v(13152)
  or u15343 (Zrpow6, Ppfow6, H70iu6);  // ../RTL/cortexm0ds_logic.v(13153)
  and u15344 (Lrpow6, Nspow6, Uspow6);  // ../RTL/cortexm0ds_logic.v(13154)
  or u15345 (Uspow6, Kqfow6, A70iu6);  // ../RTL/cortexm0ds_logic.v(13155)
  or u15346 (Nspow6, Rqfow6, T60iu6);  // ../RTL/cortexm0ds_logic.v(13156)
  and u15347 (F84ju6, Btpow6, Jqpow6);  // ../RTL/cortexm0ds_logic.v(13157)
  and u15348 (n4235, Itpow6, Jbjow6);  // ../RTL/cortexm0ds_logic.v(13158)
  not u15349 (Jqpow6, n4235);  // ../RTL/cortexm0ds_logic.v(13158)
  not u1535 (No0iu6, n116);  // ../RTL/cortexm0ds_logic.v(3482)
  and u15350 (Jbjow6, Ptpow6, Cyfpw6[3]);  // ../RTL/cortexm0ds_logic.v(13159)
  and u15351 (Ptpow6, Wtpow6, Azfow6);  // ../RTL/cortexm0ds_logic.v(13160)
  not u15352 (Azfow6, Lveow6);  // ../RTL/cortexm0ds_logic.v(13161)
  and u15353 (Lveow6, J2eow6, Uieow6);  // ../RTL/cortexm0ds_logic.v(13162)
  or u15354 (Wtpow6, Ppfow6, V2kow6);  // ../RTL/cortexm0ds_logic.v(13164)
  AL_MUX u15355 (
    .i0(V2kow6),
    .i1(Qbjow6),
    .sel(Kqfow6),
    .o(Itpow6));  // ../RTL/cortexm0ds_logic.v(13165)
  or u15356 (Qbjow6, Hzfow6, Dupow6);  // ../RTL/cortexm0ds_logic.v(13166)
  and u15357 (n4236, V2kow6, Hv3ju6);  // ../RTL/cortexm0ds_logic.v(13167)
  not u15358 (Hzfow6, n4236);  // ../RTL/cortexm0ds_logic.v(13167)
  or u15359 (Uieow6, N7pow6, Df3ju6);  // ../RTL/cortexm0ds_logic.v(13168)
  and u1536 (Bp0iu6, Ip0iu6, Pp0iu6);  // ../RTL/cortexm0ds_logic.v(3483)
  not u15360 (V2kow6, Uieow6);  // ../RTL/cortexm0ds_logic.v(13168)
  and u15361 (Df3ju6, Vwaiu6, Mr0iu6);  // ../RTL/cortexm0ds_logic.v(13169)
  and u15362 (N7pow6, Kupow6, Rupow6);  // ../RTL/cortexm0ds_logic.v(13170)
  or u15363 (n4237, F93ju6, Oa3ju6);  // ../RTL/cortexm0ds_logic.v(13171)
  not u15364 (Rupow6, n4237);  // ../RTL/cortexm0ds_logic.v(13171)
  AL_MUX u15365 (
    .i0(X43ju6),
    .i1(Yupow6),
    .sel(H4ghu6),
    .o(Oa3ju6));  // ../RTL/cortexm0ds_logic.v(13172)
  xor u15366 (n4238, G63ju6, Sc3ju6);  // ../RTL/cortexm0ds_logic.v(13173)
  not u15367 (Yupow6, n4238);  // ../RTL/cortexm0ds_logic.v(13173)
  and u15368 (Sc3ju6, Fvpow6, Mvpow6);  // ../RTL/cortexm0ds_logic.v(13175)
  not u15369 (X43ju6, Sc3ju6);  // ../RTL/cortexm0ds_logic.v(13175)
  and u1537 (n117, Wp0iu6, Dq0iu6);  // ../RTL/cortexm0ds_logic.v(3484)
  or u15370 (Mvpow6, Yn2ju6, Nwzhu6);  // ../RTL/cortexm0ds_logic.v(13176)
  or u15371 (Fvpow6, A4oiu6, Qjoiu6);  // ../RTL/cortexm0ds_logic.v(13177)
  not u15372 (F93ju6, Ej3ju6);  // ../RTL/cortexm0ds_logic.v(13178)
  AL_MUX u15373 (
    .i0(Tvpow6),
    .i1(Awpow6),
    .sel(H4ghu6),
    .o(Ej3ju6));  // ../RTL/cortexm0ds_logic.v(13179)
  and u15374 (n4239, Hwpow6, G63ju6);  // ../RTL/cortexm0ds_logic.v(13180)
  not u15375 (Awpow6, n4239);  // ../RTL/cortexm0ds_logic.v(13180)
  or u15376 (G63ju6, Owpow6, Vwpow6);  // ../RTL/cortexm0ds_logic.v(13181)
  and u15377 (n4240, Vwpow6, Owpow6);  // ../RTL/cortexm0ds_logic.v(13182)
  not u15378 (Hwpow6, n4240);  // ../RTL/cortexm0ds_logic.v(13182)
  and u15379 (Tvpow6, Cxpow6, Jxpow6);  // ../RTL/cortexm0ds_logic.v(13184)
  not u1538 (Pp0iu6, n117);  // ../RTL/cortexm0ds_logic.v(3484)
  not u15380 (Owpow6, Tvpow6);  // ../RTL/cortexm0ds_logic.v(13184)
  or u15381 (Jxpow6, Yn2ju6, Uwzhu6);  // ../RTL/cortexm0ds_logic.v(13185)
  or u15382 (Cxpow6, Cajiu6, A4oiu6);  // ../RTL/cortexm0ds_logic.v(13186)
  not u15383 (Cajiu6, S8fpw6[3]);  // ../RTL/cortexm0ds_logic.v(13187)
  or u15384 (n4241, Hv3ju6, Ppfow6);  // ../RTL/cortexm0ds_logic.v(13188)
  not u15385 (Kupow6, n4241);  // ../RTL/cortexm0ds_logic.v(13188)
  not u15386 (Hv3ju6, J2eow6);  // ../RTL/cortexm0ds_logic.v(13189)
  or u15387 (Btpow6, Eolow6, J2eow6);  // ../RTL/cortexm0ds_logic.v(13190)
  AL_MUX u15388 (
    .i0(Qxpow6),
    .i1(Xxpow6),
    .sel(H4ghu6),
    .o(J2eow6));  // ../RTL/cortexm0ds_logic.v(13191)
  and u15389 (n4242, Eypow6, Vwpow6);  // ../RTL/cortexm0ds_logic.v(13192)
  and u1539 (n118, Kq0iu6, Rq0iu6);  // ../RTL/cortexm0ds_logic.v(3485)
  not u15390 (Xxpow6, n4242);  // ../RTL/cortexm0ds_logic.v(13192)
  or u15391 (Vwpow6, Lypow6, Sypow6);  // ../RTL/cortexm0ds_logic.v(13193)
  and u15392 (n4243, Sypow6, Lypow6);  // ../RTL/cortexm0ds_logic.v(13194)
  not u15393 (Eypow6, n4243);  // ../RTL/cortexm0ds_logic.v(13194)
  not u15394 (Lypow6, Qxpow6);  // ../RTL/cortexm0ds_logic.v(13195)
  and u15395 (Qxpow6, Zypow6, Gzpow6);  // ../RTL/cortexm0ds_logic.v(13196)
  or u15396 (Gzpow6, Yn2ju6, Pxzhu6);  // ../RTL/cortexm0ds_logic.v(13197)
  or u15397 (Zypow6, B5kiu6, A4oiu6);  // ../RTL/cortexm0ds_logic.v(13198)
  and u15398 (n4244, Nzpow6, Uzpow6);  // ../RTL/cortexm0ds_logic.v(13199)
  not u15399 (Eolow6, n4244);  // ../RTL/cortexm0ds_logic.v(13199)
  buf u154 (Yyghu6, Zdtpw6);  // ../RTL/cortexm0ds_logic.v(1984)
  not u1540 (Dq0iu6, n118);  // ../RTL/cortexm0ds_logic.v(3485)
  and u15400 (Uzpow6, B0qow6, I0qow6);  // ../RTL/cortexm0ds_logic.v(13200)
  or u15401 (I0qow6, Ipfow6, E90iu6);  // ../RTL/cortexm0ds_logic.v(13201)
  or u15402 (Ipfow6, P0qow6, W0qow6);  // ../RTL/cortexm0ds_logic.v(13202)
  or u15403 (B0qow6, Rqfow6, Dc0iu6);  // ../RTL/cortexm0ds_logic.v(13203)
  not u15404 (n6000, I5khu6);  // ../RTL/cortexm0ds_logic.v(3118)
  or u15405 (Rqfow6, D1qow6, P0qow6);  // ../RTL/cortexm0ds_logic.v(13205)
  not u15406 (Gweow6, Rqfow6);  // ../RTL/cortexm0ds_logic.v(13205)
  and u15407 (Nzpow6, K1qow6, R1qow6);  // ../RTL/cortexm0ds_logic.v(13206)
  or u15408 (R1qow6, Ppfow6, Y50iu6);  // ../RTL/cortexm0ds_logic.v(13207)
  not u15409 (Ppfow6, Dupow6);  // ../RTL/cortexm0ds_logic.v(13208)
  and u1541 (n119, Yq0iu6, Fr0iu6);  // ../RTL/cortexm0ds_logic.v(3486)
  and u15410 (Dupow6, P0qow6, W0qow6);  // ../RTL/cortexm0ds_logic.v(13209)
  or u15411 (K1qow6, Kqfow6, R50iu6);  // ../RTL/cortexm0ds_logic.v(13210)
  not u15412 (Kqfow6, C3kow6);  // ../RTL/cortexm0ds_logic.v(13211)
  and u15413 (C3kow6, P0qow6, D1qow6);  // ../RTL/cortexm0ds_logic.v(13212)
  AL_MUX u15414 (
    .i0(Y1qow6),
    .i1(F2qow6),
    .sel(H4ghu6),
    .o(P0qow6));  // ../RTL/cortexm0ds_logic.v(13213)
  and u15415 (n4245, M2qow6, Sypow6);  // ../RTL/cortexm0ds_logic.v(13214)
  not u15416 (F2qow6, n4245);  // ../RTL/cortexm0ds_logic.v(13214)
  and u15417 (n4246, Y1qow6, W0qow6);  // ../RTL/cortexm0ds_logic.v(13215)
  not u15418 (Sypow6, n4246);  // ../RTL/cortexm0ds_logic.v(13215)
  or u15419 (M2qow6, W0qow6, Y1qow6);  // ../RTL/cortexm0ds_logic.v(13216)
  not u1542 (Rq0iu6, n119);  // ../RTL/cortexm0ds_logic.v(3486)
  and u15420 (W0qow6, T2qow6, A3qow6);  // ../RTL/cortexm0ds_logic.v(13218)
  not u15421 (D1qow6, W0qow6);  // ../RTL/cortexm0ds_logic.v(13218)
  or u15422 (A3qow6, Yn2ju6, N30iu6);  // ../RTL/cortexm0ds_logic.v(13219)
  or u15423 (T2qow6, Je8iu6, A4oiu6);  // ../RTL/cortexm0ds_logic.v(13220)
  not u15424 (Je8iu6, S8fpw6[0]);  // ../RTL/cortexm0ds_logic.v(13221)
  and u15425 (Y1qow6, H3qow6, O3qow6);  // ../RTL/cortexm0ds_logic.v(13222)
  or u15426 (O3qow6, Yn2ju6, O00iu6);  // ../RTL/cortexm0ds_logic.v(13223)
  or u15427 (H3qow6, Y8biu6, A4oiu6);  // ../RTL/cortexm0ds_logic.v(13224)
  not u15428 (Y8biu6, S8fpw6[1]);  // ../RTL/cortexm0ds_logic.v(13225)
  and u15429 (C2eow6, E5ehu6, V3qow6);  // ../RTL/cortexm0ds_logic.v(13226)
  or u1543 (Tq8iu6, Mr0iu6, Tr0iu6);  // ../RTL/cortexm0ds_logic.v(3487)
  and u15430 (n4247, C4qow6, J4qow6);  // ../RTL/cortexm0ds_logic.v(13227)
  not u15431 (V3qow6, n4247);  // ../RTL/cortexm0ds_logic.v(13227)
  or u15432 (J4qow6, Tr0iu6, Gwyiu6);  // ../RTL/cortexm0ds_logic.v(13228)
  or u15433 (n4248, Bmpow6, A3aju6);  // ../RTL/cortexm0ds_logic.v(13229)
  not u15434 (C4qow6, n4248);  // ../RTL/cortexm0ds_logic.v(13229)
  and u15435 (Bmpow6, Hs0iu6, K9aiu6);  // ../RTL/cortexm0ds_logic.v(13230)
  and u15436 (n4249, HRDATA[26], Q2eow6);  // ../RTL/cortexm0ds_logic.v(13231)
  not u15437 (Appow6, n4249);  // ../RTL/cortexm0ds_logic.v(13231)
  and u15438 (Q2eow6, Ytwiu6, Hemow6);  // ../RTL/cortexm0ds_logic.v(13232)
  or u15439 (n4250, Nm1ju6, Q4qow6);  // ../RTL/cortexm0ds_logic.v(13233)
  not u1544 (Fr0iu6, Tq8iu6);  // ../RTL/cortexm0ds_logic.v(3487)
  not u15440 (Hemow6, n4250);  // ../RTL/cortexm0ds_logic.v(13233)
  or u15441 (n4251, X4qow6, E5qow6);  // ../RTL/cortexm0ds_logic.v(13234)
  not u15442 (Q4qow6, n4251);  // ../RTL/cortexm0ds_logic.v(13234)
  AL_MUX u15443 (
    .i0(L5qow6),
    .i1(Glpow6),
    .sel(Cyfpw6[1]),
    .o(E5qow6));  // ../RTL/cortexm0ds_logic.v(13235)
  and u15444 (Glpow6, Gwyiu6, Nlaiu6);  // ../RTL/cortexm0ds_logic.v(13236)
  or u15445 (n4252, S5qow6, Hs0iu6);  // ../RTL/cortexm0ds_logic.v(13237)
  not u15446 (L5qow6, n4252);  // ../RTL/cortexm0ds_logic.v(13237)
  and u15447 (n4253, Z5qow6, K9aiu6);  // ../RTL/cortexm0ds_logic.v(13238)
  not u15448 (X4qow6, n4253);  // ../RTL/cortexm0ds_logic.v(13238)
  or u15449 (Z5qow6, Xkaow6, C0ehu6);  // ../RTL/cortexm0ds_logic.v(13239)
  or u1545 (n120, As0iu6, Hs0iu6);  // ../RTL/cortexm0ds_logic.v(3488)
  not u15450 (Nm1ju6, E5ehu6);  // ../RTL/cortexm0ds_logic.v(13240)
  buf u15451 (Dkfhu6, Ozkbx6[4]);  // ../RTL/cortexm0ds_logic.v(3176)
  and u15452 (Wjyiu6, Zdpow6, Ka9iu6);  // ../RTL/cortexm0ds_logic.v(13242)
  not u15453 (Ka9iu6, Jfgpw6[2]);  // ../RTL/cortexm0ds_logic.v(13243)
  or u15454 (n4254, Jfgpw6[3], Jfgpw6[4]);  // ../RTL/cortexm0ds_logic.v(13244)
  not u15455 (Zdpow6, n4254);  // ../RTL/cortexm0ds_logic.v(13244)
  or u15456 (n4255, Jfgpw6[0], Jfgpw6[1]);  // ../RTL/cortexm0ds_logic.v(13245)
  not u15457 (Rzciu6, n4255);  // ../RTL/cortexm0ds_logic.v(13245)
  or u15458 (Ft6ow6, Jmziu6, Gu8iu6);  // ../RTL/cortexm0ds_logic.v(13246)
  not u15459 (Zgziu6, Ft6ow6);  // ../RTL/cortexm0ds_logic.v(13246)
  not u1546 (Yq0iu6, n120);  // ../RTL/cortexm0ds_logic.v(3488)
  and u15460 (A0mow6, G6qow6, N6qow6);  // ../RTL/cortexm0ds_logic.v(13247)
  and u15461 (n4256, Zsfpw6[9], Cmziu6);  // ../RTL/cortexm0ds_logic.v(13248)
  not u15462 (N6qow6, n4256);  // ../RTL/cortexm0ds_logic.v(13248)
  or u15463 (n4257, Hr8iu6, Jmziu6);  // ../RTL/cortexm0ds_logic.v(13249)
  not u15464 (Cmziu6, n4257);  // ../RTL/cortexm0ds_logic.v(13249)
  or u15465 (Hr8iu6, Et8iu6, U6qow6);  // ../RTL/cortexm0ds_logic.v(13250)
  and u15466 (n4258, vis_pc_o[9], Jmziu6);  // ../RTL/cortexm0ds_logic.v(13251)
  not u15467 (G6qow6, n4258);  // ../RTL/cortexm0ds_logic.v(13251)
  and u15468 (Ar8iu6, HREADY, B7qow6);  // ../RTL/cortexm0ds_logic.v(13252)
  not u15469 (Jmziu6, Ar8iu6);  // ../RTL/cortexm0ds_logic.v(13252)
  and u1547 (n121, C0ehu6, Os0iu6);  // ../RTL/cortexm0ds_logic.v(3489)
  and u15470 (n4259, I7qow6, P7qow6);  // ../RTL/cortexm0ds_logic.v(13253)
  not u15471 (Acohu6, n4259);  // ../RTL/cortexm0ds_logic.v(13253)
  and u15472 (n4260, Umhow6, HRDATA[19]);  // ../RTL/cortexm0ds_logic.v(13254)
  not u15473 (P7qow6, n4260);  // ../RTL/cortexm0ds_logic.v(13254)
  and u15474 (n4261, Hrfpw6[3], Qqhiu6);  // ../RTL/cortexm0ds_logic.v(13255)
  not u15475 (I7qow6, n4261);  // ../RTL/cortexm0ds_logic.v(13255)
  and u15476 (n4262, W7qow6, D8qow6);  // ../RTL/cortexm0ds_logic.v(13256)
  not u15477 (Tbohu6, n4262);  // ../RTL/cortexm0ds_logic.v(13256)
  and u15478 (n4263, Umhow6, HRDATA[18]);  // ../RTL/cortexm0ds_logic.v(13257)
  not u15479 (D8qow6, n4263);  // ../RTL/cortexm0ds_logic.v(13257)
  not u1548 (Ip0iu6, n121);  // ../RTL/cortexm0ds_logic.v(3489)
  and u15480 (n4264, Hrfpw6[2], Qqhiu6);  // ../RTL/cortexm0ds_logic.v(13258)
  not u15481 (W7qow6, n4264);  // ../RTL/cortexm0ds_logic.v(13258)
  and u15482 (n4265, K8qow6, R8qow6);  // ../RTL/cortexm0ds_logic.v(13259)
  not u15483 (Mbohu6, n4265);  // ../RTL/cortexm0ds_logic.v(13259)
  and u15484 (n4266, Umhow6, HRDATA[17]);  // ../RTL/cortexm0ds_logic.v(13260)
  not u15485 (R8qow6, n4266);  // ../RTL/cortexm0ds_logic.v(13260)
  or u15486 (n4267, Wz4iu6, Qqhiu6);  // ../RTL/cortexm0ds_logic.v(13261)
  not u15487 (Umhow6, n4267);  // ../RTL/cortexm0ds_logic.v(13261)
  not u15488 (Wz4iu6, Glhiu6);  // ../RTL/cortexm0ds_logic.v(13262)
  and u15489 (Glhiu6, Vobiu6, Hs7iu6);  // ../RTL/cortexm0ds_logic.v(13263)
  or u1549 (Os0iu6, Vs0iu6, Ct0iu6);  // ../RTL/cortexm0ds_logic.v(3490)
  and u15490 (n4268, Hrfpw6[1], Qqhiu6);  // ../RTL/cortexm0ds_logic.v(13264)
  not u15491 (K8qow6, n4268);  // ../RTL/cortexm0ds_logic.v(13264)
  AL_MUX u15492 (
    .i0(Rw8iu6),
    .i1(Hrfpw6[14]),
    .sel(Qqhiu6),
    .o(Fbohu6));  // ../RTL/cortexm0ds_logic.v(13265)
  and u15493 (n4269, Dxfhu6, HREADY);  // ../RTL/cortexm0ds_logic.v(13266)
  not u15494 (Qqhiu6, n4269);  // ../RTL/cortexm0ds_logic.v(13266)
  and u15495 (n4270, Hs7iu6, Y8qow6);  // ../RTL/cortexm0ds_logic.v(13267)
  not u15496 (Rw8iu6, n4270);  // ../RTL/cortexm0ds_logic.v(13267)
  and u15497 (n4271, HRDATA[30], Vobiu6);  // ../RTL/cortexm0ds_logic.v(13268)
  not u15498 (Y8qow6, n4271);  // ../RTL/cortexm0ds_logic.v(13268)
  or u15499 (n4272, F9qow6, N19iu6);  // ../RTL/cortexm0ds_logic.v(13269)
  buf u155 (Uthpw6[10], Gyxpw6);  // ../RTL/cortexm0ds_logic.v(1882)
  and u1550 (Ct0iu6, vis_apsr_o[1], Jt0iu6);  // ../RTL/cortexm0ds_logic.v(3491)
  not u15500 (Vobiu6, n4272);  // ../RTL/cortexm0ds_logic.v(13269)
  not u15501 (N19iu6, vis_tbit_o);  // ../RTL/cortexm0ds_logic.v(13270)
  or u15502 (F9qow6, V3xhu6, Yyfhu6);  // ../RTL/cortexm0ds_logic.v(13271)
  and u15503 (V3xhu6, HRESP, Qaxiu6);  // ../RTL/cortexm0ds_logic.v(13272)
  not u15504 (Hs7iu6, Aghhu6);  // ../RTL/cortexm0ds_logic.v(13273)
  and u15505 (n4273, Kaohu6, M9qow6);  // ../RTL/cortexm0ds_logic.v(13274)
  not u15506 (Yaohu6, n4273);  // ../RTL/cortexm0ds_logic.v(13274)
  and u15507 (n4274, T9qow6, G3eiu6);  // ../RTL/cortexm0ds_logic.v(13275)
  not u15508 (M9qow6, n4274);  // ../RTL/cortexm0ds_logic.v(13275)
  and u15509 (G3eiu6, Npdhu6, HWDATA[2]);  // ../RTL/cortexm0ds_logic.v(13276)
  and u1551 (n122, Qt0iu6, Xt0iu6);  // ../RTL/cortexm0ds_logic.v(3492)
  and u15510 (T9qow6, Uzhiu6, Nzhiu6);  // ../RTL/cortexm0ds_logic.v(13277)
  buf u15511 (Bklhu6, Nvkbx6[30]);  // ../RTL/cortexm0ds_logic.v(3137)
  and u15512 (Nzhiu6, Cznow6, K5eiu6);  // ../RTL/cortexm0ds_logic.v(13279)
  not u15513 (Yreow6, Nzhiu6);  // ../RTL/cortexm0ds_logic.v(13279)
  and u15514 (K5eiu6, Jfgpw6[1], Uh7iu6);  // ../RTL/cortexm0ds_logic.v(13280)
  not u15515 (Uh7iu6, Jfgpw6[0]);  // ../RTL/cortexm0ds_logic.v(13281)
  and u15516 (Cznow6, Aaqow6, Jfgpw6[3]);  // ../RTL/cortexm0ds_logic.v(13282)
  or u15517 (n4275, U89iu6, Jfgpw6[2]);  // ../RTL/cortexm0ds_logic.v(13283)
  not u15518 (Aaqow6, n4275);  // ../RTL/cortexm0ds_logic.v(13283)
  not u15519 (U89iu6, Jfgpw6[4]);  // ../RTL/cortexm0ds_logic.v(13284)
  not u1552 (Jt0iu6, n122);  // ../RTL/cortexm0ds_logic.v(3492)
  and u15520 (Uzhiu6, Haqow6, Oaqow6);  // ../RTL/cortexm0ds_logic.v(13285)
  and u15521 (Oaqow6, Vaqow6, Cbqow6);  // ../RTL/cortexm0ds_logic.v(13286)
  and u15522 (Cbqow6, Jbqow6, Qbqow6);  // ../RTL/cortexm0ds_logic.v(13287)
  or u15523 (n4276, HWDATA[29], HWDATA[16]);  // ../RTL/cortexm0ds_logic.v(13288)
  not u15524 (Qbqow6, n4276);  // ../RTL/cortexm0ds_logic.v(13288)
  and u15525 (n4278, Lcqow6, L35ju6);  // ../RTL/cortexm0ds_logic.v(13290)
  not u15526 (Ecqow6, n4278);  // ../RTL/cortexm0ds_logic.v(13290)
  and u15527 (Xbqow6, Scqow6, Zcqow6);  // ../RTL/cortexm0ds_logic.v(13291)
  and u15528 (n4279, Gdqow6, Xc9ju6);  // ../RTL/cortexm0ds_logic.v(13292)
  not u15529 (Zcqow6, n4279);  // ../RTL/cortexm0ds_logic.v(13292)
  or u1553 (Xt0iu6, Eu0iu6, Cyfpw6[7]);  // ../RTL/cortexm0ds_logic.v(3493)
  and u15530 (n4280, Ndqow6, Udqow6);  // ../RTL/cortexm0ds_logic.v(13293)
  not u15531 (Xc9ju6, n4280);  // ../RTL/cortexm0ds_logic.v(13293)
  and u15532 (Udqow6, Beqow6, Ieqow6);  // ../RTL/cortexm0ds_logic.v(13294)
  and u15533 (Ieqow6, Peqow6, Weqow6);  // ../RTL/cortexm0ds_logic.v(13295)
  and u15534 (n4281, Fkfpw6[16], Dfqow6);  // ../RTL/cortexm0ds_logic.v(13296)
  not u15535 (Weqow6, n4281);  // ../RTL/cortexm0ds_logic.v(13296)
  and u15536 (Peqow6, Kfqow6, Rfqow6);  // ../RTL/cortexm0ds_logic.v(13297)
  and u15537 (n4282, vis_psp_o[14], Yfqow6);  // ../RTL/cortexm0ds_logic.v(13298)
  not u15538 (Rfqow6, n4282);  // ../RTL/cortexm0ds_logic.v(13298)
  and u15539 (n4283, vis_msp_o[14], Fgqow6);  // ../RTL/cortexm0ds_logic.v(13299)
  or u1554 (Qt0iu6, Mr0iu6, Cyfpw6[3]);  // ../RTL/cortexm0ds_logic.v(3494)
  not u15540 (Kfqow6, n4283);  // ../RTL/cortexm0ds_logic.v(13299)
  and u15541 (Beqow6, Mgqow6, Tgqow6);  // ../RTL/cortexm0ds_logic.v(13300)
  and u15542 (n4284, vis_r14_o[16], Ahqow6);  // ../RTL/cortexm0ds_logic.v(13301)
  not u15543 (Tgqow6, n4284);  // ../RTL/cortexm0ds_logic.v(13301)
  and u15544 (n4285, vis_r12_o[16], Hhqow6);  // ../RTL/cortexm0ds_logic.v(13302)
  not u15545 (Mgqow6, n4285);  // ../RTL/cortexm0ds_logic.v(13302)
  and u15546 (Ndqow6, Ohqow6, Vhqow6);  // ../RTL/cortexm0ds_logic.v(13303)
  and u15547 (Vhqow6, Ciqow6, Jiqow6);  // ../RTL/cortexm0ds_logic.v(13304)
  and u15548 (n4286, vis_r9_o[16], Qiqow6);  // ../RTL/cortexm0ds_logic.v(13305)
  not u15549 (Jiqow6, n4286);  // ../RTL/cortexm0ds_logic.v(13305)
  and u1555 (Uo0iu6, Lu0iu6, Su0iu6);  // ../RTL/cortexm0ds_logic.v(3495)
  and u15550 (Ciqow6, Xiqow6, Ejqow6);  // ../RTL/cortexm0ds_logic.v(13306)
  and u15551 (n4287, vis_r11_o[16], Ljqow6);  // ../RTL/cortexm0ds_logic.v(13307)
  not u15552 (Ejqow6, n4287);  // ../RTL/cortexm0ds_logic.v(13307)
  and u15553 (n4288, vis_r10_o[16], Sjqow6);  // ../RTL/cortexm0ds_logic.v(13308)
  not u15554 (Xiqow6, n4288);  // ../RTL/cortexm0ds_logic.v(13308)
  and u15555 (Ohqow6, Q10iu6, Zjqow6);  // ../RTL/cortexm0ds_logic.v(13309)
  and u15556 (n4289, vis_r8_o[16], Gkqow6);  // ../RTL/cortexm0ds_logic.v(13310)
  not u15557 (Zjqow6, n4289);  // ../RTL/cortexm0ds_logic.v(13310)
  and u15558 (Q10iu6, Nkqow6, Ukqow6);  // ../RTL/cortexm0ds_logic.v(13311)
  and u15559 (Ukqow6, Blqow6, Ilqow6);  // ../RTL/cortexm0ds_logic.v(13312)
  or u1556 (Su0iu6, Zu0iu6, Cyfpw6[4]);  // ../RTL/cortexm0ds_logic.v(3496)
  and u15560 (Ilqow6, Plqow6, Wlqow6);  // ../RTL/cortexm0ds_logic.v(13313)
  and u15561 (n4290, vis_r2_o[16], Dmqow6);  // ../RTL/cortexm0ds_logic.v(13314)
  not u15562 (Wlqow6, n4290);  // ../RTL/cortexm0ds_logic.v(13314)
  and u15563 (n4291, vis_r6_o[16], Kmqow6);  // ../RTL/cortexm0ds_logic.v(13315)
  not u15564 (Plqow6, n4291);  // ../RTL/cortexm0ds_logic.v(13315)
  and u15565 (Blqow6, Rmqow6, Ymqow6);  // ../RTL/cortexm0ds_logic.v(13316)
  and u15566 (n4292, vis_r5_o[16], Fnqow6);  // ../RTL/cortexm0ds_logic.v(13317)
  not u15567 (Ymqow6, n4292);  // ../RTL/cortexm0ds_logic.v(13317)
  and u15568 (n4293, vis_r4_o[16], Mnqow6);  // ../RTL/cortexm0ds_logic.v(13318)
  not u15569 (Rmqow6, n4293);  // ../RTL/cortexm0ds_logic.v(13318)
  and u1557 (Eblhu6, Gv0iu6, Rrlhu6);  // ../RTL/cortexm0ds_logic.v(3497)
  and u15570 (Nkqow6, Tnqow6, Aoqow6);  // ../RTL/cortexm0ds_logic.v(13319)
  and u15571 (Aoqow6, Hoqow6, Ooqow6);  // ../RTL/cortexm0ds_logic.v(13320)
  and u15572 (n4294, vis_r1_o[16], Voqow6);  // ../RTL/cortexm0ds_logic.v(13321)
  not u15573 (Ooqow6, n4294);  // ../RTL/cortexm0ds_logic.v(13321)
  and u15574 (n4295, vis_r0_o[16], Cpqow6);  // ../RTL/cortexm0ds_logic.v(13322)
  not u15575 (Hoqow6, n4295);  // ../RTL/cortexm0ds_logic.v(13322)
  and u15576 (Tnqow6, Jpqow6, Qpqow6);  // ../RTL/cortexm0ds_logic.v(13323)
  and u15577 (n4296, vis_r3_o[16], Xpqow6);  // ../RTL/cortexm0ds_logic.v(13324)
  not u15578 (Qpqow6, n4296);  // ../RTL/cortexm0ds_logic.v(13324)
  and u15579 (n4297, vis_r7_o[16], Eqqow6);  // ../RTL/cortexm0ds_logic.v(13325)
  AL_MUX u1558 (
    .i0(vis_pc_o[23]),
    .i1(Tzdpw6),
    .sel(Nv0iu6),
    .o(Gv0iu6));  // ../RTL/cortexm0ds_logic.v(3498)
  not u15580 (Jpqow6, n4297);  // ../RTL/cortexm0ds_logic.v(13325)
  and u15581 (n4298, Z54iu6, R0nhu6);  // ../RTL/cortexm0ds_logic.v(13326)
  not u15582 (Scqow6, n4298);  // ../RTL/cortexm0ds_logic.v(13326)
  and u15583 (Z54iu6, Shhpw6[16], Iqzhu6);  // ../RTL/cortexm0ds_logic.v(13327)
  and u15584 (Sqqow6, Zqqow6, Grqow6);  // ../RTL/cortexm0ds_logic.v(13329)
  and u15585 (n4299, Gdqow6, Wh8iu6);  // ../RTL/cortexm0ds_logic.v(13330)
  not u15586 (Grqow6, n4299);  // ../RTL/cortexm0ds_logic.v(13330)
  and u15587 (n4300, Nrqow6, Urqow6);  // ../RTL/cortexm0ds_logic.v(13331)
  not u15588 (Wh8iu6, n4300);  // ../RTL/cortexm0ds_logic.v(13331)
  and u15589 (Urqow6, Bsqow6, Isqow6);  // ../RTL/cortexm0ds_logic.v(13332)
  and u1559 (Lclhu6, Uv0iu6, Kqlhu6);  // ../RTL/cortexm0ds_logic.v(3499)
  and u15590 (Isqow6, Psqow6, Wsqow6);  // ../RTL/cortexm0ds_logic.v(13333)
  and u15591 (n4301, vis_r11_o[29], Ljqow6);  // ../RTL/cortexm0ds_logic.v(13334)
  not u15592 (Wsqow6, n4301);  // ../RTL/cortexm0ds_logic.v(13334)
  and u15593 (Psqow6, Dtqow6, Ktqow6);  // ../RTL/cortexm0ds_logic.v(13335)
  and u15594 (n4302, vis_r9_o[29], Qiqow6);  // ../RTL/cortexm0ds_logic.v(13336)
  not u15595 (Ktqow6, n4302);  // ../RTL/cortexm0ds_logic.v(13336)
  and u15596 (n4303, Fkfpw6[29], Dfqow6);  // ../RTL/cortexm0ds_logic.v(13337)
  not u15597 (Dtqow6, n4303);  // ../RTL/cortexm0ds_logic.v(13337)
  and u15598 (Bsqow6, Rtqow6, Ytqow6);  // ../RTL/cortexm0ds_logic.v(13338)
  and u15599 (n4304, vis_r10_o[29], Sjqow6);  // ../RTL/cortexm0ds_logic.v(13339)
  buf u156 (V5hpw6[1], Hz9ax6);  // ../RTL/cortexm0ds_logic.v(2248)
  AL_MUX u1560 (
    .i0(vis_pc_o[24]),
    .i1(A0epw6),
    .sel(Nv0iu6),
    .o(Uv0iu6));  // ../RTL/cortexm0ds_logic.v(3500)
  not u15600 (Ytqow6, n4304);  // ../RTL/cortexm0ds_logic.v(13339)
  and u15601 (n4305, vis_psp_o[27], Yfqow6);  // ../RTL/cortexm0ds_logic.v(13340)
  not u15602 (Rtqow6, n4305);  // ../RTL/cortexm0ds_logic.v(13340)
  and u15603 (Nrqow6, Fuqow6, Muqow6);  // ../RTL/cortexm0ds_logic.v(13341)
  and u15604 (Muqow6, Tuqow6, Avqow6);  // ../RTL/cortexm0ds_logic.v(13342)
  and u15605 (n4306, vis_r12_o[29], Hhqow6);  // ../RTL/cortexm0ds_logic.v(13343)
  not u15606 (Avqow6, n4306);  // ../RTL/cortexm0ds_logic.v(13343)
  and u15607 (Tuqow6, Hvqow6, Ovqow6);  // ../RTL/cortexm0ds_logic.v(13344)
  and u15608 (n4307, vis_msp_o[27], Fgqow6);  // ../RTL/cortexm0ds_logic.v(13345)
  not u15609 (Ovqow6, n4307);  // ../RTL/cortexm0ds_logic.v(13345)
  and u1561 (Sdlhu6, Bw0iu6, Dplhu6);  // ../RTL/cortexm0ds_logic.v(3501)
  and u15610 (n4308, vis_r14_o[29], Ahqow6);  // ../RTL/cortexm0ds_logic.v(13346)
  not u15611 (Hvqow6, n4308);  // ../RTL/cortexm0ds_logic.v(13346)
  and u15612 (Fuqow6, Wxzhu6, Vvqow6);  // ../RTL/cortexm0ds_logic.v(13347)
  and u15613 (n4309, vis_r8_o[29], Gkqow6);  // ../RTL/cortexm0ds_logic.v(13348)
  not u15614 (Vvqow6, n4309);  // ../RTL/cortexm0ds_logic.v(13348)
  and u15615 (Wxzhu6, Cwqow6, Jwqow6);  // ../RTL/cortexm0ds_logic.v(13349)
  and u15616 (Jwqow6, Qwqow6, Xwqow6);  // ../RTL/cortexm0ds_logic.v(13350)
  and u15617 (Xwqow6, Exqow6, Lxqow6);  // ../RTL/cortexm0ds_logic.v(13351)
  and u15618 (n4310, vis_r2_o[29], Dmqow6);  // ../RTL/cortexm0ds_logic.v(13352)
  not u15619 (Lxqow6, n4310);  // ../RTL/cortexm0ds_logic.v(13352)
  AL_MUX u1562 (
    .i0(vis_pc_o[25]),
    .i1(H0epw6),
    .sel(Nv0iu6),
    .o(Bw0iu6));  // ../RTL/cortexm0ds_logic.v(3502)
  and u15620 (n4311, vis_r6_o[29], Kmqow6);  // ../RTL/cortexm0ds_logic.v(13353)
  not u15621 (Exqow6, n4311);  // ../RTL/cortexm0ds_logic.v(13353)
  and u15622 (Qwqow6, Sxqow6, Zxqow6);  // ../RTL/cortexm0ds_logic.v(13354)
  and u15623 (n4312, vis_r5_o[29], Fnqow6);  // ../RTL/cortexm0ds_logic.v(13355)
  not u15624 (Zxqow6, n4312);  // ../RTL/cortexm0ds_logic.v(13355)
  and u15625 (n4313, vis_r4_o[29], Mnqow6);  // ../RTL/cortexm0ds_logic.v(13356)
  not u15626 (Sxqow6, n4313);  // ../RTL/cortexm0ds_logic.v(13356)
  and u15627 (Cwqow6, Gyqow6, Nyqow6);  // ../RTL/cortexm0ds_logic.v(13357)
  and u15628 (Nyqow6, Uyqow6, Bzqow6);  // ../RTL/cortexm0ds_logic.v(13358)
  and u15629 (n4314, vis_r1_o[29], Voqow6);  // ../RTL/cortexm0ds_logic.v(13359)
  and u1563 (Zelhu6, Iw0iu6, Wnlhu6);  // ../RTL/cortexm0ds_logic.v(3503)
  not u15630 (Bzqow6, n4314);  // ../RTL/cortexm0ds_logic.v(13359)
  and u15631 (n4315, vis_r0_o[29], Cpqow6);  // ../RTL/cortexm0ds_logic.v(13360)
  not u15632 (Uyqow6, n4315);  // ../RTL/cortexm0ds_logic.v(13360)
  and u15633 (Gyqow6, Izqow6, Pzqow6);  // ../RTL/cortexm0ds_logic.v(13361)
  and u15634 (n4316, vis_r3_o[29], Xpqow6);  // ../RTL/cortexm0ds_logic.v(13362)
  not u15635 (Pzqow6, n4316);  // ../RTL/cortexm0ds_logic.v(13362)
  and u15636 (n4317, vis_r7_o[29], Eqqow6);  // ../RTL/cortexm0ds_logic.v(13363)
  not u15637 (Izqow6, n4317);  // ../RTL/cortexm0ds_logic.v(13363)
  and u15638 (Lqqow6, Wzqow6, D0row6);  // ../RTL/cortexm0ds_logic.v(13364)
  and u15639 (n4318, K0row6, Sz8ju6);  // ../RTL/cortexm0ds_logic.v(13365)
  AL_MUX u1564 (
    .i0(vis_pc_o[26]),
    .i1(O0epw6),
    .sel(Nv0iu6),
    .o(Iw0iu6));  // ../RTL/cortexm0ds_logic.v(3504)
  not u15640 (D0row6, n4318);  // ../RTL/cortexm0ds_logic.v(13365)
  and u15641 (n4319, M94iu6, R0nhu6);  // ../RTL/cortexm0ds_logic.v(13366)
  not u15642 (Wzqow6, n4319);  // ../RTL/cortexm0ds_logic.v(13366)
  and u15643 (M94iu6, Shhpw6[29], Iqzhu6);  // ../RTL/cortexm0ds_logic.v(13367)
  or u15644 (n4320, HWDATA[30], HWDATA[31]);  // ../RTL/cortexm0ds_logic.v(13368)
  not u15645 (Jbqow6, n4320);  // ../RTL/cortexm0ds_logic.v(13368)
  and u15646 (Vaqow6, R0row6, Y0row6);  // ../RTL/cortexm0ds_logic.v(13369)
  or u15647 (n4321, HWDATA[27], HWDATA[28]);  // ../RTL/cortexm0ds_logic.v(13370)
  not u15648 (Y0row6, n4321);  // ../RTL/cortexm0ds_logic.v(13370)
  or u15649 (n4322, HWDATA[18], HWDATA[25]);  // ../RTL/cortexm0ds_logic.v(13371)
  and u1565 (Gglhu6, Pw0iu6, Pmlhu6);  // ../RTL/cortexm0ds_logic.v(3505)
  not u15650 (R0row6, n4322);  // ../RTL/cortexm0ds_logic.v(13371)
  and u15651 (Haqow6, F1row6, M1row6);  // ../RTL/cortexm0ds_logic.v(13372)
  and u15652 (M1row6, T1row6, A2row6);  // ../RTL/cortexm0ds_logic.v(13373)
  and u15653 (A2row6, HWDATA[24], HWDATA[26]);  // ../RTL/cortexm0ds_logic.v(13374)
  and u15654 (T1row6, HWDATA[22], HWDATA[23]);  // ../RTL/cortexm0ds_logic.v(13375)
  and u15655 (F1row6, H2row6, O2row6);  // ../RTL/cortexm0ds_logic.v(13376)
  and u15656 (O2row6, HWDATA[20], HWDATA[21]);  // ../RTL/cortexm0ds_logic.v(13377)
  and u15657 (H2row6, HWDATA[17], HWDATA[19]);  // ../RTL/cortexm0ds_logic.v(13378)
  AL_MUX u15658 (
    .i0(V2row6),
    .i1(Qnghu6),
    .sel(Eh6iu6),
    .o(Raohu6));  // ../RTL/cortexm0ds_logic.v(13379)
  not u15659 (Eh6iu6, HREADY);  // ../RTL/cortexm0ds_logic.v(13380)
  AL_MUX u1566 (
    .i0(vis_pc_o[27]),
    .i1(V0epw6),
    .sel(Nv0iu6),
    .o(Pw0iu6));  // ../RTL/cortexm0ds_logic.v(3506)
  and u15660 (V2row6, C3row6, J3row6);  // ../RTL/cortexm0ds_logic.v(13381)
  and u15661 (J3row6, Q3row6, Udpiu6);  // ../RTL/cortexm0ds_logic.v(13382)
  not u15662 (Udpiu6, Pzwiu6);  // ../RTL/cortexm0ds_logic.v(13383)
  and u15663 (n4323, Stdhu6, Gsaiu6);  // ../RTL/cortexm0ds_logic.v(13384)
  not u15664 (Q3row6, n4323);  // ../RTL/cortexm0ds_logic.v(13384)
  and u15665 (n4324, Xe9ow6, X3row6);  // ../RTL/cortexm0ds_logic.v(13385)
  not u15666 (Gsaiu6, n4324);  // ../RTL/cortexm0ds_logic.v(13385)
  and u15667 (n4325, E4row6, Y2oiu6);  // ../RTL/cortexm0ds_logic.v(13386)
  not u15668 (X3row6, n4325);  // ../RTL/cortexm0ds_logic.v(13386)
  or u15669 (E4row6, Iugiu6, P8oiu6);  // ../RTL/cortexm0ds_logic.v(13387)
  and u1567 (Nhlhu6, Ww0iu6, Illhu6);  // ../RTL/cortexm0ds_logic.v(3507)
  or u15670 (n4326, Et0ju6, Xe8iu6);  // ../RTL/cortexm0ds_logic.v(13388)
  not u15671 (P8oiu6, n4326);  // ../RTL/cortexm0ds_logic.v(13388)
  or u15672 (Et0ju6, Nlaiu6, K9aiu6);  // ../RTL/cortexm0ds_logic.v(13389)
  and u15673 (C3row6, U6piu6, Usaiu6);  // ../RTL/cortexm0ds_logic.v(13390)
  or u15674 (n4327, Qa5iu6, L4row6);  // ../RTL/cortexm0ds_logic.v(13391)
  not u15675 (Usaiu6, n4327);  // ../RTL/cortexm0ds_logic.v(13391)
  and u15676 (L4row6, Fsdhu6, Ja5iu6);  // ../RTL/cortexm0ds_logic.v(13392)
  and u15677 (Ja5iu6, S4row6, Sf7ju6);  // ../RTL/cortexm0ds_logic.v(13393)
  and u15678 (Sf7ju6, Z4row6, F23ju6);  // ../RTL/cortexm0ds_logic.v(13394)
  or u15679 (n4328, As0iu6, H4ghu6);  // ../RTL/cortexm0ds_logic.v(13395)
  AL_MUX u1568 (
    .i0(vis_pc_o[28]),
    .i1(Dx0iu6),
    .sel(Nv0iu6),
    .o(Ww0iu6));  // ../RTL/cortexm0ds_logic.v(3508)
  not u15680 (Z4row6, n4328);  // ../RTL/cortexm0ds_logic.v(13395)
  and u15681 (S4row6, Pt2ju6, Cyfpw6[3]);  // ../RTL/cortexm0ds_logic.v(13396)
  and u15682 (Qa5iu6, Su8ow6, Xe9ow6);  // ../RTL/cortexm0ds_logic.v(13397)
  and u15683 (n4329, Iepiu6, Cyfpw6[5]);  // ../RTL/cortexm0ds_logic.v(13398)
  not u15684 (Xe9ow6, n4329);  // ../RTL/cortexm0ds_logic.v(13398)
  and u15685 (n4330, Vo3ju6, G5row6);  // ../RTL/cortexm0ds_logic.v(13399)
  not u15686 (Su8ow6, n4330);  // ../RTL/cortexm0ds_logic.v(13399)
  and u15687 (n4331, N5row6, U5row6);  // ../RTL/cortexm0ds_logic.v(13400)
  not u15688 (G5row6, n4331);  // ../RTL/cortexm0ds_logic.v(13400)
  and u15689 (n4332, B6row6, X97ow6);  // ../RTL/cortexm0ds_logic.v(13401)
  and u1569 (Uilhu6, Kx0iu6, Bklhu6);  // ../RTL/cortexm0ds_logic.v(3509)
  not u15690 (U5row6, n4332);  // ../RTL/cortexm0ds_logic.v(13401)
  and u15691 (B6row6, Qe8iu6, Tfjiu6);  // ../RTL/cortexm0ds_logic.v(13402)
  and u15692 (n4333, N4kiu6, Hs0iu6);  // ../RTL/cortexm0ds_logic.v(13403)
  not u15693 (N5row6, n4333);  // ../RTL/cortexm0ds_logic.v(13403)
  and u15694 (N4kiu6, I6row6, Frziu6);  // ../RTL/cortexm0ds_logic.v(13404)
  or u15695 (n4334, Ae0iu6, C0ehu6);  // ../RTL/cortexm0ds_logic.v(13405)
  not u15696 (I6row6, n4334);  // ../RTL/cortexm0ds_logic.v(13405)
  and u15697 (U6piu6, P6row6, Zl1ju6);  // ../RTL/cortexm0ds_logic.v(13406)
  and u15698 (n4335, Emfiu6, W6row6);  // ../RTL/cortexm0ds_logic.v(13407)
  not u15699 (Zl1ju6, n4335);  // ../RTL/cortexm0ds_logic.v(13407)
  buf u157 (vis_r0_o[28], Ednpw6);  // ../RTL/cortexm0ds_logic.v(1875)
  AL_MUX u1570 (
    .i0(vis_pc_o[29]),
    .i1(Rx0iu6),
    .sel(Nv0iu6),
    .o(Kx0iu6));  // ../RTL/cortexm0ds_logic.v(3510)
  and u15700 (n4336, D7row6, Te6iu6);  // ../RTL/cortexm0ds_logic.v(13408)
  not u15701 (W6row6, n4336);  // ../RTL/cortexm0ds_logic.v(13408)
  not u15702 (Te6iu6, Ahghu6);  // ../RTL/cortexm0ds_logic.v(13409)
  or u15703 (D7row6, X7gow6, M2biu6);  // ../RTL/cortexm0ds_logic.v(13410)
  not u15704 (X7gow6, Righu6);  // ../RTL/cortexm0ds_logic.v(13411)
  or u15705 (P6row6, K7row6, Sl1ju6);  // ../RTL/cortexm0ds_logic.v(13412)
  and u15706 (n4337, R7row6, Knbow6);  // ../RTL/cortexm0ds_logic.v(13413)
  not u15707 (Sl1ju6, n4337);  // ../RTL/cortexm0ds_logic.v(13413)
  and u15708 (Knbow6, Emfiu6, Y7row6);  // ../RTL/cortexm0ds_logic.v(13414)
  not u15709 (Y7row6, M2biu6);  // ../RTL/cortexm0ds_logic.v(13415)
  or u1571 (Knmhu6, Yx0iu6, G4hpw6[0]);  // ../RTL/cortexm0ds_logic.v(3511)
  and u15710 (M2biu6, F8row6, M8row6);  // ../RTL/cortexm0ds_logic.v(13416)
  and u15711 (Zmfiu6, T8row6, A9row6);  // ../RTL/cortexm0ds_logic.v(13417)
  not u15712 (Emfiu6, Zmfiu6);  // ../RTL/cortexm0ds_logic.v(13417)
  and u15713 (T8row6, H9row6, M8row6);  // ../RTL/cortexm0ds_logic.v(13418)
  and u15714 (R7row6, O9row6, V0fow6);  // ../RTL/cortexm0ds_logic.v(13419)
  or u15715 (V0fow6, V9row6, Carow6);  // ../RTL/cortexm0ds_logic.v(13420)
  and u15716 (n4338, Jarow6, Qarow6);  // ../RTL/cortexm0ds_logic.v(13421)
  not u15717 (V9row6, n4338);  // ../RTL/cortexm0ds_logic.v(13421)
  and u15718 (n4339, Ikghu6, Jhqiu6);  // ../RTL/cortexm0ds_logic.v(13422)
  not u15719 (Jarow6, n4339);  // ../RTL/cortexm0ds_logic.v(13422)
  or u1572 (Romhu6, Yx0iu6, G4hpw6[1]);  // ../RTL/cortexm0ds_logic.v(3512)
  and u15720 (n4340, Xarow6, Ebrow6);  // ../RTL/cortexm0ds_logic.v(13423)
  not u15721 (O9row6, n4340);  // ../RTL/cortexm0ds_logic.v(13423)
  or u15722 (Ebrow6, Lbrow6, Sbrow6);  // ../RTL/cortexm0ds_logic.v(13424)
  and u15723 (Xarow6, Zbrow6, Gcrow6);  // ../RTL/cortexm0ds_logic.v(13425)
  and u15724 (n4341, Ncrow6, Ucrow6);  // ../RTL/cortexm0ds_logic.v(13426)
  not u15725 (Zbrow6, n4341);  // ../RTL/cortexm0ds_logic.v(13426)
  and u15726 (Ucrow6, Bdrow6, Idrow6);  // ../RTL/cortexm0ds_logic.v(13427)
  or u15727 (Bdrow6, Okgow6, Pdrow6);  // ../RTL/cortexm0ds_logic.v(13428)
  not u15728 (Pdrow6, L1gpw6[0]);  // ../RTL/cortexm0ds_logic.v(13429)
  or u15729 (Okgow6, A8low6, Wdrow6);  // ../RTL/cortexm0ds_logic.v(13430)
  or u1573 (Ypmhu6, Yx0iu6, G4hpw6[2]);  // ../RTL/cortexm0ds_logic.v(3513)
  or u15730 (n4342, Derow6, Kerow6);  // ../RTL/cortexm0ds_logic.v(13431)
  not u15731 (Ncrow6, n4342);  // ../RTL/cortexm0ds_logic.v(13431)
  and u15732 (Kerow6, Sbrow6, Lbrow6);  // ../RTL/cortexm0ds_logic.v(13432)
  AL_MUX u15733 (
    .i0(Rerow6),
    .i1(Yerow6),
    .sel(A8low6),
    .o(Lbrow6));  // ../RTL/cortexm0ds_logic.v(13433)
  AL_MUX u15734 (
    .i0(Ffrow6),
    .i1(Mfrow6),
    .sel(A8low6),
    .o(Derow6));  // ../RTL/cortexm0ds_logic.v(13434)
  and u15735 (n4343, Tfrow6, Agrow6);  // ../RTL/cortexm0ds_logic.v(13435)
  not u15736 (A8low6, n4343);  // ../RTL/cortexm0ds_logic.v(13435)
  and u15737 (n4344, Carow6, Hgrow6);  // ../RTL/cortexm0ds_logic.v(13436)
  not u15738 (Agrow6, n4344);  // ../RTL/cortexm0ds_logic.v(13436)
  and u15739 (n4345, Ogrow6, Vgrow6);  // ../RTL/cortexm0ds_logic.v(13437)
  or u1574 (Frmhu6, Yx0iu6, G4hpw6[3]);  // ../RTL/cortexm0ds_logic.v(3514)
  not u15740 (Hgrow6, n4345);  // ../RTL/cortexm0ds_logic.v(13437)
  and u15741 (n4346, Chrow6, Jhrow6);  // ../RTL/cortexm0ds_logic.v(13438)
  not u15742 (Vgrow6, n4346);  // ../RTL/cortexm0ds_logic.v(13438)
  AL_MUX u15743 (
    .i0(B3gpw6[0]),
    .i1(L1gpw6[0]),
    .sel(Qarow6),
    .o(Jhrow6));  // ../RTL/cortexm0ds_logic.v(13439)
  or u15744 (n4347, Mfrow6, Qhrow6);  // ../RTL/cortexm0ds_logic.v(13440)
  not u15745 (Chrow6, n4347);  // ../RTL/cortexm0ds_logic.v(13440)
  or u15746 (n4348, Rerow6, Xhrow6);  // ../RTL/cortexm0ds_logic.v(13441)
  not u15747 (Qhrow6, n4348);  // ../RTL/cortexm0ds_logic.v(13441)
  and u15748 (n4349, Xhrow6, Rerow6);  // ../RTL/cortexm0ds_logic.v(13442)
  not u15749 (Ogrow6, n4349);  // ../RTL/cortexm0ds_logic.v(13442)
  and u1575 (Gwhhu6, Fy0iu6, A4khu6);  // ../RTL/cortexm0ds_logic.v(3515)
  AL_MUX u15750 (
    .i0(L1gpw6[1]),
    .i1(B3gpw6[1]),
    .sel(Wdrow6),
    .o(Rerow6));  // ../RTL/cortexm0ds_logic.v(13443)
  not u15751 (Xhrow6, Yerow6);  // ../RTL/cortexm0ds_logic.v(13444)
  AL_MUX u15752 (
    .i0(H8gpw6[1]),
    .i1(Eirow6),
    .sel(O8low6),
    .o(Yerow6));  // ../RTL/cortexm0ds_logic.v(13445)
  and u15753 (n4350, O8low6, Lirow6);  // ../RTL/cortexm0ds_logic.v(13446)
  not u15754 (Carow6, n4350);  // ../RTL/cortexm0ds_logic.v(13446)
  and u15755 (n4351, Sirow6, Jhqiu6);  // ../RTL/cortexm0ds_logic.v(13447)
  not u15756 (Lirow6, n4351);  // ../RTL/cortexm0ds_logic.v(13447)
  or u15757 (Tfrow6, Ikghu6, Wdrow6);  // ../RTL/cortexm0ds_logic.v(13448)
  buf u15758 (Illhu6, Nvkbx6[29]);  // ../RTL/cortexm0ds_logic.v(3137)
  AL_MUX u15759 (
    .i0(H8gpw6[0]),
    .i1(Zirow6),
    .sel(O8low6),
    .o(Mfrow6));  // ../RTL/cortexm0ds_logic.v(13450)
  and u1576 (Fy0iu6, My0iu6, Ty0iu6);  // ../RTL/cortexm0ds_logic.v(3516)
  and u15760 (n4352, Gjrow6, Yyghu6);  // ../RTL/cortexm0ds_logic.v(13451)
  not u15761 (O8low6, n4352);  // ../RTL/cortexm0ds_logic.v(13451)
  and u15762 (Gjrow6, Njrow6, Jhqiu6);  // ../RTL/cortexm0ds_logic.v(13452)
  and u15763 (n4353, Sirow6, Ujrow6);  // ../RTL/cortexm0ds_logic.v(13453)
  not u15764 (Njrow6, n4353);  // ../RTL/cortexm0ds_logic.v(13453)
  and u15765 (n4354, Bkrow6, Ikrow6);  // ../RTL/cortexm0ds_logic.v(13454)
  not u15766 (Ujrow6, n4354);  // ../RTL/cortexm0ds_logic.v(13454)
  or u15767 (Ikrow6, Pkrow6, Zirow6);  // ../RTL/cortexm0ds_logic.v(13455)
  and u15768 (n4355, H8gpw6[0], Wkrow6);  // ../RTL/cortexm0ds_logic.v(13456)
  not u15769 (Pkrow6, n4355);  // ../RTL/cortexm0ds_logic.v(13456)
  and u1577 (Oxhhu6, Az0iu6, S2khu6);  // ../RTL/cortexm0ds_logic.v(3517)
  or u15770 (Wkrow6, Dlrow6, H8gpw6[1]);  // ../RTL/cortexm0ds_logic.v(13457)
  and u15771 (n4356, H8gpw6[1], Dlrow6);  // ../RTL/cortexm0ds_logic.v(13458)
  not u15772 (Bkrow6, n4356);  // ../RTL/cortexm0ds_logic.v(13458)
  not u15773 (Dlrow6, Eirow6);  // ../RTL/cortexm0ds_logic.v(13459)
  AL_MUX u15774 (
    .i0(Klrow6),
    .i1(Rlrow6),
    .sel(E2fow6),
    .o(Eirow6));  // ../RTL/cortexm0ds_logic.v(13460)
  not u15775 (Klrow6, Ylrow6);  // ../RTL/cortexm0ds_logic.v(13461)
  and u15776 (n4357, Fmrow6, Mmrow6);  // ../RTL/cortexm0ds_logic.v(13462)
  not u15777 (Sirow6, n4357);  // ../RTL/cortexm0ds_logic.v(13462)
  or u15778 (n4358, E2fow6, H7fow6);  // ../RTL/cortexm0ds_logic.v(13463)
  not u15779 (Mmrow6, n4358);  // ../RTL/cortexm0ds_logic.v(13463)
  AL_MUX u1578 (
    .i0(vis_pc_o[0]),
    .i1(Hz0iu6),
    .sel(Ty0iu6),
    .o(Az0iu6));  // ../RTL/cortexm0ds_logic.v(3518)
  buf u15780 (Pmlhu6, Nvkbx6[28]);  // ../RTL/cortexm0ds_logic.v(3137)
  and u15781 (Fmrow6, C8fow6, Tmrow6);  // ../RTL/cortexm0ds_logic.v(13465)
  AL_MUX u15782 (
    .i0(Anrow6),
    .i1(Hnrow6),
    .sel(Meeow6),
    .o(Zirow6));  // ../RTL/cortexm0ds_logic.v(13466)
  and u15783 (E2fow6, Onrow6, Vnrow6);  // ../RTL/cortexm0ds_logic.v(13467)
  not u15784 (Meeow6, E2fow6);  // ../RTL/cortexm0ds_logic.v(13467)
  and u15785 (n4359, Corow6, Jorow6);  // ../RTL/cortexm0ds_logic.v(13468)
  not u15786 (Vnrow6, n4359);  // ../RTL/cortexm0ds_logic.v(13468)
  or u15787 (Jorow6, Ylrow6, Rlrow6);  // ../RTL/cortexm0ds_logic.v(13469)
  and u15788 (Corow6, Qorow6, Xorow6);  // ../RTL/cortexm0ds_logic.v(13470)
  and u15789 (n4360, Eprow6, C8fow6);  // ../RTL/cortexm0ds_logic.v(13471)
  and u1579 (Wyhhu6, Oz0iu6, K1khu6);  // ../RTL/cortexm0ds_logic.v(3519)
  not u15790 (Xorow6, n4360);  // ../RTL/cortexm0ds_logic.v(13471)
  and u15791 (Eprow6, Tmrow6, Lprow6);  // ../RTL/cortexm0ds_logic.v(13472)
  and u15792 (n4361, Sprow6, Zprow6);  // ../RTL/cortexm0ds_logic.v(13473)
  not u15793 (Qorow6, n4361);  // ../RTL/cortexm0ds_logic.v(13473)
  and u15794 (n4362, Rlrow6, Ylrow6);  // ../RTL/cortexm0ds_logic.v(13474)
  not u15795 (Zprow6, n4362);  // ../RTL/cortexm0ds_logic.v(13474)
  AL_MUX u15796 (
    .i0(Gqrow6),
    .i1(Nqrow6),
    .sel(H7fow6),
    .o(Ylrow6));  // ../RTL/cortexm0ds_logic.v(13475)
  not u15797 (Nqrow6, Uqrow6);  // ../RTL/cortexm0ds_logic.v(13476)
  AL_MUX u15798 (
    .i0(Brrow6),
    .i1(Irrow6),
    .sel(B4fow6),
    .o(Rlrow6));  // ../RTL/cortexm0ds_logic.v(13477)
  not u15799 (Brrow6, Prrow6);  // ../RTL/cortexm0ds_logic.v(13478)
  buf u158 (Gtgpw6[11], Rz8bx6);  // ../RTL/cortexm0ds_logic.v(2375)
  AL_MUX u1580 (
    .i0(vis_pc_o[1]),
    .i1(Tugpw6[0]),
    .sel(Ty0iu6),
    .o(Oz0iu6));  // ../RTL/cortexm0ds_logic.v(3520)
  or u15800 (Sprow6, Hnrow6, Wrrow6);  // ../RTL/cortexm0ds_logic.v(13479)
  buf u15801 (Wnlhu6, Nvkbx6[27]);  // ../RTL/cortexm0ds_logic.v(3137)
  or u15802 (Onrow6, Dsrow6, B4fow6);  // ../RTL/cortexm0ds_logic.v(13481)
  or u15803 (Hnrow6, Ksrow6, Rsrow6);  // ../RTL/cortexm0ds_logic.v(13482)
  or u15804 (n4363, F6fow6, Ysrow6);  // ../RTL/cortexm0ds_logic.v(13483)
  not u15805 (Rsrow6, n4363);  // ../RTL/cortexm0ds_logic.v(13483)
  or u15806 (F6fow6, Lprow6, Ftrow6);  // ../RTL/cortexm0ds_logic.v(13484)
  AL_MUX u15807 (
    .i0(Mtrow6),
    .i1(Ttrow6),
    .sel(H7fow6),
    .o(Ksrow6));  // ../RTL/cortexm0ds_logic.v(13485)
  buf u15808 (Dplhu6, Nvkbx6[26]);  // ../RTL/cortexm0ds_logic.v(3137)
  and u15809 (H7fow6, Aurow6, Hurow6);  // ../RTL/cortexm0ds_logic.v(13487)
  and u1581 (E0ihu6, Vz0iu6, C0khu6);  // ../RTL/cortexm0ds_logic.v(3521)
  not u15810 (Lprow6, H7fow6);  // ../RTL/cortexm0ds_logic.v(13487)
  and u15811 (n4364, Ourow6, Vurow6);  // ../RTL/cortexm0ds_logic.v(13488)
  not u15812 (Hurow6, n4364);  // ../RTL/cortexm0ds_logic.v(13488)
  and u15813 (n4365, Cvrow6, Jvrow6);  // ../RTL/cortexm0ds_logic.v(13489)
  not u15814 (Vurow6, n4365);  // ../RTL/cortexm0ds_logic.v(13489)
  and u15815 (n4366, Uqrow6, Gqrow6);  // ../RTL/cortexm0ds_logic.v(13490)
  not u15816 (Jvrow6, n4366);  // ../RTL/cortexm0ds_logic.v(13490)
  and u15817 (n4367, Qvrow6, Xvrow6);  // ../RTL/cortexm0ds_logic.v(13491)
  not u15818 (Cvrow6, n4367);  // ../RTL/cortexm0ds_logic.v(13491)
  AL_MUX u15819 (
    .i0(Ewrow6),
    .i1(Lwrow6),
    .sel(O7fow6),
    .o(Xvrow6));  // ../RTL/cortexm0ds_logic.v(13492)
  AL_MUX u1582 (
    .i0(vis_pc_o[2]),
    .i1(Tugpw6[1]),
    .sel(Ty0iu6),
    .o(Vz0iu6));  // ../RTL/cortexm0ds_logic.v(3522)
  or u15820 (n4368, Mtrow6, Swrow6);  // ../RTL/cortexm0ds_logic.v(13493)
  not u15821 (Qvrow6, n4368);  // ../RTL/cortexm0ds_logic.v(13493)
  or u15822 (n4369, Gqrow6, Uqrow6);  // ../RTL/cortexm0ds_logic.v(13494)
  not u15823 (Swrow6, n4369);  // ../RTL/cortexm0ds_logic.v(13494)
  AL_MUX u15824 (
    .i0(Zwrow6),
    .i1(Gxrow6),
    .sel(Ftrow6),
    .o(Uqrow6));  // ../RTL/cortexm0ds_logic.v(13495)
  AL_MUX u15825 (
    .i0(Nxrow6),
    .i1(Uxrow6),
    .sel(Hdgow6),
    .o(Gqrow6));  // ../RTL/cortexm0ds_logic.v(13496)
  buf u15826 (Qlfhu6, Ozkbx6[3]);  // ../RTL/cortexm0ds_logic.v(3176)
  not u15827 (Ourow6, Fmrow6);  // ../RTL/cortexm0ds_logic.v(13497)
  and u15828 (C8fow6, Q8fow6, Jegow6);  // ../RTL/cortexm0ds_logic.v(13498)
  and u15829 (n4370, Byrow6, Iyrow6);  // ../RTL/cortexm0ds_logic.v(13499)
  and u1583 (M1ihu6, C01iu6, Uyjhu6);  // ../RTL/cortexm0ds_logic.v(3523)
  not u15830 (Aurow6, n4370);  // ../RTL/cortexm0ds_logic.v(13499)
  or u15831 (n4371, Pyrow6, Ftrow6);  // ../RTL/cortexm0ds_logic.v(13500)
  not u15832 (Byrow6, n4371);  // ../RTL/cortexm0ds_logic.v(13500)
  and u15833 (Ttrow6, Ftrow6, Ewrow6);  // ../RTL/cortexm0ds_logic.v(13501)
  buf u15834 (Kqlhu6, Nvkbx6[25]);  // ../RTL/cortexm0ds_logic.v(3137)
  and u15835 (Ftrow6, Wyrow6, Dzrow6);  // ../RTL/cortexm0ds_logic.v(13503)
  not u15836 (O7fow6, Ftrow6);  // ../RTL/cortexm0ds_logic.v(13503)
  and u15837 (n4372, Kzrow6, Rzrow6);  // ../RTL/cortexm0ds_logic.v(13504)
  not u15838 (Dzrow6, n4372);  // ../RTL/cortexm0ds_logic.v(13504)
  or u15839 (Rzrow6, Yzrow6, Gxrow6);  // ../RTL/cortexm0ds_logic.v(13505)
  AL_MUX u1584 (
    .i0(vis_pc_o[3]),
    .i1(Tugpw6[2]),
    .sel(Ty0iu6),
    .o(C01iu6));  // ../RTL/cortexm0ds_logic.v(3524)
  and u15840 (Kzrow6, F0sow6, M0sow6);  // ../RTL/cortexm0ds_logic.v(13506)
  and u15841 (n4373, Iyrow6, T0sow6);  // ../RTL/cortexm0ds_logic.v(13507)
  not u15842 (M0sow6, n4373);  // ../RTL/cortexm0ds_logic.v(13507)
  not u15843 (T0sow6, Pyrow6);  // ../RTL/cortexm0ds_logic.v(13508)
  or u15844 (n4374, M6fow6, A1sow6);  // ../RTL/cortexm0ds_logic.v(13509)
  not u15845 (Iyrow6, n4374);  // ../RTL/cortexm0ds_logic.v(13509)
  and u15846 (n4375, H1sow6, O1sow6);  // ../RTL/cortexm0ds_logic.v(13510)
  not u15847 (F0sow6, n4375);  // ../RTL/cortexm0ds_logic.v(13510)
  and u15848 (n4376, Gxrow6, Yzrow6);  // ../RTL/cortexm0ds_logic.v(13511)
  not u15849 (O1sow6, n4376);  // ../RTL/cortexm0ds_logic.v(13511)
  and u1585 (U2ihu6, J01iu6, Mxjhu6);  // ../RTL/cortexm0ds_logic.v(3525)
  not u15850 (Yzrow6, Zwrow6);  // ../RTL/cortexm0ds_logic.v(13512)
  AL_MUX u15851 (
    .i0(V1sow6),
    .i1(C2sow6),
    .sel(M6fow6),
    .o(Zwrow6));  // ../RTL/cortexm0ds_logic.v(13513)
  AL_MUX u15852 (
    .i0(J2sow6),
    .i1(Q2sow6),
    .sel(X2sow6),
    .o(Gxrow6));  // ../RTL/cortexm0ds_logic.v(13514)
  and u15853 (n4377, Ysrow6, Ewrow6);  // ../RTL/cortexm0ds_logic.v(13515)
  not u15854 (H1sow6, n4377);  // ../RTL/cortexm0ds_logic.v(13515)
  AL_MUX u15855 (
    .i0(E3sow6),
    .i1(L3sow6),
    .sel(V7fow6),
    .o(Ewrow6));  // ../RTL/cortexm0ds_logic.v(13516)
  buf u15856 (Rrlhu6, Nvkbx6[24]);  // ../RTL/cortexm0ds_logic.v(3137)
  not u15857 (Ysrow6, Lwrow6);  // ../RTL/cortexm0ds_logic.v(13518)
  AL_MUX u15858 (
    .i0(S3sow6),
    .i1(Z3sow6),
    .sel(M6fow6),
    .o(Lwrow6));  // ../RTL/cortexm0ds_logic.v(13519)
  and u15859 (M6fow6, G4sow6, N4sow6);  // ../RTL/cortexm0ds_logic.v(13520)
  AL_MUX u1586 (
    .i0(vis_pc_o[4]),
    .i1(Tugpw6[3]),
    .sel(Ty0iu6),
    .o(J01iu6));  // ../RTL/cortexm0ds_logic.v(3526)
  and u15860 (n4378, U4sow6, B5sow6);  // ../RTL/cortexm0ds_logic.v(13521)
  not u15861 (N4sow6, n4378);  // ../RTL/cortexm0ds_logic.v(13521)
  and u15862 (n4379, I5sow6, P5sow6);  // ../RTL/cortexm0ds_logic.v(13522)
  not u15863 (B5sow6, n4379);  // ../RTL/cortexm0ds_logic.v(13522)
  or u15864 (P5sow6, W5sow6, D6sow6);  // ../RTL/cortexm0ds_logic.v(13523)
  AL_MUX u15865 (
    .i0(R4gpw6[44]),
    .i1(R4gpw6[46]),
    .sel(Wagow6),
    .o(D6sow6));  // ../RTL/cortexm0ds_logic.v(13524)
  and u15866 (n4380, Z3sow6, K6sow6);  // ../RTL/cortexm0ds_logic.v(13525)
  not u15867 (W5sow6, n4380);  // ../RTL/cortexm0ds_logic.v(13525)
  and u15868 (n4381, V1sow6, R6sow6);  // ../RTL/cortexm0ds_logic.v(13526)
  not u15869 (K6sow6, n4381);  // ../RTL/cortexm0ds_logic.v(13526)
  and u1587 (C4ihu6, Q01iu6, Ewjhu6);  // ../RTL/cortexm0ds_logic.v(3527)
  or u15870 (I5sow6, R6sow6, V1sow6);  // ../RTL/cortexm0ds_logic.v(13527)
  AL_MUX u15871 (
    .i0(R4gpw6[45]),
    .i1(R4gpw6[47]),
    .sel(Wagow6),
    .o(V1sow6));  // ../RTL/cortexm0ds_logic.v(13528)
  not u15872 (Wagow6, A1sow6);  // ../RTL/cortexm0ds_logic.v(13529)
  not u15873 (R6sow6, C2sow6);  // ../RTL/cortexm0ds_logic.v(13530)
  AL_MUX u15874 (
    .i0(R4gpw6[41]),
    .i1(R4gpw6[43]),
    .sel(Dbgow6),
    .o(C2sow6));  // ../RTL/cortexm0ds_logic.v(13531)
  or u15875 (U4sow6, Pyrow6, A1sow6);  // ../RTL/cortexm0ds_logic.v(13532)
  and u15876 (n4382, Dbgow6, Y6sow6);  // ../RTL/cortexm0ds_logic.v(13533)
  not u15877 (G4sow6, n4382);  // ../RTL/cortexm0ds_logic.v(13533)
  and u15878 (n4383, Vbgpw6[21], Odgpw6[21]);  // ../RTL/cortexm0ds_logic.v(13534)
  not u15879 (Y6sow6, n4383);  // ../RTL/cortexm0ds_logic.v(13534)
  AL_MUX u1588 (
    .i0(vis_pc_o[5]),
    .i1(Tugpw6[4]),
    .sel(Ty0iu6),
    .o(Q01iu6));  // ../RTL/cortexm0ds_logic.v(3528)
  AL_MUX u15880 (
    .i0(R4gpw6[40]),
    .i1(R4gpw6[42]),
    .sel(Dbgow6),
    .o(Z3sow6));  // ../RTL/cortexm0ds_logic.v(13535)
  buf u15881 (Yslhu6, Nvkbx6[23]);  // ../RTL/cortexm0ds_logic.v(3137)
  and u15882 (F7sow6, M7sow6, Vbgpw6[20]);  // ../RTL/cortexm0ds_logic.v(13537)
  not u15883 (Dbgow6, F7sow6);  // ../RTL/cortexm0ds_logic.v(13537)
  and u15884 (M7sow6, Odgpw6[20], T7sow6);  // ../RTL/cortexm0ds_logic.v(13538)
  and u15885 (n4384, A8sow6, Vbgpw6[21]);  // ../RTL/cortexm0ds_logic.v(13539)
  not u15886 (T7sow6, n4384);  // ../RTL/cortexm0ds_logic.v(13539)
  and u15887 (A8sow6, Odgpw6[21], H8sow6);  // ../RTL/cortexm0ds_logic.v(13540)
  and u15888 (n4385, O8sow6, V8sow6);  // ../RTL/cortexm0ds_logic.v(13541)
  not u15889 (H8sow6, n4385);  // ../RTL/cortexm0ds_logic.v(13541)
  and u1589 (K5ihu6, X01iu6, Wujhu6);  // ../RTL/cortexm0ds_logic.v(3529)
  and u15890 (n4386, C9sow6, R4gpw6[40]);  // ../RTL/cortexm0ds_logic.v(13542)
  not u15891 (V8sow6, n4386);  // ../RTL/cortexm0ds_logic.v(13542)
  or u15892 (n4387, J9sow6, R4gpw6[42]);  // ../RTL/cortexm0ds_logic.v(13543)
  not u15893 (C9sow6, n4387);  // ../RTL/cortexm0ds_logic.v(13543)
  or u15894 (n4388, Q9sow6, R4gpw6[41]);  // ../RTL/cortexm0ds_logic.v(13544)
  not u15895 (J9sow6, n4388);  // ../RTL/cortexm0ds_logic.v(13544)
  and u15896 (n4389, R4gpw6[41], Q9sow6);  // ../RTL/cortexm0ds_logic.v(13545)
  not u15897 (O8sow6, n4389);  // ../RTL/cortexm0ds_logic.v(13545)
  AL_MUX u15898 (
    .i0(R4gpw6[46]),
    .i1(R4gpw6[44]),
    .sel(A1sow6),
    .o(S3sow6));  // ../RTL/cortexm0ds_logic.v(13546)
  and u15899 (A1sow6, X9sow6, Vbgpw6[22]);  // ../RTL/cortexm0ds_logic.v(13547)
  buf u159 (vis_r12_o[26], F4tax6);  // ../RTL/cortexm0ds_logic.v(2599)
  AL_MUX u1590 (
    .i0(vis_pc_o[6]),
    .i1(Tugpw6[5]),
    .sel(Ty0iu6),
    .o(X01iu6));  // ../RTL/cortexm0ds_logic.v(3530)
  and u15900 (X9sow6, Odgpw6[22], Easow6);  // ../RTL/cortexm0ds_logic.v(13548)
  and u15901 (n4390, Lasow6, Pyrow6);  // ../RTL/cortexm0ds_logic.v(13549)
  not u15902 (Easow6, n4390);  // ../RTL/cortexm0ds_logic.v(13549)
  and u15903 (Pyrow6, Vbgpw6[23], Odgpw6[23]);  // ../RTL/cortexm0ds_logic.v(13550)
  and u15904 (Lasow6, Sasow6, Zasow6);  // ../RTL/cortexm0ds_logic.v(13551)
  and u15905 (n4391, Gbsow6, Nbsow6);  // ../RTL/cortexm0ds_logic.v(13552)
  not u15906 (Zasow6, n4391);  // ../RTL/cortexm0ds_logic.v(13552)
  or u15907 (Nbsow6, Ubsow6, R4gpw6[47]);  // ../RTL/cortexm0ds_logic.v(13553)
  and u15908 (n4392, R4gpw6[44], Bcsow6);  // ../RTL/cortexm0ds_logic.v(13554)
  not u15909 (Gbsow6, n4392);  // ../RTL/cortexm0ds_logic.v(13554)
  and u1591 (S6ihu6, E11iu6, Otjhu6);  // ../RTL/cortexm0ds_logic.v(3531)
  and u15910 (n4393, R4gpw6[47], Ubsow6);  // ../RTL/cortexm0ds_logic.v(13555)
  not u15911 (Sasow6, n4393);  // ../RTL/cortexm0ds_logic.v(13555)
  and u15912 (n4394, Icsow6, Pcsow6);  // ../RTL/cortexm0ds_logic.v(13556)
  not u15913 (Wyrow6, n4394);  // ../RTL/cortexm0ds_logic.v(13556)
  and u15914 (Icsow6, X2sow6, Kbgow6);  // ../RTL/cortexm0ds_logic.v(13557)
  and u15915 (V7fow6, Wcsow6, Ddsow6);  // ../RTL/cortexm0ds_logic.v(13558)
  not u15916 (X2sow6, V7fow6);  // ../RTL/cortexm0ds_logic.v(13558)
  and u15917 (n4395, Kdsow6, Rdsow6);  // ../RTL/cortexm0ds_logic.v(13559)
  not u15918 (Ddsow6, n4395);  // ../RTL/cortexm0ds_logic.v(13559)
  and u15919 (n4396, Ydsow6, Fesow6);  // ../RTL/cortexm0ds_logic.v(13560)
  AL_MUX u1592 (
    .i0(vis_pc_o[7]),
    .i1(Tugpw6[6]),
    .sel(Ty0iu6),
    .o(E11iu6));  // ../RTL/cortexm0ds_logic.v(3532)
  not u15920 (Rdsow6, n4396);  // ../RTL/cortexm0ds_logic.v(13560)
  and u15921 (n4397, Mesow6, L3sow6);  // ../RTL/cortexm0ds_logic.v(13561)
  not u15922 (Fesow6, n4397);  // ../RTL/cortexm0ds_logic.v(13561)
  AL_MUX u15923 (
    .i0(R4gpw6[32]),
    .i1(R4gpw6[34]),
    .sel(Rbgow6),
    .o(L3sow6));  // ../RTL/cortexm0ds_logic.v(13562)
  or u15924 (n4398, E3sow6, Tesow6);  // ../RTL/cortexm0ds_logic.v(13563)
  not u15925 (Mesow6, n4398);  // ../RTL/cortexm0ds_logic.v(13563)
  or u15926 (n4399, Afsow6, J2sow6);  // ../RTL/cortexm0ds_logic.v(13564)
  not u15927 (Tesow6, n4399);  // ../RTL/cortexm0ds_logic.v(13564)
  AL_MUX u15928 (
    .i0(R4gpw6[36]),
    .i1(R4gpw6[38]),
    .sel(Kbgow6),
    .o(E3sow6));  // ../RTL/cortexm0ds_logic.v(13565)
  and u15929 (n4400, J2sow6, Afsow6);  // ../RTL/cortexm0ds_logic.v(13566)
  or u1593 (Msmhu6, Yx0iu6, G4hpw6[4]);  // ../RTL/cortexm0ds_logic.v(3533)
  not u15930 (Ydsow6, n4400);  // ../RTL/cortexm0ds_logic.v(13566)
  not u15931 (Afsow6, Q2sow6);  // ../RTL/cortexm0ds_logic.v(13567)
  AL_MUX u15932 (
    .i0(R4gpw6[37]),
    .i1(R4gpw6[39]),
    .sel(Kbgow6),
    .o(Q2sow6));  // ../RTL/cortexm0ds_logic.v(13568)
  AL_MUX u15933 (
    .i0(R4gpw6[33]),
    .i1(R4gpw6[35]),
    .sel(Rbgow6),
    .o(J2sow6));  // ../RTL/cortexm0ds_logic.v(13569)
  and u15934 (n4401, Pcsow6, Kbgow6);  // ../RTL/cortexm0ds_logic.v(13570)
  not u15935 (Kdsow6, n4401);  // ../RTL/cortexm0ds_logic.v(13570)
  and u15936 (n4402, Hfsow6, Vbgpw6[18]);  // ../RTL/cortexm0ds_logic.v(13571)
  not u15937 (Kbgow6, n4402);  // ../RTL/cortexm0ds_logic.v(13571)
  and u15938 (Hfsow6, Odgpw6[18], Ofsow6);  // ../RTL/cortexm0ds_logic.v(13572)
  or u15939 (Ofsow6, Vfsow6, Pcsow6);  // ../RTL/cortexm0ds_logic.v(13573)
  and u1594 (A8ihu6, L11iu6, Gsjhu6);  // ../RTL/cortexm0ds_logic.v(3534)
  and u15940 (n4403, Cgsow6, Jgsow6);  // ../RTL/cortexm0ds_logic.v(13574)
  not u15941 (Vfsow6, n4403);  // ../RTL/cortexm0ds_logic.v(13574)
  and u15942 (n4404, Qgsow6, Xgsow6);  // ../RTL/cortexm0ds_logic.v(13575)
  not u15943 (Jgsow6, n4404);  // ../RTL/cortexm0ds_logic.v(13575)
  or u15944 (Xgsow6, Ehsow6, R4gpw6[39]);  // ../RTL/cortexm0ds_logic.v(13576)
  and u15945 (n4405, R4gpw6[36], Lhsow6);  // ../RTL/cortexm0ds_logic.v(13577)
  not u15946 (Qgsow6, n4405);  // ../RTL/cortexm0ds_logic.v(13577)
  and u15947 (n4406, R4gpw6[39], Ehsow6);  // ../RTL/cortexm0ds_logic.v(13578)
  not u15948 (Cgsow6, n4406);  // ../RTL/cortexm0ds_logic.v(13578)
  and u15949 (n4407, Vbgpw6[19], Odgpw6[19]);  // ../RTL/cortexm0ds_logic.v(13579)
  AL_MUX u1595 (
    .i0(vis_pc_o[8]),
    .i1(Tugpw6[7]),
    .sel(Ty0iu6),
    .o(L11iu6));  // ../RTL/cortexm0ds_logic.v(3535)
  not u15950 (Pcsow6, n4407);  // ../RTL/cortexm0ds_logic.v(13579)
  and u15951 (n4408, Rbgow6, Shsow6);  // ../RTL/cortexm0ds_logic.v(13580)
  not u15952 (Wcsow6, n4408);  // ../RTL/cortexm0ds_logic.v(13580)
  and u15953 (Nisow6, Vbgpw6[17], Odgpw6[17]);  // ../RTL/cortexm0ds_logic.v(13581)
  not u15954 (Shsow6, Nisow6);  // ../RTL/cortexm0ds_logic.v(13581)
  and u15955 (n4409, Zhsow6, Vbgpw6[16]);  // ../RTL/cortexm0ds_logic.v(13582)
  not u15956 (Rbgow6, n4409);  // ../RTL/cortexm0ds_logic.v(13582)
  and u15957 (Zhsow6, Odgpw6[16], Gisow6);  // ../RTL/cortexm0ds_logic.v(13583)
  and u15958 (n4410, Nisow6, Uisow6);  // ../RTL/cortexm0ds_logic.v(13584)
  not u15959 (Gisow6, n4410);  // ../RTL/cortexm0ds_logic.v(13584)
  and u1596 (I9ihu6, S11iu6, Yqjhu6);  // ../RTL/cortexm0ds_logic.v(3536)
  and u15960 (Uisow6, Bjsow6, Ijsow6);  // ../RTL/cortexm0ds_logic.v(13585)
  and u15961 (n4411, Pjsow6, Wjsow6);  // ../RTL/cortexm0ds_logic.v(13586)
  not u15962 (Ijsow6, n4411);  // ../RTL/cortexm0ds_logic.v(13586)
  and u15963 (n4412, R4gpw6[33], Dksow6);  // ../RTL/cortexm0ds_logic.v(13587)
  not u15964 (Wjsow6, n4412);  // ../RTL/cortexm0ds_logic.v(13587)
  and u15965 (n4413, R4gpw6[32], Kksow6);  // ../RTL/cortexm0ds_logic.v(13588)
  not u15966 (Pjsow6, n4413);  // ../RTL/cortexm0ds_logic.v(13588)
  not u15967 (Kksow6, R4gpw6[34]);  // ../RTL/cortexm0ds_logic.v(13589)
  or u15968 (Bjsow6, Dksow6, R4gpw6[33]);  // ../RTL/cortexm0ds_logic.v(13590)
  buf u15969 (Dnfhu6, Ozkbx6[2]);  // ../RTL/cortexm0ds_logic.v(3176)
  AL_MUX u1597 (
    .i0(vis_pc_o[9]),
    .i1(Tugpw6[8]),
    .sel(Ty0iu6),
    .o(S11iu6));  // ../RTL/cortexm0ds_logic.v(3537)
  AL_MUX u15970 (
    .i0(Rksow6),
    .i1(Yksow6),
    .sel(Hdgow6),
    .o(Mtrow6));  // ../RTL/cortexm0ds_logic.v(13592)
  buf u15971 (Fulhu6, Nvkbx6[22]);  // ../RTL/cortexm0ds_logic.v(3137)
  and u15972 (Hdgow6, Flsow6, Mlsow6);  // ../RTL/cortexm0ds_logic.v(13594)
  not u15973 (Q8fow6, Hdgow6);  // ../RTL/cortexm0ds_logic.v(13594)
  or u15974 (Mlsow6, Tlsow6, Amsow6);  // ../RTL/cortexm0ds_logic.v(13595)
  or u15975 (Tlsow6, X8fow6, Vdgow6);  // ../RTL/cortexm0ds_logic.v(13596)
  and u15976 (n4414, Hmsow6, Omsow6);  // ../RTL/cortexm0ds_logic.v(13597)
  not u15977 (Flsow6, n4414);  // ../RTL/cortexm0ds_logic.v(13597)
  and u15978 (n4415, Vmsow6, Cnsow6);  // ../RTL/cortexm0ds_logic.v(13598)
  not u15979 (Omsow6, n4415);  // ../RTL/cortexm0ds_logic.v(13598)
  and u1598 (Qaihu6, Z11iu6, Qpjhu6);  // ../RTL/cortexm0ds_logic.v(3538)
  and u15980 (n4416, Jnsow6, Qnsow6);  // ../RTL/cortexm0ds_logic.v(13599)
  not u15981 (Cnsow6, n4416);  // ../RTL/cortexm0ds_logic.v(13599)
  and u15982 (Qnsow6, Xnsow6, Eosow6);  // ../RTL/cortexm0ds_logic.v(13600)
  or u15983 (Xnsow6, Nxrow6, Losow6);  // ../RTL/cortexm0ds_logic.v(13601)
  and u15984 (Jnsow6, Yksow6, Sosow6);  // ../RTL/cortexm0ds_logic.v(13602)
  and u15985 (n4417, Losow6, Nxrow6);  // ../RTL/cortexm0ds_logic.v(13603)
  not u15986 (Vmsow6, n4417);  // ../RTL/cortexm0ds_logic.v(13603)
  AL_MUX u15987 (
    .i0(Zosow6),
    .i1(Gpsow6),
    .sel(Jegow6),
    .o(Nxrow6));  // ../RTL/cortexm0ds_logic.v(13604)
  not u15988 (Zosow6, Npsow6);  // ../RTL/cortexm0ds_logic.v(13605)
  not u15989 (Losow6, Uxrow6);  // ../RTL/cortexm0ds_logic.v(13606)
  AL_MUX u1599 (
    .i0(vis_pc_o[10]),
    .i1(Tugpw6[9]),
    .sel(Ty0iu6),
    .o(Z11iu6));  // ../RTL/cortexm0ds_logic.v(3539)
  AL_MUX u15990 (
    .i0(Upsow6),
    .i1(Bqsow6),
    .sel(X8fow6),
    .o(Uxrow6));  // ../RTL/cortexm0ds_logic.v(13607)
  buf u15991 (Mvlhu6, Nvkbx6[21]);  // ../RTL/cortexm0ds_logic.v(3137)
  and u15992 (n4418, Tmrow6, Jegow6);  // ../RTL/cortexm0ds_logic.v(13609)
  not u15993 (Hmsow6, n4418);  // ../RTL/cortexm0ds_logic.v(13609)
  AL_MUX u15994 (
    .i0(Iqsow6),
    .i1(Pqsow6),
    .sel(Cegow6),
    .o(Yksow6));  // ../RTL/cortexm0ds_logic.v(13610)
  and u15995 (X8fow6, Wqsow6, Drsow6);  // ../RTL/cortexm0ds_logic.v(13611)
  not u15996 (Cegow6, X8fow6);  // ../RTL/cortexm0ds_logic.v(13611)
  and u15997 (n4419, Krsow6, Rrsow6);  // ../RTL/cortexm0ds_logic.v(13612)
  not u15998 (Drsow6, n4419);  // ../RTL/cortexm0ds_logic.v(13612)
  and u15999 (n4420, Yrsow6, Fssow6);  // ../RTL/cortexm0ds_logic.v(13613)
  buf u16 (O5ohu6, Nyhpw6);  // ../RTL/cortexm0ds_logic.v(1772)
  buf u160 (Uthpw6[3], Xu2qw6);  // ../RTL/cortexm0ds_logic.v(1882)
  and u1600 (Ybihu6, G21iu6, Iojhu6);  // ../RTL/cortexm0ds_logic.v(3540)
  not u16000 (Rrsow6, n4420);  // ../RTL/cortexm0ds_logic.v(13613)
  and u16001 (n4421, Mssow6, Iqsow6);  // ../RTL/cortexm0ds_logic.v(13614)
  not u16002 (Fssow6, n4421);  // ../RTL/cortexm0ds_logic.v(13614)
  or u16003 (n4422, Pqsow6, Tssow6);  // ../RTL/cortexm0ds_logic.v(13615)
  not u16004 (Mssow6, n4422);  // ../RTL/cortexm0ds_logic.v(13615)
  or u16005 (n4423, Atsow6, Upsow6);  // ../RTL/cortexm0ds_logic.v(13616)
  not u16006 (Tssow6, n4423);  // ../RTL/cortexm0ds_logic.v(13616)
  and u16007 (n4424, Upsow6, Atsow6);  // ../RTL/cortexm0ds_logic.v(13617)
  not u16008 (Yrsow6, n4424);  // ../RTL/cortexm0ds_logic.v(13617)
  not u16009 (Atsow6, Bqsow6);  // ../RTL/cortexm0ds_logic.v(13618)
  AL_MUX u1601 (
    .i0(vis_pc_o[11]),
    .i1(Ixdpw6),
    .sel(Ty0iu6),
    .o(G21iu6));  // ../RTL/cortexm0ds_logic.v(3541)
  AL_MUX u16010 (
    .i0(Htsow6),
    .i1(Otsow6),
    .sel(Odgow6),
    .o(Bqsow6));  // ../RTL/cortexm0ds_logic.v(13619)
  AL_MUX u16011 (
    .i0(Vtsow6),
    .i1(Cusow6),
    .sel(Jusow6),
    .o(Upsow6));  // ../RTL/cortexm0ds_logic.v(13620)
  or u16012 (Krsow6, Amsow6, Vdgow6);  // ../RTL/cortexm0ds_logic.v(13621)
  or u16013 (Wqsow6, Odgow6, Qusow6);  // ../RTL/cortexm0ds_logic.v(13622)
  AL_MUX u16014 (
    .i0(R4gpw6[52]),
    .i1(R4gpw6[54]),
    .sel(Jusow6),
    .o(Pqsow6));  // ../RTL/cortexm0ds_logic.v(13623)
  not u16015 (Jusow6, Vdgow6);  // ../RTL/cortexm0ds_logic.v(13624)
  and u16016 (Vdgow6, Xusow6, Vbgpw6[26]);  // ../RTL/cortexm0ds_logic.v(13625)
  and u16017 (Xusow6, Odgpw6[26], Evsow6);  // ../RTL/cortexm0ds_logic.v(13626)
  and u16018 (n4425, Lvsow6, Amsow6);  // ../RTL/cortexm0ds_logic.v(13627)
  not u16019 (Evsow6, n4425);  // ../RTL/cortexm0ds_logic.v(13627)
  and u1602 (Gdihu6, N21iu6, Anjhu6);  // ../RTL/cortexm0ds_logic.v(3542)
  and u16020 (Amsow6, Vbgpw6[27], Odgpw6[27]);  // ../RTL/cortexm0ds_logic.v(13628)
  and u16021 (Lvsow6, Svsow6, Zvsow6);  // ../RTL/cortexm0ds_logic.v(13629)
  and u16022 (n4426, Gwsow6, Nwsow6);  // ../RTL/cortexm0ds_logic.v(13630)
  not u16023 (Zvsow6, n4426);  // ../RTL/cortexm0ds_logic.v(13630)
  or u16024 (Nwsow6, Vtsow6, R4gpw6[55]);  // ../RTL/cortexm0ds_logic.v(13631)
  or u16025 (Gwsow6, Uwsow6, R4gpw6[54]);  // ../RTL/cortexm0ds_logic.v(13632)
  or u16026 (Svsow6, Cusow6, R4gpw6[53]);  // ../RTL/cortexm0ds_logic.v(13633)
  AL_MUX u16027 (
    .i0(R4gpw6[50]),
    .i1(R4gpw6[48]),
    .sel(Odgow6),
    .o(Iqsow6));  // ../RTL/cortexm0ds_logic.v(13634)
  and u16028 (Odgow6, Bxsow6, Vbgpw6[24]);  // ../RTL/cortexm0ds_logic.v(13635)
  and u16029 (Bxsow6, Odgpw6[24], Ixsow6);  // ../RTL/cortexm0ds_logic.v(13636)
  AL_MUX u1603 (
    .i0(vis_pc_o[12]),
    .i1(Tugpw6[11]),
    .sel(Ty0iu6),
    .o(N21iu6));  // ../RTL/cortexm0ds_logic.v(3543)
  and u16030 (n4427, Qusow6, Pxsow6);  // ../RTL/cortexm0ds_logic.v(13637)
  not u16031 (Ixsow6, n4427);  // ../RTL/cortexm0ds_logic.v(13637)
  and u16032 (Pxsow6, Wxsow6, Dysow6);  // ../RTL/cortexm0ds_logic.v(13638)
  and u16033 (n4428, Kysow6, Rysow6);  // ../RTL/cortexm0ds_logic.v(13639)
  not u16034 (Dysow6, n4428);  // ../RTL/cortexm0ds_logic.v(13639)
  or u16035 (Rysow6, Otsow6, R4gpw6[51]);  // ../RTL/cortexm0ds_logic.v(13640)
  or u16036 (Kysow6, Yysow6, R4gpw6[50]);  // ../RTL/cortexm0ds_logic.v(13641)
  or u16037 (Wxsow6, Htsow6, R4gpw6[49]);  // ../RTL/cortexm0ds_logic.v(13642)
  and u16038 (Qusow6, Vbgpw6[25], Odgpw6[25]);  // ../RTL/cortexm0ds_logic.v(13643)
  and u16039 (n4429, Eosow6, Sosow6);  // ../RTL/cortexm0ds_logic.v(13644)
  and u1604 (Oeihu6, U21iu6, Sljhu6);  // ../RTL/cortexm0ds_logic.v(3544)
  not u16040 (Rksow6, n4429);  // ../RTL/cortexm0ds_logic.v(13644)
  and u16041 (n4430, Fzsow6, Jegow6);  // ../RTL/cortexm0ds_logic.v(13645)
  not u16042 (Sosow6, n4430);  // ../RTL/cortexm0ds_logic.v(13645)
  and u16043 (n4431, Mzsow6, Tzsow6);  // ../RTL/cortexm0ds_logic.v(13646)
  not u16044 (Eosow6, n4431);  // ../RTL/cortexm0ds_logic.v(13646)
  buf u16045 (Twlhu6, Nvkbx6[20]);  // ../RTL/cortexm0ds_logic.v(3137)
  and u16046 (Mzsow6, A0tow6, H0tow6);  // ../RTL/cortexm0ds_logic.v(13648)
  not u16047 (Jegow6, Mzsow6);  // ../RTL/cortexm0ds_logic.v(13648)
  or u16048 (H0tow6, Tmrow6, O0tow6);  // ../RTL/cortexm0ds_logic.v(13649)
  and u16049 (O0tow6, V0tow6, C1tow6);  // ../RTL/cortexm0ds_logic.v(13650)
  AL_MUX u1605 (
    .i0(vis_pc_o[13]),
    .i1(Tugpw6[12]),
    .sel(Ty0iu6),
    .o(U21iu6));  // ../RTL/cortexm0ds_logic.v(3545)
  and u16050 (n4432, J1tow6, Tzsow6);  // ../RTL/cortexm0ds_logic.v(13651)
  not u16051 (C1tow6, n4432);  // ../RTL/cortexm0ds_logic.v(13651)
  AL_MUX u16052 (
    .i0(R4gpw6[56]),
    .i1(R4gpw6[58]),
    .sel(Q1tow6),
    .o(Tzsow6));  // ../RTL/cortexm0ds_logic.v(13652)
  or u16053 (n4433, Fzsow6, X1tow6);  // ../RTL/cortexm0ds_logic.v(13653)
  not u16054 (J1tow6, n4433);  // ../RTL/cortexm0ds_logic.v(13653)
  or u16055 (n4434, Npsow6, Gpsow6);  // ../RTL/cortexm0ds_logic.v(13654)
  not u16056 (X1tow6, n4434);  // ../RTL/cortexm0ds_logic.v(13654)
  AL_MUX u16057 (
    .i0(R4gpw6[60]),
    .i1(R4gpw6[62]),
    .sel(Mcgow6),
    .o(Fzsow6));  // ../RTL/cortexm0ds_logic.v(13655)
  and u16058 (n4435, Gpsow6, Npsow6);  // ../RTL/cortexm0ds_logic.v(13656)
  not u16059 (V0tow6, n4435);  // ../RTL/cortexm0ds_logic.v(13656)
  and u1606 (Wfihu6, B31iu6, Kkjhu6);  // ../RTL/cortexm0ds_logic.v(3546)
  AL_MUX u16060 (
    .i0(R4gpw6[59]),
    .i1(R4gpw6[57]),
    .sel(Qegow6),
    .o(Npsow6));  // ../RTL/cortexm0ds_logic.v(13657)
  buf u16061 (Aylhu6, Nvkbx6[19]);  // ../RTL/cortexm0ds_logic.v(3137)
  AL_MUX u16062 (
    .i0(E2tow6),
    .i1(L2tow6),
    .sel(Mcgow6),
    .o(Gpsow6));  // ../RTL/cortexm0ds_logic.v(13659)
  and u16063 (Tmrow6, Mcgow6, S2tow6);  // ../RTL/cortexm0ds_logic.v(13660)
  and u16064 (N3tow6, Vbgpw6[31], Odgpw6[31]);  // ../RTL/cortexm0ds_logic.v(13661)
  not u16065 (S2tow6, N3tow6);  // ../RTL/cortexm0ds_logic.v(13661)
  and u16066 (n4436, Z2tow6, Vbgpw6[30]);  // ../RTL/cortexm0ds_logic.v(13662)
  not u16067 (Mcgow6, n4436);  // ../RTL/cortexm0ds_logic.v(13662)
  and u16068 (Z2tow6, Odgpw6[30], G3tow6);  // ../RTL/cortexm0ds_logic.v(13663)
  and u16069 (n4437, N3tow6, U3tow6);  // ../RTL/cortexm0ds_logic.v(13664)
  AL_MUX u1607 (
    .i0(vis_pc_o[14]),
    .i1(Tugpw6[13]),
    .sel(Ty0iu6),
    .o(B31iu6));  // ../RTL/cortexm0ds_logic.v(3547)
  not u16070 (G3tow6, n4437);  // ../RTL/cortexm0ds_logic.v(13664)
  and u16071 (U3tow6, B4tow6, I4tow6);  // ../RTL/cortexm0ds_logic.v(13665)
  and u16072 (n4438, P4tow6, W4tow6);  // ../RTL/cortexm0ds_logic.v(13666)
  not u16073 (I4tow6, n4438);  // ../RTL/cortexm0ds_logic.v(13666)
  or u16074 (W4tow6, E2tow6, R4gpw6[63]);  // ../RTL/cortexm0ds_logic.v(13667)
  and u16075 (n4439, R4gpw6[60], D5tow6);  // ../RTL/cortexm0ds_logic.v(13668)
  not u16076 (P4tow6, n4439);  // ../RTL/cortexm0ds_logic.v(13668)
  not u16077 (D5tow6, R4gpw6[62]);  // ../RTL/cortexm0ds_logic.v(13669)
  or u16078 (B4tow6, L2tow6, R4gpw6[61]);  // ../RTL/cortexm0ds_logic.v(13670)
  not u16079 (L2tow6, R4gpw6[63]);  // ../RTL/cortexm0ds_logic.v(13671)
  and u1608 (Ehihu6, I31iu6, Cjjhu6);  // ../RTL/cortexm0ds_logic.v(3548)
  buf u16080 (Ighpw6[5], Pmlpw6);  // ../RTL/cortexm0ds_logic.v(1840)
  and u16081 (n4440, Q1tow6, K5tow6);  // ../RTL/cortexm0ds_logic.v(13673)
  not u16082 (A0tow6, n4440);  // ../RTL/cortexm0ds_logic.v(13673)
  and u16083 (n4441, Vbgpw6[29], Odgpw6[29]);  // ../RTL/cortexm0ds_logic.v(13674)
  not u16084 (K5tow6, n4441);  // ../RTL/cortexm0ds_logic.v(13674)
  and u16085 (Qegow6, R5tow6, Vbgpw6[28]);  // ../RTL/cortexm0ds_logic.v(13675)
  not u16086 (Q1tow6, Qegow6);  // ../RTL/cortexm0ds_logic.v(13675)
  and u16087 (R5tow6, Odgpw6[28], Y5tow6);  // ../RTL/cortexm0ds_logic.v(13676)
  and u16088 (n4442, F6tow6, Vbgpw6[29]);  // ../RTL/cortexm0ds_logic.v(13677)
  not u16089 (Y5tow6, n4442);  // ../RTL/cortexm0ds_logic.v(13677)
  AL_MUX u1609 (
    .i0(vis_pc_o[15]),
    .i1(Pxdpw6),
    .sel(Ty0iu6),
    .o(I31iu6));  // ../RTL/cortexm0ds_logic.v(3549)
  and u16090 (F6tow6, Odgpw6[29], M6tow6);  // ../RTL/cortexm0ds_logic.v(13678)
  and u16091 (n4443, T6tow6, A7tow6);  // ../RTL/cortexm0ds_logic.v(13679)
  not u16092 (M6tow6, n4443);  // ../RTL/cortexm0ds_logic.v(13679)
  and u16093 (n4444, H7tow6, R4gpw6[56]);  // ../RTL/cortexm0ds_logic.v(13680)
  not u16094 (A7tow6, n4444);  // ../RTL/cortexm0ds_logic.v(13680)
  or u16095 (n4445, O7tow6, R4gpw6[58]);  // ../RTL/cortexm0ds_logic.v(13681)
  not u16096 (H7tow6, n4445);  // ../RTL/cortexm0ds_logic.v(13681)
  or u16097 (n4446, V7tow6, R4gpw6[57]);  // ../RTL/cortexm0ds_logic.v(13682)
  not u16098 (O7tow6, n4446);  // ../RTL/cortexm0ds_logic.v(13682)
  and u16099 (n4447, R4gpw6[57], V7tow6);  // ../RTL/cortexm0ds_logic.v(13683)
  buf u161 (Jshpw6[27], Q4dbx6);  // ../RTL/cortexm0ds_logic.v(2372)
  and u1610 (Miihu6, P31iu6, Uhjhu6);  // ../RTL/cortexm0ds_logic.v(3550)
  not u16100 (T6tow6, n4447);  // ../RTL/cortexm0ds_logic.v(13683)
  and u16101 (Wrrow6, C8tow6, J8tow6);  // ../RTL/cortexm0ds_logic.v(13684)
  not u16102 (Anrow6, Wrrow6);  // ../RTL/cortexm0ds_logic.v(13684)
  and u16103 (n4448, Z2fow6, Q8tow6);  // ../RTL/cortexm0ds_logic.v(13685)
  not u16104 (J8tow6, n4448);  // ../RTL/cortexm0ds_logic.v(13685)
  and u16105 (Fdtow6, X8tow6, E9tow6);  // ../RTL/cortexm0ds_logic.v(13686)
  not u16106 (Q8tow6, Fdtow6);  // ../RTL/cortexm0ds_logic.v(13686)
  and u16107 (Z2fow6, B4fow6, I4fow6);  // ../RTL/cortexm0ds_logic.v(13687)
  AL_MUX u16108 (
    .i0(L9tow6),
    .i1(S9tow6),
    .sel(B4fow6),
    .o(C8tow6));  // ../RTL/cortexm0ds_logic.v(13688)
  buf u16109 (Hzlhu6, Nvkbx6[18]);  // ../RTL/cortexm0ds_logic.v(3137)
  AL_MUX u1611 (
    .i0(vis_pc_o[16]),
    .i1(Wxdpw6),
    .sel(Ty0iu6),
    .o(P31iu6));  // ../RTL/cortexm0ds_logic.v(3551)
  and u16110 (B4fow6, Z9tow6, Gatow6);  // ../RTL/cortexm0ds_logic.v(13690)
  buf u16111 (Qbehu6, Ozkbx6[33]);  // ../RTL/cortexm0ds_logic.v(3176)
  and u16112 (n4449, Dsrow6, Natow6);  // ../RTL/cortexm0ds_logic.v(13691)
  not u16113 (Gatow6, n4449);  // ../RTL/cortexm0ds_logic.v(13691)
  and u16114 (n4450, Uatow6, Bbtow6);  // ../RTL/cortexm0ds_logic.v(13692)
  not u16115 (Natow6, n4450);  // ../RTL/cortexm0ds_logic.v(13692)
  and u16116 (n4451, Ibtow6, Pbtow6);  // ../RTL/cortexm0ds_logic.v(13693)
  not u16117 (Bbtow6, n4451);  // ../RTL/cortexm0ds_logic.v(13693)
  and u16118 (Pbtow6, Wbtow6, Dctow6);  // ../RTL/cortexm0ds_logic.v(13694)
  or u16119 (Wbtow6, Prrow6, Irrow6);  // ../RTL/cortexm0ds_logic.v(13695)
  and u1612 (Ujihu6, W31iu6, Mgjhu6);  // ../RTL/cortexm0ds_logic.v(3552)
  or u16120 (n4452, Kctow6, Rctow6);  // ../RTL/cortexm0ds_logic.v(13696)
  not u16121 (Ibtow6, n4452);  // ../RTL/cortexm0ds_logic.v(13696)
  and u16122 (Rctow6, Nggow6, Yctow6);  // ../RTL/cortexm0ds_logic.v(13697)
  AL_MUX u16123 (
    .i0(Fdtow6),
    .i1(Mdtow6),
    .sel(Yigow6),
    .o(Kctow6));  // ../RTL/cortexm0ds_logic.v(13698)
  and u16124 (n4453, Irrow6, Prrow6);  // ../RTL/cortexm0ds_logic.v(13699)
  not u16125 (Uatow6, n4453);  // ../RTL/cortexm0ds_logic.v(13699)
  AL_MUX u16126 (
    .i0(Tdtow6),
    .i1(Aetow6),
    .sel(Nggow6),
    .o(Prrow6));  // ../RTL/cortexm0ds_logic.v(13700)
  AL_MUX u16127 (
    .i0(Hetow6),
    .i1(Oetow6),
    .sel(Yigow6),
    .o(Irrow6));  // ../RTL/cortexm0ds_logic.v(13701)
  and u16128 (n4454, Vetow6, Cftow6);  // ../RTL/cortexm0ds_logic.v(13702)
  not u16129 (Dsrow6, n4454);  // ../RTL/cortexm0ds_logic.v(13702)
  AL_MUX u1613 (
    .i0(vis_pc_o[17]),
    .i1(Dydpw6),
    .sel(Ty0iu6),
    .o(W31iu6));  // ../RTL/cortexm0ds_logic.v(3553)
  or u16130 (n4455, Jftow6, Nggow6);  // ../RTL/cortexm0ds_logic.v(13703)
  not u16131 (Vetow6, n4455);  // ../RTL/cortexm0ds_logic.v(13703)
  and u16132 (n4456, Qftow6, Xftow6);  // ../RTL/cortexm0ds_logic.v(13704)
  not u16133 (Z9tow6, n4456);  // ../RTL/cortexm0ds_logic.v(13704)
  or u16134 (n4457, Egtow6, Yigow6);  // ../RTL/cortexm0ds_logic.v(13705)
  not u16135 (Qftow6, n4457);  // ../RTL/cortexm0ds_logic.v(13705)
  buf u16136 (O0mhu6, Nvkbx6[17]);  // ../RTL/cortexm0ds_logic.v(3137)
  or u16137 (S9tow6, I4fow6, Mdtow6);  // ../RTL/cortexm0ds_logic.v(13707)
  not u16138 (Mdtow6, Lgtow6);  // ../RTL/cortexm0ds_logic.v(13708)
  and u16139 (Yigow6, Sgtow6, Zgtow6);  // ../RTL/cortexm0ds_logic.v(13709)
  and u1614 (Clihu6, D41iu6, Efjhu6);  // ../RTL/cortexm0ds_logic.v(3554)
  not u16140 (I4fow6, Yigow6);  // ../RTL/cortexm0ds_logic.v(13709)
  or u16141 (Zgtow6, Ghtow6, Nhtow6);  // ../RTL/cortexm0ds_logic.v(13710)
  or u16142 (Ghtow6, P4fow6, Mjgow6);  // ../RTL/cortexm0ds_logic.v(13711)
  and u16143 (n4458, Uhtow6, Bitow6);  // ../RTL/cortexm0ds_logic.v(13712)
  not u16144 (Sgtow6, n4458);  // ../RTL/cortexm0ds_logic.v(13712)
  and u16145 (n4459, Xftow6, Iitow6);  // ../RTL/cortexm0ds_logic.v(13713)
  not u16146 (Bitow6, n4459);  // ../RTL/cortexm0ds_logic.v(13713)
  not u16147 (Iitow6, Egtow6);  // ../RTL/cortexm0ds_logic.v(13714)
  or u16148 (n4460, Pitow6, Hkgow6);  // ../RTL/cortexm0ds_logic.v(13715)
  not u16149 (Xftow6, n4460);  // ../RTL/cortexm0ds_logic.v(13715)
  AL_MUX u1615 (
    .i0(vis_pc_o[18]),
    .i1(Kydpw6),
    .sel(Ty0iu6),
    .o(D41iu6));  // ../RTL/cortexm0ds_logic.v(3555)
  and u16150 (n4461, Witow6, Djtow6);  // ../RTL/cortexm0ds_logic.v(13716)
  not u16151 (Uhtow6, n4461);  // ../RTL/cortexm0ds_logic.v(13716)
  and u16152 (n4462, Kjtow6, Fdtow6);  // ../RTL/cortexm0ds_logic.v(13717)
  not u16153 (Djtow6, n4462);  // ../RTL/cortexm0ds_logic.v(13717)
  buf u16154 (Ighpw6[4], Yklpw6);  // ../RTL/cortexm0ds_logic.v(1840)
  and u16155 (n4463, Pitow6, Rjtow6);  // ../RTL/cortexm0ds_logic.v(13719)
  not u16156 (E9tow6, n4463);  // ../RTL/cortexm0ds_logic.v(13719)
  and u16157 (n4464, Yjtow6, G3fow6);  // ../RTL/cortexm0ds_logic.v(13720)
  not u16158 (X8tow6, n4464);  // ../RTL/cortexm0ds_logic.v(13720)
  and u16159 (Kjtow6, Lgtow6, Fktow6);  // ../RTL/cortexm0ds_logic.v(13721)
  and u1616 (Kmihu6, K41iu6, Wdjhu6);  // ../RTL/cortexm0ds_logic.v(3556)
  or u16160 (Fktow6, Mktow6, Oetow6);  // ../RTL/cortexm0ds_logic.v(13722)
  AL_MUX u16161 (
    .i0(Tktow6),
    .i1(Altow6),
    .sel(P4fow6),
    .o(Lgtow6));  // ../RTL/cortexm0ds_logic.v(13723)
  buf u16162 (V1mhu6, Nvkbx6[16]);  // ../RTL/cortexm0ds_logic.v(3137)
  AL_MUX u16163 (
    .i0(R4gpw6[2]),
    .i1(R4gpw6[0]),
    .sel(Fjgow6),
    .o(Altow6));  // ../RTL/cortexm0ds_logic.v(13725)
  and u16164 (n4465, Oetow6, Mktow6);  // ../RTL/cortexm0ds_logic.v(13726)
  not u16165 (Witow6, n4465);  // ../RTL/cortexm0ds_logic.v(13726)
  not u16166 (Mktow6, Hetow6);  // ../RTL/cortexm0ds_logic.v(13727)
  AL_MUX u16167 (
    .i0(Hltow6),
    .i1(Oltow6),
    .sel(Pitow6),
    .o(Hetow6));  // ../RTL/cortexm0ds_logic.v(13728)
  buf u16168 (C3mhu6, Nvkbx6[15]);  // ../RTL/cortexm0ds_logic.v(3137)
  and u16169 (Pitow6, Vltow6, Cmtow6);  // ../RTL/cortexm0ds_logic.v(13730)
  AL_MUX u1617 (
    .i0(vis_pc_o[19]),
    .i1(Rydpw6),
    .sel(Ty0iu6),
    .o(K41iu6));  // ../RTL/cortexm0ds_logic.v(3557)
  not u16170 (G3fow6, Pitow6);  // ../RTL/cortexm0ds_logic.v(13730)
  and u16171 (n4466, Jmtow6, Qmtow6);  // ../RTL/cortexm0ds_logic.v(13731)
  not u16172 (Cmtow6, n4466);  // ../RTL/cortexm0ds_logic.v(13731)
  and u16173 (n4467, Xmtow6, Entow6);  // ../RTL/cortexm0ds_logic.v(13732)
  not u16174 (Qmtow6, n4467);  // ../RTL/cortexm0ds_logic.v(13732)
  and u16175 (n4468, Lntow6, Rjtow6);  // ../RTL/cortexm0ds_logic.v(13733)
  not u16176 (Entow6, n4468);  // ../RTL/cortexm0ds_logic.v(13733)
  AL_MUX u16177 (
    .i0(R4gpw6[10]),
    .i1(R4gpw6[8]),
    .sel(Akgow6),
    .o(Rjtow6));  // ../RTL/cortexm0ds_logic.v(13734)
  or u16178 (n4469, Yjtow6, Sntow6);  // ../RTL/cortexm0ds_logic.v(13735)
  not u16179 (Lntow6, n4469);  // ../RTL/cortexm0ds_logic.v(13735)
  and u1618 (Snihu6, R41iu6, Ocjhu6);  // ../RTL/cortexm0ds_logic.v(3558)
  or u16180 (n4470, Zntow6, Oltow6);  // ../RTL/cortexm0ds_logic.v(13736)
  not u16181 (Sntow6, n4470);  // ../RTL/cortexm0ds_logic.v(13736)
  AL_MUX u16182 (
    .i0(R4gpw6[14]),
    .i1(R4gpw6[12]),
    .sel(Hkgow6),
    .o(Yjtow6));  // ../RTL/cortexm0ds_logic.v(13737)
  and u16183 (n4471, Oltow6, Zntow6);  // ../RTL/cortexm0ds_logic.v(13738)
  not u16184 (Xmtow6, n4471);  // ../RTL/cortexm0ds_logic.v(13738)
  or u16185 (Jmtow6, Egtow6, Hkgow6);  // ../RTL/cortexm0ds_logic.v(13739)
  and u16186 (n4472, Gotow6, Notow6);  // ../RTL/cortexm0ds_logic.v(13740)
  not u16187 (Vltow6, n4472);  // ../RTL/cortexm0ds_logic.v(13740)
  and u16188 (n4473, Vbgpw6[5], Odgpw6[5]);  // ../RTL/cortexm0ds_logic.v(13741)
  not u16189 (Notow6, n4473);  // ../RTL/cortexm0ds_logic.v(13741)
  AL_MUX u1619 (
    .i0(vis_pc_o[20]),
    .i1(Yydpw6),
    .sel(Ty0iu6),
    .o(R41iu6));  // ../RTL/cortexm0ds_logic.v(3559)
  AL_MUX u16190 (
    .i0(R4gpw6[11]),
    .i1(R4gpw6[9]),
    .sel(Akgow6),
    .o(Oltow6));  // ../RTL/cortexm0ds_logic.v(13742)
  buf u16191 (J4mhu6, Nvkbx6[14]);  // ../RTL/cortexm0ds_logic.v(3137)
  and u16192 (Akgow6, Uotow6, Vbgpw6[4]);  // ../RTL/cortexm0ds_logic.v(13744)
  not u16193 (Gotow6, Akgow6);  // ../RTL/cortexm0ds_logic.v(13744)
  and u16194 (Uotow6, Odgpw6[4], Bptow6);  // ../RTL/cortexm0ds_logic.v(13745)
  and u16195 (n4474, Iptow6, Vbgpw6[5]);  // ../RTL/cortexm0ds_logic.v(13746)
  not u16196 (Bptow6, n4474);  // ../RTL/cortexm0ds_logic.v(13746)
  and u16197 (Iptow6, Odgpw6[5], Pptow6);  // ../RTL/cortexm0ds_logic.v(13747)
  and u16198 (n4475, Wptow6, Dqtow6);  // ../RTL/cortexm0ds_logic.v(13748)
  not u16199 (Pptow6, n4475);  // ../RTL/cortexm0ds_logic.v(13748)
  buf u162 (Cjhpw6[0], Gpqpw6);  // ../RTL/cortexm0ds_logic.v(2365)
  and u1620 (Apihu6, Y41iu6, Gbjhu6);  // ../RTL/cortexm0ds_logic.v(3560)
  and u16200 (n4476, Kqtow6, R4gpw6[8]);  // ../RTL/cortexm0ds_logic.v(13749)
  not u16201 (Dqtow6, n4476);  // ../RTL/cortexm0ds_logic.v(13749)
  or u16202 (n4477, Rqtow6, R4gpw6[10]);  // ../RTL/cortexm0ds_logic.v(13750)
  not u16203 (Kqtow6, n4477);  // ../RTL/cortexm0ds_logic.v(13750)
  or u16204 (n4478, Yqtow6, R4gpw6[9]);  // ../RTL/cortexm0ds_logic.v(13751)
  not u16205 (Rqtow6, n4478);  // ../RTL/cortexm0ds_logic.v(13751)
  and u16206 (n4479, R4gpw6[9], Yqtow6);  // ../RTL/cortexm0ds_logic.v(13752)
  not u16207 (Wptow6, n4479);  // ../RTL/cortexm0ds_logic.v(13752)
  not u16208 (Hltow6, Zntow6);  // ../RTL/cortexm0ds_logic.v(13753)
  AL_MUX u16209 (
    .i0(Frtow6),
    .i1(Mrtow6),
    .sel(Hkgow6),
    .o(Zntow6));  // ../RTL/cortexm0ds_logic.v(13754)
  AL_MUX u1621 (
    .i0(vis_pc_o[21]),
    .i1(Fzdpw6),
    .sel(Ty0iu6),
    .o(Y41iu6));  // ../RTL/cortexm0ds_logic.v(3561)
  and u16210 (Hkgow6, Trtow6, Vbgpw6[6]);  // ../RTL/cortexm0ds_logic.v(13755)
  and u16211 (Trtow6, Odgpw6[6], Astow6);  // ../RTL/cortexm0ds_logic.v(13756)
  and u16212 (n4480, Hstow6, Egtow6);  // ../RTL/cortexm0ds_logic.v(13757)
  not u16213 (Astow6, n4480);  // ../RTL/cortexm0ds_logic.v(13757)
  and u16214 (Egtow6, Vbgpw6[7], Odgpw6[7]);  // ../RTL/cortexm0ds_logic.v(13758)
  and u16215 (Hstow6, Ostow6, Vstow6);  // ../RTL/cortexm0ds_logic.v(13759)
  and u16216 (n4481, Cttow6, Jttow6);  // ../RTL/cortexm0ds_logic.v(13760)
  not u16217 (Vstow6, n4481);  // ../RTL/cortexm0ds_logic.v(13760)
  or u16218 (Jttow6, Mrtow6, R4gpw6[15]);  // ../RTL/cortexm0ds_logic.v(13761)
  and u16219 (n4482, R4gpw6[12], Qttow6);  // ../RTL/cortexm0ds_logic.v(13762)
  and u1622 (Iqihu6, F51iu6, Y9jhu6);  // ../RTL/cortexm0ds_logic.v(3562)
  not u16220 (Cttow6, n4482);  // ../RTL/cortexm0ds_logic.v(13762)
  or u16221 (Ostow6, Frtow6, R4gpw6[13]);  // ../RTL/cortexm0ds_logic.v(13763)
  AL_MUX u16222 (
    .i0(Xttow6),
    .i1(Eutow6),
    .sel(Tjgow6),
    .o(Oetow6));  // ../RTL/cortexm0ds_logic.v(13764)
  and u16223 (P4fow6, Lutow6, Sutow6);  // ../RTL/cortexm0ds_logic.v(13765)
  not u16224 (Tjgow6, P4fow6);  // ../RTL/cortexm0ds_logic.v(13765)
  and u16225 (n4483, Zutow6, Gvtow6);  // ../RTL/cortexm0ds_logic.v(13766)
  not u16226 (Sutow6, n4483);  // ../RTL/cortexm0ds_logic.v(13766)
  and u16227 (n4484, Nvtow6, Uvtow6);  // ../RTL/cortexm0ds_logic.v(13767)
  not u16228 (Gvtow6, n4484);  // ../RTL/cortexm0ds_logic.v(13767)
  and u16229 (n4485, Bwtow6, Iwtow6);  // ../RTL/cortexm0ds_logic.v(13768)
  AL_MUX u1623 (
    .i0(vis_pc_o[22]),
    .i1(Mzdpw6),
    .sel(Ty0iu6),
    .o(F51iu6));  // ../RTL/cortexm0ds_logic.v(3563)
  not u16230 (Uvtow6, n4485);  // ../RTL/cortexm0ds_logic.v(13768)
  AL_MUX u16231 (
    .i0(R4gpw6[0]),
    .i1(R4gpw6[2]),
    .sel(Pwtow6),
    .o(Iwtow6));  // ../RTL/cortexm0ds_logic.v(13769)
  or u16232 (n4486, Tktow6, Wwtow6);  // ../RTL/cortexm0ds_logic.v(13770)
  not u16233 (Bwtow6, n4486);  // ../RTL/cortexm0ds_logic.v(13770)
  or u16234 (n4487, Dxtow6, Xttow6);  // ../RTL/cortexm0ds_logic.v(13771)
  not u16235 (Wwtow6, n4487);  // ../RTL/cortexm0ds_logic.v(13771)
  AL_MUX u16236 (
    .i0(R4gpw6[6]),
    .i1(R4gpw6[4]),
    .sel(Mjgow6),
    .o(Tktow6));  // ../RTL/cortexm0ds_logic.v(13772)
  buf u16237 (Edehu6, Ozkbx6[32]);  // ../RTL/cortexm0ds_logic.v(3176)
  and u16238 (n4488, Xttow6, Dxtow6);  // ../RTL/cortexm0ds_logic.v(13774)
  not u16239 (Nvtow6, n4488);  // ../RTL/cortexm0ds_logic.v(13774)
  and u1624 (Qrihu6, M51iu6, Q8jhu6);  // ../RTL/cortexm0ds_logic.v(3564)
  or u16240 (Zutow6, Nhtow6, Mjgow6);  // ../RTL/cortexm0ds_logic.v(13775)
  and u16241 (n4489, Pwtow6, Rxtow6);  // ../RTL/cortexm0ds_logic.v(13776)
  not u16242 (Lutow6, n4489);  // ../RTL/cortexm0ds_logic.v(13776)
  and u16243 (E1uow6, Vbgpw6[1], Odgpw6[1]);  // ../RTL/cortexm0ds_logic.v(13777)
  not u16244 (Rxtow6, E1uow6);  // ../RTL/cortexm0ds_logic.v(13777)
  not u16245 (Eutow6, Dxtow6);  // ../RTL/cortexm0ds_logic.v(13778)
  AL_MUX u16246 (
    .i0(Yxtow6),
    .i1(Fytow6),
    .sel(Mjgow6),
    .o(Dxtow6));  // ../RTL/cortexm0ds_logic.v(13779)
  and u16247 (Mjgow6, Mytow6, Vbgpw6[2]);  // ../RTL/cortexm0ds_logic.v(13780)
  and u16248 (Mytow6, Odgpw6[2], Tytow6);  // ../RTL/cortexm0ds_logic.v(13781)
  and u16249 (n4490, Aztow6, Nhtow6);  // ../RTL/cortexm0ds_logic.v(13782)
  AL_MUX u1625 (
    .i0(vis_pc_o[23]),
    .i1(Tzdpw6),
    .sel(Ty0iu6),
    .o(M51iu6));  // ../RTL/cortexm0ds_logic.v(3565)
  not u16250 (Tytow6, n4490);  // ../RTL/cortexm0ds_logic.v(13782)
  and u16251 (Nhtow6, Vbgpw6[3], Odgpw6[3]);  // ../RTL/cortexm0ds_logic.v(13783)
  and u16252 (Aztow6, Hztow6, Oztow6);  // ../RTL/cortexm0ds_logic.v(13784)
  and u16253 (n4491, Vztow6, C0uow6);  // ../RTL/cortexm0ds_logic.v(13785)
  not u16254 (Oztow6, n4491);  // ../RTL/cortexm0ds_logic.v(13785)
  or u16255 (C0uow6, Fytow6, R4gpw6[7]);  // ../RTL/cortexm0ds_logic.v(13786)
  or u16256 (Vztow6, J0uow6, R4gpw6[6]);  // ../RTL/cortexm0ds_logic.v(13787)
  or u16257 (Hztow6, Yxtow6, R4gpw6[5]);  // ../RTL/cortexm0ds_logic.v(13788)
  AL_MUX u16258 (
    .i0(R4gpw6[3]),
    .i1(R4gpw6[1]),
    .sel(Fjgow6),
    .o(Xttow6));  // ../RTL/cortexm0ds_logic.v(13789)
  buf u16259 (Q5mhu6, Nvkbx6[13]);  // ../RTL/cortexm0ds_logic.v(3137)
  and u1626 (Ysihu6, T51iu6, I7jhu6);  // ../RTL/cortexm0ds_logic.v(3566)
  and u16260 (Fjgow6, Q0uow6, Vbgpw6[0]);  // ../RTL/cortexm0ds_logic.v(13791)
  not u16261 (Pwtow6, Fjgow6);  // ../RTL/cortexm0ds_logic.v(13791)
  and u16262 (Q0uow6, Odgpw6[0], X0uow6);  // ../RTL/cortexm0ds_logic.v(13792)
  and u16263 (n4492, E1uow6, L1uow6);  // ../RTL/cortexm0ds_logic.v(13793)
  not u16264 (X0uow6, n4492);  // ../RTL/cortexm0ds_logic.v(13793)
  and u16265 (L1uow6, S1uow6, Z1uow6);  // ../RTL/cortexm0ds_logic.v(13794)
  and u16266 (n4493, G2uow6, N2uow6);  // ../RTL/cortexm0ds_logic.v(13795)
  not u16267 (Z1uow6, n4493);  // ../RTL/cortexm0ds_logic.v(13795)
  or u16268 (N2uow6, U2uow6, R4gpw6[3]);  // ../RTL/cortexm0ds_logic.v(13796)
  or u16269 (G2uow6, B3uow6, R4gpw6[2]);  // ../RTL/cortexm0ds_logic.v(13797)
  AL_MUX u1627 (
    .i0(vis_pc_o[24]),
    .i1(A0epw6),
    .sel(Ty0iu6),
    .o(T51iu6));  // ../RTL/cortexm0ds_logic.v(3567)
  and u16270 (n4494, R4gpw6[3], U2uow6);  // ../RTL/cortexm0ds_logic.v(13798)
  not u16271 (S1uow6, n4494);  // ../RTL/cortexm0ds_logic.v(13798)
  buf u16272 (Ighpw6[3], Jflpw6);  // ../RTL/cortexm0ds_logic.v(1840)
  and u16273 (L9tow6, I3uow6, Dctow6);  // ../RTL/cortexm0ds_logic.v(13800)
  and u16274 (n4495, K5fow6, P3uow6);  // ../RTL/cortexm0ds_logic.v(13801)
  not u16275 (Dctow6, n4495);  // ../RTL/cortexm0ds_logic.v(13801)
  and u16276 (n4496, W3uow6, D4uow6);  // ../RTL/cortexm0ds_logic.v(13802)
  not u16277 (P3uow6, n4496);  // ../RTL/cortexm0ds_logic.v(13802)
  buf u16278 (Ighpw6[2], Kalpw6);  // ../RTL/cortexm0ds_logic.v(1840)
  not u16279 (I3uow6, Rctow6);  // ../RTL/cortexm0ds_logic.v(13803)
  and u1628 (Guihu6, A61iu6, A6jhu6);  // ../RTL/cortexm0ds_logic.v(3568)
  buf u16280 (X6mhu6, Nvkbx6[12]);  // ../RTL/cortexm0ds_logic.v(3137)
  and u16281 (Nggow6, K4uow6, R4uow6);  // ../RTL/cortexm0ds_logic.v(13805)
  not u16282 (K5fow6, Nggow6);  // ../RTL/cortexm0ds_logic.v(13805)
  or u16283 (R4uow6, Y4uow6, F5uow6);  // ../RTL/cortexm0ds_logic.v(13806)
  or u16284 (Y4uow6, W4fow6, Bhgow6);  // ../RTL/cortexm0ds_logic.v(13807)
  and u16285 (n4497, M5uow6, T5uow6);  // ../RTL/cortexm0ds_logic.v(13808)
  not u16286 (K4uow6, n4497);  // ../RTL/cortexm0ds_logic.v(13808)
  and u16287 (n4498, Cftow6, A6uow6);  // ../RTL/cortexm0ds_logic.v(13809)
  not u16288 (T5uow6, n4498);  // ../RTL/cortexm0ds_logic.v(13809)
  not u16289 (A6uow6, Jftow6);  // ../RTL/cortexm0ds_logic.v(13810)
  AL_MUX u1629 (
    .i0(vis_pc_o[25]),
    .i1(H0epw6),
    .sel(Ty0iu6),
    .o(A61iu6));  // ../RTL/cortexm0ds_logic.v(3569)
  or u16290 (n4499, D5fow6, Whgow6);  // ../RTL/cortexm0ds_logic.v(13811)
  not u16291 (Cftow6, n4499);  // ../RTL/cortexm0ds_logic.v(13811)
  and u16292 (n4500, H6uow6, O6uow6);  // ../RTL/cortexm0ds_logic.v(13812)
  not u16293 (M5uow6, n4500);  // ../RTL/cortexm0ds_logic.v(13812)
  and u16294 (n4501, V6uow6, C7uow6);  // ../RTL/cortexm0ds_logic.v(13813)
  not u16295 (O6uow6, n4501);  // ../RTL/cortexm0ds_logic.v(13813)
  and u16296 (C7uow6, J7uow6, D4uow6);  // ../RTL/cortexm0ds_logic.v(13814)
  and u16297 (n4502, D5fow6, Q7uow6);  // ../RTL/cortexm0ds_logic.v(13815)
  not u16298 (D4uow6, n4502);  // ../RTL/cortexm0ds_logic.v(13815)
  buf u16299 (E8mhu6, Nvkbx6[11]);  // ../RTL/cortexm0ds_logic.v(3137)
  buf u163 (vis_r12_o[6], Hysax6);  // ../RTL/cortexm0ds_logic.v(2599)
  and u1630 (Ovihu6, H61iu6, S4jhu6);  // ../RTL/cortexm0ds_logic.v(3570)
  or u16300 (J7uow6, Tdtow6, X7uow6);  // ../RTL/cortexm0ds_logic.v(13817)
  and u16301 (V6uow6, Yctow6, W3uow6);  // ../RTL/cortexm0ds_logic.v(13818)
  and u16302 (n4503, E8uow6, Digow6);  // ../RTL/cortexm0ds_logic.v(13819)
  not u16303 (W3uow6, n4503);  // ../RTL/cortexm0ds_logic.v(13819)
  AL_MUX u16304 (
    .i0(L8uow6),
    .i1(S8uow6),
    .sel(W4fow6),
    .o(Yctow6));  // ../RTL/cortexm0ds_logic.v(13820)
  AL_MUX u16305 (
    .i0(R4gpw6[18]),
    .i1(R4gpw6[16]),
    .sel(Uggow6),
    .o(S8uow6));  // ../RTL/cortexm0ds_logic.v(13821)
  and u16306 (n4504, X7uow6, Tdtow6);  // ../RTL/cortexm0ds_logic.v(13822)
  not u16307 (H6uow6, n4504);  // ../RTL/cortexm0ds_logic.v(13822)
  AL_MUX u16308 (
    .i0(Z8uow6),
    .i1(G9uow6),
    .sel(Digow6),
    .o(Tdtow6));  // ../RTL/cortexm0ds_logic.v(13823)
  and u16309 (D5fow6, N9uow6, U9uow6);  // ../RTL/cortexm0ds_logic.v(13824)
  AL_MUX u1631 (
    .i0(vis_pc_o[26]),
    .i1(O0epw6),
    .sel(Ty0iu6),
    .o(H61iu6));  // ../RTL/cortexm0ds_logic.v(3571)
  not u16310 (Digow6, D5fow6);  // ../RTL/cortexm0ds_logic.v(13824)
  and u16311 (n4505, Bauow6, Iauow6);  // ../RTL/cortexm0ds_logic.v(13825)
  not u16312 (U9uow6, n4505);  // ../RTL/cortexm0ds_logic.v(13825)
  and u16313 (n4506, Pauow6, Wauow6);  // ../RTL/cortexm0ds_logic.v(13826)
  not u16314 (Iauow6, n4506);  // ../RTL/cortexm0ds_logic.v(13826)
  and u16315 (n4507, Dbuow6, Q7uow6);  // ../RTL/cortexm0ds_logic.v(13827)
  not u16316 (Wauow6, n4507);  // ../RTL/cortexm0ds_logic.v(13827)
  AL_MUX u16317 (
    .i0(R4gpw6[26]),
    .i1(R4gpw6[24]),
    .sel(Phgow6),
    .o(Q7uow6));  // ../RTL/cortexm0ds_logic.v(13828)
  or u16318 (n4508, E8uow6, Kbuow6);  // ../RTL/cortexm0ds_logic.v(13829)
  not u16319 (Dbuow6, n4508);  // ../RTL/cortexm0ds_logic.v(13829)
  and u1632 (Wwihu6, O61iu6, K3jhu6);  // ../RTL/cortexm0ds_logic.v(3572)
  or u16320 (n4509, G9uow6, Rbuow6);  // ../RTL/cortexm0ds_logic.v(13830)
  not u16321 (Kbuow6, n4509);  // ../RTL/cortexm0ds_logic.v(13830)
  AL_MUX u16322 (
    .i0(R4gpw6[30]),
    .i1(R4gpw6[28]),
    .sel(Whgow6),
    .o(E8uow6));  // ../RTL/cortexm0ds_logic.v(13831)
  and u16323 (n4510, Rbuow6, G9uow6);  // ../RTL/cortexm0ds_logic.v(13832)
  not u16324 (Pauow6, n4510);  // ../RTL/cortexm0ds_logic.v(13832)
  or u16325 (Bauow6, Jftow6, Whgow6);  // ../RTL/cortexm0ds_logic.v(13833)
  and u16326 (n4511, Ybuow6, Fcuow6);  // ../RTL/cortexm0ds_logic.v(13834)
  not u16327 (N9uow6, n4511);  // ../RTL/cortexm0ds_logic.v(13834)
  and u16328 (n4512, Vbgpw6[13], Odgpw6[13]);  // ../RTL/cortexm0ds_logic.v(13835)
  not u16329 (Fcuow6, n4512);  // ../RTL/cortexm0ds_logic.v(13835)
  AL_MUX u1633 (
    .i0(vis_pc_o[27]),
    .i1(V0epw6),
    .sel(Ty0iu6),
    .o(O61iu6));  // ../RTL/cortexm0ds_logic.v(3573)
  AL_MUX u16330 (
    .i0(Mcuow6),
    .i1(Tcuow6),
    .sel(Whgow6),
    .o(G9uow6));  // ../RTL/cortexm0ds_logic.v(13836)
  and u16331 (Whgow6, Aduow6, Vbgpw6[14]);  // ../RTL/cortexm0ds_logic.v(13837)
  and u16332 (Aduow6, Odgpw6[14], Hduow6);  // ../RTL/cortexm0ds_logic.v(13838)
  and u16333 (n4513, Oduow6, Jftow6);  // ../RTL/cortexm0ds_logic.v(13839)
  not u16334 (Hduow6, n4513);  // ../RTL/cortexm0ds_logic.v(13839)
  and u16335 (Jftow6, Vbgpw6[15], Odgpw6[15]);  // ../RTL/cortexm0ds_logic.v(13840)
  and u16336 (Oduow6, Vduow6, Ceuow6);  // ../RTL/cortexm0ds_logic.v(13841)
  and u16337 (n4514, Jeuow6, Qeuow6);  // ../RTL/cortexm0ds_logic.v(13842)
  not u16338 (Ceuow6, n4514);  // ../RTL/cortexm0ds_logic.v(13842)
  or u16339 (Qeuow6, Tcuow6, R4gpw6[31]);  // ../RTL/cortexm0ds_logic.v(13843)
  and u1634 (Eyihu6, V61iu6, C2jhu6);  // ../RTL/cortexm0ds_logic.v(3574)
  and u16340 (n4515, R4gpw6[28], Xeuow6);  // ../RTL/cortexm0ds_logic.v(13844)
  not u16341 (Jeuow6, n4515);  // ../RTL/cortexm0ds_logic.v(13844)
  not u16342 (Xeuow6, R4gpw6[30]);  // ../RTL/cortexm0ds_logic.v(13845)
  or u16343 (Vduow6, Mcuow6, R4gpw6[29]);  // ../RTL/cortexm0ds_logic.v(13846)
  not u16344 (Tcuow6, R4gpw6[29]);  // ../RTL/cortexm0ds_logic.v(13847)
  not u16345 (Z8uow6, Rbuow6);  // ../RTL/cortexm0ds_logic.v(13848)
  AL_MUX u16346 (
    .i0(R4gpw6[27]),
    .i1(R4gpw6[25]),
    .sel(Phgow6),
    .o(Rbuow6));  // ../RTL/cortexm0ds_logic.v(13849)
  buf u16347 (L9mhu6, Nvkbx6[10]);  // ../RTL/cortexm0ds_logic.v(3137)
  and u16348 (Phgow6, Efuow6, Vbgpw6[12]);  // ../RTL/cortexm0ds_logic.v(13851)
  not u16349 (Ybuow6, Phgow6);  // ../RTL/cortexm0ds_logic.v(13851)
  AL_MUX u1635 (
    .i0(vis_pc_o[28]),
    .i1(Dx0iu6),
    .sel(Ty0iu6),
    .o(V61iu6));  // ../RTL/cortexm0ds_logic.v(3575)
  and u16350 (Efuow6, Odgpw6[12], Lfuow6);  // ../RTL/cortexm0ds_logic.v(13852)
  and u16351 (n4516, Sfuow6, Vbgpw6[13]);  // ../RTL/cortexm0ds_logic.v(13853)
  not u16352 (Lfuow6, n4516);  // ../RTL/cortexm0ds_logic.v(13853)
  and u16353 (Sfuow6, Odgpw6[13], Zfuow6);  // ../RTL/cortexm0ds_logic.v(13854)
  and u16354 (n4517, Gguow6, Nguow6);  // ../RTL/cortexm0ds_logic.v(13855)
  not u16355 (Zfuow6, n4517);  // ../RTL/cortexm0ds_logic.v(13855)
  and u16356 (n4518, Uguow6, R4gpw6[24]);  // ../RTL/cortexm0ds_logic.v(13856)
  not u16357 (Nguow6, n4518);  // ../RTL/cortexm0ds_logic.v(13856)
  or u16358 (n4519, Bhuow6, R4gpw6[26]);  // ../RTL/cortexm0ds_logic.v(13857)
  not u16359 (Uguow6, n4519);  // ../RTL/cortexm0ds_logic.v(13857)
  and u1636 (Mzihu6, C71iu6, U0jhu6);  // ../RTL/cortexm0ds_logic.v(3576)
  or u16360 (n4520, Ihuow6, R4gpw6[25]);  // ../RTL/cortexm0ds_logic.v(13858)
  not u16361 (Bhuow6, n4520);  // ../RTL/cortexm0ds_logic.v(13858)
  and u16362 (n4521, R4gpw6[25], Ihuow6);  // ../RTL/cortexm0ds_logic.v(13859)
  not u16363 (Gguow6, n4521);  // ../RTL/cortexm0ds_logic.v(13859)
  not u16364 (X7uow6, Aetow6);  // ../RTL/cortexm0ds_logic.v(13860)
  AL_MUX u16365 (
    .i0(Phuow6),
    .i1(Whuow6),
    .sel(W4fow6),
    .o(Aetow6));  // ../RTL/cortexm0ds_logic.v(13861)
  buf u16366 (Samhu6, Nvkbx6[9]);  // ../RTL/cortexm0ds_logic.v(3137)
  and u16367 (W4fow6, Diuow6, Kiuow6);  // ../RTL/cortexm0ds_logic.v(13863)
  buf u16368 (Seehu6, Ozkbx6[31]);  // ../RTL/cortexm0ds_logic.v(3176)
  and u16369 (n4522, Riuow6, Yiuow6);  // ../RTL/cortexm0ds_logic.v(13864)
  AL_MUX u1637 (
    .i0(vis_pc_o[29]),
    .i1(Rx0iu6),
    .sel(Ty0iu6),
    .o(C71iu6));  // ../RTL/cortexm0ds_logic.v(3577)
  not u16370 (Kiuow6, n4522);  // ../RTL/cortexm0ds_logic.v(13864)
  and u16371 (n4523, Fjuow6, Mjuow6);  // ../RTL/cortexm0ds_logic.v(13865)
  not u16372 (Yiuow6, n4523);  // ../RTL/cortexm0ds_logic.v(13865)
  and u16373 (n4524, Tjuow6, Akuow6);  // ../RTL/cortexm0ds_logic.v(13866)
  not u16374 (Mjuow6, n4524);  // ../RTL/cortexm0ds_logic.v(13866)
  AL_MUX u16375 (
    .i0(R4gpw6[16]),
    .i1(R4gpw6[18]),
    .sel(Hkuow6),
    .o(Akuow6));  // ../RTL/cortexm0ds_logic.v(13867)
  or u16376 (n4525, L8uow6, Okuow6);  // ../RTL/cortexm0ds_logic.v(13868)
  not u16377 (Tjuow6, n4525);  // ../RTL/cortexm0ds_logic.v(13868)
  or u16378 (n4526, Vkuow6, Phuow6);  // ../RTL/cortexm0ds_logic.v(13869)
  not u16379 (Okuow6, n4526);  // ../RTL/cortexm0ds_logic.v(13869)
  and u1638 (Ttmhu6, V5hpw6[0], J71iu6);  // ../RTL/cortexm0ds_logic.v(3578)
  AL_MUX u16380 (
    .i0(R4gpw6[20]),
    .i1(R4gpw6[22]),
    .sel(Cluow6),
    .o(L8uow6));  // ../RTL/cortexm0ds_logic.v(13870)
  and u16381 (n4527, Phuow6, Vkuow6);  // ../RTL/cortexm0ds_logic.v(13871)
  not u16382 (Fjuow6, n4527);  // ../RTL/cortexm0ds_logic.v(13871)
  not u16383 (Vkuow6, Whuow6);  // ../RTL/cortexm0ds_logic.v(13872)
  or u16384 (Riuow6, F5uow6, Bhgow6);  // ../RTL/cortexm0ds_logic.v(13873)
  and u16385 (n4528, Hkuow6, Jluow6);  // ../RTL/cortexm0ds_logic.v(13874)
  not u16386 (Diuow6, n4528);  // ../RTL/cortexm0ds_logic.v(13874)
  and u16387 (Smuow6, Vbgpw6[9], Odgpw6[9]);  // ../RTL/cortexm0ds_logic.v(13875)
  not u16388 (Jluow6, Smuow6);  // ../RTL/cortexm0ds_logic.v(13875)
  AL_MUX u16389 (
    .i0(Qluow6),
    .i1(Xluow6),
    .sel(Uggow6),
    .o(Whuow6));  // ../RTL/cortexm0ds_logic.v(13876)
  and u1639 (Avmhu6, V5hpw6[1], Q71iu6);  // ../RTL/cortexm0ds_logic.v(3579)
  buf u16390 (Zbmhu6, Nvkbx6[8]);  // ../RTL/cortexm0ds_logic.v(3137)
  and u16391 (Uggow6, Emuow6, Vbgpw6[8]);  // ../RTL/cortexm0ds_logic.v(13878)
  not u16392 (Hkuow6, Uggow6);  // ../RTL/cortexm0ds_logic.v(13878)
  and u16393 (Emuow6, Odgpw6[8], Lmuow6);  // ../RTL/cortexm0ds_logic.v(13879)
  and u16394 (n4529, Smuow6, Zmuow6);  // ../RTL/cortexm0ds_logic.v(13880)
  not u16395 (Lmuow6, n4529);  // ../RTL/cortexm0ds_logic.v(13880)
  and u16396 (Zmuow6, Gnuow6, Nnuow6);  // ../RTL/cortexm0ds_logic.v(13881)
  and u16397 (n4530, Unuow6, Bouow6);  // ../RTL/cortexm0ds_logic.v(13882)
  not u16398 (Nnuow6, n4530);  // ../RTL/cortexm0ds_logic.v(13882)
  or u16399 (Bouow6, Xluow6, R4gpw6[19]);  // ../RTL/cortexm0ds_logic.v(13883)
  buf u164 (vis_psp_o[10], Bdjpw6);  // ../RTL/cortexm0ds_logic.v(2085)
  and u1640 (n123, X71iu6, Nv0iu6);  // ../RTL/cortexm0ds_logic.v(3580)
  or u16400 (Unuow6, Iouow6, R4gpw6[18]);  // ../RTL/cortexm0ds_logic.v(13884)
  or u16401 (Gnuow6, Qluow6, R4gpw6[17]);  // ../RTL/cortexm0ds_logic.v(13885)
  buf u16402 (Ighpw6[1], Sdlpw6);  // ../RTL/cortexm0ds_logic.v(1840)
  AL_MUX u16403 (
    .i0(Pouow6),
    .i1(Wouow6),
    .sel(Cluow6),
    .o(Phuow6));  // ../RTL/cortexm0ds_logic.v(13887)
  not u16404 (Cluow6, Bhgow6);  // ../RTL/cortexm0ds_logic.v(13888)
  and u16405 (Bhgow6, Dpuow6, Vbgpw6[10]);  // ../RTL/cortexm0ds_logic.v(13889)
  and u16406 (Dpuow6, Odgpw6[10], Kpuow6);  // ../RTL/cortexm0ds_logic.v(13890)
  and u16407 (n4531, Rpuow6, F5uow6);  // ../RTL/cortexm0ds_logic.v(13891)
  not u16408 (Kpuow6, n4531);  // ../RTL/cortexm0ds_logic.v(13891)
  and u16409 (F5uow6, Vbgpw6[11], Odgpw6[11]);  // ../RTL/cortexm0ds_logic.v(13892)
  not u1641 (Q71iu6, n123);  // ../RTL/cortexm0ds_logic.v(3580)
  and u16410 (Rpuow6, Ypuow6, Fquow6);  // ../RTL/cortexm0ds_logic.v(13893)
  and u16411 (n4532, Mquow6, Tquow6);  // ../RTL/cortexm0ds_logic.v(13894)
  not u16412 (Fquow6, n4532);  // ../RTL/cortexm0ds_logic.v(13894)
  or u16413 (Tquow6, Pouow6, R4gpw6[23]);  // ../RTL/cortexm0ds_logic.v(13895)
  or u16414 (Mquow6, Aruow6, R4gpw6[22]);  // ../RTL/cortexm0ds_logic.v(13896)
  or u16415 (Ypuow6, Wouow6, R4gpw6[21]);  // ../RTL/cortexm0ds_logic.v(13897)
  or u16416 (n4533, Qarow6, Xglow6);  // ../RTL/cortexm0ds_logic.v(13898)
  not u16417 (Ffrow6, n4533);  // ../RTL/cortexm0ds_logic.v(13898)
  and u16418 (Wdrow6, Zlghu6, Hruow6);  // ../RTL/cortexm0ds_logic.v(13899)
  not u16419 (Qarow6, Wdrow6);  // ../RTL/cortexm0ds_logic.v(13899)
  or u1642 (I5khu6, E81iu6, Aygpw6[0]);  // ../RTL/cortexm0ds_logic.v(3581)
  and u16420 (n4534, Oruow6, Vruow6);  // ../RTL/cortexm0ds_logic.v(13900)
  not u16421 (Hruow6, n4534);  // ../RTL/cortexm0ds_logic.v(13900)
  and u16422 (Vruow6, Csuow6, Jhqiu6);  // ../RTL/cortexm0ds_logic.v(13901)
  and u16423 (n4535, P9hhu6, Jehhu6);  // ../RTL/cortexm0ds_logic.v(13902)
  not u16424 (Jhqiu6, n4535);  // ../RTL/cortexm0ds_logic.v(13902)
  and u16425 (n4536, Jsuow6, Qsuow6);  // ../RTL/cortexm0ds_logic.v(13903)
  not u16426 (Csuow6, n4536);  // ../RTL/cortexm0ds_logic.v(13903)
  or u16427 (Qsuow6, F4oow6, L1gpw6[1]);  // ../RTL/cortexm0ds_logic.v(13904)
  or u16428 (Jsuow6, Xglow6, L1gpw6[0]);  // ../RTL/cortexm0ds_logic.v(13905)
  and u16429 (Oruow6, Ikghu6, Xsuow6);  // ../RTL/cortexm0ds_logic.v(13906)
  or u1643 (Q6khu6, E81iu6, Aygpw6[1]);  // ../RTL/cortexm0ds_logic.v(3582)
  and u16430 (n4537, L1gpw6[1], F4oow6);  // ../RTL/cortexm0ds_logic.v(13907)
  not u16431 (Xsuow6, n4537);  // ../RTL/cortexm0ds_logic.v(13907)
  not u16432 (F4oow6, B3gpw6[1]);  // ../RTL/cortexm0ds_logic.v(13908)
  AL_MUX u16433 (
    .i0(Oy8iu6),
    .i1(vis_primask_o),
    .sel(Cz8iu6),
    .o(K7row6));  // ../RTL/cortexm0ds_logic.v(13909)
  and u16434 (Cz8iu6, Etuow6, Ltuow6);  // ../RTL/cortexm0ds_logic.v(13910)
  and u16435 (n4538, Stuow6, Ztuow6);  // ../RTL/cortexm0ds_logic.v(13911)
  not u16436 (Ltuow6, n4538);  // ../RTL/cortexm0ds_logic.v(13911)
  and u16437 (Ztuow6, Cyfpw6[4], Gmniu6);  // ../RTL/cortexm0ds_logic.v(13912)
  and u16438 (n4539, Guuow6, Nuuow6);  // ../RTL/cortexm0ds_logic.v(13913)
  not u16439 (Gmniu6, n4539);  // ../RTL/cortexm0ds_logic.v(13913)
  or u1644 (Y7khu6, E81iu6, Aygpw6[2]);  // ../RTL/cortexm0ds_logic.v(3583)
  and u16440 (Nuuow6, Uuuow6, Bvuow6);  // ../RTL/cortexm0ds_logic.v(13914)
  or u16441 (Bvuow6, Ivuow6, Yoniu6);  // ../RTL/cortexm0ds_logic.v(13915)
  and u16442 (Yoniu6, Pvuow6, Wvuow6);  // ../RTL/cortexm0ds_logic.v(13916)
  and u16443 (n4540, Dwuow6, Kwuow6);  // ../RTL/cortexm0ds_logic.v(13917)
  not u16444 (Wvuow6, n4540);  // ../RTL/cortexm0ds_logic.v(13917)
  or u16445 (n4541, C0ehu6, H4ghu6);  // ../RTL/cortexm0ds_logic.v(13918)
  not u16446 (Dwuow6, n4541);  // ../RTL/cortexm0ds_logic.v(13918)
  or u16447 (n4542, Glaiu6, Rwuow6);  // ../RTL/cortexm0ds_logic.v(13919)
  not u16448 (Pvuow6, n4542);  // ../RTL/cortexm0ds_logic.v(13919)
  and u16449 (Rwuow6, Ywuow6, Fxuow6);  // ../RTL/cortexm0ds_logic.v(13920)
  or u1645 (G9khu6, E81iu6, Aygpw6[3]);  // ../RTL/cortexm0ds_logic.v(3584)
  or u16450 (n4543, Nlaiu6, Hs0iu6);  // ../RTL/cortexm0ds_logic.v(13921)
  not u16451 (Fxuow6, n4543);  // ../RTL/cortexm0ds_logic.v(13921)
  and u16452 (Ywuow6, Jf6ju6, Imaiu6);  // ../RTL/cortexm0ds_logic.v(13922)
  or u16453 (Uuuow6, Mxuow6, Mpniu6);  // ../RTL/cortexm0ds_logic.v(13923)
  and u16454 (Mpniu6, Txuow6, Ayuow6);  // ../RTL/cortexm0ds_logic.v(13924)
  and u16455 (Ayuow6, Hyuow6, Xiaju6);  // ../RTL/cortexm0ds_logic.v(13925)
  and u16456 (Xiaju6, Oyuow6, W8oiu6);  // ../RTL/cortexm0ds_logic.v(13926)
  and u16457 (n4544, Vyuow6, Ae0iu6);  // ../RTL/cortexm0ds_logic.v(13927)
  not u16458 (Oyuow6, n4544);  // ../RTL/cortexm0ds_logic.v(13927)
  and u16459 (Vyuow6, U4kiu6, Yljiu6);  // ../RTL/cortexm0ds_logic.v(13928)
  or u1646 (Oakhu6, E81iu6, Aygpw6[4]);  // ../RTL/cortexm0ds_logic.v(3585)
  and u16460 (Hyuow6, Czuow6, Jzuow6);  // ../RTL/cortexm0ds_logic.v(13929)
  or u16461 (Jzuow6, Z6oiu6, E4jiu6);  // ../RTL/cortexm0ds_logic.v(13930)
  not u16462 (Z6oiu6, Fhaiu6);  // ../RTL/cortexm0ds_logic.v(13931)
  and u16463 (n4545, Qzuow6, Cyfpw6[7]);  // ../RTL/cortexm0ds_logic.v(13932)
  not u16464 (Czuow6, n4545);  // ../RTL/cortexm0ds_logic.v(13932)
  and u16465 (Qzuow6, Cyfpw6[1], Xzuow6);  // ../RTL/cortexm0ds_logic.v(13933)
  and u16466 (n4546, E0vow6, Vwaiu6);  // ../RTL/cortexm0ds_logic.v(13934)
  not u16467 (Xzuow6, n4546);  // ../RTL/cortexm0ds_logic.v(13934)
  or u16468 (E0vow6, Y7ghu6, Cyfpw6[4]);  // ../RTL/cortexm0ds_logic.v(13935)
  and u16469 (Txuow6, L0vow6, S0vow6);  // ../RTL/cortexm0ds_logic.v(13936)
  and u1647 (Wbkhu6, Pzgpw6[0], J71iu6);  // ../RTL/cortexm0ds_logic.v(3586)
  AL_MUX u16470 (
    .i0(Z0vow6),
    .i1(G1vow6),
    .sel(Cyfpw6[4]),
    .o(S0vow6));  // ../RTL/cortexm0ds_logic.v(13937)
  or u16471 (G1vow6, Nlaiu6, Mr0iu6);  // ../RTL/cortexm0ds_logic.v(13938)
  or u16472 (Z0vow6, Qxaiu6, Cyfpw6[6]);  // ../RTL/cortexm0ds_logic.v(13939)
  and u16473 (L0vow6, N1vow6, U1vow6);  // ../RTL/cortexm0ds_logic.v(13940)
  and u16474 (n4547, Xe8iu6, B2vow6);  // ../RTL/cortexm0ds_logic.v(13941)
  not u16475 (U1vow6, n4547);  // ../RTL/cortexm0ds_logic.v(13941)
  or u16476 (B2vow6, U4kiu6, Vboiu6);  // ../RTL/cortexm0ds_logic.v(13942)
  or u16477 (N1vow6, Yn2ju6, Ii0iu6);  // ../RTL/cortexm0ds_logic.v(13943)
  and u16478 (Guuow6, Utniu6, I2vow6);  // ../RTL/cortexm0ds_logic.v(13944)
  and u16479 (n4548, S8fpw6[9], Wnniu6);  // ../RTL/cortexm0ds_logic.v(13945)
  and u1648 (Edkhu6, Pzgpw6[1], L81iu6);  // ../RTL/cortexm0ds_logic.v(3587)
  not u16480 (I2vow6, n4548);  // ../RTL/cortexm0ds_logic.v(13945)
  and u16481 (n4549, P2vow6, W2vow6);  // ../RTL/cortexm0ds_logic.v(13946)
  not u16482 (Wnniu6, n4549);  // ../RTL/cortexm0ds_logic.v(13946)
  or u16483 (n4550, Gz2ju6, Iugiu6);  // ../RTL/cortexm0ds_logic.v(13947)
  not u16484 (W2vow6, n4550);  // ../RTL/cortexm0ds_logic.v(13947)
  or u16485 (n4551, X5oiu6, Yn2ju6);  // ../RTL/cortexm0ds_logic.v(13948)
  not u16486 (Gz2ju6, n4551);  // ../RTL/cortexm0ds_logic.v(13948)
  not u16487 (Yn2ju6, Pfoiu6);  // ../RTL/cortexm0ds_logic.v(13949)
  not u16488 (X5oiu6, F9aju6);  // ../RTL/cortexm0ds_logic.v(13950)
  and u16489 (P2vow6, D3vow6, K3vow6);  // ../RTL/cortexm0ds_logic.v(13951)
  and u1649 (n124, X71iu6, Ty0iu6);  // ../RTL/cortexm0ds_logic.v(3588)
  and u16490 (n4552, R3vow6, Cyfpw6[4]);  // ../RTL/cortexm0ds_logic.v(13952)
  not u16491 (K3vow6, n4552);  // ../RTL/cortexm0ds_logic.v(13952)
  or u16492 (n4553, Lkaiu6, Tr0iu6);  // ../RTL/cortexm0ds_logic.v(13953)
  not u16493 (R3vow6, n4553);  // ../RTL/cortexm0ds_logic.v(13953)
  and u16494 (n4554, C0ehu6, Y3vow6);  // ../RTL/cortexm0ds_logic.v(13954)
  not u16495 (D3vow6, n4554);  // ../RTL/cortexm0ds_logic.v(13954)
  and u16496 (n4555, F4vow6, M4vow6);  // ../RTL/cortexm0ds_logic.v(13955)
  not u16497 (Y3vow6, n4555);  // ../RTL/cortexm0ds_logic.v(13955)
  or u16498 (M4vow6, G7oiu6, Hs0iu6);  // ../RTL/cortexm0ds_logic.v(13956)
  and u16499 (F4vow6, T4vow6, Ekaiu6);  // ../RTL/cortexm0ds_logic.v(13957)
  buf u165 (L1gpw6[0], Vpgbx6);  // ../RTL/cortexm0ds_logic.v(2191)
  not u1650 (L81iu6, n124);  // ../RTL/cortexm0ds_logic.v(3588)
  or u16500 (Ekaiu6, A4oiu6, Cyfpw6[0]);  // ../RTL/cortexm0ds_logic.v(13958)
  or u16501 (T4vow6, M32ju6, Tfjiu6);  // ../RTL/cortexm0ds_logic.v(13959)
  or u16502 (n4556, A5vow6, Fq8iu6);  // ../RTL/cortexm0ds_logic.v(13960)
  not u16503 (Utniu6, n4556);  // ../RTL/cortexm0ds_logic.v(13960)
  or u16504 (n4557, Mzlow6, C0ehu6);  // ../RTL/cortexm0ds_logic.v(13961)
  not u16505 (A5vow6, n4557);  // ../RTL/cortexm0ds_logic.v(13961)
  and u16506 (Etuow6, Vlliu6, H5vow6);  // ../RTL/cortexm0ds_logic.v(13962)
  and u16507 (n4558, O5vow6, Jjoiu6);  // ../RTL/cortexm0ds_logic.v(13963)
  not u16508 (H5vow6, n4558);  // ../RTL/cortexm0ds_logic.v(13963)
  and u16509 (Jjoiu6, B5kiu6, Qmliu6);  // ../RTL/cortexm0ds_logic.v(13964)
  and u1651 (Ufkhu6, S81iu6, Dmmhu6);  // ../RTL/cortexm0ds_logic.v(3589)
  not u16510 (B5kiu6, S8fpw6[2]);  // ../RTL/cortexm0ds_logic.v(13965)
  or u16511 (n4559, Wofiu6, Qjoiu6);  // ../RTL/cortexm0ds_logic.v(13966)
  not u16512 (O5vow6, n4559);  // ../RTL/cortexm0ds_logic.v(13966)
  and u16513 (n4560, V5vow6, S8fpw6[2]);  // ../RTL/cortexm0ds_logic.v(13967)
  not u16514 (Vlliu6, n4560);  // ../RTL/cortexm0ds_logic.v(13967)
  and u16515 (V5vow6, Qmliu6, Wofiu6);  // ../RTL/cortexm0ds_logic.v(13968)
  and u16516 (n4561, C6vow6, J6vow6);  // ../RTL/cortexm0ds_logic.v(13969)
  not u16517 (Oy8iu6, n4561);  // ../RTL/cortexm0ds_logic.v(13969)
  and u16518 (n4562, Stuow6, X3fpw6[1]);  // ../RTL/cortexm0ds_logic.v(13970)
  not u16519 (J6vow6, n4562);  // ../RTL/cortexm0ds_logic.v(13970)
  and u1652 (S81iu6, My0iu6, Nv0iu6);  // ../RTL/cortexm0ds_logic.v(3590)
  or u16520 (n4563, M32ju6, P1bow6);  // ../RTL/cortexm0ds_logic.v(13971)
  not u16521 (Stuow6, n4563);  // ../RTL/cortexm0ds_logic.v(13971)
  not u16522 (M32ju6, W2aow6);  // ../RTL/cortexm0ds_logic.v(13972)
  and u16523 (n4564, Qmliu6, L35ju6);  // ../RTL/cortexm0ds_logic.v(13973)
  not u16524 (C6vow6, n4564);  // ../RTL/cortexm0ds_logic.v(13973)
  and u16525 (n4565, Q6vow6, X6vow6);  // ../RTL/cortexm0ds_logic.v(13974)
  not u16526 (Qmliu6, n4565);  // ../RTL/cortexm0ds_logic.v(13974)
  and u16527 (n4566, E7vow6, Obbow6);  // ../RTL/cortexm0ds_logic.v(13975)
  not u16528 (X6vow6, n4566);  // ../RTL/cortexm0ds_logic.v(13975)
  or u16529 (n4567, A4oiu6, Cyfpw6[6]);  // ../RTL/cortexm0ds_logic.v(13976)
  and u1653 (Chkhu6, Z81iu6, Wkmhu6);  // ../RTL/cortexm0ds_logic.v(3591)
  not u16530 (E7vow6, n4567);  // ../RTL/cortexm0ds_logic.v(13976)
  not u16531 (A4oiu6, Pugiu6);  // ../RTL/cortexm0ds_logic.v(13977)
  or u16532 (Q6vow6, Kgaiu6, Ii0iu6);  // ../RTL/cortexm0ds_logic.v(13978)
  AL_MUX u16533 (
    .i0(Oodhu6),
    .i1(PORESETn),
    .sel(RSTBYPASS),
    .o(Fmdhu6));  // ../RTL/cortexm0ds_logic.v(13979)
  and u16534 (TXEV, L7vow6, Iugiu6);  // ../RTL/cortexm0ds_logic.v(13980)
  and u16535 (Iugiu6, S7vow6, Vo3ju6);  // ../RTL/cortexm0ds_logic.v(13981)
  or u16536 (n4568, Knaiu6, Cyfpw6[6]);  // ../RTL/cortexm0ds_logic.v(13982)
  not u16537 (S7vow6, n4568);  // ../RTL/cortexm0ds_logic.v(13982)
  and u16538 (L7vow6, Pt2ju6, Cyfpw6[4]);  // ../RTL/cortexm0ds_logic.v(13983)
  AL_MUX u16539 (
    .i0(Tonhu6),
    .i1(Hknhu6),
    .sel(Ujyhu6),
    .o(SWDO));  // ../RTL/cortexm0ds_logic.v(13984)
  AL_MUX u1654 (
    .i0(vis_pc_o[0]),
    .i1(Hz0iu6),
    .sel(Nv0iu6),
    .o(Z81iu6));  // ../RTL/cortexm0ds_logic.v(3592)
  not u16540 (Ujyhu6, Ighpw6[5]);  // ../RTL/cortexm0ds_logic.v(13985)
  and u16541 (n4569, HMASTER, Z7vow6);  // ../RTL/cortexm0ds_logic.v(13986)
  not u16542 (SPECHTRANS, n4569);  // ../RTL/cortexm0ds_logic.v(13986)
  and u16543 (n4570, Krzhu6, Ebxiu6);  // ../RTL/cortexm0ds_logic.v(13987)
  not u16544 (Z7vow6, n4570);  // ../RTL/cortexm0ds_logic.v(13987)
  and u16545 (SLEEPDEEP, SLEEPING, Ndghu6);  // ../RTL/cortexm0ds_logic.v(13988)
  not u16546 (HWRITE, G8vow6);  // ../RTL/cortexm0ds_logic.v(13989)
  AL_MUX u16547 (
    .i0(Ejpiu6),
    .i1(Sq4iu6),
    .sel(Xg6iu6),
    .o(G8vow6));  // ../RTL/cortexm0ds_logic.v(13990)
  and u16548 (Sq4iu6, Iqnhu6, Iqzhu6);  // ../RTL/cortexm0ds_logic.v(13991)
  and u16549 (Ejpiu6, N8vow6, U8vow6);  // ../RTL/cortexm0ds_logic.v(13992)
  and u1655 (Kikhu6, G91iu6, Pjmhu6);  // ../RTL/cortexm0ds_logic.v(3593)
  and u16550 (U8vow6, B9vow6, I9vow6);  // ../RTL/cortexm0ds_logic.v(13993)
  and u16551 (n4571, Xzmiu6, P9vow6);  // ../RTL/cortexm0ds_logic.v(13994)
  not u16552 (I9vow6, n4571);  // ../RTL/cortexm0ds_logic.v(13994)
  or u16553 (P9vow6, W9vow6, Bi0iu6);  // ../RTL/cortexm0ds_logic.v(13995)
  and u16554 (Bi0iu6, Wp0iu6, Y7ghu6);  // ../RTL/cortexm0ds_logic.v(13996)
  and u16555 (W9vow6, Kwuow6, Wp0iu6);  // ../RTL/cortexm0ds_logic.v(13997)
  or u16556 (n4572, Qjaiu6, Xkaow6);  // ../RTL/cortexm0ds_logic.v(13998)
  not u16557 (Kwuow6, n4572);  // ../RTL/cortexm0ds_logic.v(13998)
  and u16558 (n4573, Us2ju6, Davow6);  // ../RTL/cortexm0ds_logic.v(13999)
  not u16559 (B9vow6, n4573);  // ../RTL/cortexm0ds_logic.v(13999)
  AL_MUX u1656 (
    .i0(vis_pc_o[1]),
    .i1(Tugpw6[0]),
    .sel(Nv0iu6),
    .o(G91iu6));  // ../RTL/cortexm0ds_logic.v(3594)
  or u16560 (Davow6, Kavow6, Moaiu6);  // ../RTL/cortexm0ds_logic.v(14000)
  and u16561 (Moaiu6, D6kiu6, Y2oiu6);  // ../RTL/cortexm0ds_logic.v(14001)
  and u16562 (Kavow6, Ravow6, Ldoiu6);  // ../RTL/cortexm0ds_logic.v(14002)
  or u16563 (n4574, P1bow6, Sbghu6);  // ../RTL/cortexm0ds_logic.v(14003)
  not u16564 (Ravow6, n4574);  // ../RTL/cortexm0ds_logic.v(14003)
  and u16565 (Us2ju6, Cyfpw6[7], Gwyiu6);  // ../RTL/cortexm0ds_logic.v(14004)
  and u16566 (N8vow6, Lv7ow6, Yavow6);  // ../RTL/cortexm0ds_logic.v(14005)
  and u16567 (Lv7ow6, Fbvow6, Oe8ow6);  // ../RTL/cortexm0ds_logic.v(14006)
  and u16568 (n4575, Mbvow6, Ldoiu6);  // ../RTL/cortexm0ds_logic.v(14007)
  not u16569 (Fbvow6, n4575);  // ../RTL/cortexm0ds_logic.v(14007)
  and u1657 (Sjkhu6, N91iu6, Iimhu6);  // ../RTL/cortexm0ds_logic.v(3595)
  and u16570 (Mbvow6, Qe8iu6, H4ghu6);  // ../RTL/cortexm0ds_logic.v(14008)
  and u16571 (Tbvow6, Hcvow6, Ocvow6);  // ../RTL/cortexm0ds_logic.v(14010)
  and u16572 (n4576, Ym4iu6, R0nhu6);  // ../RTL/cortexm0ds_logic.v(14011)
  not u16573 (Ocvow6, n4576);  // ../RTL/cortexm0ds_logic.v(14011)
  and u16574 (Ym4iu6, Shhpw6[9], Iqzhu6);  // ../RTL/cortexm0ds_logic.v(14012)
  or u16575 (Hcvow6, Vcvow6, I28ju6);  // ../RTL/cortexm0ds_logic.v(14013)
  and u16576 (Cdvow6, Qdvow6, Xdvow6);  // ../RTL/cortexm0ds_logic.v(14015)
  and u16577 (n4577, Pl4iu6, R0nhu6);  // ../RTL/cortexm0ds_logic.v(14016)
  not u16578 (Xdvow6, n4577);  // ../RTL/cortexm0ds_logic.v(14016)
  and u16579 (Pl4iu6, Shhpw6[8], Iqzhu6);  // ../RTL/cortexm0ds_logic.v(14017)
  AL_MUX u1658 (
    .i0(vis_pc_o[2]),
    .i1(Tugpw6[1]),
    .sel(Nv0iu6),
    .o(N91iu6));  // ../RTL/cortexm0ds_logic.v(3596)
  or u16580 (Qdvow6, Vcvow6, Cz7ju6);  // ../RTL/cortexm0ds_logic.v(14018)
  and u16581 (n4578, Gk4iu6, R0nhu6);  // ../RTL/cortexm0ds_logic.v(14020)
  not u16582 (Levow6, n4578);  // ../RTL/cortexm0ds_logic.v(14020)
  and u16583 (Gk4iu6, Shhpw6[7], Iqzhu6);  // ../RTL/cortexm0ds_logic.v(14021)
  and u16584 (n4579, Sevow6, Uo6ju6);  // ../RTL/cortexm0ds_logic.v(14022)
  not u16585 (Eevow6, n4579);  // ../RTL/cortexm0ds_logic.v(14022)
  and u16586 (n4580, Xi4iu6, R0nhu6);  // ../RTL/cortexm0ds_logic.v(14024)
  not u16587 (Gfvow6, n4580);  // ../RTL/cortexm0ds_logic.v(14024)
  and u16588 (Xi4iu6, Shhpw6[6], Iqzhu6);  // ../RTL/cortexm0ds_logic.v(14025)
  and u16589 (n4581, Sevow6, Kj6ju6);  // ../RTL/cortexm0ds_logic.v(14026)
  and u1659 (Alkhu6, U91iu6, Bhmhu6);  // ../RTL/cortexm0ds_logic.v(3597)
  not u16590 (Zevow6, n4581);  // ../RTL/cortexm0ds_logic.v(14026)
  and u16591 (n4582, Oh4iu6, R0nhu6);  // ../RTL/cortexm0ds_logic.v(14028)
  not u16592 (Ufvow6, n4582);  // ../RTL/cortexm0ds_logic.v(14028)
  and u16593 (Oh4iu6, Shhpw6[5], Iqzhu6);  // ../RTL/cortexm0ds_logic.v(14029)
  and u16594 (n4583, Sevow6, Eg6ju6);  // ../RTL/cortexm0ds_logic.v(14030)
  not u16595 (Nfvow6, n4583);  // ../RTL/cortexm0ds_logic.v(14030)
  and u16596 (n4584, H34iu6, R0nhu6);  // ../RTL/cortexm0ds_logic.v(14032)
  not u16597 (Igvow6, n4584);  // ../RTL/cortexm0ds_logic.v(14032)
  and u16598 (H34iu6, Shhpw6[4], Iqzhu6);  // ../RTL/cortexm0ds_logic.v(14033)
  and u16599 (n4585, Sevow6, Zw4ju6);  // ../RTL/cortexm0ds_logic.v(14034)
  buf u166 (Dhgpw6[0], Lmkbx6);  // ../RTL/cortexm0ds_logic.v(2280)
  AL_MUX u1660 (
    .i0(vis_pc_o[3]),
    .i1(Tugpw6[2]),
    .sel(Nv0iu6),
    .o(U91iu6));  // ../RTL/cortexm0ds_logic.v(3598)
  not u16600 (Bgvow6, n4585);  // ../RTL/cortexm0ds_logic.v(14034)
  and u16601 (n4586, Df4iu6, R0nhu6);  // ../RTL/cortexm0ds_logic.v(14036)
  not u16602 (Wgvow6, n4586);  // ../RTL/cortexm0ds_logic.v(14036)
  and u16603 (Df4iu6, Shhpw6[3], Iqzhu6);  // ../RTL/cortexm0ds_logic.v(14037)
  and u16604 (n4587, Sevow6, G36ju6);  // ../RTL/cortexm0ds_logic.v(14038)
  not u16605 (Pgvow6, n4587);  // ../RTL/cortexm0ds_logic.v(14038)
  xor u16606 (n2661[0], J25ju6, Hu4ju6);  // ../RTL/cortexm0ds_logic.v(9500)
  not u16607 (CODEHINTDE[0], n5968[0]);  // ../RTL/cortexm0ds_logic.v(16977)
  and u16608 (Khvow6, Rhvow6, Yhvow6);  // ../RTL/cortexm0ds_logic.v(14040)
  and u16609 (n4588, Gdqow6, Aioiu6);  // ../RTL/cortexm0ds_logic.v(14041)
  and u1661 (Imkhu6, Ba1iu6, Ufmhu6);  // ../RTL/cortexm0ds_logic.v(3599)
  not u16610 (Yhvow6, n4588);  // ../RTL/cortexm0ds_logic.v(14041)
  and u16611 (n4589, Fivow6, Mivow6);  // ../RTL/cortexm0ds_logic.v(14042)
  not u16612 (Aioiu6, n4589);  // ../RTL/cortexm0ds_logic.v(14042)
  and u16613 (Mivow6, Tivow6, Ajvow6);  // ../RTL/cortexm0ds_logic.v(14043)
  and u16614 (Ajvow6, Hjvow6, Ojvow6);  // ../RTL/cortexm0ds_logic.v(14044)
  and u16615 (n4590, vis_r11_o[31], Ljqow6);  // ../RTL/cortexm0ds_logic.v(14045)
  not u16616 (Ojvow6, n4590);  // ../RTL/cortexm0ds_logic.v(14045)
  and u16617 (Hjvow6, Vjvow6, Ckvow6);  // ../RTL/cortexm0ds_logic.v(14046)
  and u16618 (n4591, vis_r9_o[31], Qiqow6);  // ../RTL/cortexm0ds_logic.v(14047)
  not u16619 (Ckvow6, n4591);  // ../RTL/cortexm0ds_logic.v(14047)
  AL_MUX u1662 (
    .i0(vis_pc_o[4]),
    .i1(Tugpw6[3]),
    .sel(Nv0iu6),
    .o(Ba1iu6));  // ../RTL/cortexm0ds_logic.v(3600)
  and u16620 (n4592, Fkfpw6[31], Dfqow6);  // ../RTL/cortexm0ds_logic.v(14048)
  not u16621 (Vjvow6, n4592);  // ../RTL/cortexm0ds_logic.v(14048)
  and u16622 (Tivow6, Jkvow6, Qkvow6);  // ../RTL/cortexm0ds_logic.v(14049)
  and u16623 (n4593, vis_r10_o[31], Sjqow6);  // ../RTL/cortexm0ds_logic.v(14050)
  not u16624 (Qkvow6, n4593);  // ../RTL/cortexm0ds_logic.v(14050)
  and u16625 (n4594, vis_psp_o[29], Yfqow6);  // ../RTL/cortexm0ds_logic.v(14051)
  not u16626 (Jkvow6, n4594);  // ../RTL/cortexm0ds_logic.v(14051)
  and u16627 (Fivow6, Xkvow6, Elvow6);  // ../RTL/cortexm0ds_logic.v(14052)
  and u16628 (Elvow6, Llvow6, Slvow6);  // ../RTL/cortexm0ds_logic.v(14053)
  and u16629 (n4595, vis_r12_o[31], Hhqow6);  // ../RTL/cortexm0ds_logic.v(14054)
  and u1663 (Qnkhu6, Ia1iu6, Nemhu6);  // ../RTL/cortexm0ds_logic.v(3601)
  not u16630 (Slvow6, n4595);  // ../RTL/cortexm0ds_logic.v(14054)
  and u16631 (Llvow6, Zlvow6, Gmvow6);  // ../RTL/cortexm0ds_logic.v(14055)
  and u16632 (n4596, vis_msp_o[29], Fgqow6);  // ../RTL/cortexm0ds_logic.v(14056)
  not u16633 (Gmvow6, n4596);  // ../RTL/cortexm0ds_logic.v(14056)
  and u16634 (n4597, vis_r14_o[31], Ahqow6);  // ../RTL/cortexm0ds_logic.v(14057)
  not u16635 (Zlvow6, n4597);  // ../RTL/cortexm0ds_logic.v(14057)
  and u16636 (Xkvow6, Bxzhu6, Nmvow6);  // ../RTL/cortexm0ds_logic.v(14058)
  and u16637 (n4598, vis_r8_o[31], Gkqow6);  // ../RTL/cortexm0ds_logic.v(14059)
  not u16638 (Nmvow6, n4598);  // ../RTL/cortexm0ds_logic.v(14059)
  and u16639 (Bxzhu6, Umvow6, Bnvow6);  // ../RTL/cortexm0ds_logic.v(14060)
  AL_MUX u1664 (
    .i0(vis_pc_o[5]),
    .i1(Tugpw6[4]),
    .sel(Nv0iu6),
    .o(Ia1iu6));  // ../RTL/cortexm0ds_logic.v(3602)
  and u16640 (Bnvow6, Invow6, Pnvow6);  // ../RTL/cortexm0ds_logic.v(14061)
  and u16641 (Pnvow6, Wnvow6, Dovow6);  // ../RTL/cortexm0ds_logic.v(14062)
  and u16642 (n4599, vis_r2_o[31], Dmqow6);  // ../RTL/cortexm0ds_logic.v(14063)
  not u16643 (Dovow6, n4599);  // ../RTL/cortexm0ds_logic.v(14063)
  and u16644 (n4600, vis_r6_o[31], Kmqow6);  // ../RTL/cortexm0ds_logic.v(14064)
  not u16645 (Wnvow6, n4600);  // ../RTL/cortexm0ds_logic.v(14064)
  and u16646 (Invow6, Kovow6, Rovow6);  // ../RTL/cortexm0ds_logic.v(14065)
  and u16647 (n4601, vis_r5_o[31], Fnqow6);  // ../RTL/cortexm0ds_logic.v(14066)
  not u16648 (Rovow6, n4601);  // ../RTL/cortexm0ds_logic.v(14066)
  and u16649 (n4602, vis_r4_o[31], Mnqow6);  // ../RTL/cortexm0ds_logic.v(14067)
  and u1665 (Yokhu6, Pa1iu6, Gdmhu6);  // ../RTL/cortexm0ds_logic.v(3603)
  not u16650 (Kovow6, n4602);  // ../RTL/cortexm0ds_logic.v(14067)
  and u16651 (Umvow6, Yovow6, Fpvow6);  // ../RTL/cortexm0ds_logic.v(14068)
  and u16652 (Fpvow6, Mpvow6, Tpvow6);  // ../RTL/cortexm0ds_logic.v(14069)
  and u16653 (n4603, vis_r1_o[31], Voqow6);  // ../RTL/cortexm0ds_logic.v(14070)
  not u16654 (Tpvow6, n4603);  // ../RTL/cortexm0ds_logic.v(14070)
  and u16655 (n4604, vis_r0_o[31], Cpqow6);  // ../RTL/cortexm0ds_logic.v(14071)
  not u16656 (Mpvow6, n4604);  // ../RTL/cortexm0ds_logic.v(14071)
  and u16657 (Yovow6, Aqvow6, Hqvow6);  // ../RTL/cortexm0ds_logic.v(14072)
  and u16658 (n4605, vis_r3_o[31], Xpqow6);  // ../RTL/cortexm0ds_logic.v(14073)
  not u16659 (Hqvow6, n4605);  // ../RTL/cortexm0ds_logic.v(14073)
  AL_MUX u1666 (
    .i0(vis_pc_o[6]),
    .i1(Tugpw6[5]),
    .sel(Nv0iu6),
    .o(Pa1iu6));  // ../RTL/cortexm0ds_logic.v(3604)
  and u16660 (n4606, vis_r7_o[31], Eqqow6);  // ../RTL/cortexm0ds_logic.v(14074)
  not u16661 (Aqvow6, n4606);  // ../RTL/cortexm0ds_logic.v(14074)
  and u16662 (n4607, R0nhu6, Lm1iu6);  // ../RTL/cortexm0ds_logic.v(14075)
  not u16663 (Rhvow6, n4607);  // ../RTL/cortexm0ds_logic.v(14075)
  and u16664 (Lm1iu6, Shhpw6[31], Iqzhu6);  // ../RTL/cortexm0ds_logic.v(14076)
  and u16665 (Dhvow6, Oqvow6, Vqvow6);  // ../RTL/cortexm0ds_logic.v(14077)
  and u16666 (n4608, K0row6, W89ju6);  // ../RTL/cortexm0ds_logic.v(14078)
  not u16667 (Vqvow6, n4608);  // ../RTL/cortexm0ds_logic.v(14078)
  and u16668 (Jrvow6, Qrvow6, Xrvow6);  // ../RTL/cortexm0ds_logic.v(14080)
  and u16669 (n4609, Gdqow6, T6liu6);  // ../RTL/cortexm0ds_logic.v(14081)
  and u1667 (Gqkhu6, Wa1iu6, Zbmhu6);  // ../RTL/cortexm0ds_logic.v(3605)
  not u16670 (Xrvow6, n4609);  // ../RTL/cortexm0ds_logic.v(14081)
  and u16671 (n4610, Esvow6, Lsvow6);  // ../RTL/cortexm0ds_logic.v(14082)
  not u16672 (T6liu6, n4610);  // ../RTL/cortexm0ds_logic.v(14082)
  and u16673 (Lsvow6, Ssvow6, Zsvow6);  // ../RTL/cortexm0ds_logic.v(14083)
  and u16674 (Zsvow6, Gtvow6, Ntvow6);  // ../RTL/cortexm0ds_logic.v(14084)
  and u16675 (n4611, vis_r11_o[30], Ljqow6);  // ../RTL/cortexm0ds_logic.v(14085)
  not u16676 (Ntvow6, n4611);  // ../RTL/cortexm0ds_logic.v(14085)
  and u16677 (Gtvow6, Utvow6, Buvow6);  // ../RTL/cortexm0ds_logic.v(14086)
  and u16678 (n4612, vis_r10_o[30], Sjqow6);  // ../RTL/cortexm0ds_logic.v(14087)
  not u16679 (Buvow6, n4612);  // ../RTL/cortexm0ds_logic.v(14087)
  AL_MUX u1668 (
    .i0(vis_pc_o[7]),
    .i1(Tugpw6[6]),
    .sel(Nv0iu6),
    .o(Wa1iu6));  // ../RTL/cortexm0ds_logic.v(3606)
  and u16680 (n4613, vis_r9_o[30], Qiqow6);  // ../RTL/cortexm0ds_logic.v(14088)
  not u16681 (Utvow6, n4613);  // ../RTL/cortexm0ds_logic.v(14088)
  and u16682 (Ssvow6, Iuvow6, Puvow6);  // ../RTL/cortexm0ds_logic.v(14089)
  and u16683 (n4614, Fkfpw6[30], Dfqow6);  // ../RTL/cortexm0ds_logic.v(14090)
  not u16684 (Puvow6, n4614);  // ../RTL/cortexm0ds_logic.v(14090)
  and u16685 (n4615, vis_r12_o[30], Hhqow6);  // ../RTL/cortexm0ds_logic.v(14091)
  not u16686 (Iuvow6, n4615);  // ../RTL/cortexm0ds_logic.v(14091)
  and u16687 (Esvow6, Wuvow6, Dvvow6);  // ../RTL/cortexm0ds_logic.v(14092)
  and u16688 (Dvvow6, Kvvow6, Rvvow6);  // ../RTL/cortexm0ds_logic.v(14093)
  and u16689 (n4616, vis_r14_o[30], Ahqow6);  // ../RTL/cortexm0ds_logic.v(14094)
  and u1669 (Orkhu6, Db1iu6, Samhu6);  // ../RTL/cortexm0ds_logic.v(3607)
  not u16690 (Rvvow6, n4616);  // ../RTL/cortexm0ds_logic.v(14094)
  and u16691 (Kvvow6, Yvvow6, Fwvow6);  // ../RTL/cortexm0ds_logic.v(14095)
  and u16692 (n4617, vis_psp_o[28], Yfqow6);  // ../RTL/cortexm0ds_logic.v(14096)
  not u16693 (Fwvow6, n4617);  // ../RTL/cortexm0ds_logic.v(14096)
  and u16694 (n4618, vis_r8_o[30], Gkqow6);  // ../RTL/cortexm0ds_logic.v(14097)
  not u16695 (Yvvow6, n4618);  // ../RTL/cortexm0ds_logic.v(14097)
  and u16696 (Wuvow6, Ixzhu6, Mwvow6);  // ../RTL/cortexm0ds_logic.v(14098)
  and u16697 (n4619, vis_msp_o[28], Fgqow6);  // ../RTL/cortexm0ds_logic.v(14099)
  not u16698 (Mwvow6, n4619);  // ../RTL/cortexm0ds_logic.v(14099)
  and u16699 (Ixzhu6, Twvow6, Axvow6);  // ../RTL/cortexm0ds_logic.v(14100)
  buf u167 (E1hpw6[13], Egaax6);  // ../RTL/cortexm0ds_logic.v(2367)
  AL_MUX u1670 (
    .i0(vis_pc_o[8]),
    .i1(Tugpw6[7]),
    .sel(Nv0iu6),
    .o(Db1iu6));  // ../RTL/cortexm0ds_logic.v(3608)
  and u16700 (Axvow6, Hxvow6, Oxvow6);  // ../RTL/cortexm0ds_logic.v(14101)
  and u16701 (Oxvow6, Vxvow6, Cyvow6);  // ../RTL/cortexm0ds_logic.v(14102)
  and u16702 (n4620, vis_r0_o[30], Cpqow6);  // ../RTL/cortexm0ds_logic.v(14103)
  not u16703 (Cyvow6, n4620);  // ../RTL/cortexm0ds_logic.v(14103)
  and u16704 (n4621, vis_r2_o[30], Dmqow6);  // ../RTL/cortexm0ds_logic.v(14104)
  not u16705 (Vxvow6, n4621);  // ../RTL/cortexm0ds_logic.v(14104)
  and u16706 (Hxvow6, Jyvow6, Qyvow6);  // ../RTL/cortexm0ds_logic.v(14105)
  and u16707 (n4622, vis_r5_o[30], Fnqow6);  // ../RTL/cortexm0ds_logic.v(14106)
  not u16708 (Qyvow6, n4622);  // ../RTL/cortexm0ds_logic.v(14106)
  and u16709 (n4623, vis_r4_o[30], Mnqow6);  // ../RTL/cortexm0ds_logic.v(14107)
  and u1671 (Wskhu6, Kb1iu6, L9mhu6);  // ../RTL/cortexm0ds_logic.v(3609)
  not u16710 (Jyvow6, n4623);  // ../RTL/cortexm0ds_logic.v(14107)
  and u16711 (Twvow6, Xyvow6, Ezvow6);  // ../RTL/cortexm0ds_logic.v(14108)
  and u16712 (Ezvow6, Lzvow6, Szvow6);  // ../RTL/cortexm0ds_logic.v(14109)
  and u16713 (n4624, vis_r7_o[30], Eqqow6);  // ../RTL/cortexm0ds_logic.v(14110)
  not u16714 (Szvow6, n4624);  // ../RTL/cortexm0ds_logic.v(14110)
  and u16715 (n4625, vis_r3_o[30], Xpqow6);  // ../RTL/cortexm0ds_logic.v(14111)
  not u16716 (Lzvow6, n4625);  // ../RTL/cortexm0ds_logic.v(14111)
  and u16717 (Xyvow6, Zzvow6, G0wow6);  // ../RTL/cortexm0ds_logic.v(14112)
  and u16718 (n4626, vis_r1_o[30], Voqow6);  // ../RTL/cortexm0ds_logic.v(14113)
  not u16719 (G0wow6, n4626);  // ../RTL/cortexm0ds_logic.v(14113)
  AL_MUX u1672 (
    .i0(vis_pc_o[9]),
    .i1(Tugpw6[8]),
    .sel(Nv0iu6),
    .o(Kb1iu6));  // ../RTL/cortexm0ds_logic.v(3610)
  and u16720 (n4627, vis_r6_o[30], Kmqow6);  // ../RTL/cortexm0ds_logic.v(14114)
  not u16721 (Zzvow6, n4627);  // ../RTL/cortexm0ds_logic.v(14114)
  or u16722 (Qrvow6, Naliu6, Qaxiu6);  // ../RTL/cortexm0ds_logic.v(14115)
  not u16723 (Naliu6, T94iu6);  // ../RTL/cortexm0ds_logic.v(14116)
  and u16724 (T94iu6, Shhpw6[30], Iqzhu6);  // ../RTL/cortexm0ds_logic.v(14117)
  and u16725 (Crvow6, N0wow6, U0wow6);  // ../RTL/cortexm0ds_logic.v(14118)
  and u16726 (n4628, K0row6, T39ju6);  // ../RTL/cortexm0ds_logic.v(14119)
  not u16727 (U0wow6, n4628);  // ../RTL/cortexm0ds_logic.v(14119)
  and u16728 (n4629, Ud4iu6, R0nhu6);  // ../RTL/cortexm0ds_logic.v(14121)
  not u16729 (I1wow6, n4629);  // ../RTL/cortexm0ds_logic.v(14121)
  and u1673 (Eukhu6, Rb1iu6, E8mhu6);  // ../RTL/cortexm0ds_logic.v(3611)
  and u16730 (Ud4iu6, Shhpw6[2], Iqzhu6);  // ../RTL/cortexm0ds_logic.v(14122)
  and u16731 (n4630, Sevow6, Ot5ju6);  // ../RTL/cortexm0ds_logic.v(14123)
  not u16732 (B1wow6, n4630);  // ../RTL/cortexm0ds_logic.v(14123)
  and u16733 (W1wow6, D2wow6, K2wow6);  // ../RTL/cortexm0ds_logic.v(14125)
  and u16734 (n4631, Gdqow6, Po7ju6);  // ../RTL/cortexm0ds_logic.v(14126)
  not u16735 (K2wow6, n4631);  // ../RTL/cortexm0ds_logic.v(14126)
  and u16736 (Mbniu6, R2wow6, Y2wow6);  // ../RTL/cortexm0ds_logic.v(14127)
  not u16737 (Po7ju6, Mbniu6);  // ../RTL/cortexm0ds_logic.v(14127)
  and u16738 (Y2wow6, F3wow6, M3wow6);  // ../RTL/cortexm0ds_logic.v(14128)
  and u16739 (M3wow6, T3wow6, A4wow6);  // ../RTL/cortexm0ds_logic.v(14129)
  AL_MUX u1674 (
    .i0(vis_pc_o[10]),
    .i1(Tugpw6[9]),
    .sel(Nv0iu6),
    .o(Rb1iu6));  // ../RTL/cortexm0ds_logic.v(3612)
  and u16740 (n4632, vis_r11_o[28], Ljqow6);  // ../RTL/cortexm0ds_logic.v(14130)
  not u16741 (A4wow6, n4632);  // ../RTL/cortexm0ds_logic.v(14130)
  and u16742 (T3wow6, H4wow6, O4wow6);  // ../RTL/cortexm0ds_logic.v(14131)
  and u16743 (n4633, vis_r10_o[28], Sjqow6);  // ../RTL/cortexm0ds_logic.v(14132)
  not u16744 (O4wow6, n4633);  // ../RTL/cortexm0ds_logic.v(14132)
  and u16745 (n4634, vis_r9_o[28], Qiqow6);  // ../RTL/cortexm0ds_logic.v(14133)
  not u16746 (H4wow6, n4634);  // ../RTL/cortexm0ds_logic.v(14133)
  and u16747 (F3wow6, V4wow6, C5wow6);  // ../RTL/cortexm0ds_logic.v(14134)
  and u16748 (n4635, Fkfpw6[28], Dfqow6);  // ../RTL/cortexm0ds_logic.v(14135)
  not u16749 (C5wow6, n4635);  // ../RTL/cortexm0ds_logic.v(14135)
  and u1675 (Mvkhu6, Yb1iu6, X6mhu6);  // ../RTL/cortexm0ds_logic.v(3613)
  and u16750 (n4636, vis_r12_o[28], Hhqow6);  // ../RTL/cortexm0ds_logic.v(14136)
  not u16751 (V4wow6, n4636);  // ../RTL/cortexm0ds_logic.v(14136)
  and u16752 (R2wow6, J5wow6, Q5wow6);  // ../RTL/cortexm0ds_logic.v(14137)
  and u16753 (Q5wow6, X5wow6, E6wow6);  // ../RTL/cortexm0ds_logic.v(14138)
  and u16754 (n4637, vis_r14_o[28], Ahqow6);  // ../RTL/cortexm0ds_logic.v(14139)
  not u16755 (E6wow6, n4637);  // ../RTL/cortexm0ds_logic.v(14139)
  and u16756 (X5wow6, L6wow6, S6wow6);  // ../RTL/cortexm0ds_logic.v(14140)
  and u16757 (n4638, vis_psp_o[26], Yfqow6);  // ../RTL/cortexm0ds_logic.v(14141)
  not u16758 (S6wow6, n4638);  // ../RTL/cortexm0ds_logic.v(14141)
  and u16759 (n4639, vis_r8_o[28], Gkqow6);  // ../RTL/cortexm0ds_logic.v(14142)
  AL_MUX u1676 (
    .i0(vis_pc_o[11]),
    .i1(Ixdpw6),
    .sel(Nv0iu6),
    .o(Yb1iu6));  // ../RTL/cortexm0ds_logic.v(3614)
  not u16760 (L6wow6, n4639);  // ../RTL/cortexm0ds_logic.v(14142)
  and u16761 (J5wow6, Dyzhu6, Z6wow6);  // ../RTL/cortexm0ds_logic.v(14143)
  and u16762 (n4640, vis_msp_o[26], Fgqow6);  // ../RTL/cortexm0ds_logic.v(14144)
  not u16763 (Z6wow6, n4640);  // ../RTL/cortexm0ds_logic.v(14144)
  and u16764 (Dyzhu6, G7wow6, N7wow6);  // ../RTL/cortexm0ds_logic.v(14145)
  and u16765 (N7wow6, U7wow6, B8wow6);  // ../RTL/cortexm0ds_logic.v(14146)
  and u16766 (B8wow6, I8wow6, P8wow6);  // ../RTL/cortexm0ds_logic.v(14147)
  and u16767 (n4641, vis_r0_o[28], Cpqow6);  // ../RTL/cortexm0ds_logic.v(14148)
  not u16768 (P8wow6, n4641);  // ../RTL/cortexm0ds_logic.v(14148)
  and u16769 (n4642, vis_r2_o[28], Dmqow6);  // ../RTL/cortexm0ds_logic.v(14149)
  and u1677 (Uwkhu6, Fc1iu6, Q5mhu6);  // ../RTL/cortexm0ds_logic.v(3615)
  not u16770 (I8wow6, n4642);  // ../RTL/cortexm0ds_logic.v(14149)
  and u16771 (U7wow6, W8wow6, D9wow6);  // ../RTL/cortexm0ds_logic.v(14150)
  and u16772 (n4643, vis_r5_o[28], Fnqow6);  // ../RTL/cortexm0ds_logic.v(14151)
  not u16773 (D9wow6, n4643);  // ../RTL/cortexm0ds_logic.v(14151)
  and u16774 (n4644, vis_r4_o[28], Mnqow6);  // ../RTL/cortexm0ds_logic.v(14152)
  not u16775 (W8wow6, n4644);  // ../RTL/cortexm0ds_logic.v(14152)
  and u16776 (G7wow6, K9wow6, R9wow6);  // ../RTL/cortexm0ds_logic.v(14153)
  and u16777 (R9wow6, Y9wow6, Fawow6);  // ../RTL/cortexm0ds_logic.v(14154)
  and u16778 (n4645, vis_r7_o[28], Eqqow6);  // ../RTL/cortexm0ds_logic.v(14155)
  not u16779 (Fawow6, n4645);  // ../RTL/cortexm0ds_logic.v(14155)
  AL_MUX u1678 (
    .i0(vis_pc_o[12]),
    .i1(Tugpw6[11]),
    .sel(Nv0iu6),
    .o(Fc1iu6));  // ../RTL/cortexm0ds_logic.v(3616)
  and u16780 (n4646, vis_r3_o[28], Xpqow6);  // ../RTL/cortexm0ds_logic.v(14156)
  not u16781 (Y9wow6, n4646);  // ../RTL/cortexm0ds_logic.v(14156)
  and u16782 (K9wow6, Mawow6, Tawow6);  // ../RTL/cortexm0ds_logic.v(14157)
  and u16783 (n4647, vis_r1_o[28], Voqow6);  // ../RTL/cortexm0ds_logic.v(14158)
  not u16784 (Tawow6, n4647);  // ../RTL/cortexm0ds_logic.v(14158)
  and u16785 (n4648, vis_r6_o[28], Kmqow6);  // ../RTL/cortexm0ds_logic.v(14159)
  not u16786 (Mawow6, n4648);  // ../RTL/cortexm0ds_logic.v(14159)
  or u16787 (D2wow6, Zeniu6, Qaxiu6);  // ../RTL/cortexm0ds_logic.v(14160)
  not u16788 (Zeniu6, F94iu6);  // ../RTL/cortexm0ds_logic.v(14161)
  and u16789 (F94iu6, Shhpw6[28], Iqzhu6);  // ../RTL/cortexm0ds_logic.v(14162)
  and u1679 (Cykhu6, Mc1iu6, J4mhu6);  // ../RTL/cortexm0ds_logic.v(3617)
  and u16790 (P1wow6, Abwow6, Hbwow6);  // ../RTL/cortexm0ds_logic.v(14163)
  and u16791 (n4649, K0row6, Rv8ju6);  // ../RTL/cortexm0ds_logic.v(14164)
  not u16792 (Hbwow6, n4649);  // ../RTL/cortexm0ds_logic.v(14164)
  and u16793 (Vbwow6, Ccwow6, Jcwow6);  // ../RTL/cortexm0ds_logic.v(14166)
  and u16794 (n4650, Gdqow6, A67ju6);  // ../RTL/cortexm0ds_logic.v(14167)
  not u16795 (Jcwow6, n4650);  // ../RTL/cortexm0ds_logic.v(14167)
  and u16796 (n4651, Qcwow6, Xcwow6);  // ../RTL/cortexm0ds_logic.v(14168)
  not u16797 (A67ju6, n4651);  // ../RTL/cortexm0ds_logic.v(14168)
  and u16798 (Xcwow6, Edwow6, Ldwow6);  // ../RTL/cortexm0ds_logic.v(14169)
  and u16799 (Ldwow6, Sdwow6, Zdwow6);  // ../RTL/cortexm0ds_logic.v(14170)
  buf u168 (E1hpw6[14], Nmabx6);  // ../RTL/cortexm0ds_logic.v(2367)
  AL_MUX u1680 (
    .i0(vis_pc_o[13]),
    .i1(Tugpw6[12]),
    .sel(Nv0iu6),
    .o(Mc1iu6));  // ../RTL/cortexm0ds_logic.v(3618)
  and u16800 (n4652, Fkfpw6[27], Dfqow6);  // ../RTL/cortexm0ds_logic.v(14171)
  not u16801 (Zdwow6, n4652);  // ../RTL/cortexm0ds_logic.v(14171)
  and u16802 (Sdwow6, Gewow6, Newow6);  // ../RTL/cortexm0ds_logic.v(14172)
  and u16803 (n4653, vis_psp_o[25], Yfqow6);  // ../RTL/cortexm0ds_logic.v(14173)
  not u16804 (Newow6, n4653);  // ../RTL/cortexm0ds_logic.v(14173)
  and u16805 (n4654, vis_msp_o[25], Fgqow6);  // ../RTL/cortexm0ds_logic.v(14174)
  not u16806 (Gewow6, n4654);  // ../RTL/cortexm0ds_logic.v(14174)
  and u16807 (Edwow6, Uewow6, Bfwow6);  // ../RTL/cortexm0ds_logic.v(14175)
  and u16808 (n4655, vis_r14_o[27], Ahqow6);  // ../RTL/cortexm0ds_logic.v(14176)
  not u16809 (Bfwow6, n4655);  // ../RTL/cortexm0ds_logic.v(14176)
  and u1681 (Kzkhu6, Tc1iu6, C3mhu6);  // ../RTL/cortexm0ds_logic.v(3619)
  and u16810 (n4656, vis_r12_o[27], Hhqow6);  // ../RTL/cortexm0ds_logic.v(14177)
  not u16811 (Uewow6, n4656);  // ../RTL/cortexm0ds_logic.v(14177)
  and u16812 (Qcwow6, Ifwow6, Pfwow6);  // ../RTL/cortexm0ds_logic.v(14178)
  and u16813 (Pfwow6, Wfwow6, Dgwow6);  // ../RTL/cortexm0ds_logic.v(14179)
  and u16814 (n4657, vis_r9_o[27], Qiqow6);  // ../RTL/cortexm0ds_logic.v(14180)
  not u16815 (Dgwow6, n4657);  // ../RTL/cortexm0ds_logic.v(14180)
  and u16816 (Wfwow6, Kgwow6, Rgwow6);  // ../RTL/cortexm0ds_logic.v(14181)
  and u16817 (n4658, vis_r11_o[27], Ljqow6);  // ../RTL/cortexm0ds_logic.v(14182)
  not u16818 (Rgwow6, n4658);  // ../RTL/cortexm0ds_logic.v(14182)
  and u16819 (n4659, vis_r10_o[27], Sjqow6);  // ../RTL/cortexm0ds_logic.v(14183)
  AL_MUX u1682 (
    .i0(vis_pc_o[14]),
    .i1(Tugpw6[13]),
    .sel(Nv0iu6),
    .o(Tc1iu6));  // ../RTL/cortexm0ds_logic.v(3620)
  not u16820 (Kgwow6, n4659);  // ../RTL/cortexm0ds_logic.v(14183)
  and u16821 (Ifwow6, Kyzhu6, Ygwow6);  // ../RTL/cortexm0ds_logic.v(14184)
  and u16822 (n4660, vis_r8_o[27], Gkqow6);  // ../RTL/cortexm0ds_logic.v(14185)
  not u16823 (Ygwow6, n4660);  // ../RTL/cortexm0ds_logic.v(14185)
  and u16824 (Kyzhu6, Fhwow6, Mhwow6);  // ../RTL/cortexm0ds_logic.v(14186)
  and u16825 (Mhwow6, Thwow6, Aiwow6);  // ../RTL/cortexm0ds_logic.v(14187)
  and u16826 (Aiwow6, Hiwow6, Oiwow6);  // ../RTL/cortexm0ds_logic.v(14188)
  and u16827 (n4661, vis_r2_o[27], Dmqow6);  // ../RTL/cortexm0ds_logic.v(14189)
  not u16828 (Oiwow6, n4661);  // ../RTL/cortexm0ds_logic.v(14189)
  and u16829 (n4662, vis_r6_o[27], Kmqow6);  // ../RTL/cortexm0ds_logic.v(14190)
  and u1683 (S0lhu6, Ad1iu6, V1mhu6);  // ../RTL/cortexm0ds_logic.v(3621)
  not u16830 (Hiwow6, n4662);  // ../RTL/cortexm0ds_logic.v(14190)
  and u16831 (Thwow6, Viwow6, Cjwow6);  // ../RTL/cortexm0ds_logic.v(14191)
  and u16832 (n4663, vis_r5_o[27], Fnqow6);  // ../RTL/cortexm0ds_logic.v(14192)
  not u16833 (Cjwow6, n4663);  // ../RTL/cortexm0ds_logic.v(14192)
  and u16834 (n4664, vis_r4_o[27], Mnqow6);  // ../RTL/cortexm0ds_logic.v(14193)
  not u16835 (Viwow6, n4664);  // ../RTL/cortexm0ds_logic.v(14193)
  and u16836 (Fhwow6, Jjwow6, Qjwow6);  // ../RTL/cortexm0ds_logic.v(14194)
  and u16837 (Qjwow6, Xjwow6, Ekwow6);  // ../RTL/cortexm0ds_logic.v(14195)
  and u16838 (n4665, vis_r1_o[27], Voqow6);  // ../RTL/cortexm0ds_logic.v(14196)
  not u16839 (Ekwow6, n4665);  // ../RTL/cortexm0ds_logic.v(14196)
  AL_MUX u1684 (
    .i0(vis_pc_o[15]),
    .i1(Pxdpw6),
    .sel(Nv0iu6),
    .o(Ad1iu6));  // ../RTL/cortexm0ds_logic.v(3622)
  and u16840 (n4666, vis_r0_o[27], Cpqow6);  // ../RTL/cortexm0ds_logic.v(14197)
  not u16841 (Xjwow6, n4666);  // ../RTL/cortexm0ds_logic.v(14197)
  and u16842 (Jjwow6, Lkwow6, Skwow6);  // ../RTL/cortexm0ds_logic.v(14198)
  and u16843 (n4667, vis_r3_o[27], Xpqow6);  // ../RTL/cortexm0ds_logic.v(14199)
  not u16844 (Skwow6, n4667);  // ../RTL/cortexm0ds_logic.v(14199)
  and u16845 (n4668, vis_r7_o[27], Eqqow6);  // ../RTL/cortexm0ds_logic.v(14200)
  not u16846 (Lkwow6, n4668);  // ../RTL/cortexm0ds_logic.v(14200)
  or u16847 (Ccwow6, U3liu6, Qaxiu6);  // ../RTL/cortexm0ds_logic.v(14201)
  not u16848 (U3liu6, Y84iu6);  // ../RTL/cortexm0ds_logic.v(14202)
  and u16849 (Y84iu6, Shhpw6[27], Iqzhu6);  // ../RTL/cortexm0ds_logic.v(14203)
  and u1685 (A2lhu6, Hd1iu6, O0mhu6);  // ../RTL/cortexm0ds_logic.v(3623)
  and u16850 (Obwow6, Zkwow6, Glwow6);  // ../RTL/cortexm0ds_logic.v(14204)
  and u16851 (n4669, K0row6, In8ju6);  // ../RTL/cortexm0ds_logic.v(14205)
  not u16852 (Glwow6, n4669);  // ../RTL/cortexm0ds_logic.v(14205)
  buf u16853 (Gdmhu6, Nvkbx6[7]);  // ../RTL/cortexm0ds_logic.v(3137)
  and u16854 (Bmwow6, Imwow6, Pmwow6);  // ../RTL/cortexm0ds_logic.v(14208)
  and u16855 (n4670, Gdqow6, Z17ju6);  // ../RTL/cortexm0ds_logic.v(14209)
  not u16856 (Pmwow6, n4670);  // ../RTL/cortexm0ds_logic.v(14209)
  and u16857 (n4671, Wmwow6, Dnwow6);  // ../RTL/cortexm0ds_logic.v(14210)
  not u16858 (Z17ju6, n4671);  // ../RTL/cortexm0ds_logic.v(14210)
  and u16859 (Dnwow6, Knwow6, Rnwow6);  // ../RTL/cortexm0ds_logic.v(14211)
  AL_MUX u1686 (
    .i0(vis_pc_o[16]),
    .i1(Wxdpw6),
    .sel(Nv0iu6),
    .o(Hd1iu6));  // ../RTL/cortexm0ds_logic.v(3624)
  and u16860 (Rnwow6, Ynwow6, Fowow6);  // ../RTL/cortexm0ds_logic.v(14212)
  and u16861 (n4672, Fkfpw6[26], Dfqow6);  // ../RTL/cortexm0ds_logic.v(14213)
  not u16862 (Fowow6, n4672);  // ../RTL/cortexm0ds_logic.v(14213)
  and u16863 (Ynwow6, Mowow6, Towow6);  // ../RTL/cortexm0ds_logic.v(14214)
  and u16864 (n4673, vis_psp_o[24], Yfqow6);  // ../RTL/cortexm0ds_logic.v(14215)
  not u16865 (Towow6, n4673);  // ../RTL/cortexm0ds_logic.v(14215)
  and u16866 (n4674, vis_msp_o[24], Fgqow6);  // ../RTL/cortexm0ds_logic.v(14216)
  not u16867 (Mowow6, n4674);  // ../RTL/cortexm0ds_logic.v(14216)
  and u16868 (Knwow6, Apwow6, Hpwow6);  // ../RTL/cortexm0ds_logic.v(14217)
  and u16869 (n4675, vis_r14_o[26], Ahqow6);  // ../RTL/cortexm0ds_logic.v(14218)
  and u1687 (I3lhu6, Od1iu6, Hzlhu6);  // ../RTL/cortexm0ds_logic.v(3625)
  not u16870 (Hpwow6, n4675);  // ../RTL/cortexm0ds_logic.v(14218)
  and u16871 (n4676, vis_r12_o[26], Hhqow6);  // ../RTL/cortexm0ds_logic.v(14219)
  not u16872 (Apwow6, n4676);  // ../RTL/cortexm0ds_logic.v(14219)
  and u16873 (Wmwow6, Opwow6, Vpwow6);  // ../RTL/cortexm0ds_logic.v(14220)
  and u16874 (Vpwow6, Cqwow6, Jqwow6);  // ../RTL/cortexm0ds_logic.v(14221)
  and u16875 (n4677, vis_r9_o[26], Qiqow6);  // ../RTL/cortexm0ds_logic.v(14222)
  not u16876 (Jqwow6, n4677);  // ../RTL/cortexm0ds_logic.v(14222)
  and u16877 (Cqwow6, Qqwow6, Xqwow6);  // ../RTL/cortexm0ds_logic.v(14223)
  and u16878 (n4678, vis_r11_o[26], Ljqow6);  // ../RTL/cortexm0ds_logic.v(14224)
  not u16879 (Xqwow6, n4678);  // ../RTL/cortexm0ds_logic.v(14224)
  AL_MUX u1688 (
    .i0(vis_pc_o[17]),
    .i1(Dydpw6),
    .sel(Nv0iu6),
    .o(Od1iu6));  // ../RTL/cortexm0ds_logic.v(3626)
  and u16880 (n4679, vis_r10_o[26], Sjqow6);  // ../RTL/cortexm0ds_logic.v(14225)
  not u16881 (Qqwow6, n4679);  // ../RTL/cortexm0ds_logic.v(14225)
  and u16882 (Opwow6, Ryzhu6, Erwow6);  // ../RTL/cortexm0ds_logic.v(14226)
  and u16883 (n4680, vis_r8_o[26], Gkqow6);  // ../RTL/cortexm0ds_logic.v(14227)
  not u16884 (Erwow6, n4680);  // ../RTL/cortexm0ds_logic.v(14227)
  and u16885 (Ryzhu6, Lrwow6, Srwow6);  // ../RTL/cortexm0ds_logic.v(14228)
  and u16886 (Srwow6, Zrwow6, Gswow6);  // ../RTL/cortexm0ds_logic.v(14229)
  and u16887 (Gswow6, Nswow6, Uswow6);  // ../RTL/cortexm0ds_logic.v(14230)
  and u16888 (n4681, vis_r2_o[26], Dmqow6);  // ../RTL/cortexm0ds_logic.v(14231)
  not u16889 (Uswow6, n4681);  // ../RTL/cortexm0ds_logic.v(14231)
  and u1689 (Q4lhu6, Vd1iu6, Aylhu6);  // ../RTL/cortexm0ds_logic.v(3627)
  and u16890 (n4682, vis_r6_o[26], Kmqow6);  // ../RTL/cortexm0ds_logic.v(14232)
  not u16891 (Nswow6, n4682);  // ../RTL/cortexm0ds_logic.v(14232)
  and u16892 (Zrwow6, Btwow6, Itwow6);  // ../RTL/cortexm0ds_logic.v(14233)
  and u16893 (n4683, vis_r5_o[26], Fnqow6);  // ../RTL/cortexm0ds_logic.v(14234)
  not u16894 (Itwow6, n4683);  // ../RTL/cortexm0ds_logic.v(14234)
  and u16895 (n4684, vis_r4_o[26], Mnqow6);  // ../RTL/cortexm0ds_logic.v(14235)
  not u16896 (Btwow6, n4684);  // ../RTL/cortexm0ds_logic.v(14235)
  and u16897 (Lrwow6, Ptwow6, Wtwow6);  // ../RTL/cortexm0ds_logic.v(14236)
  and u16898 (Wtwow6, Duwow6, Kuwow6);  // ../RTL/cortexm0ds_logic.v(14237)
  and u16899 (n4685, vis_r1_o[26], Voqow6);  // ../RTL/cortexm0ds_logic.v(14238)
  buf u169 (E1hpw6[11], Ux8bx6);  // ../RTL/cortexm0ds_logic.v(2367)
  AL_MUX u1690 (
    .i0(vis_pc_o[18]),
    .i1(Kydpw6),
    .sel(Nv0iu6),
    .o(Vd1iu6));  // ../RTL/cortexm0ds_logic.v(3628)
  not u16900 (Kuwow6, n4685);  // ../RTL/cortexm0ds_logic.v(14238)
  and u16901 (n4686, vis_r0_o[26], Cpqow6);  // ../RTL/cortexm0ds_logic.v(14239)
  not u16902 (Duwow6, n4686);  // ../RTL/cortexm0ds_logic.v(14239)
  and u16903 (Ptwow6, Ruwow6, Yuwow6);  // ../RTL/cortexm0ds_logic.v(14240)
  and u16904 (n4687, vis_r3_o[26], Xpqow6);  // ../RTL/cortexm0ds_logic.v(14241)
  not u16905 (Yuwow6, n4687);  // ../RTL/cortexm0ds_logic.v(14241)
  and u16906 (n4688, vis_r7_o[26], Eqqow6);  // ../RTL/cortexm0ds_logic.v(14242)
  not u16907 (Ruwow6, n4688);  // ../RTL/cortexm0ds_logic.v(14242)
  or u16908 (Imwow6, C1liu6, Qaxiu6);  // ../RTL/cortexm0ds_logic.v(14243)
  not u16909 (C1liu6, R84iu6);  // ../RTL/cortexm0ds_logic.v(14244)
  and u1691 (Y5lhu6, Ce1iu6, Twlhu6);  // ../RTL/cortexm0ds_logic.v(3629)
  and u16910 (R84iu6, Shhpw6[26], Iqzhu6);  // ../RTL/cortexm0ds_logic.v(14245)
  and u16911 (Ulwow6, Fvwow6, Mvwow6);  // ../RTL/cortexm0ds_logic.v(14246)
  or u16912 (Mvwow6, Nlwow6, Ka8ju6);  // ../RTL/cortexm0ds_logic.v(14247)
  and u16913 (Awwow6, Hwwow6, Owwow6);  // ../RTL/cortexm0ds_logic.v(14249)
  or u16914 (Owwow6, Nlwow6, I28ju6);  // ../RTL/cortexm0ds_logic.v(14250)
  and u16915 (I28ju6, Vwwow6, Cxwow6);  // ../RTL/cortexm0ds_logic.v(14251)
  and u16916 (Cxwow6, Jxwow6, Qxwow6);  // ../RTL/cortexm0ds_logic.v(14252)
  and u16917 (Qxwow6, Xxwow6, Eywow6);  // ../RTL/cortexm0ds_logic.v(14253)
  and u16918 (n4689, vis_r11_o[9], Ljqow6);  // ../RTL/cortexm0ds_logic.v(14254)
  not u16919 (Eywow6, n4689);  // ../RTL/cortexm0ds_logic.v(14254)
  AL_MUX u1692 (
    .i0(vis_pc_o[19]),
    .i1(Rydpw6),
    .sel(Nv0iu6),
    .o(Ce1iu6));  // ../RTL/cortexm0ds_logic.v(3630)
  and u16920 (Xxwow6, Lywow6, Sywow6);  // ../RTL/cortexm0ds_logic.v(14255)
  and u16921 (n4690, vis_r10_o[9], Sjqow6);  // ../RTL/cortexm0ds_logic.v(14256)
  not u16922 (Sywow6, n4690);  // ../RTL/cortexm0ds_logic.v(14256)
  and u16923 (n4691, vis_r9_o[9], Qiqow6);  // ../RTL/cortexm0ds_logic.v(14257)
  not u16924 (Lywow6, n4691);  // ../RTL/cortexm0ds_logic.v(14257)
  and u16925 (Jxwow6, Zywow6, Gzwow6);  // ../RTL/cortexm0ds_logic.v(14258)
  and u16926 (n4692, Fkfpw6[9], Dfqow6);  // ../RTL/cortexm0ds_logic.v(14259)
  not u16927 (Gzwow6, n4692);  // ../RTL/cortexm0ds_logic.v(14259)
  and u16928 (n4693, vis_r12_o[9], Hhqow6);  // ../RTL/cortexm0ds_logic.v(14260)
  not u16929 (Zywow6, n4693);  // ../RTL/cortexm0ds_logic.v(14260)
  and u1693 (G7lhu6, Je1iu6, Mvlhu6);  // ../RTL/cortexm0ds_logic.v(3631)
  and u16930 (Vwwow6, Nzwow6, Uzwow6);  // ../RTL/cortexm0ds_logic.v(14261)
  and u16931 (Uzwow6, B0xow6, I0xow6);  // ../RTL/cortexm0ds_logic.v(14262)
  and u16932 (n4694, vis_r14_o[9], Ahqow6);  // ../RTL/cortexm0ds_logic.v(14263)
  not u16933 (I0xow6, n4694);  // ../RTL/cortexm0ds_logic.v(14263)
  and u16934 (B0xow6, P0xow6, W0xow6);  // ../RTL/cortexm0ds_logic.v(14264)
  and u16935 (n4695, vis_psp_o[7], Yfqow6);  // ../RTL/cortexm0ds_logic.v(14265)
  not u16936 (W0xow6, n4695);  // ../RTL/cortexm0ds_logic.v(14265)
  and u16937 (n4696, vis_r8_o[9], Gkqow6);  // ../RTL/cortexm0ds_logic.v(14266)
  not u16938 (P0xow6, n4696);  // ../RTL/cortexm0ds_logic.v(14266)
  and u16939 (Nzwow6, Evzhu6, D1xow6);  // ../RTL/cortexm0ds_logic.v(14267)
  AL_MUX u1694 (
    .i0(vis_pc_o[20]),
    .i1(Yydpw6),
    .sel(Nv0iu6),
    .o(Je1iu6));  // ../RTL/cortexm0ds_logic.v(3632)
  and u16940 (n4697, vis_msp_o[7], Fgqow6);  // ../RTL/cortexm0ds_logic.v(14268)
  not u16941 (D1xow6, n4697);  // ../RTL/cortexm0ds_logic.v(14268)
  and u16942 (Evzhu6, K1xow6, R1xow6);  // ../RTL/cortexm0ds_logic.v(14269)
  and u16943 (R1xow6, Y1xow6, F2xow6);  // ../RTL/cortexm0ds_logic.v(14270)
  and u16944 (F2xow6, M2xow6, T2xow6);  // ../RTL/cortexm0ds_logic.v(14271)
  and u16945 (n4698, vis_r0_o[9], Cpqow6);  // ../RTL/cortexm0ds_logic.v(14272)
  not u16946 (T2xow6, n4698);  // ../RTL/cortexm0ds_logic.v(14272)
  and u16947 (n4699, vis_r2_o[9], Dmqow6);  // ../RTL/cortexm0ds_logic.v(14273)
  not u16948 (M2xow6, n4699);  // ../RTL/cortexm0ds_logic.v(14273)
  and u16949 (Y1xow6, A3xow6, H3xow6);  // ../RTL/cortexm0ds_logic.v(14274)
  and u1695 (O8lhu6, Qe1iu6, Fulhu6);  // ../RTL/cortexm0ds_logic.v(3633)
  and u16950 (n4700, vis_r5_o[9], Fnqow6);  // ../RTL/cortexm0ds_logic.v(14275)
  not u16951 (H3xow6, n4700);  // ../RTL/cortexm0ds_logic.v(14275)
  and u16952 (n4701, vis_r4_o[9], Mnqow6);  // ../RTL/cortexm0ds_logic.v(14276)
  not u16953 (A3xow6, n4701);  // ../RTL/cortexm0ds_logic.v(14276)
  and u16954 (K1xow6, O3xow6, V3xow6);  // ../RTL/cortexm0ds_logic.v(14277)
  and u16955 (V3xow6, C4xow6, J4xow6);  // ../RTL/cortexm0ds_logic.v(14278)
  and u16956 (n4702, vis_r7_o[9], Eqqow6);  // ../RTL/cortexm0ds_logic.v(14279)
  not u16957 (J4xow6, n4702);  // ../RTL/cortexm0ds_logic.v(14279)
  and u16958 (n4703, vis_r3_o[9], Xpqow6);  // ../RTL/cortexm0ds_logic.v(14280)
  not u16959 (C4xow6, n4703);  // ../RTL/cortexm0ds_logic.v(14280)
  AL_MUX u1696 (
    .i0(vis_pc_o[21]),
    .i1(Fzdpw6),
    .sel(Nv0iu6),
    .o(Qe1iu6));  // ../RTL/cortexm0ds_logic.v(3634)
  and u16960 (O3xow6, Q4xow6, X4xow6);  // ../RTL/cortexm0ds_logic.v(14281)
  and u16961 (n4704, vis_r1_o[9], Voqow6);  // ../RTL/cortexm0ds_logic.v(14282)
  not u16962 (X4xow6, n4704);  // ../RTL/cortexm0ds_logic.v(14282)
  and u16963 (n4705, vis_r6_o[9], Kmqow6);  // ../RTL/cortexm0ds_logic.v(14283)
  not u16964 (Q4xow6, n4705);  // ../RTL/cortexm0ds_logic.v(14283)
  and u16965 (n4706, Gdqow6, Goliu6);  // ../RTL/cortexm0ds_logic.v(14284)
  not u16966 (Hwwow6, n4706);  // ../RTL/cortexm0ds_logic.v(14284)
  and u16967 (n4707, E5xow6, L5xow6);  // ../RTL/cortexm0ds_logic.v(14285)
  not u16968 (Goliu6, n4707);  // ../RTL/cortexm0ds_logic.v(14285)
  and u16969 (L5xow6, S5xow6, Z5xow6);  // ../RTL/cortexm0ds_logic.v(14286)
  and u1697 (W9lhu6, Xe1iu6, Yslhu6);  // ../RTL/cortexm0ds_logic.v(3635)
  and u16970 (Z5xow6, G6xow6, N6xow6);  // ../RTL/cortexm0ds_logic.v(14287)
  and u16971 (n4708, Fkfpw6[25], Dfqow6);  // ../RTL/cortexm0ds_logic.v(14288)
  not u16972 (N6xow6, n4708);  // ../RTL/cortexm0ds_logic.v(14288)
  and u16973 (G6xow6, U6xow6, B7xow6);  // ../RTL/cortexm0ds_logic.v(14289)
  and u16974 (n4709, vis_psp_o[23], Yfqow6);  // ../RTL/cortexm0ds_logic.v(14290)
  not u16975 (B7xow6, n4709);  // ../RTL/cortexm0ds_logic.v(14290)
  and u16976 (n4710, vis_msp_o[23], Fgqow6);  // ../RTL/cortexm0ds_logic.v(14291)
  not u16977 (U6xow6, n4710);  // ../RTL/cortexm0ds_logic.v(14291)
  and u16978 (S5xow6, I7xow6, P7xow6);  // ../RTL/cortexm0ds_logic.v(14292)
  and u16979 (n4711, vis_r14_o[25], Ahqow6);  // ../RTL/cortexm0ds_logic.v(14293)
  AL_MUX u1698 (
    .i0(vis_pc_o[22]),
    .i1(Mzdpw6),
    .sel(Nv0iu6),
    .o(Xe1iu6));  // ../RTL/cortexm0ds_logic.v(3636)
  not u16980 (P7xow6, n4711);  // ../RTL/cortexm0ds_logic.v(14293)
  and u16981 (n4712, vis_r12_o[25], Hhqow6);  // ../RTL/cortexm0ds_logic.v(14294)
  not u16982 (I7xow6, n4712);  // ../RTL/cortexm0ds_logic.v(14294)
  and u16983 (E5xow6, W7xow6, D8xow6);  // ../RTL/cortexm0ds_logic.v(14295)
  and u16984 (D8xow6, K8xow6, R8xow6);  // ../RTL/cortexm0ds_logic.v(14296)
  and u16985 (n4713, vis_r9_o[25], Qiqow6);  // ../RTL/cortexm0ds_logic.v(14297)
  not u16986 (R8xow6, n4713);  // ../RTL/cortexm0ds_logic.v(14297)
  and u16987 (K8xow6, Y8xow6, F9xow6);  // ../RTL/cortexm0ds_logic.v(14298)
  and u16988 (n4714, vis_r11_o[25], Ljqow6);  // ../RTL/cortexm0ds_logic.v(14299)
  not u16989 (F9xow6, n4714);  // ../RTL/cortexm0ds_logic.v(14299)
  AL_MUX u1699 (
    .i0(vis_pc_o[30]),
    .i1(Ef1iu6),
    .sel(Ty0iu6),
    .o(R9ohu6));  // ../RTL/cortexm0ds_logic.v(3637)
  and u16990 (n4715, vis_r10_o[25], Sjqow6);  // ../RTL/cortexm0ds_logic.v(14300)
  not u16991 (Y8xow6, n4715);  // ../RTL/cortexm0ds_logic.v(14300)
  and u16992 (W7xow6, Yyzhu6, M9xow6);  // ../RTL/cortexm0ds_logic.v(14301)
  and u16993 (n4716, vis_r8_o[25], Gkqow6);  // ../RTL/cortexm0ds_logic.v(14302)
  not u16994 (M9xow6, n4716);  // ../RTL/cortexm0ds_logic.v(14302)
  and u16995 (Yyzhu6, T9xow6, Aaxow6);  // ../RTL/cortexm0ds_logic.v(14303)
  and u16996 (Aaxow6, Haxow6, Oaxow6);  // ../RTL/cortexm0ds_logic.v(14304)
  and u16997 (Oaxow6, Vaxow6, Cbxow6);  // ../RTL/cortexm0ds_logic.v(14305)
  and u16998 (n4717, vis_r2_o[25], Dmqow6);  // ../RTL/cortexm0ds_logic.v(14306)
  not u16999 (Cbxow6, n4717);  // ../RTL/cortexm0ds_logic.v(14306)
  buf u17 (Gwnhu6, T0ipw6);  // ../RTL/cortexm0ds_logic.v(1773)
  buf u170 (E1hpw6[10], Yjaax6);  // ../RTL/cortexm0ds_logic.v(2367)
  AL_MUX u1700 (
    .i0(vis_pc_o[30]),
    .i1(Ef1iu6),
    .sel(Nv0iu6),
    .o(M9ohu6));  // ../RTL/cortexm0ds_logic.v(3638)
  and u17000 (n4718, vis_r6_o[25], Kmqow6);  // ../RTL/cortexm0ds_logic.v(14307)
  not u17001 (Vaxow6, n4718);  // ../RTL/cortexm0ds_logic.v(14307)
  and u17002 (Haxow6, Jbxow6, Qbxow6);  // ../RTL/cortexm0ds_logic.v(14308)
  and u17003 (n4719, vis_r5_o[25], Fnqow6);  // ../RTL/cortexm0ds_logic.v(14309)
  not u17004 (Qbxow6, n4719);  // ../RTL/cortexm0ds_logic.v(14309)
  and u17005 (n4720, vis_r4_o[25], Mnqow6);  // ../RTL/cortexm0ds_logic.v(14310)
  not u17006 (Jbxow6, n4720);  // ../RTL/cortexm0ds_logic.v(14310)
  and u17007 (T9xow6, Xbxow6, Ecxow6);  // ../RTL/cortexm0ds_logic.v(14311)
  and u17008 (Ecxow6, Lcxow6, Scxow6);  // ../RTL/cortexm0ds_logic.v(14312)
  and u17009 (n4721, vis_r1_o[25], Voqow6);  // ../RTL/cortexm0ds_logic.v(14313)
  AL_MUX u1701 (
    .i0(Lf1iu6),
    .i1(X0ohu6),
    .sel(Sf1iu6),
    .o(X3yhu6));  // ../RTL/cortexm0ds_logic.v(3639)
  not u17010 (Scxow6, n4721);  // ../RTL/cortexm0ds_logic.v(14313)
  and u17011 (n4722, vis_r0_o[25], Cpqow6);  // ../RTL/cortexm0ds_logic.v(14314)
  not u17012 (Lcxow6, n4722);  // ../RTL/cortexm0ds_logic.v(14314)
  and u17013 (Xbxow6, Zcxow6, Gdxow6);  // ../RTL/cortexm0ds_logic.v(14315)
  and u17014 (n4723, vis_r3_o[25], Xpqow6);  // ../RTL/cortexm0ds_logic.v(14316)
  not u17015 (Gdxow6, n4723);  // ../RTL/cortexm0ds_logic.v(14316)
  and u17016 (n4724, vis_r7_o[25], Eqqow6);  // ../RTL/cortexm0ds_logic.v(14317)
  not u17017 (Zcxow6, n4724);  // ../RTL/cortexm0ds_logic.v(14317)
  and u17018 (Tvwow6, Acvow6, Ndxow6);  // ../RTL/cortexm0ds_logic.v(14318)
  or u17019 (Ndxow6, Asliu6, Qaxiu6);  // ../RTL/cortexm0ds_logic.v(14319)
  and u1702 (n125, Zf1iu6, Gg1iu6);  // ../RTL/cortexm0ds_logic.v(3640)
  not u17020 (Asliu6, K84iu6);  // ../RTL/cortexm0ds_logic.v(14320)
  and u17021 (K84iu6, Shhpw6[25], Iqzhu6);  // ../RTL/cortexm0ds_logic.v(14321)
  and u17022 (n4725, Udxow6, Znliu6);  // ../RTL/cortexm0ds_logic.v(14322)
  not u17023 (Acvow6, n4725);  // ../RTL/cortexm0ds_logic.v(14322)
  and u17024 (Iexow6, Pexow6, Wexow6);  // ../RTL/cortexm0ds_logic.v(14324)
  or u17025 (Wexow6, Nlwow6, Cz7ju6);  // ../RTL/cortexm0ds_logic.v(14325)
  and u17026 (Cz7ju6, Dfxow6, Kfxow6);  // ../RTL/cortexm0ds_logic.v(14326)
  and u17027 (Kfxow6, Rfxow6, Yfxow6);  // ../RTL/cortexm0ds_logic.v(14327)
  and u17028 (Yfxow6, Fgxow6, Mgxow6);  // ../RTL/cortexm0ds_logic.v(14328)
  and u17029 (n4726, vis_r11_o[8], Ljqow6);  // ../RTL/cortexm0ds_logic.v(14329)
  not u1703 (Q3yhu6, n125);  // ../RTL/cortexm0ds_logic.v(3640)
  not u17030 (Mgxow6, n4726);  // ../RTL/cortexm0ds_logic.v(14329)
  and u17031 (Fgxow6, Tgxow6, Ahxow6);  // ../RTL/cortexm0ds_logic.v(14330)
  and u17032 (n4727, vis_r9_o[8], Qiqow6);  // ../RTL/cortexm0ds_logic.v(14331)
  not u17033 (Ahxow6, n4727);  // ../RTL/cortexm0ds_logic.v(14331)
  and u17034 (n4728, Fkfpw6[8], Dfqow6);  // ../RTL/cortexm0ds_logic.v(14332)
  not u17035 (Tgxow6, n4728);  // ../RTL/cortexm0ds_logic.v(14332)
  and u17036 (Rfxow6, Hhxow6, Ohxow6);  // ../RTL/cortexm0ds_logic.v(14333)
  and u17037 (n4729, vis_r10_o[8], Sjqow6);  // ../RTL/cortexm0ds_logic.v(14334)
  not u17038 (Ohxow6, n4729);  // ../RTL/cortexm0ds_logic.v(14334)
  and u17039 (n4730, vis_psp_o[6], Yfqow6);  // ../RTL/cortexm0ds_logic.v(14335)
  or u1704 (Gg1iu6, Ng1iu6, Ug1iu6);  // ../RTL/cortexm0ds_logic.v(3641)
  not u17040 (Hhxow6, n4730);  // ../RTL/cortexm0ds_logic.v(14335)
  and u17041 (Dfxow6, Vhxow6, Cixow6);  // ../RTL/cortexm0ds_logic.v(14336)
  and u17042 (Cixow6, Jixow6, Qixow6);  // ../RTL/cortexm0ds_logic.v(14337)
  and u17043 (n4731, vis_r12_o[8], Hhqow6);  // ../RTL/cortexm0ds_logic.v(14338)
  not u17044 (Qixow6, n4731);  // ../RTL/cortexm0ds_logic.v(14338)
  and u17045 (Jixow6, Xixow6, Ejxow6);  // ../RTL/cortexm0ds_logic.v(14339)
  and u17046 (n4732, vis_msp_o[6], Fgqow6);  // ../RTL/cortexm0ds_logic.v(14340)
  not u17047 (Ejxow6, n4732);  // ../RTL/cortexm0ds_logic.v(14340)
  and u17048 (n4733, vis_r14_o[8], Ahqow6);  // ../RTL/cortexm0ds_logic.v(14341)
  not u17049 (Xixow6, n4733);  // ../RTL/cortexm0ds_logic.v(14341)
  or u1705 (n126, Ih1iu6, Ph1iu6);  // ../RTL/cortexm0ds_logic.v(3643)
  and u17050 (Vhxow6, Lvzhu6, Ljxow6);  // ../RTL/cortexm0ds_logic.v(14342)
  and u17051 (n4734, vis_r8_o[8], Gkqow6);  // ../RTL/cortexm0ds_logic.v(14343)
  not u17052 (Ljxow6, n4734);  // ../RTL/cortexm0ds_logic.v(14343)
  and u17053 (Lvzhu6, Sjxow6, Zjxow6);  // ../RTL/cortexm0ds_logic.v(14344)
  and u17054 (Zjxow6, Gkxow6, Nkxow6);  // ../RTL/cortexm0ds_logic.v(14345)
  and u17055 (Nkxow6, Ukxow6, Blxow6);  // ../RTL/cortexm0ds_logic.v(14346)
  and u17056 (n4735, vis_r2_o[8], Dmqow6);  // ../RTL/cortexm0ds_logic.v(14347)
  not u17057 (Blxow6, n4735);  // ../RTL/cortexm0ds_logic.v(14347)
  and u17058 (n4736, vis_r6_o[8], Kmqow6);  // ../RTL/cortexm0ds_logic.v(14348)
  not u17059 (Ukxow6, n4736);  // ../RTL/cortexm0ds_logic.v(14348)
  not u1706 (Zf1iu6, n126);  // ../RTL/cortexm0ds_logic.v(3643)
  and u17060 (Gkxow6, Ilxow6, Plxow6);  // ../RTL/cortexm0ds_logic.v(14349)
  and u17061 (n4737, vis_r5_o[8], Fnqow6);  // ../RTL/cortexm0ds_logic.v(14350)
  not u17062 (Plxow6, n4737);  // ../RTL/cortexm0ds_logic.v(14350)
  and u17063 (n4738, vis_r4_o[8], Mnqow6);  // ../RTL/cortexm0ds_logic.v(14351)
  not u17064 (Ilxow6, n4738);  // ../RTL/cortexm0ds_logic.v(14351)
  and u17065 (Sjxow6, Wlxow6, Dmxow6);  // ../RTL/cortexm0ds_logic.v(14352)
  and u17066 (Dmxow6, Kmxow6, Rmxow6);  // ../RTL/cortexm0ds_logic.v(14353)
  and u17067 (n4739, vis_r1_o[8], Voqow6);  // ../RTL/cortexm0ds_logic.v(14354)
  not u17068 (Rmxow6, n4739);  // ../RTL/cortexm0ds_logic.v(14354)
  and u17069 (n4740, vis_r0_o[8], Cpqow6);  // ../RTL/cortexm0ds_logic.v(14355)
  and u1707 (Ih1iu6, Fanhu6, Wh1iu6);  // ../RTL/cortexm0ds_logic.v(3644)
  not u17070 (Kmxow6, n4740);  // ../RTL/cortexm0ds_logic.v(14355)
  and u17071 (Wlxow6, Ymxow6, Fnxow6);  // ../RTL/cortexm0ds_logic.v(14356)
  and u17072 (n4741, vis_r3_o[8], Xpqow6);  // ../RTL/cortexm0ds_logic.v(14357)
  not u17073 (Fnxow6, n4741);  // ../RTL/cortexm0ds_logic.v(14357)
  and u17074 (n4742, vis_r7_o[8], Eqqow6);  // ../RTL/cortexm0ds_logic.v(14358)
  not u17075 (Ymxow6, n4742);  // ../RTL/cortexm0ds_logic.v(14358)
  and u17076 (K0row6, Mnxow6, Sevow6);  // ../RTL/cortexm0ds_logic.v(14359)
  not u17077 (Nlwow6, K0row6);  // ../RTL/cortexm0ds_logic.v(14359)
  and u17078 (n4743, Gdqow6, Fy6ju6);  // ../RTL/cortexm0ds_logic.v(14360)
  not u17079 (Pexow6, n4743);  // ../RTL/cortexm0ds_logic.v(14360)
  and u1708 (n127, Iahpw6[1], Di1iu6);  // ../RTL/cortexm0ds_logic.v(3645)
  and u17080 (n4744, Tnxow6, Aoxow6);  // ../RTL/cortexm0ds_logic.v(14361)
  not u17081 (Fy6ju6, n4744);  // ../RTL/cortexm0ds_logic.v(14361)
  and u17082 (Aoxow6, Hoxow6, Ooxow6);  // ../RTL/cortexm0ds_logic.v(14362)
  and u17083 (Ooxow6, Voxow6, Cpxow6);  // ../RTL/cortexm0ds_logic.v(14363)
  and u17084 (n4745, Fkfpw6[24], Dfqow6);  // ../RTL/cortexm0ds_logic.v(14364)
  not u17085 (Cpxow6, n4745);  // ../RTL/cortexm0ds_logic.v(14364)
  and u17086 (Voxow6, Jpxow6, Qpxow6);  // ../RTL/cortexm0ds_logic.v(14365)
  and u17087 (n4746, vis_psp_o[22], Yfqow6);  // ../RTL/cortexm0ds_logic.v(14366)
  not u17088 (Qpxow6, n4746);  // ../RTL/cortexm0ds_logic.v(14366)
  and u17089 (n4747, vis_msp_o[22], Fgqow6);  // ../RTL/cortexm0ds_logic.v(14367)
  not u1709 (Wh1iu6, n127);  // ../RTL/cortexm0ds_logic.v(3645)
  not u17090 (Jpxow6, n4747);  // ../RTL/cortexm0ds_logic.v(14367)
  and u17091 (Hoxow6, Xpxow6, Eqxow6);  // ../RTL/cortexm0ds_logic.v(14368)
  and u17092 (n4748, vis_r14_o[24], Ahqow6);  // ../RTL/cortexm0ds_logic.v(14369)
  not u17093 (Eqxow6, n4748);  // ../RTL/cortexm0ds_logic.v(14369)
  and u17094 (n4749, vis_r12_o[24], Hhqow6);  // ../RTL/cortexm0ds_logic.v(14370)
  not u17095 (Xpxow6, n4749);  // ../RTL/cortexm0ds_logic.v(14370)
  and u17096 (Tnxow6, Lqxow6, Sqxow6);  // ../RTL/cortexm0ds_logic.v(14371)
  and u17097 (Sqxow6, Zqxow6, Grxow6);  // ../RTL/cortexm0ds_logic.v(14372)
  and u17098 (n4750, vis_r9_o[24], Qiqow6);  // ../RTL/cortexm0ds_logic.v(14373)
  not u17099 (Grxow6, n4750);  // ../RTL/cortexm0ds_logic.v(14373)
  buf u171 (Y7ghu6, P5vpw6);  // ../RTL/cortexm0ds_logic.v(2016)
  and u1710 (n128, Ki1iu6, Ri1iu6);  // ../RTL/cortexm0ds_logic.v(3646)
  and u17100 (Zqxow6, Nrxow6, Urxow6);  // ../RTL/cortexm0ds_logic.v(14374)
  and u17101 (n4751, vis_r11_o[24], Ljqow6);  // ../RTL/cortexm0ds_logic.v(14375)
  not u17102 (Urxow6, n4751);  // ../RTL/cortexm0ds_logic.v(14375)
  and u17103 (n4752, vis_r10_o[24], Sjqow6);  // ../RTL/cortexm0ds_logic.v(14376)
  not u17104 (Nrxow6, n4752);  // ../RTL/cortexm0ds_logic.v(14376)
  and u17105 (Lqxow6, Fzzhu6, Bsxow6);  // ../RTL/cortexm0ds_logic.v(14377)
  and u17106 (n4753, vis_r8_o[24], Gkqow6);  // ../RTL/cortexm0ds_logic.v(14378)
  not u17107 (Bsxow6, n4753);  // ../RTL/cortexm0ds_logic.v(14378)
  and u17108 (Fzzhu6, Isxow6, Psxow6);  // ../RTL/cortexm0ds_logic.v(14379)
  and u17109 (Psxow6, Wsxow6, Dtxow6);  // ../RTL/cortexm0ds_logic.v(14380)
  not u1711 (J3yhu6, n128);  // ../RTL/cortexm0ds_logic.v(3646)
  and u17110 (Dtxow6, Ktxow6, Rtxow6);  // ../RTL/cortexm0ds_logic.v(14381)
  and u17111 (n4754, vis_r2_o[24], Dmqow6);  // ../RTL/cortexm0ds_logic.v(14382)
  not u17112 (Rtxow6, n4754);  // ../RTL/cortexm0ds_logic.v(14382)
  and u17113 (n4755, vis_r6_o[24], Kmqow6);  // ../RTL/cortexm0ds_logic.v(14383)
  not u17114 (Ktxow6, n4755);  // ../RTL/cortexm0ds_logic.v(14383)
  and u17115 (Wsxow6, Ytxow6, Fuxow6);  // ../RTL/cortexm0ds_logic.v(14384)
  and u17116 (n4756, vis_r5_o[24], Fnqow6);  // ../RTL/cortexm0ds_logic.v(14385)
  not u17117 (Fuxow6, n4756);  // ../RTL/cortexm0ds_logic.v(14385)
  and u17118 (n4757, vis_r4_o[24], Mnqow6);  // ../RTL/cortexm0ds_logic.v(14386)
  not u17119 (Ytxow6, n4757);  // ../RTL/cortexm0ds_logic.v(14386)
  and u1712 (n129, Yi1iu6, Fj1iu6);  // ../RTL/cortexm0ds_logic.v(3647)
  and u17120 (Isxow6, Muxow6, Tuxow6);  // ../RTL/cortexm0ds_logic.v(14387)
  and u17121 (Tuxow6, Avxow6, Hvxow6);  // ../RTL/cortexm0ds_logic.v(14388)
  and u17122 (n4758, vis_r1_o[24], Voqow6);  // ../RTL/cortexm0ds_logic.v(14389)
  not u17123 (Hvxow6, n4758);  // ../RTL/cortexm0ds_logic.v(14389)
  and u17124 (n4759, vis_r0_o[24], Cpqow6);  // ../RTL/cortexm0ds_logic.v(14390)
  not u17125 (Avxow6, n4759);  // ../RTL/cortexm0ds_logic.v(14390)
  and u17126 (Muxow6, Ovxow6, Vvxow6);  // ../RTL/cortexm0ds_logic.v(14391)
  and u17127 (n4760, vis_r3_o[24], Xpqow6);  // ../RTL/cortexm0ds_logic.v(14392)
  not u17128 (Vvxow6, n4760);  // ../RTL/cortexm0ds_logic.v(14392)
  and u17129 (n4761, vis_r7_o[24], Eqqow6);  // ../RTL/cortexm0ds_logic.v(14393)
  not u1713 (Ri1iu6, n129);  // ../RTL/cortexm0ds_logic.v(3647)
  not u17130 (Ovxow6, n4761);  // ../RTL/cortexm0ds_logic.v(14393)
  and u17131 (Bexow6, Jdvow6, Cwxow6);  // ../RTL/cortexm0ds_logic.v(14394)
  or u17132 (Cwxow6, Rykiu6, Qaxiu6);  // ../RTL/cortexm0ds_logic.v(14395)
  not u17133 (Rykiu6, D84iu6);  // ../RTL/cortexm0ds_logic.v(14396)
  and u17134 (D84iu6, Shhpw6[24], Iqzhu6);  // ../RTL/cortexm0ds_logic.v(14397)
  and u17135 (n4762, Udxow6, L35ju6);  // ../RTL/cortexm0ds_logic.v(14398)
  not u17136 (Jdvow6, n4762);  // ../RTL/cortexm0ds_logic.v(14398)
  and u17137 (n4763, Lcqow6, Uo6ju6);  // ../RTL/cortexm0ds_logic.v(14400)
  not u17138 (Qwxow6, n4763);  // ../RTL/cortexm0ds_logic.v(14400)
  and u17139 (Jwxow6, Xwxow6, Exxow6);  // ../RTL/cortexm0ds_logic.v(14401)
  or u1714 (Sr3iu6, Ofzhu6, Mdhpw6[0]);  // ../RTL/cortexm0ds_logic.v(3648)
  or u17140 (Exxow6, Ox9iu6, Qaxiu6);  // ../RTL/cortexm0ds_logic.v(14402)
  not u17141 (Ox9iu6, W74iu6);  // ../RTL/cortexm0ds_logic.v(14403)
  and u17142 (W74iu6, Shhpw6[23], Iqzhu6);  // ../RTL/cortexm0ds_logic.v(14404)
  and u17143 (n4764, Gdqow6, Xg5ju6);  // ../RTL/cortexm0ds_logic.v(14405)
  not u17144 (Xwxow6, n4764);  // ../RTL/cortexm0ds_logic.v(14405)
  and u17145 (n4765, Lxxow6, Sxxow6);  // ../RTL/cortexm0ds_logic.v(14406)
  not u17146 (Xg5ju6, n4765);  // ../RTL/cortexm0ds_logic.v(14406)
  and u17147 (Sxxow6, Zxxow6, Gyxow6);  // ../RTL/cortexm0ds_logic.v(14407)
  and u17148 (Gyxow6, Nyxow6, Uyxow6);  // ../RTL/cortexm0ds_logic.v(14408)
  and u17149 (n4766, Fkfpw6[23], Dfqow6);  // ../RTL/cortexm0ds_logic.v(14409)
  not u1715 (Yi1iu6, Sr3iu6);  // ../RTL/cortexm0ds_logic.v(3648)
  not u17150 (Uyxow6, n4766);  // ../RTL/cortexm0ds_logic.v(14409)
  and u17151 (Nyxow6, Bzxow6, Izxow6);  // ../RTL/cortexm0ds_logic.v(14410)
  and u17152 (n4767, vis_psp_o[21], Yfqow6);  // ../RTL/cortexm0ds_logic.v(14411)
  not u17153 (Izxow6, n4767);  // ../RTL/cortexm0ds_logic.v(14411)
  and u17154 (n4768, vis_msp_o[21], Fgqow6);  // ../RTL/cortexm0ds_logic.v(14412)
  not u17155 (Bzxow6, n4768);  // ../RTL/cortexm0ds_logic.v(14412)
  and u17156 (Zxxow6, Pzxow6, Wzxow6);  // ../RTL/cortexm0ds_logic.v(14413)
  and u17157 (n4769, vis_r14_o[23], Ahqow6);  // ../RTL/cortexm0ds_logic.v(14414)
  not u17158 (Wzxow6, n4769);  // ../RTL/cortexm0ds_logic.v(14414)
  and u17159 (n4770, vis_r12_o[23], Hhqow6);  // ../RTL/cortexm0ds_logic.v(14415)
  and u1716 (n130, Jdnhu6, Mj1iu6);  // ../RTL/cortexm0ds_logic.v(3649)
  not u17160 (Pzxow6, n4770);  // ../RTL/cortexm0ds_logic.v(14415)
  and u17161 (Lxxow6, D0yow6, K0yow6);  // ../RTL/cortexm0ds_logic.v(14416)
  and u17162 (K0yow6, R0yow6, Y0yow6);  // ../RTL/cortexm0ds_logic.v(14417)
  and u17163 (n4771, vis_r9_o[23], Qiqow6);  // ../RTL/cortexm0ds_logic.v(14418)
  not u17164 (Y0yow6, n4771);  // ../RTL/cortexm0ds_logic.v(14418)
  and u17165 (R0yow6, F1yow6, M1yow6);  // ../RTL/cortexm0ds_logic.v(14419)
  and u17166 (n4772, vis_r11_o[23], Ljqow6);  // ../RTL/cortexm0ds_logic.v(14420)
  not u17167 (M1yow6, n4772);  // ../RTL/cortexm0ds_logic.v(14420)
  and u17168 (n4773, vis_r10_o[23], Sjqow6);  // ../RTL/cortexm0ds_logic.v(14421)
  not u17169 (F1yow6, n4773);  // ../RTL/cortexm0ds_logic.v(14421)
  not u1717 (Ki1iu6, n130);  // ../RTL/cortexm0ds_logic.v(3649)
  and u17170 (D0yow6, Mzzhu6, T1yow6);  // ../RTL/cortexm0ds_logic.v(14422)
  and u17171 (n4774, vis_r8_o[23], Gkqow6);  // ../RTL/cortexm0ds_logic.v(14423)
  not u17172 (T1yow6, n4774);  // ../RTL/cortexm0ds_logic.v(14423)
  and u17173 (Mzzhu6, A2yow6, H2yow6);  // ../RTL/cortexm0ds_logic.v(14424)
  and u17174 (H2yow6, O2yow6, V2yow6);  // ../RTL/cortexm0ds_logic.v(14425)
  and u17175 (V2yow6, C3yow6, J3yow6);  // ../RTL/cortexm0ds_logic.v(14426)
  and u17176 (n4775, vis_r2_o[23], Dmqow6);  // ../RTL/cortexm0ds_logic.v(14427)
  not u17177 (J3yow6, n4775);  // ../RTL/cortexm0ds_logic.v(14427)
  and u17178 (n4776, vis_r6_o[23], Kmqow6);  // ../RTL/cortexm0ds_logic.v(14428)
  not u17179 (C3yow6, n4776);  // ../RTL/cortexm0ds_logic.v(14428)
  and u1718 (n131, Iahpw6[2], Di1iu6);  // ../RTL/cortexm0ds_logic.v(3650)
  and u17180 (O2yow6, Q3yow6, X3yow6);  // ../RTL/cortexm0ds_logic.v(14429)
  and u17181 (n4777, vis_r5_o[23], Fnqow6);  // ../RTL/cortexm0ds_logic.v(14430)
  not u17182 (X3yow6, n4777);  // ../RTL/cortexm0ds_logic.v(14430)
  and u17183 (n4778, vis_r4_o[23], Mnqow6);  // ../RTL/cortexm0ds_logic.v(14431)
  not u17184 (Q3yow6, n4778);  // ../RTL/cortexm0ds_logic.v(14431)
  and u17185 (A2yow6, E4yow6, L4yow6);  // ../RTL/cortexm0ds_logic.v(14432)
  and u17186 (L4yow6, S4yow6, Z4yow6);  // ../RTL/cortexm0ds_logic.v(14433)
  and u17187 (n4779, vis_r1_o[23], Voqow6);  // ../RTL/cortexm0ds_logic.v(14434)
  not u17188 (Z4yow6, n4779);  // ../RTL/cortexm0ds_logic.v(14434)
  and u17189 (n4780, vis_r0_o[23], Cpqow6);  // ../RTL/cortexm0ds_logic.v(14435)
  not u1719 (Mj1iu6, n131);  // ../RTL/cortexm0ds_logic.v(3650)
  not u17190 (S4yow6, n4780);  // ../RTL/cortexm0ds_logic.v(14435)
  and u17191 (E4yow6, G5yow6, N5yow6);  // ../RTL/cortexm0ds_logic.v(14436)
  and u17192 (n4781, vis_r3_o[23], Xpqow6);  // ../RTL/cortexm0ds_logic.v(14437)
  not u17193 (N5yow6, n4781);  // ../RTL/cortexm0ds_logic.v(14437)
  and u17194 (n4782, vis_r7_o[23], Eqqow6);  // ../RTL/cortexm0ds_logic.v(14438)
  not u17195 (G5yow6, n4782);  // ../RTL/cortexm0ds_logic.v(14438)
  and u17196 (n4783, Lcqow6, Kj6ju6);  // ../RTL/cortexm0ds_logic.v(14440)
  not u17197 (B6yow6, n4783);  // ../RTL/cortexm0ds_logic.v(14440)
  and u17198 (U5yow6, I6yow6, P6yow6);  // ../RTL/cortexm0ds_logic.v(14441)
  and u17199 (n4784, P74iu6, R0nhu6);  // ../RTL/cortexm0ds_logic.v(14442)
  buf u172 (DBGRESTARTED, K7vpw6);  // ../RTL/cortexm0ds_logic.v(2017)
  and u1720 (n132, Tj1iu6, Ak1iu6);  // ../RTL/cortexm0ds_logic.v(3651)
  not u17200 (P6yow6, n4784);  // ../RTL/cortexm0ds_logic.v(14442)
  and u17201 (P74iu6, Shhpw6[22], Iqzhu6);  // ../RTL/cortexm0ds_logic.v(14443)
  and u17202 (n4785, Gdqow6, V3aju6);  // ../RTL/cortexm0ds_logic.v(14444)
  not u17203 (I6yow6, n4785);  // ../RTL/cortexm0ds_logic.v(14444)
  and u17204 (n4786, W6yow6, D7yow6);  // ../RTL/cortexm0ds_logic.v(14445)
  not u17205 (V3aju6, n4786);  // ../RTL/cortexm0ds_logic.v(14445)
  and u17206 (D7yow6, K7yow6, R7yow6);  // ../RTL/cortexm0ds_logic.v(14446)
  and u17207 (R7yow6, Y7yow6, F8yow6);  // ../RTL/cortexm0ds_logic.v(14447)
  and u17208 (n4787, Fkfpw6[22], Dfqow6);  // ../RTL/cortexm0ds_logic.v(14448)
  not u17209 (F8yow6, n4787);  // ../RTL/cortexm0ds_logic.v(14448)
  not u1721 (C3yhu6, n132);  // ../RTL/cortexm0ds_logic.v(3651)
  and u17210 (Y7yow6, M8yow6, T8yow6);  // ../RTL/cortexm0ds_logic.v(14449)
  and u17211 (n4788, vis_psp_o[20], Yfqow6);  // ../RTL/cortexm0ds_logic.v(14450)
  not u17212 (T8yow6, n4788);  // ../RTL/cortexm0ds_logic.v(14450)
  and u17213 (n4789, vis_msp_o[20], Fgqow6);  // ../RTL/cortexm0ds_logic.v(14451)
  not u17214 (M8yow6, n4789);  // ../RTL/cortexm0ds_logic.v(14451)
  and u17215 (K7yow6, A9yow6, H9yow6);  // ../RTL/cortexm0ds_logic.v(14452)
  and u17216 (n4790, vis_r14_o[22], Ahqow6);  // ../RTL/cortexm0ds_logic.v(14453)
  not u17217 (H9yow6, n4790);  // ../RTL/cortexm0ds_logic.v(14453)
  and u17218 (n4791, vis_r12_o[22], Hhqow6);  // ../RTL/cortexm0ds_logic.v(14454)
  not u17219 (A9yow6, n4791);  // ../RTL/cortexm0ds_logic.v(14454)
  and u1722 (Ak1iu6, Hk1iu6, Ok1iu6);  // ../RTL/cortexm0ds_logic.v(3652)
  and u17220 (W6yow6, O9yow6, V9yow6);  // ../RTL/cortexm0ds_logic.v(14455)
  and u17221 (V9yow6, Cayow6, Jayow6);  // ../RTL/cortexm0ds_logic.v(14456)
  and u17222 (n4792, vis_r9_o[22], Qiqow6);  // ../RTL/cortexm0ds_logic.v(14457)
  not u17223 (Jayow6, n4792);  // ../RTL/cortexm0ds_logic.v(14457)
  and u17224 (Cayow6, Qayow6, Xayow6);  // ../RTL/cortexm0ds_logic.v(14458)
  and u17225 (n4793, vis_r11_o[22], Ljqow6);  // ../RTL/cortexm0ds_logic.v(14459)
  not u17226 (Xayow6, n4793);  // ../RTL/cortexm0ds_logic.v(14459)
  and u17227 (n4794, vis_r10_o[22], Sjqow6);  // ../RTL/cortexm0ds_logic.v(14460)
  not u17228 (Qayow6, n4794);  // ../RTL/cortexm0ds_logic.v(14460)
  and u17229 (O9yow6, Tzzhu6, Ebyow6);  // ../RTL/cortexm0ds_logic.v(14461)
  and u1723 (n133, Uthpw6[7], Vk1iu6);  // ../RTL/cortexm0ds_logic.v(3653)
  and u17230 (n4795, vis_r8_o[22], Gkqow6);  // ../RTL/cortexm0ds_logic.v(14462)
  not u17231 (Ebyow6, n4795);  // ../RTL/cortexm0ds_logic.v(14462)
  and u17232 (Tzzhu6, Lbyow6, Sbyow6);  // ../RTL/cortexm0ds_logic.v(14463)
  and u17233 (Sbyow6, Zbyow6, Gcyow6);  // ../RTL/cortexm0ds_logic.v(14464)
  and u17234 (Gcyow6, Ncyow6, Ucyow6);  // ../RTL/cortexm0ds_logic.v(14465)
  and u17235 (n4796, vis_r2_o[22], Dmqow6);  // ../RTL/cortexm0ds_logic.v(14466)
  not u17236 (Ucyow6, n4796);  // ../RTL/cortexm0ds_logic.v(14466)
  and u17237 (n4797, vis_r6_o[22], Kmqow6);  // ../RTL/cortexm0ds_logic.v(14467)
  not u17238 (Ncyow6, n4797);  // ../RTL/cortexm0ds_logic.v(14467)
  and u17239 (Zbyow6, Bdyow6, Idyow6);  // ../RTL/cortexm0ds_logic.v(14468)
  not u1724 (Ok1iu6, n133);  // ../RTL/cortexm0ds_logic.v(3653)
  and u17240 (n4798, vis_r5_o[22], Fnqow6);  // ../RTL/cortexm0ds_logic.v(14469)
  not u17241 (Idyow6, n4798);  // ../RTL/cortexm0ds_logic.v(14469)
  and u17242 (n4799, vis_r4_o[22], Mnqow6);  // ../RTL/cortexm0ds_logic.v(14470)
  not u17243 (Bdyow6, n4799);  // ../RTL/cortexm0ds_logic.v(14470)
  and u17244 (Lbyow6, Pdyow6, Wdyow6);  // ../RTL/cortexm0ds_logic.v(14471)
  and u17245 (Wdyow6, Deyow6, Keyow6);  // ../RTL/cortexm0ds_logic.v(14472)
  and u17246 (n4800, vis_r1_o[22], Voqow6);  // ../RTL/cortexm0ds_logic.v(14473)
  not u17247 (Keyow6, n4800);  // ../RTL/cortexm0ds_logic.v(14473)
  and u17248 (n4801, vis_r0_o[22], Cpqow6);  // ../RTL/cortexm0ds_logic.v(14474)
  not u17249 (Deyow6, n4801);  // ../RTL/cortexm0ds_logic.v(14474)
  and u1725 (n134, Cl1iu6, Jdnhu6);  // ../RTL/cortexm0ds_logic.v(3654)
  and u17250 (Pdyow6, Reyow6, Yeyow6);  // ../RTL/cortexm0ds_logic.v(14475)
  and u17251 (n4802, vis_r3_o[22], Xpqow6);  // ../RTL/cortexm0ds_logic.v(14476)
  not u17252 (Yeyow6, n4802);  // ../RTL/cortexm0ds_logic.v(14476)
  and u17253 (n4803, vis_r7_o[22], Eqqow6);  // ../RTL/cortexm0ds_logic.v(14477)
  not u17254 (Reyow6, n4803);  // ../RTL/cortexm0ds_logic.v(14477)
  and u17255 (n4804, Lcqow6, Eg6ju6);  // ../RTL/cortexm0ds_logic.v(14479)
  not u17256 (Mfyow6, n4804);  // ../RTL/cortexm0ds_logic.v(14479)
  and u17257 (Ffyow6, Tfyow6, Agyow6);  // ../RTL/cortexm0ds_logic.v(14480)
  or u17258 (Agyow6, Yxliu6, Qaxiu6);  // ../RTL/cortexm0ds_logic.v(14481)
  not u17259 (Yxliu6, I74iu6);  // ../RTL/cortexm0ds_logic.v(14482)
  not u1726 (Hk1iu6, n134);  // ../RTL/cortexm0ds_logic.v(3654)
  and u17260 (I74iu6, Shhpw6[21], Iqzhu6);  // ../RTL/cortexm0ds_logic.v(14483)
  and u17261 (n4805, Gdqow6, Xx9ju6);  // ../RTL/cortexm0ds_logic.v(14484)
  not u17262 (Tfyow6, n4805);  // ../RTL/cortexm0ds_logic.v(14484)
  and u17263 (n4806, Hgyow6, Ogyow6);  // ../RTL/cortexm0ds_logic.v(14485)
  not u17264 (Xx9ju6, n4806);  // ../RTL/cortexm0ds_logic.v(14485)
  and u17265 (Ogyow6, Vgyow6, Chyow6);  // ../RTL/cortexm0ds_logic.v(14486)
  and u17266 (Chyow6, Jhyow6, Qhyow6);  // ../RTL/cortexm0ds_logic.v(14487)
  and u17267 (n4807, Fkfpw6[21], Dfqow6);  // ../RTL/cortexm0ds_logic.v(14488)
  not u17268 (Qhyow6, n4807);  // ../RTL/cortexm0ds_logic.v(14488)
  and u17269 (Jhyow6, Xhyow6, Eiyow6);  // ../RTL/cortexm0ds_logic.v(14489)
  and u1727 (Tj1iu6, Jl1iu6, Ql1iu6);  // ../RTL/cortexm0ds_logic.v(3655)
  and u17270 (n4808, vis_psp_o[19], Yfqow6);  // ../RTL/cortexm0ds_logic.v(14490)
  not u17271 (Eiyow6, n4808);  // ../RTL/cortexm0ds_logic.v(14490)
  and u17272 (n4809, vis_msp_o[19], Fgqow6);  // ../RTL/cortexm0ds_logic.v(14491)
  not u17273 (Xhyow6, n4809);  // ../RTL/cortexm0ds_logic.v(14491)
  and u17274 (Vgyow6, Liyow6, Siyow6);  // ../RTL/cortexm0ds_logic.v(14492)
  and u17275 (n4810, vis_r14_o[21], Ahqow6);  // ../RTL/cortexm0ds_logic.v(14493)
  not u17276 (Siyow6, n4810);  // ../RTL/cortexm0ds_logic.v(14493)
  and u17277 (n4811, vis_r12_o[21], Hhqow6);  // ../RTL/cortexm0ds_logic.v(14494)
  not u17278 (Liyow6, n4811);  // ../RTL/cortexm0ds_logic.v(14494)
  and u17279 (Hgyow6, Ziyow6, Gjyow6);  // ../RTL/cortexm0ds_logic.v(14495)
  and u1728 (n135, Iahpw6[6], Xl1iu6);  // ../RTL/cortexm0ds_logic.v(3656)
  and u17280 (Gjyow6, Njyow6, Ujyow6);  // ../RTL/cortexm0ds_logic.v(14496)
  and u17281 (n4812, vis_r9_o[21], Qiqow6);  // ../RTL/cortexm0ds_logic.v(14497)
  not u17282 (Ujyow6, n4812);  // ../RTL/cortexm0ds_logic.v(14497)
  and u17283 (Njyow6, Bkyow6, Ikyow6);  // ../RTL/cortexm0ds_logic.v(14498)
  and u17284 (n4813, vis_r11_o[21], Ljqow6);  // ../RTL/cortexm0ds_logic.v(14499)
  not u17285 (Ikyow6, n4813);  // ../RTL/cortexm0ds_logic.v(14499)
  and u17286 (n4814, vis_r10_o[21], Sjqow6);  // ../RTL/cortexm0ds_logic.v(14500)
  not u17287 (Bkyow6, n4814);  // ../RTL/cortexm0ds_logic.v(14500)
  and u17288 (Ziyow6, A00iu6, Pkyow6);  // ../RTL/cortexm0ds_logic.v(14501)
  and u17289 (n4815, vis_r8_o[21], Gkqow6);  // ../RTL/cortexm0ds_logic.v(14502)
  not u1729 (Ql1iu6, n135);  // ../RTL/cortexm0ds_logic.v(3656)
  not u17290 (Pkyow6, n4815);  // ../RTL/cortexm0ds_logic.v(14502)
  and u17291 (A00iu6, Wkyow6, Dlyow6);  // ../RTL/cortexm0ds_logic.v(14503)
  and u17292 (Dlyow6, Klyow6, Rlyow6);  // ../RTL/cortexm0ds_logic.v(14504)
  and u17293 (Rlyow6, Ylyow6, Fmyow6);  // ../RTL/cortexm0ds_logic.v(14505)
  and u17294 (n4816, vis_r2_o[21], Dmqow6);  // ../RTL/cortexm0ds_logic.v(14506)
  not u17295 (Fmyow6, n4816);  // ../RTL/cortexm0ds_logic.v(14506)
  and u17296 (n4817, vis_r6_o[21], Kmqow6);  // ../RTL/cortexm0ds_logic.v(14507)
  not u17297 (Ylyow6, n4817);  // ../RTL/cortexm0ds_logic.v(14507)
  and u17298 (Klyow6, Mmyow6, Tmyow6);  // ../RTL/cortexm0ds_logic.v(14508)
  and u17299 (n4818, vis_r5_o[21], Fnqow6);  // ../RTL/cortexm0ds_logic.v(14509)
  buf u173 (Eafpw6[6], Nxkbx6[7]);  // ../RTL/cortexm0ds_logic.v(3167)
  and u1730 (n136, Iahpw6[7], Z4yhu6);  // ../RTL/cortexm0ds_logic.v(3657)
  not u17300 (Tmyow6, n4818);  // ../RTL/cortexm0ds_logic.v(14509)
  and u17301 (n4819, vis_r4_o[21], Mnqow6);  // ../RTL/cortexm0ds_logic.v(14510)
  not u17302 (Mmyow6, n4819);  // ../RTL/cortexm0ds_logic.v(14510)
  and u17303 (Wkyow6, Anyow6, Hnyow6);  // ../RTL/cortexm0ds_logic.v(14511)
  and u17304 (Hnyow6, Onyow6, Vnyow6);  // ../RTL/cortexm0ds_logic.v(14512)
  and u17305 (n4820, vis_r1_o[21], Voqow6);  // ../RTL/cortexm0ds_logic.v(14513)
  not u17306 (Vnyow6, n4820);  // ../RTL/cortexm0ds_logic.v(14513)
  and u17307 (n4821, vis_r0_o[21], Cpqow6);  // ../RTL/cortexm0ds_logic.v(14514)
  not u17308 (Onyow6, n4821);  // ../RTL/cortexm0ds_logic.v(14514)
  and u17309 (Anyow6, Coyow6, Joyow6);  // ../RTL/cortexm0ds_logic.v(14515)
  not u1731 (Jl1iu6, n136);  // ../RTL/cortexm0ds_logic.v(3657)
  and u17310 (n4822, vis_r3_o[21], Xpqow6);  // ../RTL/cortexm0ds_logic.v(14516)
  not u17311 (Joyow6, n4822);  // ../RTL/cortexm0ds_logic.v(14516)
  and u17312 (n4823, vis_r7_o[21], Eqqow6);  // ../RTL/cortexm0ds_logic.v(14517)
  not u17313 (Coyow6, n4823);  // ../RTL/cortexm0ds_logic.v(14517)
  and u17314 (n4824, Lcqow6, Zw4ju6);  // ../RTL/cortexm0ds_logic.v(14519)
  not u17315 (Xoyow6, n4824);  // ../RTL/cortexm0ds_logic.v(14519)
  and u17316 (Qoyow6, Epyow6, Lpyow6);  // ../RTL/cortexm0ds_logic.v(14520)
  and u17317 (n4825, B74iu6, R0nhu6);  // ../RTL/cortexm0ds_logic.v(14521)
  not u17318 (Lpyow6, n4825);  // ../RTL/cortexm0ds_logic.v(14521)
  and u17319 (B74iu6, Shhpw6[20], Iqzhu6);  // ../RTL/cortexm0ds_logic.v(14522)
  AL_MUX u1732 (
    .i0(Shhpw6[31]),
    .i1(Iahpw6[30]),
    .sel(Em1iu6),
    .o(V2yhu6));  // ../RTL/cortexm0ds_logic.v(3658)
  and u17320 (n4826, Gdqow6, Wt9ju6);  // ../RTL/cortexm0ds_logic.v(14523)
  not u17321 (Epyow6, n4826);  // ../RTL/cortexm0ds_logic.v(14523)
  and u17322 (n4827, Spyow6, Zpyow6);  // ../RTL/cortexm0ds_logic.v(14524)
  not u17323 (Wt9ju6, n4827);  // ../RTL/cortexm0ds_logic.v(14524)
  and u17324 (Zpyow6, Gqyow6, Nqyow6);  // ../RTL/cortexm0ds_logic.v(14525)
  and u17325 (Nqyow6, Uqyow6, Bryow6);  // ../RTL/cortexm0ds_logic.v(14526)
  and u17326 (n4828, Fkfpw6[20], Dfqow6);  // ../RTL/cortexm0ds_logic.v(14527)
  not u17327 (Bryow6, n4828);  // ../RTL/cortexm0ds_logic.v(14527)
  and u17328 (Uqyow6, Iryow6, Pryow6);  // ../RTL/cortexm0ds_logic.v(14528)
  and u17329 (n4829, vis_psp_o[18], Yfqow6);  // ../RTL/cortexm0ds_logic.v(14529)
  AL_MUX u1733 (
    .i0(Jshpw6[31]),
    .i1(Lm1iu6),
    .sel(Sm1iu6),
    .o(O2yhu6));  // ../RTL/cortexm0ds_logic.v(3659)
  not u17330 (Pryow6, n4829);  // ../RTL/cortexm0ds_logic.v(14529)
  and u17331 (n4830, vis_msp_o[18], Fgqow6);  // ../RTL/cortexm0ds_logic.v(14530)
  not u17332 (Iryow6, n4830);  // ../RTL/cortexm0ds_logic.v(14530)
  and u17333 (Gqyow6, Wryow6, Dsyow6);  // ../RTL/cortexm0ds_logic.v(14531)
  and u17334 (n4831, vis_r14_o[20], Ahqow6);  // ../RTL/cortexm0ds_logic.v(14532)
  not u17335 (Dsyow6, n4831);  // ../RTL/cortexm0ds_logic.v(14532)
  and u17336 (n4832, vis_r12_o[20], Hhqow6);  // ../RTL/cortexm0ds_logic.v(14533)
  not u17337 (Wryow6, n4832);  // ../RTL/cortexm0ds_logic.v(14533)
  and u17338 (Spyow6, Ksyow6, Rsyow6);  // ../RTL/cortexm0ds_logic.v(14534)
  and u17339 (Rsyow6, Ysyow6, Ftyow6);  // ../RTL/cortexm0ds_logic.v(14535)
  and u1734 (n137, Zm1iu6, Gn1iu6);  // ../RTL/cortexm0ds_logic.v(3660)
  and u17340 (n4833, vis_r9_o[20], Qiqow6);  // ../RTL/cortexm0ds_logic.v(14536)
  not u17341 (Ftyow6, n4833);  // ../RTL/cortexm0ds_logic.v(14536)
  and u17342 (Ysyow6, Mtyow6, Ttyow6);  // ../RTL/cortexm0ds_logic.v(14537)
  and u17343 (n4834, vis_r11_o[20], Ljqow6);  // ../RTL/cortexm0ds_logic.v(14538)
  not u17344 (Ttyow6, n4834);  // ../RTL/cortexm0ds_logic.v(14538)
  and u17345 (n4835, vis_r10_o[20], Sjqow6);  // ../RTL/cortexm0ds_logic.v(14539)
  not u17346 (Mtyow6, n4835);  // ../RTL/cortexm0ds_logic.v(14539)
  and u17347 (Ksyow6, H00iu6, Auyow6);  // ../RTL/cortexm0ds_logic.v(14540)
  and u17348 (n4836, vis_r8_o[20], Gkqow6);  // ../RTL/cortexm0ds_logic.v(14541)
  not u17349 (Auyow6, n4836);  // ../RTL/cortexm0ds_logic.v(14541)
  not u1735 (H2yhu6, n137);  // ../RTL/cortexm0ds_logic.v(3660)
  and u17350 (H00iu6, Huyow6, Ouyow6);  // ../RTL/cortexm0ds_logic.v(14542)
  and u17351 (Ouyow6, Vuyow6, Cvyow6);  // ../RTL/cortexm0ds_logic.v(14543)
  and u17352 (Cvyow6, Jvyow6, Qvyow6);  // ../RTL/cortexm0ds_logic.v(14544)
  and u17353 (n4837, vis_r2_o[20], Dmqow6);  // ../RTL/cortexm0ds_logic.v(14545)
  not u17354 (Qvyow6, n4837);  // ../RTL/cortexm0ds_logic.v(14545)
  and u17355 (n4838, vis_r6_o[20], Kmqow6);  // ../RTL/cortexm0ds_logic.v(14546)
  not u17356 (Jvyow6, n4838);  // ../RTL/cortexm0ds_logic.v(14546)
  and u17357 (Vuyow6, Xvyow6, Ewyow6);  // ../RTL/cortexm0ds_logic.v(14547)
  and u17358 (n4839, vis_r5_o[20], Fnqow6);  // ../RTL/cortexm0ds_logic.v(14548)
  not u17359 (Ewyow6, n4839);  // ../RTL/cortexm0ds_logic.v(14548)
  and u1736 (Gn1iu6, Nn1iu6, Un1iu6);  // ../RTL/cortexm0ds_logic.v(3661)
  and u17360 (n4840, vis_r4_o[20], Mnqow6);  // ../RTL/cortexm0ds_logic.v(14549)
  not u17361 (Xvyow6, n4840);  // ../RTL/cortexm0ds_logic.v(14549)
  and u17362 (Huyow6, Lwyow6, Swyow6);  // ../RTL/cortexm0ds_logic.v(14550)
  and u17363 (Swyow6, Zwyow6, Gxyow6);  // ../RTL/cortexm0ds_logic.v(14551)
  and u17364 (n4841, vis_r1_o[20], Voqow6);  // ../RTL/cortexm0ds_logic.v(14552)
  not u17365 (Gxyow6, n4841);  // ../RTL/cortexm0ds_logic.v(14552)
  and u17366 (n4842, vis_r0_o[20], Cpqow6);  // ../RTL/cortexm0ds_logic.v(14553)
  not u17367 (Zwyow6, n4842);  // ../RTL/cortexm0ds_logic.v(14553)
  and u17368 (Lwyow6, Nxyow6, Uxyow6);  // ../RTL/cortexm0ds_logic.v(14554)
  and u17369 (n4843, vis_r3_o[20], Xpqow6);  // ../RTL/cortexm0ds_logic.v(14555)
  and u1737 (n138, Bo1iu6, Jshpw6[31]);  // ../RTL/cortexm0ds_logic.v(3662)
  not u17370 (Uxyow6, n4843);  // ../RTL/cortexm0ds_logic.v(14555)
  and u17371 (n4844, vis_r7_o[20], Eqqow6);  // ../RTL/cortexm0ds_logic.v(14556)
  not u17372 (Nxyow6, n4844);  // ../RTL/cortexm0ds_logic.v(14556)
  or u17373 (Iyyow6, A34iu6, Qaxiu6);  // ../RTL/cortexm0ds_logic.v(14558)
  not u17374 (A34iu6, O34iu6);  // ../RTL/cortexm0ds_logic.v(14559)
  and u17375 (O34iu6, Shhpw6[1], Iqzhu6);  // ../RTL/cortexm0ds_logic.v(14560)
  and u17376 (n4845, Sevow6, Znliu6);  // ../RTL/cortexm0ds_logic.v(14561)
  not u17377 (Byyow6, n4845);  // ../RTL/cortexm0ds_logic.v(14561)
  and u17378 (n4846, Lcqow6, G36ju6);  // ../RTL/cortexm0ds_logic.v(14563)
  not u17379 (Wyyow6, n4846);  // ../RTL/cortexm0ds_logic.v(14563)
  not u1738 (Un1iu6, n138);  // ../RTL/cortexm0ds_logic.v(3662)
  and u17380 (Pyyow6, Dzyow6, Kzyow6);  // ../RTL/cortexm0ds_logic.v(14564)
  and u17381 (n4847, U64iu6, R0nhu6);  // ../RTL/cortexm0ds_logic.v(14565)
  not u17382 (Kzyow6, n4847);  // ../RTL/cortexm0ds_logic.v(14565)
  and u17383 (U64iu6, Shhpw6[19], Iqzhu6);  // ../RTL/cortexm0ds_logic.v(14566)
  and u17384 (n4848, Gdqow6, Vp9ju6);  // ../RTL/cortexm0ds_logic.v(14567)
  not u17385 (Dzyow6, n4848);  // ../RTL/cortexm0ds_logic.v(14567)
  and u17386 (n4849, Rzyow6, Yzyow6);  // ../RTL/cortexm0ds_logic.v(14568)
  not u17387 (Vp9ju6, n4849);  // ../RTL/cortexm0ds_logic.v(14568)
  and u17388 (Yzyow6, F0zow6, M0zow6);  // ../RTL/cortexm0ds_logic.v(14569)
  and u17389 (M0zow6, T0zow6, A1zow6);  // ../RTL/cortexm0ds_logic.v(14570)
  and u1739 (Nn1iu6, Io1iu6, Po1iu6);  // ../RTL/cortexm0ds_logic.v(3663)
  and u17390 (n4850, Fkfpw6[19], Dfqow6);  // ../RTL/cortexm0ds_logic.v(14571)
  not u17391 (A1zow6, n4850);  // ../RTL/cortexm0ds_logic.v(14571)
  and u17392 (T0zow6, H1zow6, O1zow6);  // ../RTL/cortexm0ds_logic.v(14572)
  and u17393 (n4851, vis_psp_o[17], Yfqow6);  // ../RTL/cortexm0ds_logic.v(14573)
  not u17394 (O1zow6, n4851);  // ../RTL/cortexm0ds_logic.v(14573)
  and u17395 (n4852, vis_msp_o[17], Fgqow6);  // ../RTL/cortexm0ds_logic.v(14574)
  not u17396 (H1zow6, n4852);  // ../RTL/cortexm0ds_logic.v(14574)
  and u17397 (F0zow6, V1zow6, C2zow6);  // ../RTL/cortexm0ds_logic.v(14575)
  and u17398 (n4853, vis_r14_o[19], Ahqow6);  // ../RTL/cortexm0ds_logic.v(14576)
  not u17399 (C2zow6, n4853);  // ../RTL/cortexm0ds_logic.v(14576)
  buf u174 (V9ghu6, F9vpw6);  // ../RTL/cortexm0ds_logic.v(2019)
  and u1740 (n139, Wo1iu6, Dp1iu6);  // ../RTL/cortexm0ds_logic.v(3664)
  and u17400 (n4854, vis_r12_o[19], Hhqow6);  // ../RTL/cortexm0ds_logic.v(14577)
  not u17401 (V1zow6, n4854);  // ../RTL/cortexm0ds_logic.v(14577)
  and u17402 (Rzyow6, J2zow6, Q2zow6);  // ../RTL/cortexm0ds_logic.v(14578)
  and u17403 (Q2zow6, X2zow6, E3zow6);  // ../RTL/cortexm0ds_logic.v(14579)
  and u17404 (n4855, vis_r9_o[19], Qiqow6);  // ../RTL/cortexm0ds_logic.v(14580)
  not u17405 (E3zow6, n4855);  // ../RTL/cortexm0ds_logic.v(14580)
  and u17406 (X2zow6, L3zow6, S3zow6);  // ../RTL/cortexm0ds_logic.v(14581)
  and u17407 (n4856, vis_r11_o[19], Ljqow6);  // ../RTL/cortexm0ds_logic.v(14582)
  not u17408 (S3zow6, n4856);  // ../RTL/cortexm0ds_logic.v(14582)
  and u17409 (n4857, vis_r10_o[19], Sjqow6);  // ../RTL/cortexm0ds_logic.v(14583)
  not u1741 (Io1iu6, n139);  // ../RTL/cortexm0ds_logic.v(3664)
  not u17410 (L3zow6, n4857);  // ../RTL/cortexm0ds_logic.v(14583)
  and u17411 (J2zow6, V00iu6, Z3zow6);  // ../RTL/cortexm0ds_logic.v(14584)
  and u17412 (n4858, vis_r8_o[19], Gkqow6);  // ../RTL/cortexm0ds_logic.v(14585)
  not u17413 (Z3zow6, n4858);  // ../RTL/cortexm0ds_logic.v(14585)
  and u17414 (V00iu6, G4zow6, N4zow6);  // ../RTL/cortexm0ds_logic.v(14586)
  and u17415 (N4zow6, U4zow6, B5zow6);  // ../RTL/cortexm0ds_logic.v(14587)
  and u17416 (B5zow6, I5zow6, P5zow6);  // ../RTL/cortexm0ds_logic.v(14588)
  and u17417 (n4859, vis_r2_o[19], Dmqow6);  // ../RTL/cortexm0ds_logic.v(14589)
  not u17418 (P5zow6, n4859);  // ../RTL/cortexm0ds_logic.v(14589)
  and u17419 (n4860, vis_r6_o[19], Kmqow6);  // ../RTL/cortexm0ds_logic.v(14590)
  and u1742 (n140, Kp1iu6, Rp1iu6);  // ../RTL/cortexm0ds_logic.v(3665)
  not u17420 (I5zow6, n4860);  // ../RTL/cortexm0ds_logic.v(14590)
  and u17421 (U4zow6, W5zow6, D6zow6);  // ../RTL/cortexm0ds_logic.v(14591)
  and u17422 (n4861, vis_r5_o[19], Fnqow6);  // ../RTL/cortexm0ds_logic.v(14592)
  not u17423 (D6zow6, n4861);  // ../RTL/cortexm0ds_logic.v(14592)
  and u17424 (n4862, vis_r4_o[19], Mnqow6);  // ../RTL/cortexm0ds_logic.v(14593)
  not u17425 (W5zow6, n4862);  // ../RTL/cortexm0ds_logic.v(14593)
  and u17426 (G4zow6, K6zow6, R6zow6);  // ../RTL/cortexm0ds_logic.v(14594)
  and u17427 (R6zow6, Y6zow6, F7zow6);  // ../RTL/cortexm0ds_logic.v(14595)
  and u17428 (n4863, vis_r1_o[19], Voqow6);  // ../RTL/cortexm0ds_logic.v(14596)
  not u17429 (F7zow6, n4863);  // ../RTL/cortexm0ds_logic.v(14596)
  not u1743 (Dp1iu6, n140);  // ../RTL/cortexm0ds_logic.v(3665)
  and u17430 (n4864, vis_r0_o[19], Cpqow6);  // ../RTL/cortexm0ds_logic.v(14597)
  not u17431 (Y6zow6, n4864);  // ../RTL/cortexm0ds_logic.v(14597)
  and u17432 (K6zow6, M7zow6, T7zow6);  // ../RTL/cortexm0ds_logic.v(14598)
  and u17433 (n4865, vis_r3_o[19], Xpqow6);  // ../RTL/cortexm0ds_logic.v(14599)
  not u17434 (T7zow6, n4865);  // ../RTL/cortexm0ds_logic.v(14599)
  and u17435 (n4866, vis_r7_o[19], Eqqow6);  // ../RTL/cortexm0ds_logic.v(14600)
  not u17436 (M7zow6, n4866);  // ../RTL/cortexm0ds_logic.v(14600)
  and u17437 (n4867, Lcqow6, Ot5ju6);  // ../RTL/cortexm0ds_logic.v(14602)
  not u17438 (H8zow6, n4867);  // ../RTL/cortexm0ds_logic.v(14602)
  and u17439 (A8zow6, O8zow6, V8zow6);  // ../RTL/cortexm0ds_logic.v(14603)
  and u1744 (Rp1iu6, Yp1iu6, Fq1iu6);  // ../RTL/cortexm0ds_logic.v(3666)
  and u17440 (n4868, N64iu6, R0nhu6);  // ../RTL/cortexm0ds_logic.v(14604)
  not u17441 (V8zow6, n4868);  // ../RTL/cortexm0ds_logic.v(14604)
  and u17442 (N64iu6, Shhpw6[18], Iqzhu6);  // ../RTL/cortexm0ds_logic.v(14605)
  and u17443 (n4869, Gdqow6, Gl9ju6);  // ../RTL/cortexm0ds_logic.v(14606)
  not u17444 (O8zow6, n4869);  // ../RTL/cortexm0ds_logic.v(14606)
  and u17445 (n4870, C9zow6, J9zow6);  // ../RTL/cortexm0ds_logic.v(14607)
  not u17446 (Gl9ju6, n4870);  // ../RTL/cortexm0ds_logic.v(14607)
  and u17447 (J9zow6, Q9zow6, X9zow6);  // ../RTL/cortexm0ds_logic.v(14608)
  and u17448 (X9zow6, Eazow6, Lazow6);  // ../RTL/cortexm0ds_logic.v(14609)
  and u17449 (n4871, Fkfpw6[18], Dfqow6);  // ../RTL/cortexm0ds_logic.v(14610)
  and u1745 (Fq1iu6, Mq1iu6, Tq1iu6);  // ../RTL/cortexm0ds_logic.v(3667)
  not u17450 (Lazow6, n4871);  // ../RTL/cortexm0ds_logic.v(14610)
  and u17451 (Eazow6, Sazow6, Zazow6);  // ../RTL/cortexm0ds_logic.v(14611)
  and u17452 (n4872, vis_psp_o[16], Yfqow6);  // ../RTL/cortexm0ds_logic.v(14612)
  not u17453 (Zazow6, n4872);  // ../RTL/cortexm0ds_logic.v(14612)
  and u17454 (n4873, vis_msp_o[16], Fgqow6);  // ../RTL/cortexm0ds_logic.v(14613)
  not u17455 (Sazow6, n4873);  // ../RTL/cortexm0ds_logic.v(14613)
  and u17456 (Q9zow6, Gbzow6, Nbzow6);  // ../RTL/cortexm0ds_logic.v(14614)
  and u17457 (n4874, vis_r14_o[18], Ahqow6);  // ../RTL/cortexm0ds_logic.v(14615)
  not u17458 (Nbzow6, n4874);  // ../RTL/cortexm0ds_logic.v(14615)
  and u17459 (n4875, vis_r12_o[18], Hhqow6);  // ../RTL/cortexm0ds_logic.v(14616)
  and u1746 (n141, Ar1iu6, Fkfpw6[31]);  // ../RTL/cortexm0ds_logic.v(3668)
  not u17460 (Gbzow6, n4875);  // ../RTL/cortexm0ds_logic.v(14616)
  and u17461 (C9zow6, Ubzow6, Bczow6);  // ../RTL/cortexm0ds_logic.v(14617)
  and u17462 (Bczow6, Iczow6, Pczow6);  // ../RTL/cortexm0ds_logic.v(14618)
  and u17463 (n4876, vis_r9_o[18], Qiqow6);  // ../RTL/cortexm0ds_logic.v(14619)
  not u17464 (Pczow6, n4876);  // ../RTL/cortexm0ds_logic.v(14619)
  and u17465 (Iczow6, Wczow6, Ddzow6);  // ../RTL/cortexm0ds_logic.v(14620)
  and u17466 (n4877, vis_r11_o[18], Ljqow6);  // ../RTL/cortexm0ds_logic.v(14621)
  not u17467 (Ddzow6, n4877);  // ../RTL/cortexm0ds_logic.v(14621)
  and u17468 (n4878, vis_r10_o[18], Sjqow6);  // ../RTL/cortexm0ds_logic.v(14622)
  not u17469 (Wczow6, n4878);  // ../RTL/cortexm0ds_logic.v(14622)
  not u1747 (Tq1iu6, n141);  // ../RTL/cortexm0ds_logic.v(3668)
  and u17470 (Ubzow6, C10iu6, Kdzow6);  // ../RTL/cortexm0ds_logic.v(14623)
  and u17471 (n4879, vis_r8_o[18], Gkqow6);  // ../RTL/cortexm0ds_logic.v(14624)
  not u17472 (Kdzow6, n4879);  // ../RTL/cortexm0ds_logic.v(14624)
  and u17473 (C10iu6, Rdzow6, Ydzow6);  // ../RTL/cortexm0ds_logic.v(14625)
  and u17474 (Ydzow6, Fezow6, Mezow6);  // ../RTL/cortexm0ds_logic.v(14626)
  and u17475 (Mezow6, Tezow6, Afzow6);  // ../RTL/cortexm0ds_logic.v(14627)
  and u17476 (n4880, vis_r2_o[18], Dmqow6);  // ../RTL/cortexm0ds_logic.v(14628)
  not u17477 (Afzow6, n4880);  // ../RTL/cortexm0ds_logic.v(14628)
  and u17478 (n4881, vis_r6_o[18], Kmqow6);  // ../RTL/cortexm0ds_logic.v(14629)
  not u17479 (Tezow6, n4881);  // ../RTL/cortexm0ds_logic.v(14629)
  and u1748 (Mq1iu6, Hr1iu6, Or1iu6);  // ../RTL/cortexm0ds_logic.v(3669)
  and u17480 (Fezow6, Hfzow6, Ofzow6);  // ../RTL/cortexm0ds_logic.v(14630)
  and u17481 (n4882, vis_r5_o[18], Fnqow6);  // ../RTL/cortexm0ds_logic.v(14631)
  not u17482 (Ofzow6, n4882);  // ../RTL/cortexm0ds_logic.v(14631)
  and u17483 (n4883, vis_r4_o[18], Mnqow6);  // ../RTL/cortexm0ds_logic.v(14632)
  not u17484 (Hfzow6, n4883);  // ../RTL/cortexm0ds_logic.v(14632)
  and u17485 (Rdzow6, Vfzow6, Cgzow6);  // ../RTL/cortexm0ds_logic.v(14633)
  and u17486 (Cgzow6, Jgzow6, Qgzow6);  // ../RTL/cortexm0ds_logic.v(14634)
  and u17487 (n4884, vis_r1_o[18], Voqow6);  // ../RTL/cortexm0ds_logic.v(14635)
  not u17488 (Qgzow6, n4884);  // ../RTL/cortexm0ds_logic.v(14635)
  and u17489 (n4885, vis_r0_o[18], Cpqow6);  // ../RTL/cortexm0ds_logic.v(14636)
  and u1749 (n142, Ligpw6[28], Vr1iu6);  // ../RTL/cortexm0ds_logic.v(3670)
  not u17490 (Jgzow6, n4885);  // ../RTL/cortexm0ds_logic.v(14636)
  and u17491 (Vfzow6, Xgzow6, Ehzow6);  // ../RTL/cortexm0ds_logic.v(14637)
  and u17492 (n4886, vis_r3_o[18], Xpqow6);  // ../RTL/cortexm0ds_logic.v(14638)
  not u17493 (Ehzow6, n4886);  // ../RTL/cortexm0ds_logic.v(14638)
  and u17494 (n4887, vis_r7_o[18], Eqqow6);  // ../RTL/cortexm0ds_logic.v(14639)
  not u17495 (Xgzow6, n4887);  // ../RTL/cortexm0ds_logic.v(14639)
  and u17496 (n4888, Lcqow6, Znliu6);  // ../RTL/cortexm0ds_logic.v(14641)
  not u17497 (Shzow6, n4888);  // ../RTL/cortexm0ds_logic.v(14641)
  and u17498 (n4889, Zhzow6, Gizow6);  // ../RTL/cortexm0ds_logic.v(14642)
  not u17499 (Znliu6, n4889);  // ../RTL/cortexm0ds_logic.v(14642)
  buf u175 (vis_r4_o[4], C2uax6);  // ../RTL/cortexm0ds_logic.v(2626)
  not u1750 (Or1iu6, n142);  // ../RTL/cortexm0ds_logic.v(3670)
  and u17500 (Gizow6, Nizow6, Uizow6);  // ../RTL/cortexm0ds_logic.v(14643)
  and u17501 (Uizow6, Bjzow6, Ijzow6);  // ../RTL/cortexm0ds_logic.v(14644)
  and u17502 (n4890, Fkfpw6[1], Dfqow6);  // ../RTL/cortexm0ds_logic.v(14645)
  not u17503 (Ijzow6, n4890);  // ../RTL/cortexm0ds_logic.v(14645)
  and u17504 (n4891, vis_r14_o[1], Ahqow6);  // ../RTL/cortexm0ds_logic.v(14646)
  not u17505 (Bjzow6, n4891);  // ../RTL/cortexm0ds_logic.v(14646)
  and u17506 (Nizow6, Pjzow6, Wjzow6);  // ../RTL/cortexm0ds_logic.v(14647)
  and u17507 (n4892, vis_r12_o[1], Hhqow6);  // ../RTL/cortexm0ds_logic.v(14648)
  not u17508 (Wjzow6, n4892);  // ../RTL/cortexm0ds_logic.v(14648)
  and u17509 (n4893, vis_r11_o[1], Ljqow6);  // ../RTL/cortexm0ds_logic.v(14649)
  and u1751 (n143, Engpw6[28], Cs1iu6);  // ../RTL/cortexm0ds_logic.v(3671)
  not u17510 (Pjzow6, n4893);  // ../RTL/cortexm0ds_logic.v(14649)
  and u17511 (Zhzow6, Dkzow6, Kkzow6);  // ../RTL/cortexm0ds_logic.v(14650)
  and u17512 (Kkzow6, Rkzow6, Ykzow6);  // ../RTL/cortexm0ds_logic.v(14651)
  and u17513 (n4894, vis_r10_o[1], Sjqow6);  // ../RTL/cortexm0ds_logic.v(14652)
  not u17514 (Ykzow6, n4894);  // ../RTL/cortexm0ds_logic.v(14652)
  and u17515 (n4895, vis_r9_o[1], Qiqow6);  // ../RTL/cortexm0ds_logic.v(14653)
  not u17516 (Rkzow6, n4895);  // ../RTL/cortexm0ds_logic.v(14653)
  and u17517 (Dkzow6, O00iu6, Flzow6);  // ../RTL/cortexm0ds_logic.v(14654)
  and u17518 (n4896, vis_r8_o[1], Gkqow6);  // ../RTL/cortexm0ds_logic.v(14655)
  not u17519 (Flzow6, n4896);  // ../RTL/cortexm0ds_logic.v(14655)
  not u1752 (Hr1iu6, n143);  // ../RTL/cortexm0ds_logic.v(3671)
  and u17520 (O00iu6, Mlzow6, Tlzow6);  // ../RTL/cortexm0ds_logic.v(14656)
  and u17521 (Tlzow6, Amzow6, Hmzow6);  // ../RTL/cortexm0ds_logic.v(14657)
  and u17522 (Hmzow6, Omzow6, Vmzow6);  // ../RTL/cortexm0ds_logic.v(14658)
  and u17523 (n4897, vis_r0_o[1], Cpqow6);  // ../RTL/cortexm0ds_logic.v(14659)
  not u17524 (Vmzow6, n4897);  // ../RTL/cortexm0ds_logic.v(14659)
  and u17525 (n4898, vis_r2_o[1], Dmqow6);  // ../RTL/cortexm0ds_logic.v(14660)
  not u17526 (Omzow6, n4898);  // ../RTL/cortexm0ds_logic.v(14660)
  and u17527 (Amzow6, Cnzow6, Jnzow6);  // ../RTL/cortexm0ds_logic.v(14661)
  and u17528 (n4899, vis_r5_o[1], Fnqow6);  // ../RTL/cortexm0ds_logic.v(14662)
  not u17529 (Jnzow6, n4899);  // ../RTL/cortexm0ds_logic.v(14662)
  and u1753 (Yp1iu6, Js1iu6, Qs1iu6);  // ../RTL/cortexm0ds_logic.v(3672)
  and u17530 (n4900, vis_r4_o[1], Mnqow6);  // ../RTL/cortexm0ds_logic.v(14663)
  not u17531 (Cnzow6, n4900);  // ../RTL/cortexm0ds_logic.v(14663)
  and u17532 (Mlzow6, Qnzow6, Xnzow6);  // ../RTL/cortexm0ds_logic.v(14664)
  and u17533 (Xnzow6, Eozow6, Lozow6);  // ../RTL/cortexm0ds_logic.v(14665)
  and u17534 (n4901, vis_r7_o[1], Eqqow6);  // ../RTL/cortexm0ds_logic.v(14666)
  not u17535 (Lozow6, n4901);  // ../RTL/cortexm0ds_logic.v(14666)
  and u17536 (n4902, vis_r3_o[1], Xpqow6);  // ../RTL/cortexm0ds_logic.v(14667)
  not u17537 (Eozow6, n4902);  // ../RTL/cortexm0ds_logic.v(14667)
  and u17538 (Qnzow6, Sozow6, Zozow6);  // ../RTL/cortexm0ds_logic.v(14668)
  and u17539 (n4903, vis_r1_o[1], Voqow6);  // ../RTL/cortexm0ds_logic.v(14669)
  and u1754 (n144, Akgpw6[28], Xs1iu6);  // ../RTL/cortexm0ds_logic.v(3673)
  not u17540 (Zozow6, n4903);  // ../RTL/cortexm0ds_logic.v(14669)
  and u17541 (n4904, vis_r6_o[1], Kmqow6);  // ../RTL/cortexm0ds_logic.v(14670)
  not u17542 (Sozow6, n4904);  // ../RTL/cortexm0ds_logic.v(14670)
  and u17543 (Lcqow6, Gpzow6, Qaxiu6);  // ../RTL/cortexm0ds_logic.v(14671)
  and u17544 (n4905, L3ehu6, X71iu6);  // ../RTL/cortexm0ds_logic.v(14672)
  not u17545 (Gpzow6, n4905);  // ../RTL/cortexm0ds_logic.v(14672)
  and u17546 (Lhzow6, Npzow6, Upzow6);  // ../RTL/cortexm0ds_logic.v(14673)
  and u17547 (n4906, Gdqow6, Fh9ju6);  // ../RTL/cortexm0ds_logic.v(14674)
  not u17548 (Upzow6, n4906);  // ../RTL/cortexm0ds_logic.v(14674)
  and u17549 (n4907, Bqzow6, Iqzow6);  // ../RTL/cortexm0ds_logic.v(14675)
  not u1755 (Qs1iu6, n144);  // ../RTL/cortexm0ds_logic.v(3673)
  not u17550 (Fh9ju6, n4907);  // ../RTL/cortexm0ds_logic.v(14675)
  and u17551 (Iqzow6, Pqzow6, Wqzow6);  // ../RTL/cortexm0ds_logic.v(14676)
  and u17552 (Wqzow6, Drzow6, Krzow6);  // ../RTL/cortexm0ds_logic.v(14677)
  and u17553 (n4908, Fkfpw6[17], Dfqow6);  // ../RTL/cortexm0ds_logic.v(14678)
  not u17554 (Krzow6, n4908);  // ../RTL/cortexm0ds_logic.v(14678)
  and u17555 (Drzow6, Rrzow6, Yrzow6);  // ../RTL/cortexm0ds_logic.v(14679)
  and u17556 (n4909, vis_psp_o[15], Yfqow6);  // ../RTL/cortexm0ds_logic.v(14680)
  not u17557 (Yrzow6, n4909);  // ../RTL/cortexm0ds_logic.v(14680)
  and u17558 (n4910, vis_msp_o[15], Fgqow6);  // ../RTL/cortexm0ds_logic.v(14681)
  not u17559 (Rrzow6, n4910);  // ../RTL/cortexm0ds_logic.v(14681)
  and u1756 (Js1iu6, Et1iu6, Lt1iu6);  // ../RTL/cortexm0ds_logic.v(3674)
  and u17560 (Pqzow6, Fszow6, Mszow6);  // ../RTL/cortexm0ds_logic.v(14682)
  and u17561 (n4911, vis_r14_o[17], Ahqow6);  // ../RTL/cortexm0ds_logic.v(14683)
  not u17562 (Mszow6, n4911);  // ../RTL/cortexm0ds_logic.v(14683)
  and u17563 (n4912, vis_r12_o[17], Hhqow6);  // ../RTL/cortexm0ds_logic.v(14684)
  not u17564 (Fszow6, n4912);  // ../RTL/cortexm0ds_logic.v(14684)
  and u17565 (Bqzow6, Tszow6, Atzow6);  // ../RTL/cortexm0ds_logic.v(14685)
  and u17566 (Atzow6, Htzow6, Otzow6);  // ../RTL/cortexm0ds_logic.v(14686)
  and u17567 (n4913, vis_r9_o[17], Qiqow6);  // ../RTL/cortexm0ds_logic.v(14687)
  not u17568 (Otzow6, n4913);  // ../RTL/cortexm0ds_logic.v(14687)
  and u17569 (Htzow6, Vtzow6, Cuzow6);  // ../RTL/cortexm0ds_logic.v(14688)
  and u1757 (n145, HRDATA[31], St1iu6);  // ../RTL/cortexm0ds_logic.v(3675)
  and u17570 (n4914, vis_r11_o[17], Ljqow6);  // ../RTL/cortexm0ds_logic.v(14689)
  not u17571 (Cuzow6, n4914);  // ../RTL/cortexm0ds_logic.v(14689)
  and u17572 (n4915, vis_r10_o[17], Sjqow6);  // ../RTL/cortexm0ds_logic.v(14690)
  not u17573 (Vtzow6, n4915);  // ../RTL/cortexm0ds_logic.v(14690)
  and u17574 (Tszow6, J10iu6, Juzow6);  // ../RTL/cortexm0ds_logic.v(14691)
  and u17575 (n4916, vis_r8_o[17], Gkqow6);  // ../RTL/cortexm0ds_logic.v(14692)
  not u17576 (Juzow6, n4916);  // ../RTL/cortexm0ds_logic.v(14692)
  and u17577 (J10iu6, Quzow6, Xuzow6);  // ../RTL/cortexm0ds_logic.v(14693)
  and u17578 (Xuzow6, Evzow6, Lvzow6);  // ../RTL/cortexm0ds_logic.v(14694)
  and u17579 (Lvzow6, Svzow6, Zvzow6);  // ../RTL/cortexm0ds_logic.v(14695)
  not u1758 (Lt1iu6, n145);  // ../RTL/cortexm0ds_logic.v(3675)
  and u17580 (n4917, vis_r2_o[17], Dmqow6);  // ../RTL/cortexm0ds_logic.v(14696)
  not u17581 (Zvzow6, n4917);  // ../RTL/cortexm0ds_logic.v(14696)
  and u17582 (n4918, vis_r6_o[17], Kmqow6);  // ../RTL/cortexm0ds_logic.v(14697)
  not u17583 (Svzow6, n4918);  // ../RTL/cortexm0ds_logic.v(14697)
  and u17584 (Evzow6, Gwzow6, Nwzow6);  // ../RTL/cortexm0ds_logic.v(14698)
  and u17585 (n4919, vis_r5_o[17], Fnqow6);  // ../RTL/cortexm0ds_logic.v(14699)
  not u17586 (Nwzow6, n4919);  // ../RTL/cortexm0ds_logic.v(14699)
  and u17587 (n4920, vis_r4_o[17], Mnqow6);  // ../RTL/cortexm0ds_logic.v(14700)
  not u17588 (Gwzow6, n4920);  // ../RTL/cortexm0ds_logic.v(14700)
  and u17589 (Quzow6, Uwzow6, Bxzow6);  // ../RTL/cortexm0ds_logic.v(14701)
  and u1759 (n146, E1hpw6[31], Zt1iu6);  // ../RTL/cortexm0ds_logic.v(3676)
  and u17590 (Bxzow6, Ixzow6, Pxzow6);  // ../RTL/cortexm0ds_logic.v(14702)
  and u17591 (n4921, vis_r1_o[17], Voqow6);  // ../RTL/cortexm0ds_logic.v(14703)
  not u17592 (Pxzow6, n4921);  // ../RTL/cortexm0ds_logic.v(14703)
  and u17593 (n4922, vis_r0_o[17], Cpqow6);  // ../RTL/cortexm0ds_logic.v(14704)
  not u17594 (Ixzow6, n4922);  // ../RTL/cortexm0ds_logic.v(14704)
  and u17595 (Uwzow6, Wxzow6, Dyzow6);  // ../RTL/cortexm0ds_logic.v(14705)
  and u17596 (n4923, vis_r3_o[17], Xpqow6);  // ../RTL/cortexm0ds_logic.v(14706)
  not u17597 (Dyzow6, n4923);  // ../RTL/cortexm0ds_logic.v(14706)
  and u17598 (n4924, vis_r7_o[17], Eqqow6);  // ../RTL/cortexm0ds_logic.v(14707)
  not u17599 (Wxzow6, n4924);  // ../RTL/cortexm0ds_logic.v(14707)
  buf u176 (vis_r14_o[1], Onypw6);  // ../RTL/cortexm0ds_logic.v(2497)
  not u1760 (Et1iu6, n146);  // ../RTL/cortexm0ds_logic.v(3676)
  and u17600 (Gdqow6, Sevow6, X71iu6);  // ../RTL/cortexm0ds_logic.v(14708)
  and u17601 (n4925, G64iu6, R0nhu6);  // ../RTL/cortexm0ds_logic.v(14709)
  not u17602 (Npzow6, n4925);  // ../RTL/cortexm0ds_logic.v(14709)
  and u17603 (G64iu6, Shhpw6[17], Iqzhu6);  // ../RTL/cortexm0ds_logic.v(14710)
  and u17604 (n4926, Yyzow6, W89ju6);  // ../RTL/cortexm0ds_logic.v(14712)
  not u17605 (Ryzow6, n4926);  // ../RTL/cortexm0ds_logic.v(14712)
  and u17606 (n4927, Fzzow6, Mzzow6);  // ../RTL/cortexm0ds_logic.v(14713)
  not u17607 (W89ju6, n4927);  // ../RTL/cortexm0ds_logic.v(14713)
  and u17608 (Mzzow6, Tzzow6, A00pw6);  // ../RTL/cortexm0ds_logic.v(14714)
  and u17609 (A00pw6, H00pw6, O00pw6);  // ../RTL/cortexm0ds_logic.v(14715)
  and u1761 (Kp1iu6, Gu1iu6, Nu1iu6);  // ../RTL/cortexm0ds_logic.v(3677)
  and u17610 (n4928, Fkfpw6[15], Dfqow6);  // ../RTL/cortexm0ds_logic.v(14716)
  not u17611 (O00pw6, n4928);  // ../RTL/cortexm0ds_logic.v(14716)
  and u17612 (H00pw6, V00pw6, C10pw6);  // ../RTL/cortexm0ds_logic.v(14717)
  and u17613 (n4929, vis_psp_o[13], Yfqow6);  // ../RTL/cortexm0ds_logic.v(14718)
  not u17614 (C10pw6, n4929);  // ../RTL/cortexm0ds_logic.v(14718)
  and u17615 (n4930, vis_msp_o[13], Fgqow6);  // ../RTL/cortexm0ds_logic.v(14719)
  not u17616 (V00pw6, n4930);  // ../RTL/cortexm0ds_logic.v(14719)
  and u17617 (Tzzow6, J10pw6, Q10pw6);  // ../RTL/cortexm0ds_logic.v(14720)
  and u17618 (n4931, vis_r14_o[15], Ahqow6);  // ../RTL/cortexm0ds_logic.v(14721)
  not u17619 (Q10pw6, n4931);  // ../RTL/cortexm0ds_logic.v(14721)
  and u1762 (Nu1iu6, Uu1iu6, Bv1iu6);  // ../RTL/cortexm0ds_logic.v(3678)
  and u17620 (n4932, vis_r12_o[15], Hhqow6);  // ../RTL/cortexm0ds_logic.v(14722)
  not u17621 (J10pw6, n4932);  // ../RTL/cortexm0ds_logic.v(14722)
  and u17622 (Fzzow6, X10pw6, E20pw6);  // ../RTL/cortexm0ds_logic.v(14723)
  and u17623 (E20pw6, L20pw6, S20pw6);  // ../RTL/cortexm0ds_logic.v(14724)
  and u17624 (n4933, vis_r9_o[15], Qiqow6);  // ../RTL/cortexm0ds_logic.v(14725)
  not u17625 (S20pw6, n4933);  // ../RTL/cortexm0ds_logic.v(14725)
  and u17626 (L20pw6, Z20pw6, G30pw6);  // ../RTL/cortexm0ds_logic.v(14726)
  and u17627 (n4934, vis_r11_o[15], Ljqow6);  // ../RTL/cortexm0ds_logic.v(14727)
  not u17628 (G30pw6, n4934);  // ../RTL/cortexm0ds_logic.v(14727)
  and u17629 (n4935, vis_r10_o[15], Sjqow6);  // ../RTL/cortexm0ds_logic.v(14728)
  and u1763 (n147, Iv1iu6, vis_pc_o[30]);  // ../RTL/cortexm0ds_logic.v(3679)
  not u17630 (Z20pw6, n4935);  // ../RTL/cortexm0ds_logic.v(14728)
  and u17631 (X10pw6, X10iu6, N30pw6);  // ../RTL/cortexm0ds_logic.v(14729)
  and u17632 (n4936, vis_r8_o[15], Gkqow6);  // ../RTL/cortexm0ds_logic.v(14730)
  not u17633 (N30pw6, n4936);  // ../RTL/cortexm0ds_logic.v(14730)
  and u17634 (X10iu6, U30pw6, B40pw6);  // ../RTL/cortexm0ds_logic.v(14731)
  and u17635 (B40pw6, I40pw6, P40pw6);  // ../RTL/cortexm0ds_logic.v(14732)
  and u17636 (P40pw6, W40pw6, D50pw6);  // ../RTL/cortexm0ds_logic.v(14733)
  and u17637 (n4937, vis_r2_o[15], Dmqow6);  // ../RTL/cortexm0ds_logic.v(14734)
  not u17638 (D50pw6, n4937);  // ../RTL/cortexm0ds_logic.v(14734)
  and u17639 (n4938, vis_r6_o[15], Kmqow6);  // ../RTL/cortexm0ds_logic.v(14735)
  not u1764 (Bv1iu6, n147);  // ../RTL/cortexm0ds_logic.v(3679)
  not u17640 (W40pw6, n4938);  // ../RTL/cortexm0ds_logic.v(14735)
  and u17641 (I40pw6, K50pw6, R50pw6);  // ../RTL/cortexm0ds_logic.v(14736)
  and u17642 (n4939, vis_r5_o[15], Fnqow6);  // ../RTL/cortexm0ds_logic.v(14737)
  not u17643 (R50pw6, n4939);  // ../RTL/cortexm0ds_logic.v(14737)
  and u17644 (n4940, vis_r4_o[15], Mnqow6);  // ../RTL/cortexm0ds_logic.v(14738)
  not u17645 (K50pw6, n4940);  // ../RTL/cortexm0ds_logic.v(14738)
  and u17646 (U30pw6, Y50pw6, F60pw6);  // ../RTL/cortexm0ds_logic.v(14739)
  and u17647 (F60pw6, M60pw6, T60pw6);  // ../RTL/cortexm0ds_logic.v(14740)
  and u17648 (n4941, vis_r1_o[15], Voqow6);  // ../RTL/cortexm0ds_logic.v(14741)
  not u17649 (T60pw6, n4941);  // ../RTL/cortexm0ds_logic.v(14741)
  and u1765 (Uu1iu6, Pv1iu6, Wv1iu6);  // ../RTL/cortexm0ds_logic.v(3680)
  and u17650 (n4942, vis_r0_o[15], Cpqow6);  // ../RTL/cortexm0ds_logic.v(14742)
  not u17651 (M60pw6, n4942);  // ../RTL/cortexm0ds_logic.v(14742)
  and u17652 (Y50pw6, A70pw6, H70pw6);  // ../RTL/cortexm0ds_logic.v(14743)
  and u17653 (n4943, vis_r3_o[15], Xpqow6);  // ../RTL/cortexm0ds_logic.v(14744)
  not u17654 (H70pw6, n4943);  // ../RTL/cortexm0ds_logic.v(14744)
  and u17655 (n4944, vis_r7_o[15], Eqqow6);  // ../RTL/cortexm0ds_logic.v(14745)
  not u17656 (A70pw6, n4944);  // ../RTL/cortexm0ds_logic.v(14745)
  and u17657 (Kyzow6, O70pw6, Oqvow6);  // ../RTL/cortexm0ds_logic.v(14746)
  and u17658 (n4945, Udxow6, Uo6ju6);  // ../RTL/cortexm0ds_logic.v(14747)
  not u17659 (Oqvow6, n4945);  // ../RTL/cortexm0ds_logic.v(14747)
  and u1766 (n148, Plgpw6[28], Dw1iu6);  // ../RTL/cortexm0ds_logic.v(3681)
  and u17660 (n4946, V70pw6, C80pw6);  // ../RTL/cortexm0ds_logic.v(14748)
  not u17661 (Uo6ju6, n4946);  // ../RTL/cortexm0ds_logic.v(14748)
  and u17662 (C80pw6, J80pw6, Q80pw6);  // ../RTL/cortexm0ds_logic.v(14749)
  and u17663 (Q80pw6, X80pw6, E90pw6);  // ../RTL/cortexm0ds_logic.v(14750)
  and u17664 (n4947, Fkfpw6[7], Dfqow6);  // ../RTL/cortexm0ds_logic.v(14751)
  not u17665 (E90pw6, n4947);  // ../RTL/cortexm0ds_logic.v(14751)
  and u17666 (X80pw6, L90pw6, S90pw6);  // ../RTL/cortexm0ds_logic.v(14752)
  and u17667 (n4948, vis_psp_o[5], Yfqow6);  // ../RTL/cortexm0ds_logic.v(14753)
  not u17668 (S90pw6, n4948);  // ../RTL/cortexm0ds_logic.v(14753)
  and u17669 (n4949, vis_msp_o[5], Fgqow6);  // ../RTL/cortexm0ds_logic.v(14754)
  not u1767 (Wv1iu6, n148);  // ../RTL/cortexm0ds_logic.v(3681)
  not u17670 (L90pw6, n4949);  // ../RTL/cortexm0ds_logic.v(14754)
  and u17671 (J80pw6, Z90pw6, Ga0pw6);  // ../RTL/cortexm0ds_logic.v(14755)
  and u17672 (n4950, vis_r14_o[7], Ahqow6);  // ../RTL/cortexm0ds_logic.v(14756)
  not u17673 (Ga0pw6, n4950);  // ../RTL/cortexm0ds_logic.v(14756)
  and u17674 (n4951, vis_r12_o[7], Hhqow6);  // ../RTL/cortexm0ds_logic.v(14757)
  not u17675 (Z90pw6, n4951);  // ../RTL/cortexm0ds_logic.v(14757)
  and u17676 (V70pw6, Na0pw6, Ua0pw6);  // ../RTL/cortexm0ds_logic.v(14758)
  and u17677 (Ua0pw6, Bb0pw6, Ib0pw6);  // ../RTL/cortexm0ds_logic.v(14759)
  and u17678 (n4952, vis_r9_o[7], Qiqow6);  // ../RTL/cortexm0ds_logic.v(14760)
  not u17679 (Ib0pw6, n4952);  // ../RTL/cortexm0ds_logic.v(14760)
  and u1768 (n149, K7hpw6[31], Kw1iu6);  // ../RTL/cortexm0ds_logic.v(3682)
  and u17680 (Bb0pw6, Pb0pw6, Wb0pw6);  // ../RTL/cortexm0ds_logic.v(14761)
  and u17681 (n4953, vis_r11_o[7], Ljqow6);  // ../RTL/cortexm0ds_logic.v(14762)
  not u17682 (Wb0pw6, n4953);  // ../RTL/cortexm0ds_logic.v(14762)
  and u17683 (n4954, vis_r10_o[7], Sjqow6);  // ../RTL/cortexm0ds_logic.v(14763)
  not u17684 (Pb0pw6, n4954);  // ../RTL/cortexm0ds_logic.v(14763)
  and u17685 (Na0pw6, Svzhu6, Dc0pw6);  // ../RTL/cortexm0ds_logic.v(14764)
  and u17686 (n4955, vis_r8_o[7], Gkqow6);  // ../RTL/cortexm0ds_logic.v(14765)
  not u17687 (Dc0pw6, n4955);  // ../RTL/cortexm0ds_logic.v(14765)
  and u17688 (Svzhu6, Kc0pw6, Rc0pw6);  // ../RTL/cortexm0ds_logic.v(14766)
  and u17689 (Rc0pw6, Yc0pw6, Fd0pw6);  // ../RTL/cortexm0ds_logic.v(14767)
  not u1769 (Pv1iu6, n149);  // ../RTL/cortexm0ds_logic.v(3682)
  and u17690 (Fd0pw6, Md0pw6, Td0pw6);  // ../RTL/cortexm0ds_logic.v(14768)
  and u17691 (n4956, vis_r0_o[7], Cpqow6);  // ../RTL/cortexm0ds_logic.v(14769)
  not u17692 (Td0pw6, n4956);  // ../RTL/cortexm0ds_logic.v(14769)
  and u17693 (n4957, vis_r2_o[7], Dmqow6);  // ../RTL/cortexm0ds_logic.v(14770)
  not u17694 (Md0pw6, n4957);  // ../RTL/cortexm0ds_logic.v(14770)
  and u17695 (Yc0pw6, Ae0pw6, He0pw6);  // ../RTL/cortexm0ds_logic.v(14771)
  and u17696 (n4958, vis_r5_o[7], Fnqow6);  // ../RTL/cortexm0ds_logic.v(14772)
  not u17697 (He0pw6, n4958);  // ../RTL/cortexm0ds_logic.v(14772)
  and u17698 (n4959, vis_r4_o[7], Mnqow6);  // ../RTL/cortexm0ds_logic.v(14773)
  not u17699 (Ae0pw6, n4959);  // ../RTL/cortexm0ds_logic.v(14773)
  buf u177 (vis_r8_o[10], Ocsax6);  // ../RTL/cortexm0ds_logic.v(2579)
  and u1770 (Gu1iu6, Rw1iu6, Yw1iu6);  // ../RTL/cortexm0ds_logic.v(3683)
  and u17700 (Kc0pw6, Oe0pw6, Ve0pw6);  // ../RTL/cortexm0ds_logic.v(14774)
  and u17701 (Ve0pw6, Cf0pw6, Jf0pw6);  // ../RTL/cortexm0ds_logic.v(14775)
  and u17702 (n4960, vis_r7_o[7], Eqqow6);  // ../RTL/cortexm0ds_logic.v(14776)
  not u17703 (Jf0pw6, n4960);  // ../RTL/cortexm0ds_logic.v(14776)
  and u17704 (n4961, vis_r3_o[7], Xpqow6);  // ../RTL/cortexm0ds_logic.v(14777)
  not u17705 (Cf0pw6, n4961);  // ../RTL/cortexm0ds_logic.v(14777)
  and u17706 (Oe0pw6, Qf0pw6, Xf0pw6);  // ../RTL/cortexm0ds_logic.v(14778)
  and u17707 (n4962, vis_r1_o[7], Voqow6);  // ../RTL/cortexm0ds_logic.v(14779)
  not u17708 (Xf0pw6, n4962);  // ../RTL/cortexm0ds_logic.v(14779)
  and u17709 (n4963, vis_r6_o[7], Kmqow6);  // ../RTL/cortexm0ds_logic.v(14780)
  and u1771 (Zm1iu6, Fx1iu6, Mx1iu6);  // ../RTL/cortexm0ds_logic.v(3684)
  not u17710 (Qf0pw6, n4963);  // ../RTL/cortexm0ds_logic.v(14780)
  and u17711 (n4964, S54iu6, R0nhu6);  // ../RTL/cortexm0ds_logic.v(14781)
  not u17712 (O70pw6, n4964);  // ../RTL/cortexm0ds_logic.v(14781)
  and u17713 (S54iu6, Shhpw6[15], Iqzhu6);  // ../RTL/cortexm0ds_logic.v(14782)
  and u17714 (n4965, Yyzow6, T39ju6);  // ../RTL/cortexm0ds_logic.v(14784)
  not u17715 (Lg0pw6, n4965);  // ../RTL/cortexm0ds_logic.v(14784)
  and u17716 (n4966, Sg0pw6, Zg0pw6);  // ../RTL/cortexm0ds_logic.v(14785)
  not u17717 (T39ju6, n4966);  // ../RTL/cortexm0ds_logic.v(14785)
  and u17718 (Zg0pw6, Gh0pw6, Nh0pw6);  // ../RTL/cortexm0ds_logic.v(14786)
  and u17719 (Nh0pw6, Uh0pw6, Bi0pw6);  // ../RTL/cortexm0ds_logic.v(14787)
  and u1772 (n150, ECOREVNUM[23], Tx1iu6);  // ../RTL/cortexm0ds_logic.v(3685)
  and u17720 (n4967, vis_r11_o[14], Ljqow6);  // ../RTL/cortexm0ds_logic.v(14788)
  not u17721 (Bi0pw6, n4967);  // ../RTL/cortexm0ds_logic.v(14788)
  and u17722 (Uh0pw6, Ii0pw6, Pi0pw6);  // ../RTL/cortexm0ds_logic.v(14789)
  and u17723 (n4968, vis_r9_o[14], Qiqow6);  // ../RTL/cortexm0ds_logic.v(14790)
  not u17724 (Pi0pw6, n4968);  // ../RTL/cortexm0ds_logic.v(14790)
  and u17725 (n4969, Fkfpw6[14], Dfqow6);  // ../RTL/cortexm0ds_logic.v(14791)
  not u17726 (Ii0pw6, n4969);  // ../RTL/cortexm0ds_logic.v(14791)
  and u17727 (Gh0pw6, Wi0pw6, Dj0pw6);  // ../RTL/cortexm0ds_logic.v(14792)
  and u17728 (n4970, vis_r10_o[14], Sjqow6);  // ../RTL/cortexm0ds_logic.v(14793)
  not u17729 (Dj0pw6, n4970);  // ../RTL/cortexm0ds_logic.v(14793)
  not u1773 (Mx1iu6, n150);  // ../RTL/cortexm0ds_logic.v(3685)
  and u17730 (n4971, vis_psp_o[12], Yfqow6);  // ../RTL/cortexm0ds_logic.v(14794)
  not u17731 (Wi0pw6, n4971);  // ../RTL/cortexm0ds_logic.v(14794)
  and u17732 (Sg0pw6, Kj0pw6, Rj0pw6);  // ../RTL/cortexm0ds_logic.v(14795)
  and u17733 (Rj0pw6, Yj0pw6, Fk0pw6);  // ../RTL/cortexm0ds_logic.v(14796)
  and u17734 (n4972, vis_r12_o[14], Hhqow6);  // ../RTL/cortexm0ds_logic.v(14797)
  not u17735 (Fk0pw6, n4972);  // ../RTL/cortexm0ds_logic.v(14797)
  and u17736 (Yj0pw6, Mk0pw6, Tk0pw6);  // ../RTL/cortexm0ds_logic.v(14798)
  and u17737 (n4973, vis_msp_o[12], Fgqow6);  // ../RTL/cortexm0ds_logic.v(14799)
  not u17738 (Tk0pw6, n4973);  // ../RTL/cortexm0ds_logic.v(14799)
  and u17739 (n4974, vis_r14_o[14], Ahqow6);  // ../RTL/cortexm0ds_logic.v(14800)
  and u1774 (n151, Uthpw6[31], Sf1iu6);  // ../RTL/cortexm0ds_logic.v(3686)
  not u17740 (Mk0pw6, n4974);  // ../RTL/cortexm0ds_logic.v(14800)
  and u17741 (Kj0pw6, E20iu6, Al0pw6);  // ../RTL/cortexm0ds_logic.v(14801)
  and u17742 (n4975, vis_r8_o[14], Gkqow6);  // ../RTL/cortexm0ds_logic.v(14802)
  not u17743 (Al0pw6, n4975);  // ../RTL/cortexm0ds_logic.v(14802)
  and u17744 (E20iu6, Hl0pw6, Ol0pw6);  // ../RTL/cortexm0ds_logic.v(14803)
  and u17745 (Ol0pw6, Vl0pw6, Cm0pw6);  // ../RTL/cortexm0ds_logic.v(14804)
  and u17746 (Cm0pw6, Jm0pw6, Qm0pw6);  // ../RTL/cortexm0ds_logic.v(14805)
  and u17747 (n4976, vis_r2_o[14], Dmqow6);  // ../RTL/cortexm0ds_logic.v(14806)
  not u17748 (Qm0pw6, n4976);  // ../RTL/cortexm0ds_logic.v(14806)
  and u17749 (n4977, vis_r6_o[14], Kmqow6);  // ../RTL/cortexm0ds_logic.v(14807)
  not u1775 (Fx1iu6, n151);  // ../RTL/cortexm0ds_logic.v(3686)
  not u17750 (Jm0pw6, n4977);  // ../RTL/cortexm0ds_logic.v(14807)
  and u17751 (Vl0pw6, Xm0pw6, En0pw6);  // ../RTL/cortexm0ds_logic.v(14808)
  and u17752 (n4978, vis_r5_o[14], Fnqow6);  // ../RTL/cortexm0ds_logic.v(14809)
  not u17753 (En0pw6, n4978);  // ../RTL/cortexm0ds_logic.v(14809)
  and u17754 (n4979, vis_r4_o[14], Mnqow6);  // ../RTL/cortexm0ds_logic.v(14810)
  not u17755 (Xm0pw6, n4979);  // ../RTL/cortexm0ds_logic.v(14810)
  and u17756 (Hl0pw6, Ln0pw6, Sn0pw6);  // ../RTL/cortexm0ds_logic.v(14811)
  and u17757 (Sn0pw6, Zn0pw6, Go0pw6);  // ../RTL/cortexm0ds_logic.v(14812)
  and u17758 (n4980, vis_r1_o[14], Voqow6);  // ../RTL/cortexm0ds_logic.v(14813)
  not u17759 (Go0pw6, n4980);  // ../RTL/cortexm0ds_logic.v(14813)
  and u1776 (n152, Ay1iu6, Hy1iu6);  // ../RTL/cortexm0ds_logic.v(3687)
  and u17760 (n4981, vis_r0_o[14], Cpqow6);  // ../RTL/cortexm0ds_logic.v(14814)
  not u17761 (Zn0pw6, n4981);  // ../RTL/cortexm0ds_logic.v(14814)
  and u17762 (Ln0pw6, No0pw6, Uo0pw6);  // ../RTL/cortexm0ds_logic.v(14815)
  and u17763 (n4982, vis_r3_o[14], Xpqow6);  // ../RTL/cortexm0ds_logic.v(14816)
  not u17764 (Uo0pw6, n4982);  // ../RTL/cortexm0ds_logic.v(14816)
  and u17765 (n4983, vis_r7_o[14], Eqqow6);  // ../RTL/cortexm0ds_logic.v(14817)
  not u17766 (No0pw6, n4983);  // ../RTL/cortexm0ds_logic.v(14817)
  and u17767 (Eg0pw6, Bp0pw6, N0wow6);  // ../RTL/cortexm0ds_logic.v(14818)
  and u17768 (n4984, Udxow6, Kj6ju6);  // ../RTL/cortexm0ds_logic.v(14819)
  not u17769 (N0wow6, n4984);  // ../RTL/cortexm0ds_logic.v(14819)
  not u1777 (A2yhu6, n152);  // ../RTL/cortexm0ds_logic.v(3687)
  and u17770 (n4985, Ip0pw6, Pp0pw6);  // ../RTL/cortexm0ds_logic.v(14820)
  not u17771 (Kj6ju6, n4985);  // ../RTL/cortexm0ds_logic.v(14820)
  and u17772 (Pp0pw6, Wp0pw6, Dq0pw6);  // ../RTL/cortexm0ds_logic.v(14821)
  and u17773 (Dq0pw6, Kq0pw6, Rq0pw6);  // ../RTL/cortexm0ds_logic.v(14822)
  and u17774 (n4986, Fkfpw6[6], Dfqow6);  // ../RTL/cortexm0ds_logic.v(14823)
  not u17775 (Rq0pw6, n4986);  // ../RTL/cortexm0ds_logic.v(14823)
  and u17776 (Kq0pw6, Yq0pw6, Fr0pw6);  // ../RTL/cortexm0ds_logic.v(14824)
  and u17777 (n4987, vis_psp_o[4], Yfqow6);  // ../RTL/cortexm0ds_logic.v(14825)
  not u17778 (Fr0pw6, n4987);  // ../RTL/cortexm0ds_logic.v(14825)
  and u17779 (n4988, vis_msp_o[4], Fgqow6);  // ../RTL/cortexm0ds_logic.v(14826)
  and u1778 (Hy1iu6, Oy1iu6, Vy1iu6);  // ../RTL/cortexm0ds_logic.v(3688)
  not u17780 (Yq0pw6, n4988);  // ../RTL/cortexm0ds_logic.v(14826)
  and u17781 (Wp0pw6, Mr0pw6, Tr0pw6);  // ../RTL/cortexm0ds_logic.v(14827)
  and u17782 (n4989, vis_r14_o[6], Ahqow6);  // ../RTL/cortexm0ds_logic.v(14828)
  not u17783 (Tr0pw6, n4989);  // ../RTL/cortexm0ds_logic.v(14828)
  and u17784 (n4990, vis_r12_o[6], Hhqow6);  // ../RTL/cortexm0ds_logic.v(14829)
  not u17785 (Mr0pw6, n4990);  // ../RTL/cortexm0ds_logic.v(14829)
  and u17786 (Ip0pw6, As0pw6, Hs0pw6);  // ../RTL/cortexm0ds_logic.v(14830)
  and u17787 (Hs0pw6, Os0pw6, Vs0pw6);  // ../RTL/cortexm0ds_logic.v(14831)
  and u17788 (n4991, vis_r9_o[6], Qiqow6);  // ../RTL/cortexm0ds_logic.v(14832)
  not u17789 (Vs0pw6, n4991);  // ../RTL/cortexm0ds_logic.v(14832)
  and u1779 (Oy1iu6, Cz1iu6, Jz1iu6);  // ../RTL/cortexm0ds_logic.v(3689)
  and u17790 (Os0pw6, Ct0pw6, Jt0pw6);  // ../RTL/cortexm0ds_logic.v(14833)
  and u17791 (n4992, vis_r11_o[6], Ljqow6);  // ../RTL/cortexm0ds_logic.v(14834)
  not u17792 (Jt0pw6, n4992);  // ../RTL/cortexm0ds_logic.v(14834)
  and u17793 (n4993, vis_r10_o[6], Sjqow6);  // ../RTL/cortexm0ds_logic.v(14835)
  not u17794 (Ct0pw6, n4993);  // ../RTL/cortexm0ds_logic.v(14835)
  and u17795 (As0pw6, Zvzhu6, Qt0pw6);  // ../RTL/cortexm0ds_logic.v(14836)
  and u17796 (n4994, vis_r8_o[6], Gkqow6);  // ../RTL/cortexm0ds_logic.v(14837)
  not u17797 (Qt0pw6, n4994);  // ../RTL/cortexm0ds_logic.v(14837)
  and u17798 (Zvzhu6, Xt0pw6, Eu0pw6);  // ../RTL/cortexm0ds_logic.v(14838)
  and u17799 (Eu0pw6, Lu0pw6, Su0pw6);  // ../RTL/cortexm0ds_logic.v(14839)
  buf u178 (Uthpw6[1], L9bbx6);  // ../RTL/cortexm0ds_logic.v(1882)
  and u1780 (n153, Uthpw6[31], Vk1iu6);  // ../RTL/cortexm0ds_logic.v(3690)
  and u17800 (Su0pw6, Zu0pw6, Gv0pw6);  // ../RTL/cortexm0ds_logic.v(14840)
  and u17801 (n4995, vis_r0_o[6], Cpqow6);  // ../RTL/cortexm0ds_logic.v(14841)
  not u17802 (Gv0pw6, n4995);  // ../RTL/cortexm0ds_logic.v(14841)
  and u17803 (n4996, vis_r2_o[6], Dmqow6);  // ../RTL/cortexm0ds_logic.v(14842)
  not u17804 (Zu0pw6, n4996);  // ../RTL/cortexm0ds_logic.v(14842)
  and u17805 (Lu0pw6, Nv0pw6, Uv0pw6);  // ../RTL/cortexm0ds_logic.v(14843)
  and u17806 (n4997, vis_r5_o[6], Fnqow6);  // ../RTL/cortexm0ds_logic.v(14844)
  not u17807 (Uv0pw6, n4997);  // ../RTL/cortexm0ds_logic.v(14844)
  and u17808 (n4998, vis_r4_o[6], Mnqow6);  // ../RTL/cortexm0ds_logic.v(14845)
  not u17809 (Nv0pw6, n4998);  // ../RTL/cortexm0ds_logic.v(14845)
  not u1781 (Jz1iu6, n153);  // ../RTL/cortexm0ds_logic.v(3690)
  and u17810 (Xt0pw6, Bw0pw6, Iw0pw6);  // ../RTL/cortexm0ds_logic.v(14846)
  and u17811 (Iw0pw6, Pw0pw6, Ww0pw6);  // ../RTL/cortexm0ds_logic.v(14847)
  and u17812 (n4999, vis_r7_o[6], Eqqow6);  // ../RTL/cortexm0ds_logic.v(14848)
  not u17813 (Ww0pw6, n4999);  // ../RTL/cortexm0ds_logic.v(14848)
  and u17814 (n5000, vis_r3_o[6], Xpqow6);  // ../RTL/cortexm0ds_logic.v(14849)
  not u17815 (Pw0pw6, n5000);  // ../RTL/cortexm0ds_logic.v(14849)
  and u17816 (Bw0pw6, Dx0pw6, Kx0pw6);  // ../RTL/cortexm0ds_logic.v(14850)
  and u17817 (n5001, vis_r1_o[6], Voqow6);  // ../RTL/cortexm0ds_logic.v(14851)
  not u17818 (Kx0pw6, n5001);  // ../RTL/cortexm0ds_logic.v(14851)
  and u17819 (n5002, vis_r6_o[6], Kmqow6);  // ../RTL/cortexm0ds_logic.v(14852)
  and u1782 (n154, ECOREVNUM[27], Qz1iu6);  // ../RTL/cortexm0ds_logic.v(3691)
  not u17820 (Dx0pw6, n5002);  // ../RTL/cortexm0ds_logic.v(14852)
  and u17821 (n5003, L54iu6, R0nhu6);  // ../RTL/cortexm0ds_logic.v(14853)
  not u17822 (Bp0pw6, n5003);  // ../RTL/cortexm0ds_logic.v(14853)
  and u17823 (L54iu6, Shhpw6[14], Iqzhu6);  // ../RTL/cortexm0ds_logic.v(14854)
  and u17824 (n5004, Yyzow6, Sz8ju6);  // ../RTL/cortexm0ds_logic.v(14856)
  not u17825 (Yx0pw6, n5004);  // ../RTL/cortexm0ds_logic.v(14856)
  and u17826 (n5005, Fy0pw6, My0pw6);  // ../RTL/cortexm0ds_logic.v(14857)
  not u17827 (Sz8ju6, n5005);  // ../RTL/cortexm0ds_logic.v(14857)
  and u17828 (My0pw6, Ty0pw6, Az0pw6);  // ../RTL/cortexm0ds_logic.v(14858)
  and u17829 (Az0pw6, Hz0pw6, Oz0pw6);  // ../RTL/cortexm0ds_logic.v(14859)
  not u1783 (Cz1iu6, n154);  // ../RTL/cortexm0ds_logic.v(3691)
  and u17830 (n5006, Fkfpw6[13], Dfqow6);  // ../RTL/cortexm0ds_logic.v(14860)
  not u17831 (Oz0pw6, n5006);  // ../RTL/cortexm0ds_logic.v(14860)
  and u17832 (Hz0pw6, Vz0pw6, C01pw6);  // ../RTL/cortexm0ds_logic.v(14861)
  and u17833 (n5007, vis_psp_o[11], Yfqow6);  // ../RTL/cortexm0ds_logic.v(14862)
  not u17834 (C01pw6, n5007);  // ../RTL/cortexm0ds_logic.v(14862)
  and u17835 (n5008, vis_msp_o[11], Fgqow6);  // ../RTL/cortexm0ds_logic.v(14863)
  not u17836 (Vz0pw6, n5008);  // ../RTL/cortexm0ds_logic.v(14863)
  and u17837 (Ty0pw6, J01pw6, Q01pw6);  // ../RTL/cortexm0ds_logic.v(14864)
  and u17838 (n5009, vis_r14_o[13], Ahqow6);  // ../RTL/cortexm0ds_logic.v(14865)
  not u17839 (Q01pw6, n5009);  // ../RTL/cortexm0ds_logic.v(14865)
  and u1784 (Ay1iu6, Xz1iu6, E02iu6);  // ../RTL/cortexm0ds_logic.v(3692)
  and u17840 (n5010, vis_r12_o[13], Hhqow6);  // ../RTL/cortexm0ds_logic.v(14866)
  not u17841 (J01pw6, n5010);  // ../RTL/cortexm0ds_logic.v(14866)
  and u17842 (Fy0pw6, X01pw6, E11pw6);  // ../RTL/cortexm0ds_logic.v(14867)
  and u17843 (E11pw6, L11pw6, S11pw6);  // ../RTL/cortexm0ds_logic.v(14868)
  and u17844 (n5011, vis_r9_o[13], Qiqow6);  // ../RTL/cortexm0ds_logic.v(14869)
  not u17845 (S11pw6, n5011);  // ../RTL/cortexm0ds_logic.v(14869)
  and u17846 (L11pw6, Z11pw6, G21pw6);  // ../RTL/cortexm0ds_logic.v(14870)
  and u17847 (n5012, vis_r11_o[13], Ljqow6);  // ../RTL/cortexm0ds_logic.v(14871)
  not u17848 (G21pw6, n5012);  // ../RTL/cortexm0ds_logic.v(14871)
  and u17849 (n5013, vis_r10_o[13], Sjqow6);  // ../RTL/cortexm0ds_logic.v(14872)
  and u1785 (n155, Iahpw6[30], Xl1iu6);  // ../RTL/cortexm0ds_logic.v(3693)
  not u17850 (Z11pw6, n5013);  // ../RTL/cortexm0ds_logic.v(14872)
  and u17851 (X01pw6, L20iu6, N21pw6);  // ../RTL/cortexm0ds_logic.v(14873)
  and u17852 (n5014, vis_r8_o[13], Gkqow6);  // ../RTL/cortexm0ds_logic.v(14874)
  not u17853 (N21pw6, n5014);  // ../RTL/cortexm0ds_logic.v(14874)
  and u17854 (L20iu6, U21pw6, B31pw6);  // ../RTL/cortexm0ds_logic.v(14875)
  and u17855 (B31pw6, I31pw6, P31pw6);  // ../RTL/cortexm0ds_logic.v(14876)
  and u17856 (P31pw6, W31pw6, D41pw6);  // ../RTL/cortexm0ds_logic.v(14877)
  and u17857 (n5015, vis_r2_o[13], Dmqow6);  // ../RTL/cortexm0ds_logic.v(14878)
  not u17858 (D41pw6, n5015);  // ../RTL/cortexm0ds_logic.v(14878)
  and u17859 (n5016, vis_r6_o[13], Kmqow6);  // ../RTL/cortexm0ds_logic.v(14879)
  not u1786 (E02iu6, n155);  // ../RTL/cortexm0ds_logic.v(3693)
  not u17860 (W31pw6, n5016);  // ../RTL/cortexm0ds_logic.v(14879)
  and u17861 (I31pw6, K41pw6, R41pw6);  // ../RTL/cortexm0ds_logic.v(14880)
  and u17862 (n5017, vis_r5_o[13], Fnqow6);  // ../RTL/cortexm0ds_logic.v(14881)
  not u17863 (R41pw6, n5017);  // ../RTL/cortexm0ds_logic.v(14881)
  and u17864 (n5018, vis_r4_o[13], Mnqow6);  // ../RTL/cortexm0ds_logic.v(14882)
  not u17865 (K41pw6, n5018);  // ../RTL/cortexm0ds_logic.v(14882)
  and u17866 (U21pw6, Y41pw6, F51pw6);  // ../RTL/cortexm0ds_logic.v(14883)
  and u17867 (F51pw6, M51pw6, T51pw6);  // ../RTL/cortexm0ds_logic.v(14884)
  and u17868 (n5019, vis_r1_o[13], Voqow6);  // ../RTL/cortexm0ds_logic.v(14885)
  not u17869 (T51pw6, n5019);  // ../RTL/cortexm0ds_logic.v(14885)
  or u1787 (Xz1iu6, L02iu6, Jayhu6);  // ../RTL/cortexm0ds_logic.v(3694)
  and u17870 (n5020, vis_r0_o[13], Cpqow6);  // ../RTL/cortexm0ds_logic.v(14886)
  not u17871 (M51pw6, n5020);  // ../RTL/cortexm0ds_logic.v(14886)
  and u17872 (Y41pw6, A61pw6, H61pw6);  // ../RTL/cortexm0ds_logic.v(14887)
  and u17873 (n5021, vis_r3_o[13], Xpqow6);  // ../RTL/cortexm0ds_logic.v(14888)
  not u17874 (H61pw6, n5021);  // ../RTL/cortexm0ds_logic.v(14888)
  and u17875 (n5022, vis_r7_o[13], Eqqow6);  // ../RTL/cortexm0ds_logic.v(14889)
  not u17876 (A61pw6, n5022);  // ../RTL/cortexm0ds_logic.v(14889)
  and u17877 (Rx0pw6, O61pw6, Zqqow6);  // ../RTL/cortexm0ds_logic.v(14890)
  and u17878 (n5023, Udxow6, Eg6ju6);  // ../RTL/cortexm0ds_logic.v(14891)
  not u17879 (Zqqow6, n5023);  // ../RTL/cortexm0ds_logic.v(14891)
  not u1788 (Jayhu6, Mdhpw6[3]);  // ../RTL/cortexm0ds_logic.v(3695)
  and u17880 (n5024, V61pw6, C71pw6);  // ../RTL/cortexm0ds_logic.v(14892)
  not u17881 (Eg6ju6, n5024);  // ../RTL/cortexm0ds_logic.v(14892)
  and u17882 (C71pw6, J71pw6, Q71pw6);  // ../RTL/cortexm0ds_logic.v(14893)
  and u17883 (Q71pw6, X71pw6, E81pw6);  // ../RTL/cortexm0ds_logic.v(14894)
  and u17884 (n5025, Fkfpw6[5], Dfqow6);  // ../RTL/cortexm0ds_logic.v(14895)
  not u17885 (E81pw6, n5025);  // ../RTL/cortexm0ds_logic.v(14895)
  and u17886 (X71pw6, L81pw6, S81pw6);  // ../RTL/cortexm0ds_logic.v(14896)
  and u17887 (n5026, vis_psp_o[3], Yfqow6);  // ../RTL/cortexm0ds_logic.v(14897)
  not u17888 (S81pw6, n5026);  // ../RTL/cortexm0ds_logic.v(14897)
  and u17889 (n5027, vis_msp_o[3], Fgqow6);  // ../RTL/cortexm0ds_logic.v(14898)
  and u1789 (n156, S02iu6, Z02iu6);  // ../RTL/cortexm0ds_logic.v(3696)
  not u17890 (L81pw6, n5027);  // ../RTL/cortexm0ds_logic.v(14898)
  and u17891 (J71pw6, Z81pw6, G91pw6);  // ../RTL/cortexm0ds_logic.v(14899)
  and u17892 (n5028, vis_r14_o[5], Ahqow6);  // ../RTL/cortexm0ds_logic.v(14900)
  not u17893 (G91pw6, n5028);  // ../RTL/cortexm0ds_logic.v(14900)
  and u17894 (n5029, vis_r12_o[5], Hhqow6);  // ../RTL/cortexm0ds_logic.v(14901)
  not u17895 (Z81pw6, n5029);  // ../RTL/cortexm0ds_logic.v(14901)
  and u17896 (V61pw6, N91pw6, U91pw6);  // ../RTL/cortexm0ds_logic.v(14902)
  and u17897 (U91pw6, Ba1pw6, Ia1pw6);  // ../RTL/cortexm0ds_logic.v(14903)
  and u17898 (n5030, vis_r9_o[5], Qiqow6);  // ../RTL/cortexm0ds_logic.v(14904)
  not u17899 (Ia1pw6, n5030);  // ../RTL/cortexm0ds_logic.v(14904)
  buf u179 (vis_r12_o[24], F2tax6);  // ../RTL/cortexm0ds_logic.v(2599)
  not u1790 (T1yhu6, n156);  // ../RTL/cortexm0ds_logic.v(3696)
  and u17900 (Ba1pw6, Pa1pw6, Wa1pw6);  // ../RTL/cortexm0ds_logic.v(14905)
  and u17901 (n5031, vis_r11_o[5], Ljqow6);  // ../RTL/cortexm0ds_logic.v(14906)
  not u17902 (Wa1pw6, n5031);  // ../RTL/cortexm0ds_logic.v(14906)
  and u17903 (n5032, vis_r10_o[5], Sjqow6);  // ../RTL/cortexm0ds_logic.v(14907)
  not u17904 (Pa1pw6, n5032);  // ../RTL/cortexm0ds_logic.v(14907)
  and u17905 (N91pw6, Gwzhu6, Db1pw6);  // ../RTL/cortexm0ds_logic.v(14908)
  and u17906 (n5033, vis_r8_o[5], Gkqow6);  // ../RTL/cortexm0ds_logic.v(14909)
  not u17907 (Db1pw6, n5033);  // ../RTL/cortexm0ds_logic.v(14909)
  and u17908 (Gwzhu6, Kb1pw6, Rb1pw6);  // ../RTL/cortexm0ds_logic.v(14910)
  and u17909 (Rb1pw6, Yb1pw6, Fc1pw6);  // ../RTL/cortexm0ds_logic.v(14911)
  and u1791 (Z02iu6, G12iu6, Vy1iu6);  // ../RTL/cortexm0ds_logic.v(3697)
  and u17910 (Fc1pw6, Mc1pw6, Tc1pw6);  // ../RTL/cortexm0ds_logic.v(14912)
  and u17911 (n5034, vis_r0_o[5], Cpqow6);  // ../RTL/cortexm0ds_logic.v(14913)
  not u17912 (Tc1pw6, n5034);  // ../RTL/cortexm0ds_logic.v(14913)
  and u17913 (n5035, vis_r2_o[5], Dmqow6);  // ../RTL/cortexm0ds_logic.v(14914)
  not u17914 (Mc1pw6, n5035);  // ../RTL/cortexm0ds_logic.v(14914)
  and u17915 (Yb1pw6, Ad1pw6, Hd1pw6);  // ../RTL/cortexm0ds_logic.v(14915)
  and u17916 (n5036, vis_r5_o[5], Fnqow6);  // ../RTL/cortexm0ds_logic.v(14916)
  not u17917 (Hd1pw6, n5036);  // ../RTL/cortexm0ds_logic.v(14916)
  and u17918 (n5037, vis_r4_o[5], Mnqow6);  // ../RTL/cortexm0ds_logic.v(14917)
  not u17919 (Ad1pw6, n5037);  // ../RTL/cortexm0ds_logic.v(14917)
  and u1792 (n157, Zbhpw6[30], Cl1iu6);  // ../RTL/cortexm0ds_logic.v(3698)
  and u17920 (Kb1pw6, Od1pw6, Vd1pw6);  // ../RTL/cortexm0ds_logic.v(14918)
  and u17921 (Vd1pw6, Ce1pw6, Je1pw6);  // ../RTL/cortexm0ds_logic.v(14919)
  and u17922 (n5038, vis_r7_o[5], Eqqow6);  // ../RTL/cortexm0ds_logic.v(14920)
  not u17923 (Je1pw6, n5038);  // ../RTL/cortexm0ds_logic.v(14920)
  and u17924 (n5039, vis_r3_o[5], Xpqow6);  // ../RTL/cortexm0ds_logic.v(14921)
  not u17925 (Ce1pw6, n5039);  // ../RTL/cortexm0ds_logic.v(14921)
  and u17926 (Od1pw6, Qe1pw6, Xe1pw6);  // ../RTL/cortexm0ds_logic.v(14922)
  and u17927 (n5040, vis_r1_o[5], Voqow6);  // ../RTL/cortexm0ds_logic.v(14923)
  not u17928 (Xe1pw6, n5040);  // ../RTL/cortexm0ds_logic.v(14923)
  and u17929 (n5041, vis_r6_o[5], Kmqow6);  // ../RTL/cortexm0ds_logic.v(14924)
  not u1793 (Vy1iu6, n157);  // ../RTL/cortexm0ds_logic.v(3698)
  not u17930 (Qe1pw6, n5041);  // ../RTL/cortexm0ds_logic.v(14924)
  and u17931 (n5042, E54iu6, R0nhu6);  // ../RTL/cortexm0ds_logic.v(14925)
  not u17932 (O61pw6, n5042);  // ../RTL/cortexm0ds_logic.v(14925)
  and u17933 (E54iu6, Shhpw6[13], Iqzhu6);  // ../RTL/cortexm0ds_logic.v(14926)
  and u17934 (n5043, Yyzow6, Rv8ju6);  // ../RTL/cortexm0ds_logic.v(14928)
  not u17935 (Lf1pw6, n5043);  // ../RTL/cortexm0ds_logic.v(14928)
  and u17936 (n5044, Sf1pw6, Zf1pw6);  // ../RTL/cortexm0ds_logic.v(14929)
  not u17937 (Rv8ju6, n5044);  // ../RTL/cortexm0ds_logic.v(14929)
  and u17938 (Zf1pw6, Gg1pw6, Ng1pw6);  // ../RTL/cortexm0ds_logic.v(14930)
  and u17939 (Ng1pw6, Ug1pw6, Bh1pw6);  // ../RTL/cortexm0ds_logic.v(14931)
  and u1794 (G12iu6, N12iu6, U12iu6);  // ../RTL/cortexm0ds_logic.v(3699)
  and u17940 (n5045, vis_r11_o[12], Ljqow6);  // ../RTL/cortexm0ds_logic.v(14932)
  not u17941 (Bh1pw6, n5045);  // ../RTL/cortexm0ds_logic.v(14932)
  and u17942 (Ug1pw6, Ih1pw6, Ph1pw6);  // ../RTL/cortexm0ds_logic.v(14933)
  and u17943 (n5046, vis_r10_o[12], Sjqow6);  // ../RTL/cortexm0ds_logic.v(14934)
  not u17944 (Ph1pw6, n5046);  // ../RTL/cortexm0ds_logic.v(14934)
  and u17945 (n5047, vis_r9_o[12], Qiqow6);  // ../RTL/cortexm0ds_logic.v(14935)
  not u17946 (Ih1pw6, n5047);  // ../RTL/cortexm0ds_logic.v(14935)
  and u17947 (Gg1pw6, Wh1pw6, Di1pw6);  // ../RTL/cortexm0ds_logic.v(14936)
  and u17948 (n5048, Fkfpw6[12], Dfqow6);  // ../RTL/cortexm0ds_logic.v(14937)
  not u17949 (Di1pw6, n5048);  // ../RTL/cortexm0ds_logic.v(14937)
  and u1795 (n158, Uthpw6[30], Vk1iu6);  // ../RTL/cortexm0ds_logic.v(3700)
  and u17950 (n5049, vis_r12_o[12], Hhqow6);  // ../RTL/cortexm0ds_logic.v(14938)
  not u17951 (Wh1pw6, n5049);  // ../RTL/cortexm0ds_logic.v(14938)
  and u17952 (Sf1pw6, Ki1pw6, Ri1pw6);  // ../RTL/cortexm0ds_logic.v(14939)
  and u17953 (Ri1pw6, Yi1pw6, Fj1pw6);  // ../RTL/cortexm0ds_logic.v(14940)
  and u17954 (n5050, vis_r14_o[12], Ahqow6);  // ../RTL/cortexm0ds_logic.v(14941)
  not u17955 (Fj1pw6, n5050);  // ../RTL/cortexm0ds_logic.v(14941)
  and u17956 (Yi1pw6, Mj1pw6, Tj1pw6);  // ../RTL/cortexm0ds_logic.v(14942)
  and u17957 (n5051, vis_psp_o[10], Yfqow6);  // ../RTL/cortexm0ds_logic.v(14943)
  not u17958 (Tj1pw6, n5051);  // ../RTL/cortexm0ds_logic.v(14943)
  and u17959 (n5052, vis_r8_o[12], Gkqow6);  // ../RTL/cortexm0ds_logic.v(14944)
  not u1796 (U12iu6, n158);  // ../RTL/cortexm0ds_logic.v(3700)
  not u17960 (Mj1pw6, n5052);  // ../RTL/cortexm0ds_logic.v(14944)
  and u17961 (Ki1pw6, S20iu6, Ak1pw6);  // ../RTL/cortexm0ds_logic.v(14945)
  and u17962 (n5053, vis_msp_o[10], Fgqow6);  // ../RTL/cortexm0ds_logic.v(14946)
  not u17963 (Ak1pw6, n5053);  // ../RTL/cortexm0ds_logic.v(14946)
  and u17964 (S20iu6, Hk1pw6, Ok1pw6);  // ../RTL/cortexm0ds_logic.v(14947)
  and u17965 (Ok1pw6, Vk1pw6, Cl1pw6);  // ../RTL/cortexm0ds_logic.v(14948)
  and u17966 (Cl1pw6, Jl1pw6, Ql1pw6);  // ../RTL/cortexm0ds_logic.v(14949)
  and u17967 (n5054, vis_r0_o[12], Cpqow6);  // ../RTL/cortexm0ds_logic.v(14950)
  not u17968 (Ql1pw6, n5054);  // ../RTL/cortexm0ds_logic.v(14950)
  and u17969 (n5055, vis_r2_o[12], Dmqow6);  // ../RTL/cortexm0ds_logic.v(14951)
  and u1797 (n159, ECOREVNUM[26], Qz1iu6);  // ../RTL/cortexm0ds_logic.v(3701)
  not u17970 (Jl1pw6, n5055);  // ../RTL/cortexm0ds_logic.v(14951)
  and u17971 (Vk1pw6, Xl1pw6, Em1pw6);  // ../RTL/cortexm0ds_logic.v(14952)
  and u17972 (n5056, vis_r5_o[12], Fnqow6);  // ../RTL/cortexm0ds_logic.v(14953)
  not u17973 (Em1pw6, n5056);  // ../RTL/cortexm0ds_logic.v(14953)
  and u17974 (n5057, vis_r4_o[12], Mnqow6);  // ../RTL/cortexm0ds_logic.v(14954)
  not u17975 (Xl1pw6, n5057);  // ../RTL/cortexm0ds_logic.v(14954)
  and u17976 (Hk1pw6, Lm1pw6, Sm1pw6);  // ../RTL/cortexm0ds_logic.v(14955)
  and u17977 (Sm1pw6, Zm1pw6, Gn1pw6);  // ../RTL/cortexm0ds_logic.v(14956)
  and u17978 (n5058, vis_r7_o[12], Eqqow6);  // ../RTL/cortexm0ds_logic.v(14957)
  not u17979 (Gn1pw6, n5058);  // ../RTL/cortexm0ds_logic.v(14957)
  not u1798 (N12iu6, n159);  // ../RTL/cortexm0ds_logic.v(3701)
  and u17980 (n5059, vis_r3_o[12], Xpqow6);  // ../RTL/cortexm0ds_logic.v(14958)
  not u17981 (Zm1pw6, n5059);  // ../RTL/cortexm0ds_logic.v(14958)
  and u17982 (Lm1pw6, Nn1pw6, Un1pw6);  // ../RTL/cortexm0ds_logic.v(14959)
  and u17983 (n5060, vis_r1_o[12], Voqow6);  // ../RTL/cortexm0ds_logic.v(14960)
  not u17984 (Un1pw6, n5060);  // ../RTL/cortexm0ds_logic.v(14960)
  and u17985 (n5061, vis_r6_o[12], Kmqow6);  // ../RTL/cortexm0ds_logic.v(14961)
  not u17986 (Nn1pw6, n5061);  // ../RTL/cortexm0ds_logic.v(14961)
  and u17987 (Ef1pw6, Bo1pw6, Abwow6);  // ../RTL/cortexm0ds_logic.v(14962)
  and u17988 (n5062, Udxow6, Zw4ju6);  // ../RTL/cortexm0ds_logic.v(14963)
  not u17989 (Abwow6, n5062);  // ../RTL/cortexm0ds_logic.v(14963)
  and u1799 (S02iu6, B22iu6, I22iu6);  // ../RTL/cortexm0ds_logic.v(3702)
  and u17990 (n5063, Io1pw6, Po1pw6);  // ../RTL/cortexm0ds_logic.v(14964)
  not u17991 (Zw4ju6, n5063);  // ../RTL/cortexm0ds_logic.v(14964)
  and u17992 (Po1pw6, Wo1pw6, Dp1pw6);  // ../RTL/cortexm0ds_logic.v(14965)
  and u17993 (Dp1pw6, Kp1pw6, Rp1pw6);  // ../RTL/cortexm0ds_logic.v(14966)
  and u17994 (n5064, Fkfpw6[4], Dfqow6);  // ../RTL/cortexm0ds_logic.v(14967)
  not u17995 (Rp1pw6, n5064);  // ../RTL/cortexm0ds_logic.v(14967)
  and u17996 (Kp1pw6, Yp1pw6, Fq1pw6);  // ../RTL/cortexm0ds_logic.v(14968)
  and u17997 (n5065, vis_psp_o[2], Yfqow6);  // ../RTL/cortexm0ds_logic.v(14969)
  not u17998 (Fq1pw6, n5065);  // ../RTL/cortexm0ds_logic.v(14969)
  and u17999 (n5066, vis_msp_o[2], Fgqow6);  // ../RTL/cortexm0ds_logic.v(14970)
  buf u18 (X0ohu6, A3ipw6);  // ../RTL/cortexm0ds_logic.v(1774)
  not u180 (Svdpw6, Jvvpw6);  // ../RTL/cortexm0ds_logic.v(2030)
  and u1800 (n160, Iahpw6[29], Xl1iu6);  // ../RTL/cortexm0ds_logic.v(3703)
  not u18000 (Yp1pw6, n5066);  // ../RTL/cortexm0ds_logic.v(14970)
  and u18001 (Wo1pw6, Mq1pw6, Tq1pw6);  // ../RTL/cortexm0ds_logic.v(14971)
  and u18002 (n5067, vis_r14_o[4], Ahqow6);  // ../RTL/cortexm0ds_logic.v(14972)
  not u18003 (Tq1pw6, n5067);  // ../RTL/cortexm0ds_logic.v(14972)
  and u18004 (n5068, vis_r12_o[4], Hhqow6);  // ../RTL/cortexm0ds_logic.v(14973)
  not u18005 (Mq1pw6, n5068);  // ../RTL/cortexm0ds_logic.v(14973)
  and u18006 (Io1pw6, Ar1pw6, Hr1pw6);  // ../RTL/cortexm0ds_logic.v(14974)
  and u18007 (Hr1pw6, Or1pw6, Vr1pw6);  // ../RTL/cortexm0ds_logic.v(14975)
  and u18008 (n5069, vis_r9_o[4], Qiqow6);  // ../RTL/cortexm0ds_logic.v(14976)
  not u18009 (Vr1pw6, n5069);  // ../RTL/cortexm0ds_logic.v(14976)
  not u1801 (I22iu6, n160);  // ../RTL/cortexm0ds_logic.v(3703)
  and u18010 (Or1pw6, Cs1pw6, Js1pw6);  // ../RTL/cortexm0ds_logic.v(14977)
  and u18011 (n5070, vis_r11_o[4], Ljqow6);  // ../RTL/cortexm0ds_logic.v(14978)
  not u18012 (Js1pw6, n5070);  // ../RTL/cortexm0ds_logic.v(14978)
  and u18013 (n5071, vis_r10_o[4], Sjqow6);  // ../RTL/cortexm0ds_logic.v(14979)
  not u18014 (Cs1pw6, n5071);  // ../RTL/cortexm0ds_logic.v(14979)
  and u18015 (Ar1pw6, Nwzhu6, Qs1pw6);  // ../RTL/cortexm0ds_logic.v(14980)
  and u18016 (n5072, vis_r8_o[4], Gkqow6);  // ../RTL/cortexm0ds_logic.v(14981)
  not u18017 (Qs1pw6, n5072);  // ../RTL/cortexm0ds_logic.v(14981)
  and u18018 (Nwzhu6, Xs1pw6, Et1pw6);  // ../RTL/cortexm0ds_logic.v(14982)
  and u18019 (Et1pw6, Lt1pw6, St1pw6);  // ../RTL/cortexm0ds_logic.v(14983)
  and u1802 (n161, Iahpw6[30], Z4yhu6);  // ../RTL/cortexm0ds_logic.v(3704)
  and u18020 (St1pw6, Zt1pw6, Gu1pw6);  // ../RTL/cortexm0ds_logic.v(14984)
  and u18021 (n5073, vis_r0_o[4], Cpqow6);  // ../RTL/cortexm0ds_logic.v(14985)
  not u18022 (Gu1pw6, n5073);  // ../RTL/cortexm0ds_logic.v(14985)
  and u18023 (n5074, vis_r2_o[4], Dmqow6);  // ../RTL/cortexm0ds_logic.v(14986)
  not u18024 (Zt1pw6, n5074);  // ../RTL/cortexm0ds_logic.v(14986)
  and u18025 (Lt1pw6, Nu1pw6, Uu1pw6);  // ../RTL/cortexm0ds_logic.v(14987)
  and u18026 (n5075, vis_r5_o[4], Fnqow6);  // ../RTL/cortexm0ds_logic.v(14988)
  not u18027 (Uu1pw6, n5075);  // ../RTL/cortexm0ds_logic.v(14988)
  and u18028 (n5076, vis_r4_o[4], Mnqow6);  // ../RTL/cortexm0ds_logic.v(14989)
  not u18029 (Nu1pw6, n5076);  // ../RTL/cortexm0ds_logic.v(14989)
  not u1803 (B22iu6, n161);  // ../RTL/cortexm0ds_logic.v(3704)
  and u18030 (Xs1pw6, Bv1pw6, Iv1pw6);  // ../RTL/cortexm0ds_logic.v(14990)
  and u18031 (Iv1pw6, Pv1pw6, Wv1pw6);  // ../RTL/cortexm0ds_logic.v(14991)
  and u18032 (n5077, vis_r7_o[4], Eqqow6);  // ../RTL/cortexm0ds_logic.v(14992)
  not u18033 (Wv1pw6, n5077);  // ../RTL/cortexm0ds_logic.v(14992)
  and u18034 (n5078, vis_r3_o[4], Xpqow6);  // ../RTL/cortexm0ds_logic.v(14993)
  not u18035 (Pv1pw6, n5078);  // ../RTL/cortexm0ds_logic.v(14993)
  and u18036 (Bv1pw6, Dw1pw6, Kw1pw6);  // ../RTL/cortexm0ds_logic.v(14994)
  and u18037 (n5079, vis_r1_o[4], Voqow6);  // ../RTL/cortexm0ds_logic.v(14995)
  not u18038 (Kw1pw6, n5079);  // ../RTL/cortexm0ds_logic.v(14995)
  and u18039 (n5080, vis_r6_o[4], Kmqow6);  // ../RTL/cortexm0ds_logic.v(14996)
  and u1804 (n162, P22iu6, W22iu6);  // ../RTL/cortexm0ds_logic.v(3705)
  not u18040 (Dw1pw6, n5080);  // ../RTL/cortexm0ds_logic.v(14996)
  and u18041 (n5081, X44iu6, R0nhu6);  // ../RTL/cortexm0ds_logic.v(14997)
  not u18042 (Bo1pw6, n5081);  // ../RTL/cortexm0ds_logic.v(14997)
  and u18043 (X44iu6, Shhpw6[12], Iqzhu6);  // ../RTL/cortexm0ds_logic.v(14998)
  and u18044 (n5082, Yyzow6, In8ju6);  // ../RTL/cortexm0ds_logic.v(15000)
  not u18045 (Yw1pw6, n5082);  // ../RTL/cortexm0ds_logic.v(15000)
  and u18046 (n5083, Fx1pw6, Mx1pw6);  // ../RTL/cortexm0ds_logic.v(15001)
  not u18047 (In8ju6, n5083);  // ../RTL/cortexm0ds_logic.v(15001)
  and u18048 (Mx1pw6, Tx1pw6, Ay1pw6);  // ../RTL/cortexm0ds_logic.v(15002)
  and u18049 (Ay1pw6, Hy1pw6, Oy1pw6);  // ../RTL/cortexm0ds_logic.v(15003)
  not u1805 (M1yhu6, n162);  // ../RTL/cortexm0ds_logic.v(3705)
  and u18050 (n5084, vis_r11_o[11], Ljqow6);  // ../RTL/cortexm0ds_logic.v(15004)
  not u18051 (Oy1pw6, n5084);  // ../RTL/cortexm0ds_logic.v(15004)
  and u18052 (Hy1pw6, Vy1pw6, Cz1pw6);  // ../RTL/cortexm0ds_logic.v(15005)
  and u18053 (n5085, vis_r9_o[11], Qiqow6);  // ../RTL/cortexm0ds_logic.v(15006)
  not u18054 (Cz1pw6, n5085);  // ../RTL/cortexm0ds_logic.v(15006)
  and u18055 (n5086, Fkfpw6[11], Dfqow6);  // ../RTL/cortexm0ds_logic.v(15007)
  not u18056 (Vy1pw6, n5086);  // ../RTL/cortexm0ds_logic.v(15007)
  and u18057 (Tx1pw6, Jz1pw6, Qz1pw6);  // ../RTL/cortexm0ds_logic.v(15008)
  and u18058 (n5087, vis_r10_o[11], Sjqow6);  // ../RTL/cortexm0ds_logic.v(15009)
  not u18059 (Qz1pw6, n5087);  // ../RTL/cortexm0ds_logic.v(15009)
  and u1806 (W22iu6, D32iu6, K32iu6);  // ../RTL/cortexm0ds_logic.v(3706)
  and u18060 (n5088, vis_psp_o[9], Yfqow6);  // ../RTL/cortexm0ds_logic.v(15010)
  not u18061 (Jz1pw6, n5088);  // ../RTL/cortexm0ds_logic.v(15010)
  and u18062 (Fx1pw6, Xz1pw6, E02pw6);  // ../RTL/cortexm0ds_logic.v(15011)
  and u18063 (E02pw6, L02pw6, S02pw6);  // ../RTL/cortexm0ds_logic.v(15012)
  and u18064 (n5089, vis_r12_o[11], Hhqow6);  // ../RTL/cortexm0ds_logic.v(15013)
  not u18065 (S02pw6, n5089);  // ../RTL/cortexm0ds_logic.v(15013)
  and u18066 (L02pw6, Z02pw6, G12pw6);  // ../RTL/cortexm0ds_logic.v(15014)
  and u18067 (n5090, vis_msp_o[9], Fgqow6);  // ../RTL/cortexm0ds_logic.v(15015)
  not u18068 (G12pw6, n5090);  // ../RTL/cortexm0ds_logic.v(15015)
  and u18069 (n5091, vis_r14_o[11], Ahqow6);  // ../RTL/cortexm0ds_logic.v(15016)
  and u1807 (n163, ECOREVNUM[25], Qz1iu6);  // ../RTL/cortexm0ds_logic.v(3707)
  not u18070 (Z02pw6, n5091);  // ../RTL/cortexm0ds_logic.v(15016)
  and u18071 (Xz1pw6, Z20iu6, N12pw6);  // ../RTL/cortexm0ds_logic.v(15017)
  and u18072 (n5092, vis_r8_o[11], Gkqow6);  // ../RTL/cortexm0ds_logic.v(15018)
  not u18073 (N12pw6, n5092);  // ../RTL/cortexm0ds_logic.v(15018)
  and u18074 (Z20iu6, U12pw6, B22pw6);  // ../RTL/cortexm0ds_logic.v(15019)
  and u18075 (B22pw6, I22pw6, P22pw6);  // ../RTL/cortexm0ds_logic.v(15020)
  and u18076 (P22pw6, W22pw6, D32pw6);  // ../RTL/cortexm0ds_logic.v(15021)
  and u18077 (n5093, vis_r2_o[11], Dmqow6);  // ../RTL/cortexm0ds_logic.v(15022)
  not u18078 (D32pw6, n5093);  // ../RTL/cortexm0ds_logic.v(15022)
  and u18079 (n5094, vis_r6_o[11], Kmqow6);  // ../RTL/cortexm0ds_logic.v(15023)
  not u1808 (K32iu6, n163);  // ../RTL/cortexm0ds_logic.v(3707)
  not u18080 (W22pw6, n5094);  // ../RTL/cortexm0ds_logic.v(15023)
  and u18081 (I22pw6, K32pw6, R32pw6);  // ../RTL/cortexm0ds_logic.v(15024)
  and u18082 (n5095, vis_r5_o[11], Fnqow6);  // ../RTL/cortexm0ds_logic.v(15025)
  not u18083 (R32pw6, n5095);  // ../RTL/cortexm0ds_logic.v(15025)
  and u18084 (n5096, vis_r4_o[11], Mnqow6);  // ../RTL/cortexm0ds_logic.v(15026)
  not u18085 (K32pw6, n5096);  // ../RTL/cortexm0ds_logic.v(15026)
  and u18086 (U12pw6, Y32pw6, F42pw6);  // ../RTL/cortexm0ds_logic.v(15027)
  and u18087 (F42pw6, M42pw6, T42pw6);  // ../RTL/cortexm0ds_logic.v(15028)
  and u18088 (n5097, vis_r1_o[11], Voqow6);  // ../RTL/cortexm0ds_logic.v(15029)
  not u18089 (T42pw6, n5097);  // ../RTL/cortexm0ds_logic.v(15029)
  and u1809 (D32iu6, R32iu6, Y32iu6);  // ../RTL/cortexm0ds_logic.v(3708)
  and u18090 (n5098, vis_r0_o[11], Cpqow6);  // ../RTL/cortexm0ds_logic.v(15030)
  not u18091 (M42pw6, n5098);  // ../RTL/cortexm0ds_logic.v(15030)
  and u18092 (Y32pw6, A52pw6, H52pw6);  // ../RTL/cortexm0ds_logic.v(15031)
  and u18093 (n5099, vis_r3_o[11], Xpqow6);  // ../RTL/cortexm0ds_logic.v(15032)
  not u18094 (H52pw6, n5099);  // ../RTL/cortexm0ds_logic.v(15032)
  and u18095 (n5100, vis_r7_o[11], Eqqow6);  // ../RTL/cortexm0ds_logic.v(15033)
  not u18096 (A52pw6, n5100);  // ../RTL/cortexm0ds_logic.v(15033)
  and u18097 (Rw1pw6, O52pw6, Zkwow6);  // ../RTL/cortexm0ds_logic.v(15034)
  and u18098 (n5101, Udxow6, G36ju6);  // ../RTL/cortexm0ds_logic.v(15035)
  not u18099 (Zkwow6, n5101);  // ../RTL/cortexm0ds_logic.v(15035)
  buf u181 (vis_r2_o[16], U0rax6);  // ../RTL/cortexm0ds_logic.v(2551)
  and u1810 (n164, F42iu6, Cl1iu6);  // ../RTL/cortexm0ds_logic.v(3709)
  and u18100 (n5102, V52pw6, C62pw6);  // ../RTL/cortexm0ds_logic.v(15036)
  not u18101 (G36ju6, n5102);  // ../RTL/cortexm0ds_logic.v(15036)
  and u18102 (C62pw6, J62pw6, Q62pw6);  // ../RTL/cortexm0ds_logic.v(15037)
  and u18103 (Q62pw6, X62pw6, E72pw6);  // ../RTL/cortexm0ds_logic.v(15038)
  and u18104 (n5103, Fkfpw6[3], Dfqow6);  // ../RTL/cortexm0ds_logic.v(15039)
  not u18105 (E72pw6, n5103);  // ../RTL/cortexm0ds_logic.v(15039)
  and u18106 (X62pw6, L72pw6, S72pw6);  // ../RTL/cortexm0ds_logic.v(15040)
  and u18107 (n5104, vis_psp_o[1], Yfqow6);  // ../RTL/cortexm0ds_logic.v(15041)
  not u18108 (S72pw6, n5104);  // ../RTL/cortexm0ds_logic.v(15041)
  and u18109 (n5105, vis_msp_o[1], Fgqow6);  // ../RTL/cortexm0ds_logic.v(15042)
  not u1811 (Y32iu6, n164);  // ../RTL/cortexm0ds_logic.v(3709)
  not u18110 (L72pw6, n5105);  // ../RTL/cortexm0ds_logic.v(15042)
  and u18111 (J62pw6, Z72pw6, G82pw6);  // ../RTL/cortexm0ds_logic.v(15043)
  and u18112 (n5106, vis_r14_o[3], Ahqow6);  // ../RTL/cortexm0ds_logic.v(15044)
  not u18113 (G82pw6, n5106);  // ../RTL/cortexm0ds_logic.v(15044)
  and u18114 (n5107, vis_r12_o[3], Hhqow6);  // ../RTL/cortexm0ds_logic.v(15045)
  not u18115 (Z72pw6, n5107);  // ../RTL/cortexm0ds_logic.v(15045)
  and u18116 (V52pw6, N82pw6, U82pw6);  // ../RTL/cortexm0ds_logic.v(15046)
  and u18117 (U82pw6, B92pw6, I92pw6);  // ../RTL/cortexm0ds_logic.v(15047)
  and u18118 (n5108, vis_r9_o[3], Qiqow6);  // ../RTL/cortexm0ds_logic.v(15048)
  not u18119 (I92pw6, n5108);  // ../RTL/cortexm0ds_logic.v(15048)
  and u1812 (F42iu6, Gwnhu6, M42iu6);  // ../RTL/cortexm0ds_logic.v(3710)
  and u18120 (B92pw6, P92pw6, W92pw6);  // ../RTL/cortexm0ds_logic.v(15049)
  and u18121 (n5109, vis_r11_o[3], Ljqow6);  // ../RTL/cortexm0ds_logic.v(15050)
  not u18122 (W92pw6, n5109);  // ../RTL/cortexm0ds_logic.v(15050)
  and u18123 (n5110, vis_r10_o[3], Sjqow6);  // ../RTL/cortexm0ds_logic.v(15051)
  not u18124 (P92pw6, n5110);  // ../RTL/cortexm0ds_logic.v(15051)
  and u18125 (N82pw6, Uwzhu6, Da2pw6);  // ../RTL/cortexm0ds_logic.v(15052)
  and u18126 (n5111, vis_r8_o[3], Gkqow6);  // ../RTL/cortexm0ds_logic.v(15053)
  not u18127 (Da2pw6, n5111);  // ../RTL/cortexm0ds_logic.v(15053)
  and u18128 (Uwzhu6, Ka2pw6, Ra2pw6);  // ../RTL/cortexm0ds_logic.v(15054)
  and u18129 (Ra2pw6, Ya2pw6, Fb2pw6);  // ../RTL/cortexm0ds_logic.v(15055)
  and u1813 (n165, Zbhpw6[28], T42iu6);  // ../RTL/cortexm0ds_logic.v(3711)
  and u18130 (Fb2pw6, Mb2pw6, Tb2pw6);  // ../RTL/cortexm0ds_logic.v(15056)
  and u18131 (n5112, vis_r0_o[3], Cpqow6);  // ../RTL/cortexm0ds_logic.v(15057)
  not u18132 (Tb2pw6, n5112);  // ../RTL/cortexm0ds_logic.v(15057)
  and u18133 (n5113, vis_r2_o[3], Dmqow6);  // ../RTL/cortexm0ds_logic.v(15058)
  not u18134 (Mb2pw6, n5113);  // ../RTL/cortexm0ds_logic.v(15058)
  and u18135 (Ya2pw6, Ac2pw6, Hc2pw6);  // ../RTL/cortexm0ds_logic.v(15059)
  and u18136 (n5114, vis_r5_o[3], Fnqow6);  // ../RTL/cortexm0ds_logic.v(15060)
  not u18137 (Hc2pw6, n5114);  // ../RTL/cortexm0ds_logic.v(15060)
  and u18138 (n5115, vis_r4_o[3], Mnqow6);  // ../RTL/cortexm0ds_logic.v(15061)
  not u18139 (Ac2pw6, n5115);  // ../RTL/cortexm0ds_logic.v(15061)
  not u1814 (M42iu6, n165);  // ../RTL/cortexm0ds_logic.v(3711)
  and u18140 (Ka2pw6, Oc2pw6, Vc2pw6);  // ../RTL/cortexm0ds_logic.v(15062)
  and u18141 (Vc2pw6, Cd2pw6, Jd2pw6);  // ../RTL/cortexm0ds_logic.v(15063)
  and u18142 (n5116, vis_r7_o[3], Eqqow6);  // ../RTL/cortexm0ds_logic.v(15064)
  not u18143 (Jd2pw6, n5116);  // ../RTL/cortexm0ds_logic.v(15064)
  and u18144 (n5117, vis_r3_o[3], Xpqow6);  // ../RTL/cortexm0ds_logic.v(15065)
  not u18145 (Cd2pw6, n5117);  // ../RTL/cortexm0ds_logic.v(15065)
  and u18146 (Oc2pw6, Qd2pw6, Xd2pw6);  // ../RTL/cortexm0ds_logic.v(15066)
  and u18147 (n5118, vis_r1_o[3], Voqow6);  // ../RTL/cortexm0ds_logic.v(15067)
  not u18148 (Xd2pw6, n5118);  // ../RTL/cortexm0ds_logic.v(15067)
  and u18149 (n5119, vis_r6_o[3], Kmqow6);  // ../RTL/cortexm0ds_logic.v(15068)
  or u1815 (T42iu6, A52iu6, W9ohu6);  // ../RTL/cortexm0ds_logic.v(3712)
  not u18150 (Qd2pw6, n5119);  // ../RTL/cortexm0ds_logic.v(15068)
  and u18151 (n5120, Q44iu6, R0nhu6);  // ../RTL/cortexm0ds_logic.v(15069)
  not u18152 (O52pw6, n5120);  // ../RTL/cortexm0ds_logic.v(15069)
  and u18153 (Q44iu6, Shhpw6[11], Iqzhu6);  // ../RTL/cortexm0ds_logic.v(15070)
  or u18154 (Le2pw6, Vcvow6, Ka8ju6);  // ../RTL/cortexm0ds_logic.v(15072)
  and u18155 (Ka8ju6, Se2pw6, Ze2pw6);  // ../RTL/cortexm0ds_logic.v(15073)
  and u18156 (Ze2pw6, Gf2pw6, Nf2pw6);  // ../RTL/cortexm0ds_logic.v(15074)
  and u18157 (Nf2pw6, Uf2pw6, Bg2pw6);  // ../RTL/cortexm0ds_logic.v(15075)
  and u18158 (n5121, vis_r11_o[10], Ljqow6);  // ../RTL/cortexm0ds_logic.v(15076)
  not u18159 (Bg2pw6, n5121);  // ../RTL/cortexm0ds_logic.v(15076)
  and u1816 (n166, Uthpw6[29], Vk1iu6);  // ../RTL/cortexm0ds_logic.v(3713)
  and u18160 (Uf2pw6, Ig2pw6, Pg2pw6);  // ../RTL/cortexm0ds_logic.v(15077)
  and u18161 (n5122, vis_r9_o[10], Qiqow6);  // ../RTL/cortexm0ds_logic.v(15078)
  not u18162 (Pg2pw6, n5122);  // ../RTL/cortexm0ds_logic.v(15078)
  and u18163 (n5123, Fkfpw6[10], Dfqow6);  // ../RTL/cortexm0ds_logic.v(15079)
  not u18164 (Ig2pw6, n5123);  // ../RTL/cortexm0ds_logic.v(15079)
  and u18165 (Gf2pw6, Wg2pw6, Dh2pw6);  // ../RTL/cortexm0ds_logic.v(15080)
  and u18166 (n5124, vis_r10_o[10], Sjqow6);  // ../RTL/cortexm0ds_logic.v(15081)
  not u18167 (Dh2pw6, n5124);  // ../RTL/cortexm0ds_logic.v(15081)
  and u18168 (n5125, vis_psp_o[8], Yfqow6);  // ../RTL/cortexm0ds_logic.v(15082)
  not u18169 (Wg2pw6, n5125);  // ../RTL/cortexm0ds_logic.v(15082)
  not u1817 (R32iu6, n166);  // ../RTL/cortexm0ds_logic.v(3713)
  and u18170 (Se2pw6, Kh2pw6, Rh2pw6);  // ../RTL/cortexm0ds_logic.v(15083)
  and u18171 (Rh2pw6, Yh2pw6, Fi2pw6);  // ../RTL/cortexm0ds_logic.v(15084)
  and u18172 (n5126, vis_r12_o[10], Hhqow6);  // ../RTL/cortexm0ds_logic.v(15085)
  not u18173 (Fi2pw6, n5126);  // ../RTL/cortexm0ds_logic.v(15085)
  and u18174 (Yh2pw6, Mi2pw6, Ti2pw6);  // ../RTL/cortexm0ds_logic.v(15086)
  and u18175 (n5127, vis_msp_o[8], Fgqow6);  // ../RTL/cortexm0ds_logic.v(15087)
  not u18176 (Ti2pw6, n5127);  // ../RTL/cortexm0ds_logic.v(15087)
  and u18177 (n5128, vis_r14_o[10], Ahqow6);  // ../RTL/cortexm0ds_logic.v(15088)
  not u18178 (Mi2pw6, n5128);  // ../RTL/cortexm0ds_logic.v(15088)
  and u18179 (Kh2pw6, G30iu6, Aj2pw6);  // ../RTL/cortexm0ds_logic.v(15089)
  and u1818 (P22iu6, H52iu6, O52iu6);  // ../RTL/cortexm0ds_logic.v(3714)
  and u18180 (n5129, vis_r8_o[10], Gkqow6);  // ../RTL/cortexm0ds_logic.v(15090)
  not u18181 (Aj2pw6, n5129);  // ../RTL/cortexm0ds_logic.v(15090)
  and u18182 (G30iu6, Hj2pw6, Oj2pw6);  // ../RTL/cortexm0ds_logic.v(15091)
  and u18183 (Oj2pw6, Vj2pw6, Ck2pw6);  // ../RTL/cortexm0ds_logic.v(15092)
  and u18184 (Ck2pw6, Jk2pw6, Qk2pw6);  // ../RTL/cortexm0ds_logic.v(15093)
  and u18185 (n5130, vis_r2_o[10], Dmqow6);  // ../RTL/cortexm0ds_logic.v(15094)
  not u18186 (Qk2pw6, n5130);  // ../RTL/cortexm0ds_logic.v(15094)
  and u18187 (n5131, vis_r6_o[10], Kmqow6);  // ../RTL/cortexm0ds_logic.v(15095)
  not u18188 (Jk2pw6, n5131);  // ../RTL/cortexm0ds_logic.v(15095)
  and u18189 (Vj2pw6, Xk2pw6, El2pw6);  // ../RTL/cortexm0ds_logic.v(15096)
  and u1819 (n167, Iahpw6[28], Xl1iu6);  // ../RTL/cortexm0ds_logic.v(3715)
  and u18190 (n5132, vis_r5_o[10], Fnqow6);  // ../RTL/cortexm0ds_logic.v(15097)
  not u18191 (El2pw6, n5132);  // ../RTL/cortexm0ds_logic.v(15097)
  and u18192 (n5133, vis_r4_o[10], Mnqow6);  // ../RTL/cortexm0ds_logic.v(15098)
  not u18193 (Xk2pw6, n5133);  // ../RTL/cortexm0ds_logic.v(15098)
  and u18194 (Hj2pw6, Ll2pw6, Sl2pw6);  // ../RTL/cortexm0ds_logic.v(15099)
  and u18195 (Sl2pw6, Zl2pw6, Gm2pw6);  // ../RTL/cortexm0ds_logic.v(15100)
  and u18196 (n5134, vis_r1_o[10], Voqow6);  // ../RTL/cortexm0ds_logic.v(15101)
  not u18197 (Gm2pw6, n5134);  // ../RTL/cortexm0ds_logic.v(15101)
  and u18198 (n5135, vis_r0_o[10], Cpqow6);  // ../RTL/cortexm0ds_logic.v(15102)
  not u18199 (Zl2pw6, n5135);  // ../RTL/cortexm0ds_logic.v(15102)
  buf u182 (vis_r1_o[3], Ktppw6);  // ../RTL/cortexm0ds_logic.v(1876)
  not u1820 (O52iu6, n167);  // ../RTL/cortexm0ds_logic.v(3715)
  and u18200 (Ll2pw6, Nm2pw6, Um2pw6);  // ../RTL/cortexm0ds_logic.v(15103)
  and u18201 (n5136, vis_r3_o[10], Xpqow6);  // ../RTL/cortexm0ds_logic.v(15104)
  not u18202 (Um2pw6, n5136);  // ../RTL/cortexm0ds_logic.v(15104)
  and u18203 (n5137, vis_r7_o[10], Eqqow6);  // ../RTL/cortexm0ds_logic.v(15105)
  not u18204 (Nm2pw6, n5137);  // ../RTL/cortexm0ds_logic.v(15105)
  not u18205 (Vcvow6, Yyzow6);  // ../RTL/cortexm0ds_logic.v(15106)
  and u18206 (Yyzow6, Qaxiu6, Bn2pw6);  // ../RTL/cortexm0ds_logic.v(15107)
  and u18207 (n5138, J71iu6, L3ehu6);  // ../RTL/cortexm0ds_logic.v(15108)
  not u18208 (Bn2pw6, n5138);  // ../RTL/cortexm0ds_logic.v(15108)
  and u18209 (Ee2pw6, In2pw6, Fvwow6);  // ../RTL/cortexm0ds_logic.v(15109)
  and u1821 (n168, Iahpw6[29], Z4yhu6);  // ../RTL/cortexm0ds_logic.v(3716)
  and u18210 (n5139, Udxow6, Ot5ju6);  // ../RTL/cortexm0ds_logic.v(15110)
  not u18211 (Fvwow6, n5139);  // ../RTL/cortexm0ds_logic.v(15110)
  and u18212 (n5140, Pn2pw6, Wn2pw6);  // ../RTL/cortexm0ds_logic.v(15111)
  not u18213 (Ot5ju6, n5140);  // ../RTL/cortexm0ds_logic.v(15111)
  and u18214 (Wn2pw6, Do2pw6, Ko2pw6);  // ../RTL/cortexm0ds_logic.v(15112)
  and u18215 (Ko2pw6, Ro2pw6, Yo2pw6);  // ../RTL/cortexm0ds_logic.v(15113)
  and u18216 (n5141, Fkfpw6[2], Dfqow6);  // ../RTL/cortexm0ds_logic.v(15114)
  not u18217 (Yo2pw6, n5141);  // ../RTL/cortexm0ds_logic.v(15114)
  and u18218 (Ro2pw6, Fp2pw6, Mp2pw6);  // ../RTL/cortexm0ds_logic.v(15115)
  and u18219 (n5142, vis_psp_o[0], Yfqow6);  // ../RTL/cortexm0ds_logic.v(15116)
  not u1822 (H52iu6, n168);  // ../RTL/cortexm0ds_logic.v(3716)
  not u18220 (Mp2pw6, n5142);  // ../RTL/cortexm0ds_logic.v(15116)
  and u18221 (Yfqow6, Tp2pw6, Vrfhu6);  // ../RTL/cortexm0ds_logic.v(15117)
  and u18222 (Tp2pw6, Aq2pw6, Hq2pw6);  // ../RTL/cortexm0ds_logic.v(15118)
  and u18223 (n5143, vis_msp_o[0], Fgqow6);  // ../RTL/cortexm0ds_logic.v(15119)
  not u18224 (Fp2pw6, n5143);  // ../RTL/cortexm0ds_logic.v(15119)
  and u18225 (Fgqow6, Oq2pw6, Aq2pw6);  // ../RTL/cortexm0ds_logic.v(15120)
  and u18226 (Oq2pw6, Hq2pw6, Vq2pw6);  // ../RTL/cortexm0ds_logic.v(15121)
  and u18227 (Do2pw6, Cr2pw6, Jr2pw6);  // ../RTL/cortexm0ds_logic.v(15122)
  and u18228 (n5144, vis_r14_o[2], Ahqow6);  // ../RTL/cortexm0ds_logic.v(15123)
  not u18229 (Jr2pw6, n5144);  // ../RTL/cortexm0ds_logic.v(15123)
  and u1823 (n169, V52iu6, C62iu6);  // ../RTL/cortexm0ds_logic.v(3717)
  and u18230 (n5145, vis_r12_o[2], Hhqow6);  // ../RTL/cortexm0ds_logic.v(15124)
  not u18231 (Cr2pw6, n5145);  // ../RTL/cortexm0ds_logic.v(15124)
  and u18232 (Pn2pw6, Qr2pw6, Xr2pw6);  // ../RTL/cortexm0ds_logic.v(15125)
  and u18233 (Xr2pw6, Es2pw6, Ls2pw6);  // ../RTL/cortexm0ds_logic.v(15126)
  and u18234 (n5146, vis_r9_o[2], Qiqow6);  // ../RTL/cortexm0ds_logic.v(15127)
  not u18235 (Ls2pw6, n5146);  // ../RTL/cortexm0ds_logic.v(15127)
  and u18236 (Es2pw6, Ss2pw6, Zs2pw6);  // ../RTL/cortexm0ds_logic.v(15128)
  and u18237 (n5147, vis_r11_o[2], Ljqow6);  // ../RTL/cortexm0ds_logic.v(15129)
  not u18238 (Zs2pw6, n5147);  // ../RTL/cortexm0ds_logic.v(15129)
  and u18239 (n5148, vis_r10_o[2], Sjqow6);  // ../RTL/cortexm0ds_logic.v(15130)
  not u1824 (F1yhu6, n169);  // ../RTL/cortexm0ds_logic.v(3717)
  not u18240 (Ss2pw6, n5148);  // ../RTL/cortexm0ds_logic.v(15130)
  and u18241 (Qr2pw6, Pxzhu6, Gt2pw6);  // ../RTL/cortexm0ds_logic.v(15131)
  and u18242 (n5149, vis_r8_o[2], Gkqow6);  // ../RTL/cortexm0ds_logic.v(15132)
  not u18243 (Gt2pw6, n5149);  // ../RTL/cortexm0ds_logic.v(15132)
  and u18244 (Pxzhu6, Nt2pw6, Ut2pw6);  // ../RTL/cortexm0ds_logic.v(15133)
  and u18245 (Ut2pw6, Bu2pw6, Iu2pw6);  // ../RTL/cortexm0ds_logic.v(15134)
  and u18246 (Iu2pw6, Pu2pw6, Wu2pw6);  // ../RTL/cortexm0ds_logic.v(15135)
  and u18247 (n5150, vis_r0_o[2], Cpqow6);  // ../RTL/cortexm0ds_logic.v(15136)
  not u18248 (Wu2pw6, n5150);  // ../RTL/cortexm0ds_logic.v(15136)
  and u18249 (n5151, vis_r2_o[2], Dmqow6);  // ../RTL/cortexm0ds_logic.v(15137)
  and u1825 (C62iu6, J62iu6, Q62iu6);  // ../RTL/cortexm0ds_logic.v(3718)
  not u18250 (Pu2pw6, n5151);  // ../RTL/cortexm0ds_logic.v(15137)
  and u18251 (Bu2pw6, Dv2pw6, Kv2pw6);  // ../RTL/cortexm0ds_logic.v(15138)
  and u18252 (n5152, vis_r5_o[2], Fnqow6);  // ../RTL/cortexm0ds_logic.v(15139)
  not u18253 (Kv2pw6, n5152);  // ../RTL/cortexm0ds_logic.v(15139)
  and u18254 (n5153, vis_r4_o[2], Mnqow6);  // ../RTL/cortexm0ds_logic.v(15140)
  not u18255 (Dv2pw6, n5153);  // ../RTL/cortexm0ds_logic.v(15140)
  and u18256 (Nt2pw6, Rv2pw6, Yv2pw6);  // ../RTL/cortexm0ds_logic.v(15141)
  and u18257 (Yv2pw6, Fw2pw6, Mw2pw6);  // ../RTL/cortexm0ds_logic.v(15142)
  and u18258 (n5154, vis_r7_o[2], Eqqow6);  // ../RTL/cortexm0ds_logic.v(15143)
  not u18259 (Mw2pw6, n5154);  // ../RTL/cortexm0ds_logic.v(15143)
  and u1826 (n170, Cl1iu6, Zbhpw6[28]);  // ../RTL/cortexm0ds_logic.v(3719)
  and u18260 (n5155, vis_r3_o[2], Xpqow6);  // ../RTL/cortexm0ds_logic.v(15144)
  not u18261 (Fw2pw6, n5155);  // ../RTL/cortexm0ds_logic.v(15144)
  and u18262 (Rv2pw6, Tw2pw6, Ax2pw6);  // ../RTL/cortexm0ds_logic.v(15145)
  and u18263 (n5156, vis_r1_o[2], Voqow6);  // ../RTL/cortexm0ds_logic.v(15146)
  not u18264 (Ax2pw6, n5156);  // ../RTL/cortexm0ds_logic.v(15146)
  and u18265 (n5157, vis_r6_o[2], Kmqow6);  // ../RTL/cortexm0ds_logic.v(15147)
  not u18266 (Tw2pw6, n5157);  // ../RTL/cortexm0ds_logic.v(15147)
  and u18267 (Udxow6, J71iu6, Sevow6);  // ../RTL/cortexm0ds_logic.v(15148)
  and u18268 (n5158, J44iu6, R0nhu6);  // ../RTL/cortexm0ds_logic.v(15149)
  not u18269 (In2pw6, n5158);  // ../RTL/cortexm0ds_logic.v(15149)
  not u1827 (Q62iu6, n170);  // ../RTL/cortexm0ds_logic.v(3719)
  and u18270 (J44iu6, Shhpw6[10], Iqzhu6);  // ../RTL/cortexm0ds_logic.v(15150)
  and u18271 (n5159, Sevow6, L35ju6);  // ../RTL/cortexm0ds_logic.v(15152)
  not u18272 (Ox2pw6, n5159);  // ../RTL/cortexm0ds_logic.v(15152)
  and u18273 (n5160, Vx2pw6, Cy2pw6);  // ../RTL/cortexm0ds_logic.v(15153)
  not u18274 (L35ju6, n5160);  // ../RTL/cortexm0ds_logic.v(15153)
  and u18275 (Cy2pw6, Jy2pw6, Qy2pw6);  // ../RTL/cortexm0ds_logic.v(15154)
  and u18276 (Qy2pw6, Xy2pw6, Ez2pw6);  // ../RTL/cortexm0ds_logic.v(15155)
  and u18277 (n5161, Fkfpw6[0], Dfqow6);  // ../RTL/cortexm0ds_logic.v(15156)
  not u18278 (Ez2pw6, n5161);  // ../RTL/cortexm0ds_logic.v(15156)
  and u18279 (Dfqow6, Lz2pw6, Aq2pw6);  // ../RTL/cortexm0ds_logic.v(15157)
  and u1828 (J62iu6, X62iu6, E72iu6);  // ../RTL/cortexm0ds_logic.v(3720)
  and u18280 (n5162, vis_r14_o[0], Ahqow6);  // ../RTL/cortexm0ds_logic.v(15158)
  not u18281 (Xy2pw6, n5162);  // ../RTL/cortexm0ds_logic.v(15158)
  and u18282 (Ahqow6, Sz2pw6, Aq2pw6);  // ../RTL/cortexm0ds_logic.v(15159)
  and u18283 (Jy2pw6, Zz2pw6, G03pw6);  // ../RTL/cortexm0ds_logic.v(15160)
  and u18284 (n5163, vis_r12_o[0], Hhqow6);  // ../RTL/cortexm0ds_logic.v(15161)
  not u18285 (G03pw6, n5163);  // ../RTL/cortexm0ds_logic.v(15161)
  and u18286 (Hhqow6, Aq2pw6, N03pw6);  // ../RTL/cortexm0ds_logic.v(15162)
  or u18287 (n5164, Ntniu6, Roniu6);  // ../RTL/cortexm0ds_logic.v(15163)
  not u18288 (Aq2pw6, n5164);  // ../RTL/cortexm0ds_logic.v(15163)
  and u18289 (n5165, vis_r11_o[0], Ljqow6);  // ../RTL/cortexm0ds_logic.v(15164)
  and u1829 (n171, Uthpw6[28], Vk1iu6);  // ../RTL/cortexm0ds_logic.v(3721)
  not u18290 (Zz2pw6, n5165);  // ../RTL/cortexm0ds_logic.v(15164)
  and u18291 (Ljqow6, Lz2pw6, U03pw6);  // ../RTL/cortexm0ds_logic.v(15165)
  or u18292 (n5166, Qrniu6, Ivuow6);  // ../RTL/cortexm0ds_logic.v(15166)
  not u18293 (Lz2pw6, n5166);  // ../RTL/cortexm0ds_logic.v(15166)
  and u18294 (Vx2pw6, B13pw6, I13pw6);  // ../RTL/cortexm0ds_logic.v(15167)
  and u18295 (I13pw6, P13pw6, W13pw6);  // ../RTL/cortexm0ds_logic.v(15168)
  and u18296 (n5167, vis_r10_o[0], Sjqow6);  // ../RTL/cortexm0ds_logic.v(15169)
  not u18297 (W13pw6, n5167);  // ../RTL/cortexm0ds_logic.v(15169)
  and u18298 (Sjqow6, Sz2pw6, U03pw6);  // ../RTL/cortexm0ds_logic.v(15170)
  or u18299 (n5168, Ivuow6, X3fpw6[0]);  // ../RTL/cortexm0ds_logic.v(15171)
  buf u183 (Npdhu6, C1wpw6);  // ../RTL/cortexm0ds_logic.v(2033)
  not u1830 (E72iu6, n171);  // ../RTL/cortexm0ds_logic.v(3721)
  not u18300 (Sz2pw6, n5168);  // ../RTL/cortexm0ds_logic.v(15171)
  and u18301 (n5169, vis_r9_o[0], Qiqow6);  // ../RTL/cortexm0ds_logic.v(15172)
  not u18302 (P13pw6, n5169);  // ../RTL/cortexm0ds_logic.v(15172)
  and u18303 (Qiqow6, U03pw6, Hq2pw6);  // ../RTL/cortexm0ds_logic.v(15173)
  and u18304 (B13pw6, N30iu6, D23pw6);  // ../RTL/cortexm0ds_logic.v(15174)
  and u18305 (n5170, vis_r8_o[0], Gkqow6);  // ../RTL/cortexm0ds_logic.v(15175)
  not u18306 (D23pw6, n5170);  // ../RTL/cortexm0ds_logic.v(15175)
  and u18307 (Gkqow6, U03pw6, N03pw6);  // ../RTL/cortexm0ds_logic.v(15176)
  or u18308 (n5171, Ntniu6, X3fpw6[2]);  // ../RTL/cortexm0ds_logic.v(15177)
  not u18309 (U03pw6, n5171);  // ../RTL/cortexm0ds_logic.v(15177)
  and u1831 (n172, ECOREVNUM[24], Qz1iu6);  // ../RTL/cortexm0ds_logic.v(3722)
  not u18310 (Ntniu6, X3fpw6[3]);  // ../RTL/cortexm0ds_logic.v(15178)
  and u18311 (N30iu6, K23pw6, R23pw6);  // ../RTL/cortexm0ds_logic.v(15179)
  and u18312 (R23pw6, Y23pw6, F33pw6);  // ../RTL/cortexm0ds_logic.v(15180)
  and u18313 (F33pw6, M33pw6, T33pw6);  // ../RTL/cortexm0ds_logic.v(15181)
  and u18314 (n5172, vis_r0_o[0], Cpqow6);  // ../RTL/cortexm0ds_logic.v(15182)
  not u18315 (T33pw6, n5172);  // ../RTL/cortexm0ds_logic.v(15182)
  and u18316 (Cpqow6, A43pw6, N03pw6);  // ../RTL/cortexm0ds_logic.v(15183)
  and u18317 (n5173, vis_r2_o[0], Dmqow6);  // ../RTL/cortexm0ds_logic.v(15184)
  not u18318 (M33pw6, n5173);  // ../RTL/cortexm0ds_logic.v(15184)
  and u18319 (Dmqow6, H43pw6, O43pw6);  // ../RTL/cortexm0ds_logic.v(15185)
  not u1832 (X62iu6, n172);  // ../RTL/cortexm0ds_logic.v(3722)
  or u18320 (n5174, X3fpw6[0], X3fpw6[2]);  // ../RTL/cortexm0ds_logic.v(15186)
  not u18321 (H43pw6, n5174);  // ../RTL/cortexm0ds_logic.v(15186)
  and u18322 (Y23pw6, V43pw6, C53pw6);  // ../RTL/cortexm0ds_logic.v(15187)
  and u18323 (n5175, vis_r5_o[0], Fnqow6);  // ../RTL/cortexm0ds_logic.v(15188)
  not u18324 (C53pw6, n5175);  // ../RTL/cortexm0ds_logic.v(15188)
  and u18325 (Fnqow6, J53pw6, Hq2pw6);  // ../RTL/cortexm0ds_logic.v(15189)
  and u18326 (n5176, vis_r4_o[0], Mnqow6);  // ../RTL/cortexm0ds_logic.v(15190)
  not u18327 (V43pw6, n5176);  // ../RTL/cortexm0ds_logic.v(15190)
  and u18328 (Mnqow6, J53pw6, N03pw6);  // ../RTL/cortexm0ds_logic.v(15191)
  or u18329 (n5177, X3fpw6[0], X3fpw6[1]);  // ../RTL/cortexm0ds_logic.v(15192)
  and u1833 (V52iu6, S72iu6, Z72iu6);  // ../RTL/cortexm0ds_logic.v(3724)
  not u18330 (N03pw6, n5177);  // ../RTL/cortexm0ds_logic.v(15192)
  or u18331 (n5178, Roniu6, X3fpw6[3]);  // ../RTL/cortexm0ds_logic.v(15193)
  not u18332 (J53pw6, n5178);  // ../RTL/cortexm0ds_logic.v(15193)
  and u18333 (K23pw6, Q53pw6, X53pw6);  // ../RTL/cortexm0ds_logic.v(15194)
  and u18334 (X53pw6, E63pw6, L63pw6);  // ../RTL/cortexm0ds_logic.v(15195)
  and u18335 (n5179, vis_r7_o[0], Eqqow6);  // ../RTL/cortexm0ds_logic.v(15196)
  not u18336 (L63pw6, n5179);  // ../RTL/cortexm0ds_logic.v(15196)
  and u18337 (Eqqow6, S63pw6, X3fpw6[0]);  // ../RTL/cortexm0ds_logic.v(15197)
  and u18338 (S63pw6, X3fpw6[2], O43pw6);  // ../RTL/cortexm0ds_logic.v(15198)
  and u18339 (n5180, vis_r3_o[0], Xpqow6);  // ../RTL/cortexm0ds_logic.v(15199)
  and u1834 (n173, Iahpw6[27], Xl1iu6);  // ../RTL/cortexm0ds_logic.v(3725)
  not u18340 (E63pw6, n5180);  // ../RTL/cortexm0ds_logic.v(15199)
  and u18341 (Xpqow6, Z63pw6, X3fpw6[0]);  // ../RTL/cortexm0ds_logic.v(15200)
  and u18342 (Z63pw6, O43pw6, Roniu6);  // ../RTL/cortexm0ds_logic.v(15201)
  not u18343 (Roniu6, X3fpw6[2]);  // ../RTL/cortexm0ds_logic.v(15202)
  and u18344 (Q53pw6, G73pw6, N73pw6);  // ../RTL/cortexm0ds_logic.v(15203)
  and u18345 (n5181, vis_r1_o[0], Voqow6);  // ../RTL/cortexm0ds_logic.v(15204)
  not u18346 (N73pw6, n5181);  // ../RTL/cortexm0ds_logic.v(15204)
  and u18347 (Voqow6, A43pw6, Hq2pw6);  // ../RTL/cortexm0ds_logic.v(15205)
  or u18348 (n5182, Qrniu6, X3fpw6[1]);  // ../RTL/cortexm0ds_logic.v(15206)
  not u18349 (Hq2pw6, n5182);  // ../RTL/cortexm0ds_logic.v(15206)
  not u1835 (Z72iu6, n173);  // ../RTL/cortexm0ds_logic.v(3725)
  or u18350 (n5183, X3fpw6[2], X3fpw6[3]);  // ../RTL/cortexm0ds_logic.v(15207)
  not u18351 (A43pw6, n5183);  // ../RTL/cortexm0ds_logic.v(15207)
  and u18352 (n5184, vis_r6_o[0], Kmqow6);  // ../RTL/cortexm0ds_logic.v(15208)
  not u18353 (G73pw6, n5184);  // ../RTL/cortexm0ds_logic.v(15208)
  and u18354 (Kmqow6, U73pw6, X3fpw6[2]);  // ../RTL/cortexm0ds_logic.v(15209)
  and u18355 (U73pw6, O43pw6, Qrniu6);  // ../RTL/cortexm0ds_logic.v(15210)
  not u18356 (Qrniu6, X3fpw6[0]);  // ../RTL/cortexm0ds_logic.v(15211)
  or u18357 (n5185, Ivuow6, X3fpw6[3]);  // ../RTL/cortexm0ds_logic.v(15212)
  not u18358 (O43pw6, n5185);  // ../RTL/cortexm0ds_logic.v(15212)
  not u18359 (Ivuow6, X3fpw6[1]);  // ../RTL/cortexm0ds_logic.v(15213)
  and u1836 (n174, Iahpw6[28], Z4yhu6);  // ../RTL/cortexm0ds_logic.v(3726)
  and u18360 (Sevow6, L3ehu6, Qaxiu6);  // ../RTL/cortexm0ds_logic.v(15214)
  not u18361 (Qaxiu6, R0nhu6);  // ../RTL/cortexm0ds_logic.v(15215)
  and u18362 (n5186, T24iu6, R0nhu6);  // ../RTL/cortexm0ds_logic.v(15216)
  not u18363 (Hx2pw6, n5186);  // ../RTL/cortexm0ds_logic.v(15216)
  and u18364 (T24iu6, Shhpw6[0], Iqzhu6);  // ../RTL/cortexm0ds_logic.v(15217)
  and u18365 (n5187, B83pw6, I83pw6);  // ../RTL/cortexm0ds_logic.v(15218)
  not u18366 (HTRANS[1], n5187);  // ../RTL/cortexm0ds_logic.v(15218)
  and u18367 (n5188, Xg6iu6, Kzciu6);  // ../RTL/cortexm0ds_logic.v(15219)
  not u18368 (I83pw6, n5188);  // ../RTL/cortexm0ds_logic.v(15219)
  and u18369 (n5189, P83pw6, W83pw6);  // ../RTL/cortexm0ds_logic.v(15220)
  not u1837 (S72iu6, n174);  // ../RTL/cortexm0ds_logic.v(3726)
  not u18370 (Kzciu6, n5189);  // ../RTL/cortexm0ds_logic.v(15220)
  or u18371 (n5190, D93pw6, Jshpw6[28]);  // ../RTL/cortexm0ds_logic.v(15221)
  not u18372 (W83pw6, n5190);  // ../RTL/cortexm0ds_logic.v(15221)
  not u18373 (D93pw6, Jshpw6[31]);  // ../RTL/cortexm0ds_logic.v(15222)
  and u18374 (P83pw6, Jshpw6[30], Jshpw6[29]);  // ../RTL/cortexm0ds_logic.v(15223)
  AL_MUX u18375 (
    .i0(K93pw6),
    .i1(I7cow6),
    .sel(W7cow6),
    .o(B83pw6));  // ../RTL/cortexm0ds_logic.v(15224)
  and u18376 (W7cow6, Ympiu6, L18iu6);  // ../RTL/cortexm0ds_logic.v(15225)
  AL_MUX u18377 (
    .i0(Rx0iu6),
    .i1(Ef1iu6),
    .sel(Dx0iu6),
    .o(I7cow6));  // ../RTL/cortexm0ds_logic.v(15226)
  and u18378 (n5191, R93pw6, S18iu6);  // ../RTL/cortexm0ds_logic.v(15227)
  not u18379 (K93pw6, n5191);  // ../RTL/cortexm0ds_logic.v(15227)
  and u1838 (n175, G82iu6, N82iu6);  // ../RTL/cortexm0ds_logic.v(3727)
  and u18380 (R93pw6, Y93pw6, Z18iu6);  // ../RTL/cortexm0ds_logic.v(15228)
  and u18381 (Wyciu6, Fa3pw6, Ma3pw6);  // ../RTL/cortexm0ds_logic.v(15229)
  not u18382 (Z18iu6, Wyciu6);  // ../RTL/cortexm0ds_logic.v(15229)
  and u18383 (n5192, Ta3pw6, Ab3pw6);  // ../RTL/cortexm0ds_logic.v(15230)
  not u18384 (Ma3pw6, n5192);  // ../RTL/cortexm0ds_logic.v(15230)
  and u18385 (n5193, Iiliu6, Hb3pw6);  // ../RTL/cortexm0ds_logic.v(15231)
  not u18386 (Ab3pw6, n5193);  // ../RTL/cortexm0ds_logic.v(15231)
  or u18387 (Hb3pw6, X71iu6, Ympiu6);  // ../RTL/cortexm0ds_logic.v(15232)
  and u18388 (n5194, J71iu6, Ob3pw6);  // ../RTL/cortexm0ds_logic.v(15233)
  not u18389 (Fa3pw6, n5194);  // ../RTL/cortexm0ds_logic.v(15233)
  not u1839 (Y0yhu6, n175);  // ../RTL/cortexm0ds_logic.v(3727)
  or u18390 (Y93pw6, Pyciu6, V0epw6);  // ../RTL/cortexm0ds_logic.v(15234)
  and u18391 (n5195, Vb3pw6, Ef1iu6);  // ../RTL/cortexm0ds_logic.v(15235)
  not u18392 (Pyciu6, n5195);  // ../RTL/cortexm0ds_logic.v(15235)
  and u18393 (Vb3pw6, Rx0iu6, Dx0iu6);  // ../RTL/cortexm0ds_logic.v(15236)
  and u18394 (n4277[0], Hx2pw6, Ox2pw6);  // ../RTL/cortexm0ds_logic.v(14039)
  AL_MUX u18395 (
    .i0(Jc3pw6),
    .i1(Qc3pw6),
    .sel(Xg6iu6),
    .o(Cc3pw6));  // ../RTL/cortexm0ds_logic.v(15238)
  and u18396 (n7[6], F8yhu6, M8yhu6);  // ../RTL/cortexm0ds_logic.v(3185)
  not u18397 (Qc3pw6, Ht6iu6);  // ../RTL/cortexm0ds_logic.v(15239)
  and u18398 (Jc3pw6, Ob3pw6, Xc3pw6);  // ../RTL/cortexm0ds_logic.v(15240)
  or u18399 (Xc3pw6, Ed3pw6, Sdaiu6);  // ../RTL/cortexm0ds_logic.v(15241)
  not u184 (Tugpw6[9], n1272[9]);  // ../RTL/cortexm0ds_logic.v(16030)
  and u1840 (N82iu6, U82iu6, L72iu6);  // ../RTL/cortexm0ds_logic.v(3728)
  and u18400 (n5196, Ld3pw6, Sd3pw6);  // ../RTL/cortexm0ds_logic.v(15242)
  and u18401 (n5197, Zd3pw6, Ge3pw6);  // ../RTL/cortexm0ds_logic.v(15243)
  not u18402 (Sd3pw6, n5197);  // ../RTL/cortexm0ds_logic.v(15243)
  or u18403 (n5198, Ympiu6, Sdaiu6);  // ../RTL/cortexm0ds_logic.v(15244)
  not u18404 (Ge3pw6, n5198);  // ../RTL/cortexm0ds_logic.v(15244)
  and u18405 (Zd3pw6, Mnxow6, Ze9iu6);  // ../RTL/cortexm0ds_logic.v(15245)
  and u18406 (n5199, Ne3pw6, Aphpw6[1]);  // ../RTL/cortexm0ds_logic.v(15246)
  not u18407 (Ld3pw6, n5199);  // ../RTL/cortexm0ds_logic.v(15246)
  not u18408 (HWDATA[0], n4277[0]);  // ../RTL/cortexm0ds_logic.v(14039)
  not u18409 (HSIZE[0], n5196);  // ../RTL/cortexm0ds_logic.v(15237)
  and u1841 (n176, Uthpw6[27], Vk1iu6);  // ../RTL/cortexm0ds_logic.v(3729)
  and u18410 (n5201, HADDR[29], Bf3pw6);  // ../RTL/cortexm0ds_logic.v(15248)
  not u18411 (Ue3pw6, n5201);  // ../RTL/cortexm0ds_logic.v(15248)
  not u18412 (Bf3pw6, HADDR[31]);  // ../RTL/cortexm0ds_logic.v(15249)
  and u18413 (n5202, If3pw6, Pf3pw6);  // ../RTL/cortexm0ds_logic.v(15251)
  not u18414 (Ef1iu6, n5202);  // ../RTL/cortexm0ds_logic.v(15251)
  or u18415 (Pf3pw6, T2iiu6, R65ju6);  // ../RTL/cortexm0ds_logic.v(15252)
  AL_MUX u18416 (
    .i0(Wtoiu6),
    .i1(Wf3pw6),
    .sel(Mm4ju6),
    .o(R65ju6));  // ../RTL/cortexm0ds_logic.v(15253)
  and u18417 (Wf3pw6, Dg3pw6, Kg3pw6);  // ../RTL/cortexm0ds_logic.v(15254)
  and u18418 (Kg3pw6, Rg3pw6, Yg3pw6);  // ../RTL/cortexm0ds_logic.v(15255)
  and u18419 (Yg3pw6, Fh3pw6, Mh3pw6);  // ../RTL/cortexm0ds_logic.v(15256)
  not u1842 (U82iu6, n176);  // ../RTL/cortexm0ds_logic.v(3729)
  and u18420 (n5203, Jo4ju6, vis_r14_o[31]);  // ../RTL/cortexm0ds_logic.v(15257)
  not u18421 (Mh3pw6, n5203);  // ../RTL/cortexm0ds_logic.v(15257)
  and u18422 (Fh3pw6, Th3pw6, Ai3pw6);  // ../RTL/cortexm0ds_logic.v(15258)
  and u18423 (n5204, Ep4ju6, vis_psp_o[29]);  // ../RTL/cortexm0ds_logic.v(15259)
  not u18424 (Ai3pw6, n5204);  // ../RTL/cortexm0ds_logic.v(15259)
  and u18425 (n5205, Lp4ju6, vis_msp_o[29]);  // ../RTL/cortexm0ds_logic.v(15260)
  not u18426 (Th3pw6, n5205);  // ../RTL/cortexm0ds_logic.v(15260)
  and u18427 (Rg3pw6, Hi3pw6, Oi3pw6);  // ../RTL/cortexm0ds_logic.v(15261)
  and u18428 (n5206, Gq4ju6, vis_r12_o[31]);  // ../RTL/cortexm0ds_logic.v(15262)
  not u18429 (Oi3pw6, n5206);  // ../RTL/cortexm0ds_logic.v(15262)
  and u1843 (G82iu6, B92iu6, I92iu6);  // ../RTL/cortexm0ds_logic.v(3730)
  and u18430 (n5207, Nq4ju6, vis_r11_o[31]);  // ../RTL/cortexm0ds_logic.v(15263)
  not u18431 (Hi3pw6, n5207);  // ../RTL/cortexm0ds_logic.v(15263)
  and u18432 (Dg3pw6, Vi3pw6, Cj3pw6);  // ../RTL/cortexm0ds_logic.v(15264)
  and u18433 (Cj3pw6, Jj3pw6, Qj3pw6);  // ../RTL/cortexm0ds_logic.v(15265)
  and u18434 (n5208, Wr4ju6, vis_r10_o[31]);  // ../RTL/cortexm0ds_logic.v(15266)
  not u18435 (Qj3pw6, n5208);  // ../RTL/cortexm0ds_logic.v(15266)
  and u18436 (n5209, Ds4ju6, vis_r9_o[31]);  // ../RTL/cortexm0ds_logic.v(15267)
  not u18437 (Jj3pw6, n5209);  // ../RTL/cortexm0ds_logic.v(15267)
  and u18438 (Vi3pw6, R50iu6, Xj3pw6);  // ../RTL/cortexm0ds_logic.v(15268)
  and u18439 (n5210, Rs4ju6, vis_r8_o[31]);  // ../RTL/cortexm0ds_logic.v(15269)
  and u1844 (n177, Iahpw6[26], Xl1iu6);  // ../RTL/cortexm0ds_logic.v(3731)
  not u18440 (Xj3pw6, n5210);  // ../RTL/cortexm0ds_logic.v(15269)
  and u18441 (R50iu6, Ek3pw6, Lk3pw6);  // ../RTL/cortexm0ds_logic.v(15270)
  and u18442 (Lk3pw6, Sk3pw6, Zk3pw6);  // ../RTL/cortexm0ds_logic.v(15271)
  and u18443 (Zk3pw6, Gl3pw6, Nl3pw6);  // ../RTL/cortexm0ds_logic.v(15272)
  and u18444 (n5211, V6now6, vis_r2_o[31]);  // ../RTL/cortexm0ds_logic.v(15273)
  not u18445 (Nl3pw6, n5211);  // ../RTL/cortexm0ds_logic.v(15273)
  and u18446 (n5212, C7now6, vis_r6_o[31]);  // ../RTL/cortexm0ds_logic.v(15274)
  not u18447 (Gl3pw6, n5212);  // ../RTL/cortexm0ds_logic.v(15274)
  and u18448 (Sk3pw6, Ul3pw6, Bm3pw6);  // ../RTL/cortexm0ds_logic.v(15275)
  and u18449 (n5213, X7now6, vis_r5_o[31]);  // ../RTL/cortexm0ds_logic.v(15276)
  not u1845 (I92iu6, n177);  // ../RTL/cortexm0ds_logic.v(3731)
  not u18450 (Bm3pw6, n5213);  // ../RTL/cortexm0ds_logic.v(15276)
  and u18451 (n5214, E8now6, vis_r4_o[31]);  // ../RTL/cortexm0ds_logic.v(15277)
  not u18452 (Ul3pw6, n5214);  // ../RTL/cortexm0ds_logic.v(15277)
  and u18453 (Ek3pw6, Im3pw6, Pm3pw6);  // ../RTL/cortexm0ds_logic.v(15278)
  and u18454 (Pm3pw6, Wm3pw6, Dn3pw6);  // ../RTL/cortexm0ds_logic.v(15279)
  and u18455 (n5215, N9now6, vis_r1_o[31]);  // ../RTL/cortexm0ds_logic.v(15280)
  not u18456 (Dn3pw6, n5215);  // ../RTL/cortexm0ds_logic.v(15280)
  and u18457 (n5216, U9now6, vis_r0_o[31]);  // ../RTL/cortexm0ds_logic.v(15281)
  not u18458 (Wm3pw6, n5216);  // ../RTL/cortexm0ds_logic.v(15281)
  and u18459 (Im3pw6, Kn3pw6, Rn3pw6);  // ../RTL/cortexm0ds_logic.v(15282)
  and u1846 (n178, Iahpw6[27], Z4yhu6);  // ../RTL/cortexm0ds_logic.v(3732)
  and u18460 (n5217, Panow6, vis_r3_o[31]);  // ../RTL/cortexm0ds_logic.v(15283)
  not u18461 (Rn3pw6, n5217);  // ../RTL/cortexm0ds_logic.v(15283)
  and u18462 (n5218, Wanow6, vis_r7_o[31]);  // ../RTL/cortexm0ds_logic.v(15284)
  not u18463 (Kn3pw6, n5218);  // ../RTL/cortexm0ds_logic.v(15284)
  not u18464 (Wtoiu6, Fkfpw6[31]);  // ../RTL/cortexm0ds_logic.v(15285)
  and u18465 (If3pw6, Yn3pw6, Fo3pw6);  // ../RTL/cortexm0ds_logic.v(15286)
  and u18466 (n5219, Eafpw6[31], A3iiu6);  // ../RTL/cortexm0ds_logic.v(15287)
  not u18467 (Fo3pw6, n5219);  // ../RTL/cortexm0ds_logic.v(15287)
  and u18468 (n5220, N5fpw6[30], Sdaiu6);  // ../RTL/cortexm0ds_logic.v(15288)
  not u18469 (Yn3pw6, n5220);  // ../RTL/cortexm0ds_logic.v(15288)
  not u1847 (B92iu6, n178);  // ../RTL/cortexm0ds_logic.v(3732)
  or u18470 (HPROT[2], HADDR[30], HADDR[29]);  // ../RTL/cortexm0ds_logic.v(15289)
  and u18471 (L18iu6, Mo3pw6, To3pw6);  // ../RTL/cortexm0ds_logic.v(15291)
  and u18472 (To3pw6, Ap3pw6, Hp3pw6);  // ../RTL/cortexm0ds_logic.v(15292)
  and u18473 (Hp3pw6, Op3pw6, Hq1ju6);  // ../RTL/cortexm0ds_logic.v(15293)
  and u18474 (n5221, Vp3pw6, Pthiu6);  // ../RTL/cortexm0ds_logic.v(15294)
  not u18475 (Hq1ju6, n5221);  // ../RTL/cortexm0ds_logic.v(15294)
  and u18476 (Vp3pw6, Ls1ju6, Y2oiu6);  // ../RTL/cortexm0ds_logic.v(15295)
  and u18477 (Op3pw6, Cq3pw6, Oq1ju6);  // ../RTL/cortexm0ds_logic.v(15296)
  and u18478 (Ap3pw6, Jq3pw6, Qq3pw6);  // ../RTL/cortexm0ds_logic.v(15297)
  and u18479 (n5222, Xq3pw6, Glaiu6);  // ../RTL/cortexm0ds_logic.v(15298)
  and u1848 (n179, P92iu6, W92iu6);  // ../RTL/cortexm0ds_logic.v(3733)
  not u18480 (Qq3pw6, n5222);  // ../RTL/cortexm0ds_logic.v(15298)
  and u18481 (Glaiu6, M2piu6, Cyfpw6[5]);  // ../RTL/cortexm0ds_logic.v(15299)
  and u18482 (M2piu6, Xzmiu6, Y7ghu6);  // ../RTL/cortexm0ds_logic.v(15300)
  and u18483 (n7[5], Ogyhu6, Vgyhu6);  // ../RTL/cortexm0ds_logic.v(3185)
  not u18484 (Xq3pw6, Qy1ju6);  // ../RTL/cortexm0ds_logic.v(15301)
  and u18485 (Jq3pw6, Bgaow6, Er3pw6);  // ../RTL/cortexm0ds_logic.v(15302)
  and u18486 (n5223, I82ju6, Oiaiu6);  // ../RTL/cortexm0ds_logic.v(15303)
  not u18487 (Er3pw6, n5223);  // ../RTL/cortexm0ds_logic.v(15303)
  and u18488 (n5224, Lr3pw6, Whfiu6);  // ../RTL/cortexm0ds_logic.v(15304)
  not u18489 (Bgaow6, n5224);  // ../RTL/cortexm0ds_logic.v(15304)
  not u1849 (R0yhu6, n179);  // ../RTL/cortexm0ds_logic.v(3733)
  and u18490 (Lr3pw6, D6kiu6, Sijiu6);  // ../RTL/cortexm0ds_logic.v(15305)
  and u18491 (Mo3pw6, Sr3pw6, Zr3pw6);  // ../RTL/cortexm0ds_logic.v(15306)
  and u18492 (Zr3pw6, Gs3pw6, Ns3pw6);  // ../RTL/cortexm0ds_logic.v(15307)
  and u18493 (n5225, Qe8iu6, Us3pw6);  // ../RTL/cortexm0ds_logic.v(15308)
  not u18494 (Ns3pw6, n5225);  // ../RTL/cortexm0ds_logic.v(15308)
  and u18495 (n5226, S62ju6, Jc2ju6);  // ../RTL/cortexm0ds_logic.v(15309)
  not u18496 (Us3pw6, n5226);  // ../RTL/cortexm0ds_logic.v(15309)
  or u18497 (S62ju6, Mr0iu6, Cyfpw6[4]);  // ../RTL/cortexm0ds_logic.v(15310)
  and u18498 (Gs3pw6, Bt3pw6, It3pw6);  // ../RTL/cortexm0ds_logic.v(15311)
  and u18499 (n5227, Y0jiu6, Zqaju6);  // ../RTL/cortexm0ds_logic.v(15312)
  buf u185 (vis_r12_o[27], F6tax6);  // ../RTL/cortexm0ds_logic.v(2599)
  and u1850 (W92iu6, Da2iu6, Ka2iu6);  // ../RTL/cortexm0ds_logic.v(3734)
  not u18500 (It3pw6, n5227);  // ../RTL/cortexm0ds_logic.v(15312)
  and u18501 (Zqaju6, Sijiu6, Ii0iu6);  // ../RTL/cortexm0ds_logic.v(15313)
  and u18502 (n5228, Pt3pw6, O96ow6);  // ../RTL/cortexm0ds_logic.v(15314)
  not u18503 (Bt3pw6, n5228);  // ../RTL/cortexm0ds_logic.v(15314)
  and u18504 (O96ow6, Cyfpw6[4], Geaiu6);  // ../RTL/cortexm0ds_logic.v(15315)
  or u18505 (n5229, R2aiu6, Cyfpw6[6]);  // ../RTL/cortexm0ds_logic.v(15316)
  not u18506 (Pt3pw6, n5229);  // ../RTL/cortexm0ds_logic.v(15316)
  and u18507 (Sr3pw6, Yavow6, Rcziu6);  // ../RTL/cortexm0ds_logic.v(15317)
  and u18508 (Yavow6, Wt3pw6, Du3pw6);  // ../RTL/cortexm0ds_logic.v(15318)
  and u18509 (n5230, Ku3pw6, Mo2ju6);  // ../RTL/cortexm0ds_logic.v(15319)
  and u1851 (n180, Uthpw6[26], Vk1iu6);  // ../RTL/cortexm0ds_logic.v(3735)
  not u18510 (Du3pw6, n5230);  // ../RTL/cortexm0ds_logic.v(15319)
  and u18511 (Mo2ju6, Nlaiu6, Hs0iu6);  // ../RTL/cortexm0ds_logic.v(15320)
  or u18512 (n5231, P1bow6, Cyfpw6[4]);  // ../RTL/cortexm0ds_logic.v(15321)
  not u18513 (Ku3pw6, n5231);  // ../RTL/cortexm0ds_logic.v(15321)
  and u18514 (n5232, Ru3pw6, Apaiu6);  // ../RTL/cortexm0ds_logic.v(15322)
  not u18515 (Wt3pw6, n5232);  // ../RTL/cortexm0ds_logic.v(15322)
  or u18516 (Jhcpw6, Lkaiu6, Mr0iu6);  // ../RTL/cortexm0ds_logic.v(15323)
  not u18517 (Ru3pw6, Jhcpw6);  // ../RTL/cortexm0ds_logic.v(15323)
  and u18518 (HALTED, Pzwiu6, Wofiu6);  // ../RTL/cortexm0ds_logic.v(15324)
  buf u18519 (vis_r7_o[9], Ez1qw6);  // ../RTL/cortexm0ds_logic.v(2654)
  not u1852 (Ka2iu6, n180);  // ../RTL/cortexm0ds_logic.v(3735)
  buf u18520 (vis_r7_o[21], Lfwax6);  // ../RTL/cortexm0ds_logic.v(2654)
  and u18521 (n5233, N5fpw6[8], Sdaiu6);  // ../RTL/cortexm0ds_logic.v(15327)
  not u18522 (Fv3pw6, n5233);  // ../RTL/cortexm0ds_logic.v(15327)
  and u18523 (Yu3pw6, Mv3pw6, Tv3pw6);  // ../RTL/cortexm0ds_logic.v(15328)
  and u18524 (n5234, B7iiu6, He0iu6);  // ../RTL/cortexm0ds_logic.v(15329)
  not u18525 (Tv3pw6, n5234);  // ../RTL/cortexm0ds_logic.v(15329)
  AL_MUX u18526 (
    .i0(Aw3pw6),
    .i1(Fkfpw6[9]),
    .sel(Cn5ju6),
    .o(He0iu6));  // ../RTL/cortexm0ds_logic.v(15330)
  and u18527 (n5235, Hw3pw6, Ow3pw6);  // ../RTL/cortexm0ds_logic.v(15331)
  not u18528 (Aw3pw6, n5235);  // ../RTL/cortexm0ds_logic.v(15331)
  and u18529 (Ow3pw6, Vw3pw6, Cx3pw6);  // ../RTL/cortexm0ds_logic.v(15332)
  and u1853 (n181, Zbhpw6[26], Cl1iu6);  // ../RTL/cortexm0ds_logic.v(3736)
  and u18530 (Cx3pw6, Jx3pw6, Qx3pw6);  // ../RTL/cortexm0ds_logic.v(15333)
  and u18531 (n5236, Jo4ju6, vis_r14_o[9]);  // ../RTL/cortexm0ds_logic.v(15334)
  not u18532 (Qx3pw6, n5236);  // ../RTL/cortexm0ds_logic.v(15334)
  and u18533 (Jx3pw6, Xx3pw6, Ey3pw6);  // ../RTL/cortexm0ds_logic.v(15335)
  and u18534 (n5237, Ep4ju6, vis_psp_o[7]);  // ../RTL/cortexm0ds_logic.v(15336)
  not u18535 (Ey3pw6, n5237);  // ../RTL/cortexm0ds_logic.v(15336)
  and u18536 (n5238, Lp4ju6, vis_msp_o[7]);  // ../RTL/cortexm0ds_logic.v(15337)
  not u18537 (Xx3pw6, n5238);  // ../RTL/cortexm0ds_logic.v(15337)
  and u18538 (Vw3pw6, Ly3pw6, Sy3pw6);  // ../RTL/cortexm0ds_logic.v(15338)
  and u18539 (n5239, Gq4ju6, vis_r12_o[9]);  // ../RTL/cortexm0ds_logic.v(15339)
  not u1854 (Da2iu6, n181);  // ../RTL/cortexm0ds_logic.v(3736)
  not u18540 (Sy3pw6, n5239);  // ../RTL/cortexm0ds_logic.v(15339)
  and u18541 (n5240, Nq4ju6, vis_r11_o[9]);  // ../RTL/cortexm0ds_logic.v(15340)
  not u18542 (Ly3pw6, n5240);  // ../RTL/cortexm0ds_logic.v(15340)
  and u18543 (Hw3pw6, Zy3pw6, Gz3pw6);  // ../RTL/cortexm0ds_logic.v(15341)
  and u18544 (Gz3pw6, Nz3pw6, Uz3pw6);  // ../RTL/cortexm0ds_logic.v(15342)
  and u18545 (n5241, Wr4ju6, vis_r10_o[9]);  // ../RTL/cortexm0ds_logic.v(15343)
  not u18546 (Uz3pw6, n5241);  // ../RTL/cortexm0ds_logic.v(15343)
  and u18547 (n5242, Ds4ju6, vis_r9_o[9]);  // ../RTL/cortexm0ds_logic.v(15344)
  not u18548 (Nz3pw6, n5242);  // ../RTL/cortexm0ds_logic.v(15344)
  and u18549 (Zy3pw6, U30iu6, B04pw6);  // ../RTL/cortexm0ds_logic.v(15345)
  and u1855 (P92iu6, Ra2iu6, Ya2iu6);  // ../RTL/cortexm0ds_logic.v(3737)
  and u18550 (n5243, Rs4ju6, vis_r8_o[9]);  // ../RTL/cortexm0ds_logic.v(15346)
  not u18551 (B04pw6, n5243);  // ../RTL/cortexm0ds_logic.v(15346)
  and u18552 (U30iu6, I04pw6, P04pw6);  // ../RTL/cortexm0ds_logic.v(15347)
  and u18553 (P04pw6, W04pw6, D14pw6);  // ../RTL/cortexm0ds_logic.v(15348)
  and u18554 (D14pw6, K14pw6, R14pw6);  // ../RTL/cortexm0ds_logic.v(15349)
  and u18555 (n5244, V6now6, vis_r2_o[9]);  // ../RTL/cortexm0ds_logic.v(15350)
  not u18556 (R14pw6, n5244);  // ../RTL/cortexm0ds_logic.v(15350)
  and u18557 (n5245, C7now6, vis_r6_o[9]);  // ../RTL/cortexm0ds_logic.v(15351)
  not u18558 (K14pw6, n5245);  // ../RTL/cortexm0ds_logic.v(15351)
  and u18559 (W04pw6, Y14pw6, F24pw6);  // ../RTL/cortexm0ds_logic.v(15352)
  and u1856 (n182, Iahpw6[25], Xl1iu6);  // ../RTL/cortexm0ds_logic.v(3738)
  and u18560 (n5246, X7now6, vis_r5_o[9]);  // ../RTL/cortexm0ds_logic.v(15353)
  not u18561 (F24pw6, n5246);  // ../RTL/cortexm0ds_logic.v(15353)
  and u18562 (n5247, E8now6, vis_r4_o[9]);  // ../RTL/cortexm0ds_logic.v(15354)
  not u18563 (Y14pw6, n5247);  // ../RTL/cortexm0ds_logic.v(15354)
  and u18564 (I04pw6, M24pw6, T24pw6);  // ../RTL/cortexm0ds_logic.v(15355)
  and u18565 (T24pw6, A34pw6, H34pw6);  // ../RTL/cortexm0ds_logic.v(15356)
  and u18566 (n5248, N9now6, vis_r1_o[9]);  // ../RTL/cortexm0ds_logic.v(15357)
  not u18567 (H34pw6, n5248);  // ../RTL/cortexm0ds_logic.v(15357)
  and u18568 (n5249, U9now6, vis_r0_o[9]);  // ../RTL/cortexm0ds_logic.v(15358)
  not u18569 (A34pw6, n5249);  // ../RTL/cortexm0ds_logic.v(15358)
  not u1857 (Ya2iu6, n182);  // ../RTL/cortexm0ds_logic.v(3738)
  and u18570 (M24pw6, O34pw6, V34pw6);  // ../RTL/cortexm0ds_logic.v(15359)
  and u18571 (n5250, Panow6, vis_r3_o[9]);  // ../RTL/cortexm0ds_logic.v(15360)
  not u18572 (V34pw6, n5250);  // ../RTL/cortexm0ds_logic.v(15360)
  and u18573 (n5251, Wanow6, vis_r7_o[9]);  // ../RTL/cortexm0ds_logic.v(15361)
  not u18574 (O34pw6, n5251);  // ../RTL/cortexm0ds_logic.v(15361)
  and u18575 (n5252, Eafpw6[9], A3iiu6);  // ../RTL/cortexm0ds_logic.v(15362)
  not u18576 (Mv3pw6, n5252);  // ../RTL/cortexm0ds_logic.v(15362)
  buf u18577 (vis_r7_o[12], Lvwax6);  // ../RTL/cortexm0ds_logic.v(2654)
  buf u18578 (vis_r7_o[24], M3wax6);  // ../RTL/cortexm0ds_logic.v(2654)
  and u18579 (n5253, N5fpw6[5], Sdaiu6);  // ../RTL/cortexm0ds_logic.v(15365)
  and u1858 (n183, Iahpw6[26], Z4yhu6);  // ../RTL/cortexm0ds_logic.v(3739)
  not u18580 (J44pw6, n5253);  // ../RTL/cortexm0ds_logic.v(15365)
  and u18581 (C44pw6, Q44pw6, X44pw6);  // ../RTL/cortexm0ds_logic.v(15366)
  and u18582 (n5254, B7iiu6, Qf0iu6);  // ../RTL/cortexm0ds_logic.v(15367)
  not u18583 (X44pw6, n5254);  // ../RTL/cortexm0ds_logic.v(15367)
  AL_MUX u18584 (
    .i0(E54pw6),
    .i1(Fkfpw6[6]),
    .sel(Cn5ju6),
    .o(Qf0iu6));  // ../RTL/cortexm0ds_logic.v(15368)
  and u18585 (n5255, L54pw6, S54pw6);  // ../RTL/cortexm0ds_logic.v(15369)
  not u18586 (E54pw6, n5255);  // ../RTL/cortexm0ds_logic.v(15369)
  and u18587 (S54pw6, Z54pw6, G64pw6);  // ../RTL/cortexm0ds_logic.v(15370)
  and u18588 (G64pw6, N64pw6, U64pw6);  // ../RTL/cortexm0ds_logic.v(15371)
  and u18589 (n5256, Jo4ju6, vis_r14_o[6]);  // ../RTL/cortexm0ds_logic.v(15372)
  not u1859 (Ra2iu6, n183);  // ../RTL/cortexm0ds_logic.v(3739)
  not u18590 (U64pw6, n5256);  // ../RTL/cortexm0ds_logic.v(15372)
  and u18591 (N64pw6, B74pw6, I74pw6);  // ../RTL/cortexm0ds_logic.v(15373)
  and u18592 (n5257, Ep4ju6, vis_psp_o[4]);  // ../RTL/cortexm0ds_logic.v(15374)
  not u18593 (I74pw6, n5257);  // ../RTL/cortexm0ds_logic.v(15374)
  and u18594 (n5258, Lp4ju6, vis_msp_o[4]);  // ../RTL/cortexm0ds_logic.v(15375)
  not u18595 (B74pw6, n5258);  // ../RTL/cortexm0ds_logic.v(15375)
  and u18596 (Z54pw6, P74pw6, W74pw6);  // ../RTL/cortexm0ds_logic.v(15376)
  and u18597 (n5259, Gq4ju6, vis_r12_o[6]);  // ../RTL/cortexm0ds_logic.v(15377)
  not u18598 (W74pw6, n5259);  // ../RTL/cortexm0ds_logic.v(15377)
  and u18599 (n5260, Nq4ju6, vis_r11_o[6]);  // ../RTL/cortexm0ds_logic.v(15378)
  buf u186 (vis_psp_o[1], D1zpw6);  // ../RTL/cortexm0ds_logic.v(2085)
  and u1860 (n184, Fb2iu6, Mb2iu6);  // ../RTL/cortexm0ds_logic.v(3740)
  not u18600 (P74pw6, n5260);  // ../RTL/cortexm0ds_logic.v(15378)
  and u18601 (L54pw6, D84pw6, K84pw6);  // ../RTL/cortexm0ds_logic.v(15379)
  and u18602 (K84pw6, R84pw6, Y84pw6);  // ../RTL/cortexm0ds_logic.v(15380)
  and u18603 (n5261, Wr4ju6, vis_r10_o[6]);  // ../RTL/cortexm0ds_logic.v(15381)
  not u18604 (Y84pw6, n5261);  // ../RTL/cortexm0ds_logic.v(15381)
  and u18605 (n5262, Ds4ju6, vis_r9_o[6]);  // ../RTL/cortexm0ds_logic.v(15382)
  not u18606 (R84pw6, n5262);  // ../RTL/cortexm0ds_logic.v(15382)
  and u18607 (D84pw6, P40iu6, F94pw6);  // ../RTL/cortexm0ds_logic.v(15383)
  and u18608 (n5263, Rs4ju6, vis_r8_o[6]);  // ../RTL/cortexm0ds_logic.v(15384)
  not u18609 (F94pw6, n5263);  // ../RTL/cortexm0ds_logic.v(15384)
  not u1861 (K0yhu6, n184);  // ../RTL/cortexm0ds_logic.v(3740)
  and u18610 (P40iu6, M94pw6, T94pw6);  // ../RTL/cortexm0ds_logic.v(15385)
  and u18611 (T94pw6, Aa4pw6, Ha4pw6);  // ../RTL/cortexm0ds_logic.v(15386)
  and u18612 (Ha4pw6, Oa4pw6, Va4pw6);  // ../RTL/cortexm0ds_logic.v(15387)
  and u18613 (n5264, V6now6, vis_r2_o[6]);  // ../RTL/cortexm0ds_logic.v(15388)
  not u18614 (Va4pw6, n5264);  // ../RTL/cortexm0ds_logic.v(15388)
  and u18615 (n5265, C7now6, vis_r6_o[6]);  // ../RTL/cortexm0ds_logic.v(15389)
  not u18616 (Oa4pw6, n5265);  // ../RTL/cortexm0ds_logic.v(15389)
  and u18617 (Aa4pw6, Cb4pw6, Jb4pw6);  // ../RTL/cortexm0ds_logic.v(15390)
  and u18618 (n5266, X7now6, vis_r5_o[6]);  // ../RTL/cortexm0ds_logic.v(15391)
  not u18619 (Jb4pw6, n5266);  // ../RTL/cortexm0ds_logic.v(15391)
  and u1862 (Mb2iu6, Tb2iu6, L72iu6);  // ../RTL/cortexm0ds_logic.v(3741)
  and u18620 (n5267, E8now6, vis_r4_o[6]);  // ../RTL/cortexm0ds_logic.v(15392)
  not u18621 (Cb4pw6, n5267);  // ../RTL/cortexm0ds_logic.v(15392)
  and u18622 (M94pw6, Qb4pw6, Xb4pw6);  // ../RTL/cortexm0ds_logic.v(15393)
  and u18623 (Xb4pw6, Ec4pw6, Lc4pw6);  // ../RTL/cortexm0ds_logic.v(15394)
  and u18624 (n5268, N9now6, vis_r1_o[6]);  // ../RTL/cortexm0ds_logic.v(15395)
  not u18625 (Lc4pw6, n5268);  // ../RTL/cortexm0ds_logic.v(15395)
  and u18626 (n5269, U9now6, vis_r0_o[6]);  // ../RTL/cortexm0ds_logic.v(15396)
  not u18627 (Ec4pw6, n5269);  // ../RTL/cortexm0ds_logic.v(15396)
  and u18628 (Qb4pw6, Sc4pw6, Zc4pw6);  // ../RTL/cortexm0ds_logic.v(15397)
  and u18629 (n5270, Panow6, vis_r3_o[6]);  // ../RTL/cortexm0ds_logic.v(15398)
  and u1863 (n185, Uthpw6[25], Vk1iu6);  // ../RTL/cortexm0ds_logic.v(3742)
  not u18630 (Zc4pw6, n5270);  // ../RTL/cortexm0ds_logic.v(15398)
  and u18631 (n5271, Wanow6, vis_r7_o[6]);  // ../RTL/cortexm0ds_logic.v(15399)
  not u18632 (Sc4pw6, n5271);  // ../RTL/cortexm0ds_logic.v(15399)
  and u18633 (n5272, Eafpw6[6], A3iiu6);  // ../RTL/cortexm0ds_logic.v(15400)
  not u18634 (Q44pw6, n5272);  // ../RTL/cortexm0ds_logic.v(15400)
  and u18635 (n5200[0], L18iu6, Ze9iu6);  // ../RTL/cortexm0ds_logic.v(15247)
  and u18636 (n5273, Gd4pw6, Nd4pw6);  // ../RTL/cortexm0ds_logic.v(15402)
  not u18637 (Rx0iu6, n5273);  // ../RTL/cortexm0ds_logic.v(15402)
  or u18638 (Nd4pw6, T2iiu6, Sg0iu6);  // ../RTL/cortexm0ds_logic.v(15403)
  AL_MUX u18639 (
    .i0(Galiu6),
    .i1(Ud4pw6),
    .sel(Mm4ju6),
    .o(Sg0iu6));  // ../RTL/cortexm0ds_logic.v(15404)
  not u1864 (Tb2iu6, n185);  // ../RTL/cortexm0ds_logic.v(3742)
  and u18640 (Ud4pw6, Be4pw6, Ie4pw6);  // ../RTL/cortexm0ds_logic.v(15405)
  and u18641 (Ie4pw6, Pe4pw6, We4pw6);  // ../RTL/cortexm0ds_logic.v(15406)
  and u18642 (We4pw6, Df4pw6, Kf4pw6);  // ../RTL/cortexm0ds_logic.v(15407)
  and u18643 (n5274, Jo4ju6, vis_r14_o[30]);  // ../RTL/cortexm0ds_logic.v(15408)
  not u18644 (Kf4pw6, n5274);  // ../RTL/cortexm0ds_logic.v(15408)
  and u18645 (Df4pw6, Rf4pw6, Yf4pw6);  // ../RTL/cortexm0ds_logic.v(15409)
  and u18646 (n5275, Ep4ju6, vis_psp_o[28]);  // ../RTL/cortexm0ds_logic.v(15410)
  not u18647 (Yf4pw6, n5275);  // ../RTL/cortexm0ds_logic.v(15410)
  and u18648 (n5276, Lp4ju6, vis_msp_o[28]);  // ../RTL/cortexm0ds_logic.v(15411)
  not u18649 (Rf4pw6, n5276);  // ../RTL/cortexm0ds_logic.v(15411)
  and u1865 (Fb2iu6, Ac2iu6, Hc2iu6);  // ../RTL/cortexm0ds_logic.v(3743)
  and u18650 (Pe4pw6, Fg4pw6, Mg4pw6);  // ../RTL/cortexm0ds_logic.v(15412)
  and u18651 (n5277, Gq4ju6, vis_r12_o[30]);  // ../RTL/cortexm0ds_logic.v(15413)
  not u18652 (Mg4pw6, n5277);  // ../RTL/cortexm0ds_logic.v(15413)
  and u18653 (n5278, Nq4ju6, vis_r11_o[30]);  // ../RTL/cortexm0ds_logic.v(15414)
  not u18654 (Fg4pw6, n5278);  // ../RTL/cortexm0ds_logic.v(15414)
  and u18655 (Be4pw6, Tg4pw6, Ah4pw6);  // ../RTL/cortexm0ds_logic.v(15415)
  and u18656 (Ah4pw6, Hh4pw6, Oh4pw6);  // ../RTL/cortexm0ds_logic.v(15416)
  and u18657 (n5279, Wr4ju6, vis_r10_o[30]);  // ../RTL/cortexm0ds_logic.v(15417)
  not u18658 (Oh4pw6, n5279);  // ../RTL/cortexm0ds_logic.v(15417)
  and u18659 (n5280, Ds4ju6, vis_r9_o[30]);  // ../RTL/cortexm0ds_logic.v(15418)
  and u1866 (n186, Iahpw6[24], Xl1iu6);  // ../RTL/cortexm0ds_logic.v(3744)
  not u18660 (Hh4pw6, n5280);  // ../RTL/cortexm0ds_logic.v(15418)
  and u18661 (Tg4pw6, Y50iu6, Vh4pw6);  // ../RTL/cortexm0ds_logic.v(15419)
  and u18662 (n5281, Rs4ju6, vis_r8_o[30]);  // ../RTL/cortexm0ds_logic.v(15420)
  not u18663 (Vh4pw6, n5281);  // ../RTL/cortexm0ds_logic.v(15420)
  and u18664 (Y50iu6, Ci4pw6, Ji4pw6);  // ../RTL/cortexm0ds_logic.v(15421)
  and u18665 (Ji4pw6, Qi4pw6, Xi4pw6);  // ../RTL/cortexm0ds_logic.v(15422)
  and u18666 (Xi4pw6, Ej4pw6, Lj4pw6);  // ../RTL/cortexm0ds_logic.v(15423)
  and u18667 (n5282, V6now6, vis_r2_o[30]);  // ../RTL/cortexm0ds_logic.v(15424)
  not u18668 (Lj4pw6, n5282);  // ../RTL/cortexm0ds_logic.v(15424)
  and u18669 (n5283, C7now6, vis_r6_o[30]);  // ../RTL/cortexm0ds_logic.v(15425)
  not u1867 (Hc2iu6, n186);  // ../RTL/cortexm0ds_logic.v(3744)
  not u18670 (Ej4pw6, n5283);  // ../RTL/cortexm0ds_logic.v(15425)
  and u18671 (Qi4pw6, Sj4pw6, Zj4pw6);  // ../RTL/cortexm0ds_logic.v(15426)
  and u18672 (n5284, X7now6, vis_r5_o[30]);  // ../RTL/cortexm0ds_logic.v(15427)
  not u18673 (Zj4pw6, n5284);  // ../RTL/cortexm0ds_logic.v(15427)
  and u18674 (n5285, E8now6, vis_r4_o[30]);  // ../RTL/cortexm0ds_logic.v(15428)
  not u18675 (Sj4pw6, n5285);  // ../RTL/cortexm0ds_logic.v(15428)
  and u18676 (Ci4pw6, Gk4pw6, Nk4pw6);  // ../RTL/cortexm0ds_logic.v(15429)
  and u18677 (Nk4pw6, Uk4pw6, Bl4pw6);  // ../RTL/cortexm0ds_logic.v(15430)
  and u18678 (n5286, N9now6, vis_r1_o[30]);  // ../RTL/cortexm0ds_logic.v(15431)
  not u18679 (Bl4pw6, n5286);  // ../RTL/cortexm0ds_logic.v(15431)
  and u1868 (n187, Iahpw6[25], Z4yhu6);  // ../RTL/cortexm0ds_logic.v(3745)
  and u18680 (n5287, U9now6, vis_r0_o[30]);  // ../RTL/cortexm0ds_logic.v(15432)
  not u18681 (Uk4pw6, n5287);  // ../RTL/cortexm0ds_logic.v(15432)
  and u18682 (Gk4pw6, Il4pw6, Pl4pw6);  // ../RTL/cortexm0ds_logic.v(15433)
  and u18683 (n5288, Panow6, vis_r3_o[30]);  // ../RTL/cortexm0ds_logic.v(15434)
  not u18684 (Pl4pw6, n5288);  // ../RTL/cortexm0ds_logic.v(15434)
  and u18685 (n5289, Wanow6, vis_r7_o[30]);  // ../RTL/cortexm0ds_logic.v(15435)
  not u18686 (Il4pw6, n5289);  // ../RTL/cortexm0ds_logic.v(15435)
  not u18687 (Galiu6, Fkfpw6[30]);  // ../RTL/cortexm0ds_logic.v(15436)
  and u18688 (Gd4pw6, Wl4pw6, Dm4pw6);  // ../RTL/cortexm0ds_logic.v(15437)
  and u18689 (n5290, Eafpw6[30], A3iiu6);  // ../RTL/cortexm0ds_logic.v(15438)
  not u1869 (Ac2iu6, n187);  // ../RTL/cortexm0ds_logic.v(3745)
  not u18690 (Dm4pw6, n5290);  // ../RTL/cortexm0ds_logic.v(15438)
  and u18691 (n5291, N5fpw6[29], Sdaiu6);  // ../RTL/cortexm0ds_logic.v(15439)
  not u18692 (Wl4pw6, n5291);  // ../RTL/cortexm0ds_logic.v(15439)
  buf u18693 (Nemhu6, Nvkbx6[6]);  // ../RTL/cortexm0ds_logic.v(3137)
  and u18694 (n5292, Km4pw6, Rm4pw6);  // ../RTL/cortexm0ds_logic.v(15442)
  not u18695 (Dx0iu6, n5292);  // ../RTL/cortexm0ds_logic.v(15442)
  or u18696 (Rm4pw6, T2iiu6, Pi0iu6);  // ../RTL/cortexm0ds_logic.v(15443)
  AL_MUX u18697 (
    .i0(Sm8iu6),
    .i1(Ym4pw6),
    .sel(Mm4ju6),
    .o(Pi0iu6));  // ../RTL/cortexm0ds_logic.v(15444)
  and u18698 (Ym4pw6, Fn4pw6, Mn4pw6);  // ../RTL/cortexm0ds_logic.v(15445)
  and u18699 (Mn4pw6, Tn4pw6, Ao4pw6);  // ../RTL/cortexm0ds_logic.v(15446)
  buf u187 (vis_r4_o[7], Xhuax6);  // ../RTL/cortexm0ds_logic.v(2626)
  and u1870 (n188, Oc2iu6, Vc2iu6);  // ../RTL/cortexm0ds_logic.v(3746)
  and u18700 (Ao4pw6, Ho4pw6, Oo4pw6);  // ../RTL/cortexm0ds_logic.v(15447)
  and u18701 (n5293, Jo4ju6, vis_r14_o[29]);  // ../RTL/cortexm0ds_logic.v(15448)
  not u18702 (Oo4pw6, n5293);  // ../RTL/cortexm0ds_logic.v(15448)
  and u18703 (Ho4pw6, Vo4pw6, Cp4pw6);  // ../RTL/cortexm0ds_logic.v(15449)
  and u18704 (n5294, Ep4ju6, vis_psp_o[27]);  // ../RTL/cortexm0ds_logic.v(15450)
  not u18705 (Cp4pw6, n5294);  // ../RTL/cortexm0ds_logic.v(15450)
  and u18706 (n5295, Lp4ju6, vis_msp_o[27]);  // ../RTL/cortexm0ds_logic.v(15451)
  not u18707 (Vo4pw6, n5295);  // ../RTL/cortexm0ds_logic.v(15451)
  and u18708 (Tn4pw6, Jp4pw6, Qp4pw6);  // ../RTL/cortexm0ds_logic.v(15452)
  and u18709 (n5296, Gq4ju6, vis_r12_o[29]);  // ../RTL/cortexm0ds_logic.v(15453)
  not u1871 (D0yhu6, n188);  // ../RTL/cortexm0ds_logic.v(3746)
  not u18710 (Qp4pw6, n5296);  // ../RTL/cortexm0ds_logic.v(15453)
  and u18711 (n5297, Nq4ju6, vis_r11_o[29]);  // ../RTL/cortexm0ds_logic.v(15454)
  not u18712 (Jp4pw6, n5297);  // ../RTL/cortexm0ds_logic.v(15454)
  and u18713 (Fn4pw6, Xp4pw6, Eq4pw6);  // ../RTL/cortexm0ds_logic.v(15455)
  and u18714 (Eq4pw6, Lq4pw6, Sq4pw6);  // ../RTL/cortexm0ds_logic.v(15456)
  and u18715 (n5298, Wr4ju6, vis_r10_o[29]);  // ../RTL/cortexm0ds_logic.v(15457)
  not u18716 (Sq4pw6, n5298);  // ../RTL/cortexm0ds_logic.v(15457)
  and u18717 (n5299, Ds4ju6, vis_r9_o[29]);  // ../RTL/cortexm0ds_logic.v(15458)
  not u18718 (Lq4pw6, n5299);  // ../RTL/cortexm0ds_logic.v(15458)
  and u18719 (Xp4pw6, M60iu6, Zq4pw6);  // ../RTL/cortexm0ds_logic.v(15459)
  and u1872 (Vc2iu6, Cd2iu6, L72iu6);  // ../RTL/cortexm0ds_logic.v(3747)
  and u18720 (n5300, Rs4ju6, vis_r8_o[29]);  // ../RTL/cortexm0ds_logic.v(15460)
  not u18721 (Zq4pw6, n5300);  // ../RTL/cortexm0ds_logic.v(15460)
  and u18722 (M60iu6, Gr4pw6, Nr4pw6);  // ../RTL/cortexm0ds_logic.v(15461)
  and u18723 (Nr4pw6, Ur4pw6, Bs4pw6);  // ../RTL/cortexm0ds_logic.v(15462)
  and u18724 (Bs4pw6, Is4pw6, Ps4pw6);  // ../RTL/cortexm0ds_logic.v(15463)
  and u18725 (n5301, V6now6, vis_r2_o[29]);  // ../RTL/cortexm0ds_logic.v(15464)
  not u18726 (Ps4pw6, n5301);  // ../RTL/cortexm0ds_logic.v(15464)
  and u18727 (n5302, C7now6, vis_r6_o[29]);  // ../RTL/cortexm0ds_logic.v(15465)
  not u18728 (Is4pw6, n5302);  // ../RTL/cortexm0ds_logic.v(15465)
  and u18729 (Ur4pw6, Ws4pw6, Dt4pw6);  // ../RTL/cortexm0ds_logic.v(15466)
  and u1873 (n189, Uthpw6[24], Vk1iu6);  // ../RTL/cortexm0ds_logic.v(3748)
  and u18730 (n5303, X7now6, vis_r5_o[29]);  // ../RTL/cortexm0ds_logic.v(15467)
  not u18731 (Dt4pw6, n5303);  // ../RTL/cortexm0ds_logic.v(15467)
  and u18732 (n5304, E8now6, vis_r4_o[29]);  // ../RTL/cortexm0ds_logic.v(15468)
  not u18733 (Ws4pw6, n5304);  // ../RTL/cortexm0ds_logic.v(15468)
  and u18734 (Gr4pw6, Kt4pw6, Rt4pw6);  // ../RTL/cortexm0ds_logic.v(15469)
  and u18735 (Rt4pw6, Yt4pw6, Fu4pw6);  // ../RTL/cortexm0ds_logic.v(15470)
  and u18736 (n5305, N9now6, vis_r1_o[29]);  // ../RTL/cortexm0ds_logic.v(15471)
  not u18737 (Fu4pw6, n5305);  // ../RTL/cortexm0ds_logic.v(15471)
  and u18738 (n5306, U9now6, vis_r0_o[29]);  // ../RTL/cortexm0ds_logic.v(15472)
  not u18739 (Yt4pw6, n5306);  // ../RTL/cortexm0ds_logic.v(15472)
  not u1874 (Cd2iu6, n189);  // ../RTL/cortexm0ds_logic.v(3748)
  and u18740 (Kt4pw6, Mu4pw6, Tu4pw6);  // ../RTL/cortexm0ds_logic.v(15473)
  and u18741 (n5307, Panow6, vis_r3_o[29]);  // ../RTL/cortexm0ds_logic.v(15474)
  not u18742 (Tu4pw6, n5307);  // ../RTL/cortexm0ds_logic.v(15474)
  and u18743 (n5308, Wanow6, vis_r7_o[29]);  // ../RTL/cortexm0ds_logic.v(15475)
  not u18744 (Mu4pw6, n5308);  // ../RTL/cortexm0ds_logic.v(15475)
  not u18745 (Sm8iu6, Fkfpw6[29]);  // ../RTL/cortexm0ds_logic.v(15476)
  and u18746 (Km4pw6, Av4pw6, Hv4pw6);  // ../RTL/cortexm0ds_logic.v(15477)
  and u18747 (n5309, Eafpw6[29], A3iiu6);  // ../RTL/cortexm0ds_logic.v(15478)
  not u18748 (Hv4pw6, n5309);  // ../RTL/cortexm0ds_logic.v(15478)
  and u18749 (n5310, N5fpw6[28], Sdaiu6);  // ../RTL/cortexm0ds_logic.v(15479)
  and u1875 (Oc2iu6, Jd2iu6, Qd2iu6);  // ../RTL/cortexm0ds_logic.v(3749)
  not u18750 (Av4pw6, n5310);  // ../RTL/cortexm0ds_logic.v(15479)
  and u18751 (n5311, Ov4pw6, Vv4pw6);  // ../RTL/cortexm0ds_logic.v(15481)
  not u18752 (V0epw6, n5311);  // ../RTL/cortexm0ds_logic.v(15481)
  or u18753 (Vv4pw6, T2iiu6, Wi0iu6);  // ../RTL/cortexm0ds_logic.v(15482)
  AL_MUX u18754 (
    .i0(Seniu6),
    .i1(Cw4pw6),
    .sel(Mm4ju6),
    .o(Wi0iu6));  // ../RTL/cortexm0ds_logic.v(15483)
  and u18755 (Cw4pw6, Jw4pw6, Qw4pw6);  // ../RTL/cortexm0ds_logic.v(15484)
  and u18756 (Qw4pw6, Xw4pw6, Ex4pw6);  // ../RTL/cortexm0ds_logic.v(15485)
  and u18757 (Ex4pw6, Lx4pw6, Sx4pw6);  // ../RTL/cortexm0ds_logic.v(15486)
  and u18758 (n5312, Jo4ju6, vis_r14_o[28]);  // ../RTL/cortexm0ds_logic.v(15487)
  not u18759 (Sx4pw6, n5312);  // ../RTL/cortexm0ds_logic.v(15487)
  and u1876 (n190, Iahpw6[23], Xl1iu6);  // ../RTL/cortexm0ds_logic.v(3750)
  and u18760 (Lx4pw6, Zx4pw6, Gy4pw6);  // ../RTL/cortexm0ds_logic.v(15488)
  and u18761 (n5313, Ep4ju6, vis_psp_o[26]);  // ../RTL/cortexm0ds_logic.v(15489)
  not u18762 (Gy4pw6, n5313);  // ../RTL/cortexm0ds_logic.v(15489)
  and u18763 (n5314, Lp4ju6, vis_msp_o[26]);  // ../RTL/cortexm0ds_logic.v(15490)
  not u18764 (Zx4pw6, n5314);  // ../RTL/cortexm0ds_logic.v(15490)
  and u18765 (Xw4pw6, Ny4pw6, Uy4pw6);  // ../RTL/cortexm0ds_logic.v(15491)
  and u18766 (n5315, Gq4ju6, vis_r12_o[28]);  // ../RTL/cortexm0ds_logic.v(15492)
  not u18767 (Uy4pw6, n5315);  // ../RTL/cortexm0ds_logic.v(15492)
  and u18768 (n5316, Nq4ju6, vis_r11_o[28]);  // ../RTL/cortexm0ds_logic.v(15493)
  not u18769 (Ny4pw6, n5316);  // ../RTL/cortexm0ds_logic.v(15493)
  not u1877 (Qd2iu6, n190);  // ../RTL/cortexm0ds_logic.v(3750)
  and u18770 (Jw4pw6, Bz4pw6, Iz4pw6);  // ../RTL/cortexm0ds_logic.v(15494)
  and u18771 (Iz4pw6, Pz4pw6, Wz4pw6);  // ../RTL/cortexm0ds_logic.v(15495)
  and u18772 (n5317, Wr4ju6, vis_r10_o[28]);  // ../RTL/cortexm0ds_logic.v(15496)
  not u18773 (Wz4pw6, n5317);  // ../RTL/cortexm0ds_logic.v(15496)
  and u18774 (n5318, Ds4ju6, vis_r9_o[28]);  // ../RTL/cortexm0ds_logic.v(15497)
  not u18775 (Pz4pw6, n5318);  // ../RTL/cortexm0ds_logic.v(15497)
  and u18776 (Bz4pw6, T60iu6, D05pw6);  // ../RTL/cortexm0ds_logic.v(15498)
  and u18777 (n5319, Rs4ju6, vis_r8_o[28]);  // ../RTL/cortexm0ds_logic.v(15499)
  not u18778 (D05pw6, n5319);  // ../RTL/cortexm0ds_logic.v(15499)
  buf u18779 (Ufmhu6, Nvkbx6[5]);  // ../RTL/cortexm0ds_logic.v(3137)
  and u1878 (n191, Iahpw6[24], Z4yhu6);  // ../RTL/cortexm0ds_logic.v(3751)
  and u18780 (T60iu6, K05pw6, R05pw6);  // ../RTL/cortexm0ds_logic.v(15501)
  not u18781 (Ltnow6, T60iu6);  // ../RTL/cortexm0ds_logic.v(15501)
  and u18782 (R05pw6, Y05pw6, F15pw6);  // ../RTL/cortexm0ds_logic.v(15502)
  and u18783 (F15pw6, M15pw6, T15pw6);  // ../RTL/cortexm0ds_logic.v(15503)
  and u18784 (n5320, V6now6, vis_r2_o[28]);  // ../RTL/cortexm0ds_logic.v(15504)
  not u18785 (T15pw6, n5320);  // ../RTL/cortexm0ds_logic.v(15504)
  and u18786 (n5321, C7now6, vis_r6_o[28]);  // ../RTL/cortexm0ds_logic.v(15505)
  not u18787 (M15pw6, n5321);  // ../RTL/cortexm0ds_logic.v(15505)
  and u18788 (Y05pw6, A25pw6, H25pw6);  // ../RTL/cortexm0ds_logic.v(15506)
  and u18789 (n5322, X7now6, vis_r5_o[28]);  // ../RTL/cortexm0ds_logic.v(15507)
  not u1879 (Jd2iu6, n191);  // ../RTL/cortexm0ds_logic.v(3751)
  not u18790 (H25pw6, n5322);  // ../RTL/cortexm0ds_logic.v(15507)
  and u18791 (n5323, E8now6, vis_r4_o[28]);  // ../RTL/cortexm0ds_logic.v(15508)
  not u18792 (A25pw6, n5323);  // ../RTL/cortexm0ds_logic.v(15508)
  and u18793 (K05pw6, O25pw6, V25pw6);  // ../RTL/cortexm0ds_logic.v(15509)
  and u18794 (V25pw6, C35pw6, J35pw6);  // ../RTL/cortexm0ds_logic.v(15510)
  and u18795 (n5324, N9now6, vis_r1_o[28]);  // ../RTL/cortexm0ds_logic.v(15511)
  not u18796 (J35pw6, n5324);  // ../RTL/cortexm0ds_logic.v(15511)
  and u18797 (n5325, U9now6, vis_r0_o[28]);  // ../RTL/cortexm0ds_logic.v(15512)
  not u18798 (C35pw6, n5325);  // ../RTL/cortexm0ds_logic.v(15512)
  and u18799 (O25pw6, Q35pw6, X35pw6);  // ../RTL/cortexm0ds_logic.v(15513)
  buf u188 (vis_r14_o[4], Txmax6);  // ../RTL/cortexm0ds_logic.v(2497)
  and u1880 (n192, Xd2iu6, Ee2iu6);  // ../RTL/cortexm0ds_logic.v(3752)
  and u18800 (n5326, Panow6, vis_r3_o[28]);  // ../RTL/cortexm0ds_logic.v(15514)
  not u18801 (X35pw6, n5326);  // ../RTL/cortexm0ds_logic.v(15514)
  and u18802 (n5327, Wanow6, vis_r7_o[28]);  // ../RTL/cortexm0ds_logic.v(15515)
  not u18803 (Q35pw6, n5327);  // ../RTL/cortexm0ds_logic.v(15515)
  not u18804 (Seniu6, Fkfpw6[28]);  // ../RTL/cortexm0ds_logic.v(15516)
  and u18805 (Ov4pw6, E45pw6, L45pw6);  // ../RTL/cortexm0ds_logic.v(15517)
  and u18806 (n5328, N5fpw6[27], Sdaiu6);  // ../RTL/cortexm0ds_logic.v(15518)
  not u18807 (L45pw6, n5328);  // ../RTL/cortexm0ds_logic.v(15518)
  and u18808 (n5329, Eafpw6[28], A3iiu6);  // ../RTL/cortexm0ds_logic.v(15519)
  not u18809 (E45pw6, n5329);  // ../RTL/cortexm0ds_logic.v(15519)
  not u1881 (Wzxhu6, n192);  // ../RTL/cortexm0ds_logic.v(3752)
  and u18810 (n5330, S45pw6, Z45pw6);  // ../RTL/cortexm0ds_logic.v(15521)
  not u18811 (O0epw6, n5330);  // ../RTL/cortexm0ds_logic.v(15521)
  and u18812 (n5331, B7iiu6, Dj0iu6);  // ../RTL/cortexm0ds_logic.v(15522)
  not u18813 (Z45pw6, n5331);  // ../RTL/cortexm0ds_logic.v(15522)
  AL_MUX u18814 (
    .i0(G55pw6),
    .i1(Fkfpw6[27]),
    .sel(Cn5ju6),
    .o(Dj0iu6));  // ../RTL/cortexm0ds_logic.v(15523)
  and u18815 (n5332, N55pw6, U55pw6);  // ../RTL/cortexm0ds_logic.v(15524)
  not u18816 (G55pw6, n5332);  // ../RTL/cortexm0ds_logic.v(15524)
  and u18817 (U55pw6, B65pw6, I65pw6);  // ../RTL/cortexm0ds_logic.v(15525)
  and u18818 (I65pw6, P65pw6, W65pw6);  // ../RTL/cortexm0ds_logic.v(15526)
  and u18819 (n5333, Jo4ju6, vis_r14_o[27]);  // ../RTL/cortexm0ds_logic.v(15527)
  and u1882 (Ee2iu6, Le2iu6, L72iu6);  // ../RTL/cortexm0ds_logic.v(3753)
  not u18820 (W65pw6, n5333);  // ../RTL/cortexm0ds_logic.v(15527)
  and u18821 (P65pw6, D75pw6, K75pw6);  // ../RTL/cortexm0ds_logic.v(15528)
  and u18822 (n5334, Ep4ju6, vis_psp_o[25]);  // ../RTL/cortexm0ds_logic.v(15529)
  not u18823 (K75pw6, n5334);  // ../RTL/cortexm0ds_logic.v(15529)
  and u18824 (n5335, Lp4ju6, vis_msp_o[25]);  // ../RTL/cortexm0ds_logic.v(15530)
  not u18825 (D75pw6, n5335);  // ../RTL/cortexm0ds_logic.v(15530)
  and u18826 (B65pw6, R75pw6, Y75pw6);  // ../RTL/cortexm0ds_logic.v(15531)
  and u18827 (n5336, Gq4ju6, vis_r12_o[27]);  // ../RTL/cortexm0ds_logic.v(15532)
  not u18828 (Y75pw6, n5336);  // ../RTL/cortexm0ds_logic.v(15532)
  and u18829 (n5337, Nq4ju6, vis_r11_o[27]);  // ../RTL/cortexm0ds_logic.v(15533)
  and u1883 (n193, Uthpw6[23], Vk1iu6);  // ../RTL/cortexm0ds_logic.v(3754)
  not u18830 (R75pw6, n5337);  // ../RTL/cortexm0ds_logic.v(15533)
  and u18831 (N55pw6, F85pw6, M85pw6);  // ../RTL/cortexm0ds_logic.v(15534)
  and u18832 (M85pw6, T85pw6, A95pw6);  // ../RTL/cortexm0ds_logic.v(15535)
  and u18833 (n5338, Wr4ju6, vis_r10_o[27]);  // ../RTL/cortexm0ds_logic.v(15536)
  not u18834 (A95pw6, n5338);  // ../RTL/cortexm0ds_logic.v(15536)
  and u18835 (n5339, Ds4ju6, vis_r9_o[27]);  // ../RTL/cortexm0ds_logic.v(15537)
  not u18836 (T85pw6, n5339);  // ../RTL/cortexm0ds_logic.v(15537)
  and u18837 (F85pw6, A70iu6, H95pw6);  // ../RTL/cortexm0ds_logic.v(15538)
  and u18838 (n5340, Rs4ju6, vis_r8_o[27]);  // ../RTL/cortexm0ds_logic.v(15539)
  not u18839 (H95pw6, n5340);  // ../RTL/cortexm0ds_logic.v(15539)
  not u1884 (Le2iu6, n193);  // ../RTL/cortexm0ds_logic.v(3754)
  and u18840 (A70iu6, O95pw6, V95pw6);  // ../RTL/cortexm0ds_logic.v(15540)
  and u18841 (V95pw6, Ca5pw6, Ja5pw6);  // ../RTL/cortexm0ds_logic.v(15541)
  and u18842 (Ja5pw6, Qa5pw6, Xa5pw6);  // ../RTL/cortexm0ds_logic.v(15542)
  and u18843 (n5341, V6now6, vis_r2_o[27]);  // ../RTL/cortexm0ds_logic.v(15543)
  not u18844 (Xa5pw6, n5341);  // ../RTL/cortexm0ds_logic.v(15543)
  and u18845 (n5342, C7now6, vis_r6_o[27]);  // ../RTL/cortexm0ds_logic.v(15544)
  not u18846 (Qa5pw6, n5342);  // ../RTL/cortexm0ds_logic.v(15544)
  and u18847 (Ca5pw6, Eb5pw6, Lb5pw6);  // ../RTL/cortexm0ds_logic.v(15545)
  and u18848 (n5343, X7now6, vis_r5_o[27]);  // ../RTL/cortexm0ds_logic.v(15546)
  not u18849 (Lb5pw6, n5343);  // ../RTL/cortexm0ds_logic.v(15546)
  and u1885 (Xd2iu6, Se2iu6, Ze2iu6);  // ../RTL/cortexm0ds_logic.v(3755)
  and u18850 (n5344, E8now6, vis_r4_o[27]);  // ../RTL/cortexm0ds_logic.v(15547)
  not u18851 (Eb5pw6, n5344);  // ../RTL/cortexm0ds_logic.v(15547)
  and u18852 (O95pw6, Sb5pw6, Zb5pw6);  // ../RTL/cortexm0ds_logic.v(15548)
  and u18853 (Zb5pw6, Gc5pw6, Nc5pw6);  // ../RTL/cortexm0ds_logic.v(15549)
  and u18854 (n5345, N9now6, vis_r1_o[27]);  // ../RTL/cortexm0ds_logic.v(15550)
  not u18855 (Nc5pw6, n5345);  // ../RTL/cortexm0ds_logic.v(15550)
  and u18856 (n5346, U9now6, vis_r0_o[27]);  // ../RTL/cortexm0ds_logic.v(15551)
  not u18857 (Gc5pw6, n5346);  // ../RTL/cortexm0ds_logic.v(15551)
  and u18858 (Sb5pw6, Uc5pw6, Bd5pw6);  // ../RTL/cortexm0ds_logic.v(15552)
  and u18859 (n5347, Panow6, vis_r3_o[27]);  // ../RTL/cortexm0ds_logic.v(15553)
  and u1886 (n194, Iahpw6[22], Xl1iu6);  // ../RTL/cortexm0ds_logic.v(3756)
  not u18860 (Bd5pw6, n5347);  // ../RTL/cortexm0ds_logic.v(15553)
  and u18861 (n5348, Wanow6, vis_r7_o[27]);  // ../RTL/cortexm0ds_logic.v(15554)
  not u18862 (Uc5pw6, n5348);  // ../RTL/cortexm0ds_logic.v(15554)
  and u18863 (S45pw6, Id5pw6, Pd5pw6);  // ../RTL/cortexm0ds_logic.v(15555)
  and u18864 (n5349, N5fpw6[26], Sdaiu6);  // ../RTL/cortexm0ds_logic.v(15556)
  not u18865 (Pd5pw6, n5349);  // ../RTL/cortexm0ds_logic.v(15556)
  and u18866 (n5350, Eafpw6[27], A3iiu6);  // ../RTL/cortexm0ds_logic.v(15557)
  not u18867 (Id5pw6, n5350);  // ../RTL/cortexm0ds_logic.v(15557)
  and u18868 (n5351, Wd5pw6, De5pw6);  // ../RTL/cortexm0ds_logic.v(15559)
  not u18869 (H0epw6, n5351);  // ../RTL/cortexm0ds_logic.v(15559)
  not u1887 (Ze2iu6, n194);  // ../RTL/cortexm0ds_logic.v(3756)
  and u18870 (n5352, B7iiu6, Kj0iu6);  // ../RTL/cortexm0ds_logic.v(15560)
  not u18871 (De5pw6, n5352);  // ../RTL/cortexm0ds_logic.v(15560)
  AL_MUX u18872 (
    .i0(Ke5pw6),
    .i1(Fkfpw6[26]),
    .sel(Cn5ju6),
    .o(Kj0iu6));  // ../RTL/cortexm0ds_logic.v(15561)
  and u18873 (n5353, Re5pw6, Ye5pw6);  // ../RTL/cortexm0ds_logic.v(15562)
  not u18874 (Ke5pw6, n5353);  // ../RTL/cortexm0ds_logic.v(15562)
  and u18875 (Ye5pw6, Ff5pw6, Mf5pw6);  // ../RTL/cortexm0ds_logic.v(15563)
  and u18876 (Mf5pw6, Tf5pw6, Ag5pw6);  // ../RTL/cortexm0ds_logic.v(15564)
  and u18877 (n5354, Jo4ju6, vis_r14_o[26]);  // ../RTL/cortexm0ds_logic.v(15565)
  not u18878 (Ag5pw6, n5354);  // ../RTL/cortexm0ds_logic.v(15565)
  and u18879 (Tf5pw6, Hg5pw6, Og5pw6);  // ../RTL/cortexm0ds_logic.v(15566)
  and u1888 (n195, Iahpw6[23], Z4yhu6);  // ../RTL/cortexm0ds_logic.v(3757)
  and u18880 (n5355, Ep4ju6, vis_psp_o[24]);  // ../RTL/cortexm0ds_logic.v(15567)
  not u18881 (Og5pw6, n5355);  // ../RTL/cortexm0ds_logic.v(15567)
  and u18882 (n5356, Lp4ju6, vis_msp_o[24]);  // ../RTL/cortexm0ds_logic.v(15568)
  not u18883 (Hg5pw6, n5356);  // ../RTL/cortexm0ds_logic.v(15568)
  and u18884 (Ff5pw6, Vg5pw6, Ch5pw6);  // ../RTL/cortexm0ds_logic.v(15569)
  and u18885 (n5357, Gq4ju6, vis_r12_o[26]);  // ../RTL/cortexm0ds_logic.v(15570)
  not u18886 (Ch5pw6, n5357);  // ../RTL/cortexm0ds_logic.v(15570)
  and u18887 (n5358, Nq4ju6, vis_r11_o[26]);  // ../RTL/cortexm0ds_logic.v(15571)
  not u18888 (Vg5pw6, n5358);  // ../RTL/cortexm0ds_logic.v(15571)
  and u18889 (Re5pw6, Jh5pw6, Qh5pw6);  // ../RTL/cortexm0ds_logic.v(15572)
  not u1889 (Se2iu6, n195);  // ../RTL/cortexm0ds_logic.v(3757)
  and u18890 (Qh5pw6, Xh5pw6, Ei5pw6);  // ../RTL/cortexm0ds_logic.v(15573)
  and u18891 (n5359, Wr4ju6, vis_r10_o[26]);  // ../RTL/cortexm0ds_logic.v(15574)
  not u18892 (Ei5pw6, n5359);  // ../RTL/cortexm0ds_logic.v(15574)
  and u18893 (n5360, Ds4ju6, vis_r9_o[26]);  // ../RTL/cortexm0ds_logic.v(15575)
  not u18894 (Xh5pw6, n5360);  // ../RTL/cortexm0ds_logic.v(15575)
  and u18895 (Jh5pw6, H70iu6, Li5pw6);  // ../RTL/cortexm0ds_logic.v(15576)
  and u18896 (n5361, Rs4ju6, vis_r8_o[26]);  // ../RTL/cortexm0ds_logic.v(15577)
  not u18897 (Li5pw6, n5361);  // ../RTL/cortexm0ds_logic.v(15577)
  and u18898 (H70iu6, Si5pw6, Zi5pw6);  // ../RTL/cortexm0ds_logic.v(15578)
  and u18899 (Zi5pw6, Gj5pw6, Nj5pw6);  // ../RTL/cortexm0ds_logic.v(15579)
  buf u189 (vis_r8_o[13], O8sax6);  // ../RTL/cortexm0ds_logic.v(2579)
  and u1890 (n196, Gf2iu6, Nf2iu6);  // ../RTL/cortexm0ds_logic.v(3758)
  and u18900 (Nj5pw6, Uj5pw6, Bk5pw6);  // ../RTL/cortexm0ds_logic.v(15580)
  and u18901 (n5362, V6now6, vis_r2_o[26]);  // ../RTL/cortexm0ds_logic.v(15581)
  not u18902 (Bk5pw6, n5362);  // ../RTL/cortexm0ds_logic.v(15581)
  and u18903 (n5363, C7now6, vis_r6_o[26]);  // ../RTL/cortexm0ds_logic.v(15582)
  not u18904 (Uj5pw6, n5363);  // ../RTL/cortexm0ds_logic.v(15582)
  and u18905 (Gj5pw6, Ik5pw6, Pk5pw6);  // ../RTL/cortexm0ds_logic.v(15583)
  and u18906 (n5364, X7now6, vis_r5_o[26]);  // ../RTL/cortexm0ds_logic.v(15584)
  not u18907 (Pk5pw6, n5364);  // ../RTL/cortexm0ds_logic.v(15584)
  and u18908 (n5365, E8now6, vis_r4_o[26]);  // ../RTL/cortexm0ds_logic.v(15585)
  not u18909 (Ik5pw6, n5365);  // ../RTL/cortexm0ds_logic.v(15585)
  not u1891 (Pzxhu6, n196);  // ../RTL/cortexm0ds_logic.v(3758)
  and u18910 (Si5pw6, Wk5pw6, Dl5pw6);  // ../RTL/cortexm0ds_logic.v(15586)
  and u18911 (Dl5pw6, Kl5pw6, Rl5pw6);  // ../RTL/cortexm0ds_logic.v(15587)
  and u18912 (n5366, N9now6, vis_r1_o[26]);  // ../RTL/cortexm0ds_logic.v(15588)
  not u18913 (Rl5pw6, n5366);  // ../RTL/cortexm0ds_logic.v(15588)
  and u18914 (n5367, U9now6, vis_r0_o[26]);  // ../RTL/cortexm0ds_logic.v(15589)
  not u18915 (Kl5pw6, n5367);  // ../RTL/cortexm0ds_logic.v(15589)
  and u18916 (Wk5pw6, Yl5pw6, Fm5pw6);  // ../RTL/cortexm0ds_logic.v(15590)
  and u18917 (n5368, Panow6, vis_r3_o[26]);  // ../RTL/cortexm0ds_logic.v(15591)
  not u18918 (Fm5pw6, n5368);  // ../RTL/cortexm0ds_logic.v(15591)
  and u18919 (n5369, Wanow6, vis_r7_o[26]);  // ../RTL/cortexm0ds_logic.v(15592)
  and u1892 (n197, Iahpw6[22], Z4yhu6);  // ../RTL/cortexm0ds_logic.v(3759)
  not u18920 (Yl5pw6, n5369);  // ../RTL/cortexm0ds_logic.v(15592)
  and u18921 (Wd5pw6, Mm5pw6, Tm5pw6);  // ../RTL/cortexm0ds_logic.v(15593)
  and u18922 (n5370, N5fpw6[25], Sdaiu6);  // ../RTL/cortexm0ds_logic.v(15594)
  not u18923 (Tm5pw6, n5370);  // ../RTL/cortexm0ds_logic.v(15594)
  and u18924 (n5371, Eafpw6[26], A3iiu6);  // ../RTL/cortexm0ds_logic.v(15595)
  not u18925 (Mm5pw6, n5371);  // ../RTL/cortexm0ds_logic.v(15595)
  and u18926 (n5372, An5pw6, Hn5pw6);  // ../RTL/cortexm0ds_logic.v(15597)
  not u18927 (A0epw6, n5372);  // ../RTL/cortexm0ds_logic.v(15597)
  and u18928 (n5373, B7iiu6, Rj0iu6);  // ../RTL/cortexm0ds_logic.v(15598)
  not u18929 (Hn5pw6, n5373);  // ../RTL/cortexm0ds_logic.v(15598)
  not u1893 (Nf2iu6, n197);  // ../RTL/cortexm0ds_logic.v(3759)
  AL_MUX u18930 (
    .i0(On5pw6),
    .i1(Fkfpw6[25]),
    .sel(Cn5ju6),
    .o(Rj0iu6));  // ../RTL/cortexm0ds_logic.v(15599)
  and u18931 (n5374, Vn5pw6, Co5pw6);  // ../RTL/cortexm0ds_logic.v(15600)
  not u18932 (On5pw6, n5374);  // ../RTL/cortexm0ds_logic.v(15600)
  and u18933 (Co5pw6, Jo5pw6, Qo5pw6);  // ../RTL/cortexm0ds_logic.v(15601)
  and u18934 (Qo5pw6, Xo5pw6, Ep5pw6);  // ../RTL/cortexm0ds_logic.v(15602)
  and u18935 (n5375, Jo4ju6, vis_r14_o[25]);  // ../RTL/cortexm0ds_logic.v(15603)
  not u18936 (Ep5pw6, n5375);  // ../RTL/cortexm0ds_logic.v(15603)
  and u18937 (Xo5pw6, Lp5pw6, Sp5pw6);  // ../RTL/cortexm0ds_logic.v(15604)
  and u18938 (n5376, Ep4ju6, vis_psp_o[23]);  // ../RTL/cortexm0ds_logic.v(15605)
  not u18939 (Sp5pw6, n5376);  // ../RTL/cortexm0ds_logic.v(15605)
  and u1894 (Gf2iu6, Uf2iu6, Bg2iu6);  // ../RTL/cortexm0ds_logic.v(3760)
  and u18940 (n5377, Lp4ju6, vis_msp_o[23]);  // ../RTL/cortexm0ds_logic.v(15606)
  not u18941 (Lp5pw6, n5377);  // ../RTL/cortexm0ds_logic.v(15606)
  and u18942 (Jo5pw6, Zp5pw6, Gq5pw6);  // ../RTL/cortexm0ds_logic.v(15607)
  and u18943 (n5378, Gq4ju6, vis_r12_o[25]);  // ../RTL/cortexm0ds_logic.v(15608)
  not u18944 (Gq5pw6, n5378);  // ../RTL/cortexm0ds_logic.v(15608)
  and u18945 (n5379, Nq4ju6, vis_r11_o[25]);  // ../RTL/cortexm0ds_logic.v(15609)
  not u18946 (Zp5pw6, n5379);  // ../RTL/cortexm0ds_logic.v(15609)
  and u18947 (Vn5pw6, Nq5pw6, Uq5pw6);  // ../RTL/cortexm0ds_logic.v(15610)
  and u18948 (Uq5pw6, Br5pw6, Ir5pw6);  // ../RTL/cortexm0ds_logic.v(15611)
  and u18949 (n5380, Wr4ju6, vis_r10_o[25]);  // ../RTL/cortexm0ds_logic.v(15612)
  and u1895 (n198, Uthpw6[22], Vk1iu6);  // ../RTL/cortexm0ds_logic.v(3761)
  not u18950 (Ir5pw6, n5380);  // ../RTL/cortexm0ds_logic.v(15612)
  and u18951 (n5381, Ds4ju6, vis_r9_o[25]);  // ../RTL/cortexm0ds_logic.v(15613)
  not u18952 (Br5pw6, n5381);  // ../RTL/cortexm0ds_logic.v(15613)
  and u18953 (Nq5pw6, O70iu6, Pr5pw6);  // ../RTL/cortexm0ds_logic.v(15614)
  and u18954 (n5382, Rs4ju6, vis_r8_o[25]);  // ../RTL/cortexm0ds_logic.v(15615)
  not u18955 (Pr5pw6, n5382);  // ../RTL/cortexm0ds_logic.v(15615)
  and u18956 (O70iu6, Wr5pw6, Ds5pw6);  // ../RTL/cortexm0ds_logic.v(15616)
  and u18957 (Ds5pw6, Ks5pw6, Rs5pw6);  // ../RTL/cortexm0ds_logic.v(15617)
  and u18958 (Rs5pw6, Ys5pw6, Ft5pw6);  // ../RTL/cortexm0ds_logic.v(15618)
  and u18959 (n5383, V6now6, vis_r2_o[25]);  // ../RTL/cortexm0ds_logic.v(15619)
  not u1896 (Bg2iu6, n198);  // ../RTL/cortexm0ds_logic.v(3761)
  not u18960 (Ft5pw6, n5383);  // ../RTL/cortexm0ds_logic.v(15619)
  and u18961 (n5384, C7now6, vis_r6_o[25]);  // ../RTL/cortexm0ds_logic.v(15620)
  not u18962 (Ys5pw6, n5384);  // ../RTL/cortexm0ds_logic.v(15620)
  and u18963 (Ks5pw6, Mt5pw6, Tt5pw6);  // ../RTL/cortexm0ds_logic.v(15621)
  and u18964 (n5385, X7now6, vis_r5_o[25]);  // ../RTL/cortexm0ds_logic.v(15622)
  not u18965 (Tt5pw6, n5385);  // ../RTL/cortexm0ds_logic.v(15622)
  and u18966 (n5386, E8now6, vis_r4_o[25]);  // ../RTL/cortexm0ds_logic.v(15623)
  not u18967 (Mt5pw6, n5386);  // ../RTL/cortexm0ds_logic.v(15623)
  and u18968 (Wr5pw6, Au5pw6, Hu5pw6);  // ../RTL/cortexm0ds_logic.v(15624)
  and u18969 (Hu5pw6, Ou5pw6, Vu5pw6);  // ../RTL/cortexm0ds_logic.v(15625)
  and u1897 (n199, Iahpw6[21], Xl1iu6);  // ../RTL/cortexm0ds_logic.v(3762)
  and u18970 (n5387, N9now6, vis_r1_o[25]);  // ../RTL/cortexm0ds_logic.v(15626)
  not u18971 (Vu5pw6, n5387);  // ../RTL/cortexm0ds_logic.v(15626)
  and u18972 (n5388, U9now6, vis_r0_o[25]);  // ../RTL/cortexm0ds_logic.v(15627)
  not u18973 (Ou5pw6, n5388);  // ../RTL/cortexm0ds_logic.v(15627)
  and u18974 (Au5pw6, Cv5pw6, Jv5pw6);  // ../RTL/cortexm0ds_logic.v(15628)
  and u18975 (n5389, Panow6, vis_r3_o[25]);  // ../RTL/cortexm0ds_logic.v(15629)
  not u18976 (Jv5pw6, n5389);  // ../RTL/cortexm0ds_logic.v(15629)
  and u18977 (n5390, Wanow6, vis_r7_o[25]);  // ../RTL/cortexm0ds_logic.v(15630)
  not u18978 (Cv5pw6, n5390);  // ../RTL/cortexm0ds_logic.v(15630)
  and u18979 (An5pw6, Qv5pw6, Xv5pw6);  // ../RTL/cortexm0ds_logic.v(15631)
  not u1898 (Uf2iu6, n199);  // ../RTL/cortexm0ds_logic.v(3762)
  and u18980 (n5391, N5fpw6[24], Sdaiu6);  // ../RTL/cortexm0ds_logic.v(15632)
  not u18981 (Xv5pw6, n5391);  // ../RTL/cortexm0ds_logic.v(15632)
  and u18982 (n5392, Eafpw6[25], A3iiu6);  // ../RTL/cortexm0ds_logic.v(15633)
  not u18983 (Qv5pw6, n5392);  // ../RTL/cortexm0ds_logic.v(15633)
  and u18984 (n5393, Ew5pw6, Lw5pw6);  // ../RTL/cortexm0ds_logic.v(15635)
  not u18985 (Tzdpw6, n5393);  // ../RTL/cortexm0ds_logic.v(15635)
  or u18986 (Lw5pw6, T2iiu6, Yj0iu6);  // ../RTL/cortexm0ds_logic.v(15636)
  AL_MUX u18987 (
    .i0(Kykiu6),
    .i1(Sw5pw6),
    .sel(Mm4ju6),
    .o(Yj0iu6));  // ../RTL/cortexm0ds_logic.v(15637)
  and u18988 (Sw5pw6, Zw5pw6, Gx5pw6);  // ../RTL/cortexm0ds_logic.v(15638)
  and u18989 (Gx5pw6, Nx5pw6, Ux5pw6);  // ../RTL/cortexm0ds_logic.v(15639)
  and u1899 (n200, Ig2iu6, Pg2iu6);  // ../RTL/cortexm0ds_logic.v(3763)
  and u18990 (Ux5pw6, By5pw6, Iy5pw6);  // ../RTL/cortexm0ds_logic.v(15640)
  and u18991 (n5394, Jo4ju6, vis_r14_o[24]);  // ../RTL/cortexm0ds_logic.v(15641)
  not u18992 (Iy5pw6, n5394);  // ../RTL/cortexm0ds_logic.v(15641)
  and u18993 (By5pw6, Py5pw6, Wy5pw6);  // ../RTL/cortexm0ds_logic.v(15642)
  and u18994 (n5395, Ep4ju6, vis_psp_o[22]);  // ../RTL/cortexm0ds_logic.v(15643)
  not u18995 (Wy5pw6, n5395);  // ../RTL/cortexm0ds_logic.v(15643)
  and u18996 (n5396, Lp4ju6, vis_msp_o[22]);  // ../RTL/cortexm0ds_logic.v(15644)
  not u18997 (Py5pw6, n5396);  // ../RTL/cortexm0ds_logic.v(15644)
  and u18998 (Nx5pw6, Dz5pw6, Kz5pw6);  // ../RTL/cortexm0ds_logic.v(15645)
  and u18999 (n5397, Gq4ju6, vis_r12_o[24]);  // ../RTL/cortexm0ds_logic.v(15646)
  buf u19 (Q8nhu6, A5ipw6);  // ../RTL/cortexm0ds_logic.v(1775)
  buf u190 (Vbgpw6[7], C10bx6);  // ../RTL/cortexm0ds_logic.v(3092)
  not u1900 (Izxhu6, n200);  // ../RTL/cortexm0ds_logic.v(3763)
  not u19000 (Kz5pw6, n5397);  // ../RTL/cortexm0ds_logic.v(15646)
  and u19001 (n5398, Nq4ju6, vis_r11_o[24]);  // ../RTL/cortexm0ds_logic.v(15647)
  not u19002 (Dz5pw6, n5398);  // ../RTL/cortexm0ds_logic.v(15647)
  and u19003 (Zw5pw6, Rz5pw6, Yz5pw6);  // ../RTL/cortexm0ds_logic.v(15648)
  and u19004 (Yz5pw6, F06pw6, M06pw6);  // ../RTL/cortexm0ds_logic.v(15649)
  and u19005 (n5399, Wr4ju6, vis_r10_o[24]);  // ../RTL/cortexm0ds_logic.v(15650)
  not u19006 (M06pw6, n5399);  // ../RTL/cortexm0ds_logic.v(15650)
  and u19007 (n5400, Ds4ju6, vis_r9_o[24]);  // ../RTL/cortexm0ds_logic.v(15651)
  not u19008 (F06pw6, n5400);  // ../RTL/cortexm0ds_logic.v(15651)
  and u19009 (Rz5pw6, V70iu6, T06pw6);  // ../RTL/cortexm0ds_logic.v(15652)
  and u1901 (Pg2iu6, Wg2iu6, L72iu6);  // ../RTL/cortexm0ds_logic.v(3764)
  and u19010 (n5401, Rs4ju6, vis_r8_o[24]);  // ../RTL/cortexm0ds_logic.v(15653)
  not u19011 (T06pw6, n5401);  // ../RTL/cortexm0ds_logic.v(15653)
  and u19012 (V70iu6, A16pw6, H16pw6);  // ../RTL/cortexm0ds_logic.v(15654)
  and u19013 (H16pw6, O16pw6, V16pw6);  // ../RTL/cortexm0ds_logic.v(15655)
  and u19014 (V16pw6, C26pw6, J26pw6);  // ../RTL/cortexm0ds_logic.v(15656)
  and u19015 (n5402, V6now6, vis_r2_o[24]);  // ../RTL/cortexm0ds_logic.v(15657)
  not u19016 (J26pw6, n5402);  // ../RTL/cortexm0ds_logic.v(15657)
  and u19017 (n5403, C7now6, vis_r6_o[24]);  // ../RTL/cortexm0ds_logic.v(15658)
  not u19018 (C26pw6, n5403);  // ../RTL/cortexm0ds_logic.v(15658)
  and u19019 (O16pw6, Q26pw6, X26pw6);  // ../RTL/cortexm0ds_logic.v(15659)
  and u1902 (n201, Uthpw6[21], Vk1iu6);  // ../RTL/cortexm0ds_logic.v(3765)
  and u19020 (n5404, X7now6, vis_r5_o[24]);  // ../RTL/cortexm0ds_logic.v(15660)
  not u19021 (X26pw6, n5404);  // ../RTL/cortexm0ds_logic.v(15660)
  and u19022 (n5405, E8now6, vis_r4_o[24]);  // ../RTL/cortexm0ds_logic.v(15661)
  not u19023 (Q26pw6, n5405);  // ../RTL/cortexm0ds_logic.v(15661)
  and u19024 (A16pw6, E36pw6, L36pw6);  // ../RTL/cortexm0ds_logic.v(15662)
  and u19025 (L36pw6, S36pw6, Z36pw6);  // ../RTL/cortexm0ds_logic.v(15663)
  and u19026 (n5406, N9now6, vis_r1_o[24]);  // ../RTL/cortexm0ds_logic.v(15664)
  not u19027 (Z36pw6, n5406);  // ../RTL/cortexm0ds_logic.v(15664)
  and u19028 (n5407, U9now6, vis_r0_o[24]);  // ../RTL/cortexm0ds_logic.v(15665)
  not u19029 (S36pw6, n5407);  // ../RTL/cortexm0ds_logic.v(15665)
  not u1903 (Wg2iu6, n201);  // ../RTL/cortexm0ds_logic.v(3765)
  and u19030 (E36pw6, G46pw6, N46pw6);  // ../RTL/cortexm0ds_logic.v(15666)
  and u19031 (n5408, Panow6, vis_r3_o[24]);  // ../RTL/cortexm0ds_logic.v(15667)
  not u19032 (N46pw6, n5408);  // ../RTL/cortexm0ds_logic.v(15667)
  and u19033 (n5409, Wanow6, vis_r7_o[24]);  // ../RTL/cortexm0ds_logic.v(15668)
  not u19034 (G46pw6, n5409);  // ../RTL/cortexm0ds_logic.v(15668)
  not u19035 (Kykiu6, Fkfpw6[24]);  // ../RTL/cortexm0ds_logic.v(15669)
  and u19036 (Ew5pw6, U46pw6, B56pw6);  // ../RTL/cortexm0ds_logic.v(15670)
  and u19037 (n5410, N5fpw6[23], Sdaiu6);  // ../RTL/cortexm0ds_logic.v(15671)
  not u19038 (B56pw6, n5410);  // ../RTL/cortexm0ds_logic.v(15671)
  and u19039 (n5411, Eafpw6[24], A3iiu6);  // ../RTL/cortexm0ds_logic.v(15672)
  and u1904 (Ig2iu6, Dh2iu6, Kh2iu6);  // ../RTL/cortexm0ds_logic.v(3766)
  not u19040 (U46pw6, n5411);  // ../RTL/cortexm0ds_logic.v(15672)
  and u19041 (n5412, I56pw6, P56pw6);  // ../RTL/cortexm0ds_logic.v(15674)
  not u19042 (Mzdpw6, n5412);  // ../RTL/cortexm0ds_logic.v(15674)
  or u19043 (P56pw6, T2iiu6, Fk0iu6);  // ../RTL/cortexm0ds_logic.v(15675)
  AL_MUX u19044 (
    .i0(Ax9iu6),
    .i1(W56pw6),
    .sel(Mm4ju6),
    .o(Fk0iu6));  // ../RTL/cortexm0ds_logic.v(15676)
  and u19045 (W56pw6, D66pw6, K66pw6);  // ../RTL/cortexm0ds_logic.v(15677)
  and u19046 (K66pw6, R66pw6, Y66pw6);  // ../RTL/cortexm0ds_logic.v(15678)
  and u19047 (Y66pw6, F76pw6, M76pw6);  // ../RTL/cortexm0ds_logic.v(15679)
  and u19048 (n5413, Jo4ju6, vis_r14_o[23]);  // ../RTL/cortexm0ds_logic.v(15680)
  not u19049 (M76pw6, n5413);  // ../RTL/cortexm0ds_logic.v(15680)
  and u1905 (n202, Iahpw6[20], Xl1iu6);  // ../RTL/cortexm0ds_logic.v(3767)
  and u19050 (F76pw6, T76pw6, A86pw6);  // ../RTL/cortexm0ds_logic.v(15681)
  and u19051 (n5414, Ep4ju6, vis_psp_o[21]);  // ../RTL/cortexm0ds_logic.v(15682)
  not u19052 (A86pw6, n5414);  // ../RTL/cortexm0ds_logic.v(15682)
  and u19053 (n5415, Lp4ju6, vis_msp_o[21]);  // ../RTL/cortexm0ds_logic.v(15683)
  not u19054 (T76pw6, n5415);  // ../RTL/cortexm0ds_logic.v(15683)
  and u19055 (R66pw6, H86pw6, O86pw6);  // ../RTL/cortexm0ds_logic.v(15684)
  and u19056 (n5416, Gq4ju6, vis_r12_o[23]);  // ../RTL/cortexm0ds_logic.v(15685)
  not u19057 (O86pw6, n5416);  // ../RTL/cortexm0ds_logic.v(15685)
  and u19058 (n5417, Nq4ju6, vis_r11_o[23]);  // ../RTL/cortexm0ds_logic.v(15686)
  not u19059 (H86pw6, n5417);  // ../RTL/cortexm0ds_logic.v(15686)
  not u1906 (Kh2iu6, n202);  // ../RTL/cortexm0ds_logic.v(3767)
  and u19060 (D66pw6, V86pw6, C96pw6);  // ../RTL/cortexm0ds_logic.v(15687)
  and u19061 (C96pw6, J96pw6, Q96pw6);  // ../RTL/cortexm0ds_logic.v(15688)
  and u19062 (n5418, Wr4ju6, vis_r10_o[23]);  // ../RTL/cortexm0ds_logic.v(15689)
  not u19063 (Q96pw6, n5418);  // ../RTL/cortexm0ds_logic.v(15689)
  and u19064 (n5419, Ds4ju6, vis_r9_o[23]);  // ../RTL/cortexm0ds_logic.v(15690)
  not u19065 (J96pw6, n5419);  // ../RTL/cortexm0ds_logic.v(15690)
  and u19066 (V86pw6, C80iu6, X96pw6);  // ../RTL/cortexm0ds_logic.v(15691)
  and u19067 (n5420, Rs4ju6, vis_r8_o[23]);  // ../RTL/cortexm0ds_logic.v(15692)
  not u19068 (X96pw6, n5420);  // ../RTL/cortexm0ds_logic.v(15692)
  and u19069 (C80iu6, Ea6pw6, La6pw6);  // ../RTL/cortexm0ds_logic.v(15693)
  and u1907 (n203, Iahpw6[21], Z4yhu6);  // ../RTL/cortexm0ds_logic.v(3768)
  and u19070 (La6pw6, Sa6pw6, Za6pw6);  // ../RTL/cortexm0ds_logic.v(15694)
  and u19071 (Za6pw6, Gb6pw6, Nb6pw6);  // ../RTL/cortexm0ds_logic.v(15695)
  and u19072 (n5421, V6now6, vis_r2_o[23]);  // ../RTL/cortexm0ds_logic.v(15696)
  not u19073 (Nb6pw6, n5421);  // ../RTL/cortexm0ds_logic.v(15696)
  and u19074 (n5422, C7now6, vis_r6_o[23]);  // ../RTL/cortexm0ds_logic.v(15697)
  not u19075 (Gb6pw6, n5422);  // ../RTL/cortexm0ds_logic.v(15697)
  and u19076 (Sa6pw6, Ub6pw6, Bc6pw6);  // ../RTL/cortexm0ds_logic.v(15698)
  and u19077 (n5423, X7now6, vis_r5_o[23]);  // ../RTL/cortexm0ds_logic.v(15699)
  not u19078 (Bc6pw6, n5423);  // ../RTL/cortexm0ds_logic.v(15699)
  and u19079 (n5424, E8now6, vis_r4_o[23]);  // ../RTL/cortexm0ds_logic.v(15700)
  not u1908 (Dh2iu6, n203);  // ../RTL/cortexm0ds_logic.v(3768)
  not u19080 (Ub6pw6, n5424);  // ../RTL/cortexm0ds_logic.v(15700)
  and u19081 (Ea6pw6, Ic6pw6, Pc6pw6);  // ../RTL/cortexm0ds_logic.v(15701)
  and u19082 (Pc6pw6, Wc6pw6, Dd6pw6);  // ../RTL/cortexm0ds_logic.v(15702)
  and u19083 (n5425, N9now6, vis_r1_o[23]);  // ../RTL/cortexm0ds_logic.v(15703)
  not u19084 (Dd6pw6, n5425);  // ../RTL/cortexm0ds_logic.v(15703)
  and u19085 (n5426, U9now6, vis_r0_o[23]);  // ../RTL/cortexm0ds_logic.v(15704)
  not u19086 (Wc6pw6, n5426);  // ../RTL/cortexm0ds_logic.v(15704)
  and u19087 (Ic6pw6, Kd6pw6, Rd6pw6);  // ../RTL/cortexm0ds_logic.v(15705)
  and u19088 (n5427, Panow6, vis_r3_o[23]);  // ../RTL/cortexm0ds_logic.v(15706)
  not u19089 (Rd6pw6, n5427);  // ../RTL/cortexm0ds_logic.v(15706)
  and u1909 (n204, Rh2iu6, Yh2iu6);  // ../RTL/cortexm0ds_logic.v(3769)
  and u19090 (n5428, Wanow6, vis_r7_o[23]);  // ../RTL/cortexm0ds_logic.v(15707)
  not u19091 (Kd6pw6, n5428);  // ../RTL/cortexm0ds_logic.v(15707)
  not u19092 (Ax9iu6, Fkfpw6[23]);  // ../RTL/cortexm0ds_logic.v(15708)
  and u19093 (I56pw6, Yd6pw6, Fe6pw6);  // ../RTL/cortexm0ds_logic.v(15709)
  and u19094 (n5429, N5fpw6[22], Sdaiu6);  // ../RTL/cortexm0ds_logic.v(15710)
  not u19095 (Fe6pw6, n5429);  // ../RTL/cortexm0ds_logic.v(15710)
  and u19096 (n5430, Eafpw6[23], A3iiu6);  // ../RTL/cortexm0ds_logic.v(15711)
  not u19097 (Yd6pw6, n5430);  // ../RTL/cortexm0ds_logic.v(15711)
  and u19098 (n5431, Me6pw6, Te6pw6);  // ../RTL/cortexm0ds_logic.v(15713)
  not u19099 (Fzdpw6, n5431);  // ../RTL/cortexm0ds_logic.v(15713)
  buf u191 (vis_apsr_o[0], X5ibx6);  // ../RTL/cortexm0ds_logic.v(1880)
  not u1910 (Bzxhu6, n204);  // ../RTL/cortexm0ds_logic.v(3769)
  or u19100 (Te6pw6, T2iiu6, Mk0iu6);  // ../RTL/cortexm0ds_logic.v(15714)
  AL_MUX u19101 (
    .i0(Suliu6),
    .i1(Af6pw6),
    .sel(Mm4ju6),
    .o(Mk0iu6));  // ../RTL/cortexm0ds_logic.v(15715)
  and u19102 (Af6pw6, Hf6pw6, Of6pw6);  // ../RTL/cortexm0ds_logic.v(15716)
  and u19103 (Of6pw6, Vf6pw6, Cg6pw6);  // ../RTL/cortexm0ds_logic.v(15717)
  and u19104 (Cg6pw6, Jg6pw6, Qg6pw6);  // ../RTL/cortexm0ds_logic.v(15718)
  and u19105 (n5432, Jo4ju6, vis_r14_o[22]);  // ../RTL/cortexm0ds_logic.v(15719)
  not u19106 (Qg6pw6, n5432);  // ../RTL/cortexm0ds_logic.v(15719)
  and u19107 (Jg6pw6, Xg6pw6, Eh6pw6);  // ../RTL/cortexm0ds_logic.v(15720)
  and u19108 (n5433, Ep4ju6, vis_psp_o[20]);  // ../RTL/cortexm0ds_logic.v(15721)
  not u19109 (Eh6pw6, n5433);  // ../RTL/cortexm0ds_logic.v(15721)
  and u1911 (Yh2iu6, Fi2iu6, L72iu6);  // ../RTL/cortexm0ds_logic.v(3770)
  and u19110 (n5434, Lp4ju6, vis_msp_o[20]);  // ../RTL/cortexm0ds_logic.v(15722)
  not u19111 (Xg6pw6, n5434);  // ../RTL/cortexm0ds_logic.v(15722)
  and u19112 (Vf6pw6, Lh6pw6, Sh6pw6);  // ../RTL/cortexm0ds_logic.v(15723)
  and u19113 (n5435, Gq4ju6, vis_r12_o[22]);  // ../RTL/cortexm0ds_logic.v(15724)
  not u19114 (Sh6pw6, n5435);  // ../RTL/cortexm0ds_logic.v(15724)
  and u19115 (n5436, Nq4ju6, vis_r11_o[22]);  // ../RTL/cortexm0ds_logic.v(15725)
  not u19116 (Lh6pw6, n5436);  // ../RTL/cortexm0ds_logic.v(15725)
  and u19117 (Hf6pw6, Zh6pw6, Gi6pw6);  // ../RTL/cortexm0ds_logic.v(15726)
  and u19118 (Gi6pw6, Ni6pw6, Ui6pw6);  // ../RTL/cortexm0ds_logic.v(15727)
  and u19119 (n5437, Wr4ju6, vis_r10_o[22]);  // ../RTL/cortexm0ds_logic.v(15728)
  and u1912 (n205, Uthpw6[20], Vk1iu6);  // ../RTL/cortexm0ds_logic.v(3771)
  not u19120 (Ui6pw6, n5437);  // ../RTL/cortexm0ds_logic.v(15728)
  and u19121 (n5438, Ds4ju6, vis_r9_o[22]);  // ../RTL/cortexm0ds_logic.v(15729)
  not u19122 (Ni6pw6, n5438);  // ../RTL/cortexm0ds_logic.v(15729)
  and u19123 (Zh6pw6, J80iu6, Bj6pw6);  // ../RTL/cortexm0ds_logic.v(15730)
  and u19124 (n5439, Rs4ju6, vis_r8_o[22]);  // ../RTL/cortexm0ds_logic.v(15731)
  not u19125 (Bj6pw6, n5439);  // ../RTL/cortexm0ds_logic.v(15731)
  and u19126 (J80iu6, Ij6pw6, Pj6pw6);  // ../RTL/cortexm0ds_logic.v(15732)
  and u19127 (Pj6pw6, Wj6pw6, Dk6pw6);  // ../RTL/cortexm0ds_logic.v(15733)
  and u19128 (Dk6pw6, Kk6pw6, Rk6pw6);  // ../RTL/cortexm0ds_logic.v(15734)
  and u19129 (n5440, V6now6, vis_r2_o[22]);  // ../RTL/cortexm0ds_logic.v(15735)
  not u1913 (Fi2iu6, n205);  // ../RTL/cortexm0ds_logic.v(3771)
  not u19130 (Rk6pw6, n5440);  // ../RTL/cortexm0ds_logic.v(15735)
  and u19131 (n5441, C7now6, vis_r6_o[22]);  // ../RTL/cortexm0ds_logic.v(15736)
  not u19132 (Kk6pw6, n5441);  // ../RTL/cortexm0ds_logic.v(15736)
  and u19133 (Wj6pw6, Yk6pw6, Fl6pw6);  // ../RTL/cortexm0ds_logic.v(15737)
  and u19134 (n5442, X7now6, vis_r5_o[22]);  // ../RTL/cortexm0ds_logic.v(15738)
  not u19135 (Fl6pw6, n5442);  // ../RTL/cortexm0ds_logic.v(15738)
  and u19136 (n5443, E8now6, vis_r4_o[22]);  // ../RTL/cortexm0ds_logic.v(15739)
  not u19137 (Yk6pw6, n5443);  // ../RTL/cortexm0ds_logic.v(15739)
  and u19138 (Ij6pw6, Ml6pw6, Tl6pw6);  // ../RTL/cortexm0ds_logic.v(15740)
  and u19139 (Tl6pw6, Am6pw6, Hm6pw6);  // ../RTL/cortexm0ds_logic.v(15741)
  and u1914 (Rh2iu6, Mi2iu6, Ti2iu6);  // ../RTL/cortexm0ds_logic.v(3772)
  and u19140 (n5444, N9now6, vis_r1_o[22]);  // ../RTL/cortexm0ds_logic.v(15742)
  not u19141 (Hm6pw6, n5444);  // ../RTL/cortexm0ds_logic.v(15742)
  and u19142 (n5445, U9now6, vis_r0_o[22]);  // ../RTL/cortexm0ds_logic.v(15743)
  not u19143 (Am6pw6, n5445);  // ../RTL/cortexm0ds_logic.v(15743)
  and u19144 (Ml6pw6, Om6pw6, Vm6pw6);  // ../RTL/cortexm0ds_logic.v(15744)
  and u19145 (n5446, Panow6, vis_r3_o[22]);  // ../RTL/cortexm0ds_logic.v(15745)
  not u19146 (Vm6pw6, n5446);  // ../RTL/cortexm0ds_logic.v(15745)
  and u19147 (n5447, Wanow6, vis_r7_o[22]);  // ../RTL/cortexm0ds_logic.v(15746)
  not u19148 (Om6pw6, n5447);  // ../RTL/cortexm0ds_logic.v(15746)
  not u19149 (Suliu6, Fkfpw6[22]);  // ../RTL/cortexm0ds_logic.v(15747)
  and u1915 (n206, Iahpw6[19], Xl1iu6);  // ../RTL/cortexm0ds_logic.v(3773)
  and u19150 (Me6pw6, Cn6pw6, Jn6pw6);  // ../RTL/cortexm0ds_logic.v(15748)
  and u19151 (n5448, N5fpw6[21], Sdaiu6);  // ../RTL/cortexm0ds_logic.v(15749)
  not u19152 (Jn6pw6, n5448);  // ../RTL/cortexm0ds_logic.v(15749)
  and u19153 (n5449, Eafpw6[22], A3iiu6);  // ../RTL/cortexm0ds_logic.v(15750)
  not u19154 (Cn6pw6, n5449);  // ../RTL/cortexm0ds_logic.v(15750)
  and u19155 (n5450, Qn6pw6, Xn6pw6);  // ../RTL/cortexm0ds_logic.v(15752)
  not u19156 (Yydpw6, n5450);  // ../RTL/cortexm0ds_logic.v(15752)
  or u19157 (Xn6pw6, T2iiu6, Tk0iu6);  // ../RTL/cortexm0ds_logic.v(15753)
  AL_MUX u19158 (
    .i0(Rxliu6),
    .i1(Eo6pw6),
    .sel(Mm4ju6),
    .o(Tk0iu6));  // ../RTL/cortexm0ds_logic.v(15754)
  and u19159 (Eo6pw6, Lo6pw6, So6pw6);  // ../RTL/cortexm0ds_logic.v(15755)
  not u1916 (Ti2iu6, n206);  // ../RTL/cortexm0ds_logic.v(3773)
  and u19160 (So6pw6, Zo6pw6, Gp6pw6);  // ../RTL/cortexm0ds_logic.v(15756)
  and u19161 (Gp6pw6, Np6pw6, Up6pw6);  // ../RTL/cortexm0ds_logic.v(15757)
  and u19162 (n5451, Jo4ju6, vis_r14_o[21]);  // ../RTL/cortexm0ds_logic.v(15758)
  not u19163 (Up6pw6, n5451);  // ../RTL/cortexm0ds_logic.v(15758)
  and u19164 (Np6pw6, Bq6pw6, Iq6pw6);  // ../RTL/cortexm0ds_logic.v(15759)
  and u19165 (n5452, Ep4ju6, vis_psp_o[19]);  // ../RTL/cortexm0ds_logic.v(15760)
  not u19166 (Iq6pw6, n5452);  // ../RTL/cortexm0ds_logic.v(15760)
  and u19167 (n5453, Lp4ju6, vis_msp_o[19]);  // ../RTL/cortexm0ds_logic.v(15761)
  not u19168 (Bq6pw6, n5453);  // ../RTL/cortexm0ds_logic.v(15761)
  and u19169 (Zo6pw6, Pq6pw6, Wq6pw6);  // ../RTL/cortexm0ds_logic.v(15762)
  and u1917 (n207, Iahpw6[20], Z4yhu6);  // ../RTL/cortexm0ds_logic.v(3774)
  and u19170 (n5454, Gq4ju6, vis_r12_o[21]);  // ../RTL/cortexm0ds_logic.v(15763)
  not u19171 (Wq6pw6, n5454);  // ../RTL/cortexm0ds_logic.v(15763)
  and u19172 (n5455, Nq4ju6, vis_r11_o[21]);  // ../RTL/cortexm0ds_logic.v(15764)
  not u19173 (Pq6pw6, n5455);  // ../RTL/cortexm0ds_logic.v(15764)
  and u19174 (Lo6pw6, Dr6pw6, Kr6pw6);  // ../RTL/cortexm0ds_logic.v(15765)
  and u19175 (Kr6pw6, Rr6pw6, Yr6pw6);  // ../RTL/cortexm0ds_logic.v(15766)
  and u19176 (n5456, Wr4ju6, vis_r10_o[21]);  // ../RTL/cortexm0ds_logic.v(15767)
  not u19177 (Yr6pw6, n5456);  // ../RTL/cortexm0ds_logic.v(15767)
  and u19178 (n5457, Ds4ju6, vis_r9_o[21]);  // ../RTL/cortexm0ds_logic.v(15768)
  not u19179 (Rr6pw6, n5457);  // ../RTL/cortexm0ds_logic.v(15768)
  not u1918 (Mi2iu6, n207);  // ../RTL/cortexm0ds_logic.v(3774)
  and u19180 (Dr6pw6, Q80iu6, Fs6pw6);  // ../RTL/cortexm0ds_logic.v(15769)
  and u19181 (n5458, Rs4ju6, vis_r8_o[21]);  // ../RTL/cortexm0ds_logic.v(15770)
  not u19182 (Fs6pw6, n5458);  // ../RTL/cortexm0ds_logic.v(15770)
  and u19183 (Q80iu6, Ms6pw6, Ts6pw6);  // ../RTL/cortexm0ds_logic.v(15771)
  and u19184 (Ts6pw6, At6pw6, Ht6pw6);  // ../RTL/cortexm0ds_logic.v(15772)
  and u19185 (Ht6pw6, Ot6pw6, Vt6pw6);  // ../RTL/cortexm0ds_logic.v(15773)
  and u19186 (n5459, V6now6, vis_r2_o[21]);  // ../RTL/cortexm0ds_logic.v(15774)
  not u19187 (Vt6pw6, n5459);  // ../RTL/cortexm0ds_logic.v(15774)
  and u19188 (n5460, C7now6, vis_r6_o[21]);  // ../RTL/cortexm0ds_logic.v(15775)
  not u19189 (Ot6pw6, n5460);  // ../RTL/cortexm0ds_logic.v(15775)
  and u1919 (n208, Aj2iu6, Hj2iu6);  // ../RTL/cortexm0ds_logic.v(3775)
  and u19190 (At6pw6, Cu6pw6, Ju6pw6);  // ../RTL/cortexm0ds_logic.v(15776)
  and u19191 (n5461, X7now6, vis_r5_o[21]);  // ../RTL/cortexm0ds_logic.v(15777)
  not u19192 (Ju6pw6, n5461);  // ../RTL/cortexm0ds_logic.v(15777)
  and u19193 (n5462, E8now6, vis_r4_o[21]);  // ../RTL/cortexm0ds_logic.v(15778)
  not u19194 (Cu6pw6, n5462);  // ../RTL/cortexm0ds_logic.v(15778)
  and u19195 (Ms6pw6, Qu6pw6, Xu6pw6);  // ../RTL/cortexm0ds_logic.v(15779)
  and u19196 (Xu6pw6, Ev6pw6, Lv6pw6);  // ../RTL/cortexm0ds_logic.v(15780)
  and u19197 (n5463, N9now6, vis_r1_o[21]);  // ../RTL/cortexm0ds_logic.v(15781)
  not u19198 (Lv6pw6, n5463);  // ../RTL/cortexm0ds_logic.v(15781)
  and u19199 (n5464, U9now6, vis_r0_o[21]);  // ../RTL/cortexm0ds_logic.v(15782)
  buf u192 (vis_r4_o[5], Zduax6);  // ../RTL/cortexm0ds_logic.v(2626)
  not u1920 (Uyxhu6, n208);  // ../RTL/cortexm0ds_logic.v(3775)
  not u19200 (Ev6pw6, n5464);  // ../RTL/cortexm0ds_logic.v(15782)
  and u19201 (Qu6pw6, Sv6pw6, Zv6pw6);  // ../RTL/cortexm0ds_logic.v(15783)
  and u19202 (n5465, Panow6, vis_r3_o[21]);  // ../RTL/cortexm0ds_logic.v(15784)
  not u19203 (Zv6pw6, n5465);  // ../RTL/cortexm0ds_logic.v(15784)
  and u19204 (n5466, Wanow6, vis_r7_o[21]);  // ../RTL/cortexm0ds_logic.v(15785)
  not u19205 (Sv6pw6, n5466);  // ../RTL/cortexm0ds_logic.v(15785)
  not u19206 (Rxliu6, Fkfpw6[21]);  // ../RTL/cortexm0ds_logic.v(15786)
  and u19207 (Qn6pw6, Gw6pw6, Nw6pw6);  // ../RTL/cortexm0ds_logic.v(15787)
  and u19208 (n5467, N5fpw6[20], Sdaiu6);  // ../RTL/cortexm0ds_logic.v(15788)
  not u19209 (Nw6pw6, n5467);  // ../RTL/cortexm0ds_logic.v(15788)
  and u1921 (n209, Iahpw6[19], Z4yhu6);  // ../RTL/cortexm0ds_logic.v(3776)
  and u19210 (n5468, Eafpw6[21], A3iiu6);  // ../RTL/cortexm0ds_logic.v(15789)
  not u19211 (Gw6pw6, n5468);  // ../RTL/cortexm0ds_logic.v(15789)
  and u19212 (n5469, Uw6pw6, Bx6pw6);  // ../RTL/cortexm0ds_logic.v(15791)
  not u19213 (Rydpw6, n5469);  // ../RTL/cortexm0ds_logic.v(15791)
  or u19214 (Bx6pw6, T2iiu6, Al0iu6);  // ../RTL/cortexm0ds_logic.v(15792)
  AL_MUX u19215 (
    .i0(X0miu6),
    .i1(Ix6pw6),
    .sel(Mm4ju6),
    .o(Al0iu6));  // ../RTL/cortexm0ds_logic.v(15793)
  and u19216 (Ix6pw6, Px6pw6, Wx6pw6);  // ../RTL/cortexm0ds_logic.v(15794)
  and u19217 (Wx6pw6, Dy6pw6, Ky6pw6);  // ../RTL/cortexm0ds_logic.v(15795)
  and u19218 (Ky6pw6, Ry6pw6, Yy6pw6);  // ../RTL/cortexm0ds_logic.v(15796)
  and u19219 (n5470, Jo4ju6, vis_r14_o[20]);  // ../RTL/cortexm0ds_logic.v(15797)
  not u1922 (Hj2iu6, n209);  // ../RTL/cortexm0ds_logic.v(3776)
  not u19220 (Yy6pw6, n5470);  // ../RTL/cortexm0ds_logic.v(15797)
  and u19221 (Ry6pw6, Fz6pw6, Mz6pw6);  // ../RTL/cortexm0ds_logic.v(15798)
  and u19222 (n5471, Ep4ju6, vis_psp_o[18]);  // ../RTL/cortexm0ds_logic.v(15799)
  not u19223 (Mz6pw6, n5471);  // ../RTL/cortexm0ds_logic.v(15799)
  and u19224 (n5472, Lp4ju6, vis_msp_o[18]);  // ../RTL/cortexm0ds_logic.v(15800)
  not u19225 (Fz6pw6, n5472);  // ../RTL/cortexm0ds_logic.v(15800)
  and u19226 (Dy6pw6, Tz6pw6, A07pw6);  // ../RTL/cortexm0ds_logic.v(15801)
  and u19227 (n5473, Gq4ju6, vis_r12_o[20]);  // ../RTL/cortexm0ds_logic.v(15802)
  not u19228 (A07pw6, n5473);  // ../RTL/cortexm0ds_logic.v(15802)
  and u19229 (n5474, Nq4ju6, vis_r11_o[20]);  // ../RTL/cortexm0ds_logic.v(15803)
  and u1923 (Aj2iu6, Oj2iu6, Vj2iu6);  // ../RTL/cortexm0ds_logic.v(3777)
  not u19230 (Tz6pw6, n5474);  // ../RTL/cortexm0ds_logic.v(15803)
  and u19231 (Px6pw6, H07pw6, O07pw6);  // ../RTL/cortexm0ds_logic.v(15804)
  and u19232 (O07pw6, V07pw6, C17pw6);  // ../RTL/cortexm0ds_logic.v(15805)
  and u19233 (n5475, Wr4ju6, vis_r10_o[20]);  // ../RTL/cortexm0ds_logic.v(15806)
  not u19234 (C17pw6, n5475);  // ../RTL/cortexm0ds_logic.v(15806)
  and u19235 (n5476, Ds4ju6, vis_r9_o[20]);  // ../RTL/cortexm0ds_logic.v(15807)
  not u19236 (V07pw6, n5476);  // ../RTL/cortexm0ds_logic.v(15807)
  and u19237 (H07pw6, X80iu6, J17pw6);  // ../RTL/cortexm0ds_logic.v(15808)
  and u19238 (n5477, Rs4ju6, vis_r8_o[20]);  // ../RTL/cortexm0ds_logic.v(15809)
  not u19239 (J17pw6, n5477);  // ../RTL/cortexm0ds_logic.v(15809)
  and u1924 (n210, Uthpw6[19], Vk1iu6);  // ../RTL/cortexm0ds_logic.v(3778)
  and u19240 (X80iu6, Q17pw6, X17pw6);  // ../RTL/cortexm0ds_logic.v(15810)
  and u19241 (X17pw6, E27pw6, L27pw6);  // ../RTL/cortexm0ds_logic.v(15811)
  and u19242 (L27pw6, S27pw6, Z27pw6);  // ../RTL/cortexm0ds_logic.v(15812)
  and u19243 (n5478, V6now6, vis_r2_o[20]);  // ../RTL/cortexm0ds_logic.v(15813)
  not u19244 (Z27pw6, n5478);  // ../RTL/cortexm0ds_logic.v(15813)
  and u19245 (n5479, C7now6, vis_r6_o[20]);  // ../RTL/cortexm0ds_logic.v(15814)
  not u19246 (S27pw6, n5479);  // ../RTL/cortexm0ds_logic.v(15814)
  and u19247 (E27pw6, G37pw6, N37pw6);  // ../RTL/cortexm0ds_logic.v(15815)
  and u19248 (n5480, X7now6, vis_r5_o[20]);  // ../RTL/cortexm0ds_logic.v(15816)
  not u19249 (N37pw6, n5480);  // ../RTL/cortexm0ds_logic.v(15816)
  not u1925 (Vj2iu6, n210);  // ../RTL/cortexm0ds_logic.v(3778)
  and u19250 (n5481, E8now6, vis_r4_o[20]);  // ../RTL/cortexm0ds_logic.v(15817)
  not u19251 (G37pw6, n5481);  // ../RTL/cortexm0ds_logic.v(15817)
  and u19252 (Q17pw6, U37pw6, B47pw6);  // ../RTL/cortexm0ds_logic.v(15818)
  and u19253 (B47pw6, I47pw6, P47pw6);  // ../RTL/cortexm0ds_logic.v(15819)
  and u19254 (n5482, N9now6, vis_r1_o[20]);  // ../RTL/cortexm0ds_logic.v(15820)
  not u19255 (P47pw6, n5482);  // ../RTL/cortexm0ds_logic.v(15820)
  and u19256 (n5483, U9now6, vis_r0_o[20]);  // ../RTL/cortexm0ds_logic.v(15821)
  not u19257 (I47pw6, n5483);  // ../RTL/cortexm0ds_logic.v(15821)
  and u19258 (U37pw6, W47pw6, D57pw6);  // ../RTL/cortexm0ds_logic.v(15822)
  and u19259 (n5484, Panow6, vis_r3_o[20]);  // ../RTL/cortexm0ds_logic.v(15823)
  and u1926 (n211, Iahpw6[18], Xl1iu6);  // ../RTL/cortexm0ds_logic.v(3779)
  not u19260 (D57pw6, n5484);  // ../RTL/cortexm0ds_logic.v(15823)
  and u19261 (n5485, Wanow6, vis_r7_o[20]);  // ../RTL/cortexm0ds_logic.v(15824)
  not u19262 (W47pw6, n5485);  // ../RTL/cortexm0ds_logic.v(15824)
  not u19263 (X0miu6, Fkfpw6[20]);  // ../RTL/cortexm0ds_logic.v(15825)
  and u19264 (Uw6pw6, K57pw6, R57pw6);  // ../RTL/cortexm0ds_logic.v(15826)
  and u19265 (n5486, N5fpw6[19], Sdaiu6);  // ../RTL/cortexm0ds_logic.v(15827)
  not u19266 (R57pw6, n5486);  // ../RTL/cortexm0ds_logic.v(15827)
  and u19267 (n5487, Eafpw6[20], A3iiu6);  // ../RTL/cortexm0ds_logic.v(15828)
  not u19268 (K57pw6, n5487);  // ../RTL/cortexm0ds_logic.v(15828)
  not u19269 (HADDR[0], n5488[0]);  // ../RTL/cortexm0ds_logic.v(15829)
  not u1927 (Oj2iu6, n211);  // ../RTL/cortexm0ds_logic.v(3779)
  buf u19270 (HBURST[0], 1'b0);  // ../RTL/cortexm0ds_logic.v(1725)
  and u19271 (n5489, M67pw6, Ne3pw6);  // ../RTL/cortexm0ds_logic.v(15830)
  not u19272 (F67pw6, n5489);  // ../RTL/cortexm0ds_logic.v(15830)
  and u19273 (M67pw6, Tnhpw6[1], T67pw6);  // ../RTL/cortexm0ds_logic.v(15831)
  not u19274 (T67pw6, Aphpw6[2]);  // ../RTL/cortexm0ds_logic.v(15832)
  and u19275 (n5490, Hz0iu6, Ze9iu6);  // ../RTL/cortexm0ds_logic.v(15833)
  not u19276 (Y57pw6, n5490);  // ../RTL/cortexm0ds_logic.v(15833)
  and u19277 (Hz0iu6, A77pw6, Ed3pw6);  // ../RTL/cortexm0ds_logic.v(15834)
  and u19278 (A77pw6, Iiliu6, Ob3pw6);  // ../RTL/cortexm0ds_logic.v(15835)
  and u19279 (n5491, H77pw6, O77pw6);  // ../RTL/cortexm0ds_logic.v(15836)
  and u1928 (n212, Ck2iu6, Jk2iu6);  // ../RTL/cortexm0ds_logic.v(3780)
  not u19280 (Iiliu6, n5491);  // ../RTL/cortexm0ds_logic.v(15836)
  or u19281 (O77pw6, T2iiu6, Hl0iu6);  // ../RTL/cortexm0ds_logic.v(15837)
  AL_MUX u19282 (
    .i0(Rjliu6),
    .i1(V77pw6),
    .sel(Mm4ju6),
    .o(Hl0iu6));  // ../RTL/cortexm0ds_logic.v(15838)
  and u19283 (V77pw6, C87pw6, J87pw6);  // ../RTL/cortexm0ds_logic.v(15839)
  and u19284 (J87pw6, Q87pw6, X87pw6);  // ../RTL/cortexm0ds_logic.v(15840)
  and u19285 (X87pw6, E97pw6, L97pw6);  // ../RTL/cortexm0ds_logic.v(15841)
  and u19286 (n5492, Jo4ju6, vis_r14_o[1]);  // ../RTL/cortexm0ds_logic.v(15842)
  not u19287 (L97pw6, n5492);  // ../RTL/cortexm0ds_logic.v(15842)
  and u19288 (n5493, Gq4ju6, vis_r12_o[1]);  // ../RTL/cortexm0ds_logic.v(15843)
  not u19289 (E97pw6, n5493);  // ../RTL/cortexm0ds_logic.v(15843)
  not u1929 (Nyxhu6, n212);  // ../RTL/cortexm0ds_logic.v(3780)
  and u19290 (Q87pw6, S97pw6, Z97pw6);  // ../RTL/cortexm0ds_logic.v(15844)
  and u19291 (n5494, Nq4ju6, vis_r11_o[1]);  // ../RTL/cortexm0ds_logic.v(15845)
  not u19292 (Z97pw6, n5494);  // ../RTL/cortexm0ds_logic.v(15845)
  and u19293 (n5495, Wr4ju6, vis_r10_o[1]);  // ../RTL/cortexm0ds_logic.v(15846)
  not u19294 (S97pw6, n5495);  // ../RTL/cortexm0ds_logic.v(15846)
  and u19295 (C87pw6, Ga7pw6, E90iu6);  // ../RTL/cortexm0ds_logic.v(15847)
  and u19296 (E90iu6, Na7pw6, Ua7pw6);  // ../RTL/cortexm0ds_logic.v(15848)
  and u19297 (Ua7pw6, Bb7pw6, Ib7pw6);  // ../RTL/cortexm0ds_logic.v(15849)
  and u19298 (Ib7pw6, Pb7pw6, Wb7pw6);  // ../RTL/cortexm0ds_logic.v(15850)
  and u19299 (n5496, V6now6, vis_r2_o[1]);  // ../RTL/cortexm0ds_logic.v(15851)
  buf u193 (vis_r14_o[2], Uvmax6);  // ../RTL/cortexm0ds_logic.v(2497)
  and u1930 (n213, Iahpw6[18], Z4yhu6);  // ../RTL/cortexm0ds_logic.v(3781)
  not u19300 (Wb7pw6, n5496);  // ../RTL/cortexm0ds_logic.v(15851)
  and u19301 (n5497, C7now6, vis_r6_o[1]);  // ../RTL/cortexm0ds_logic.v(15852)
  not u19302 (Pb7pw6, n5497);  // ../RTL/cortexm0ds_logic.v(15852)
  and u19303 (Bb7pw6, Dc7pw6, Kc7pw6);  // ../RTL/cortexm0ds_logic.v(15853)
  and u19304 (n5498, X7now6, vis_r5_o[1]);  // ../RTL/cortexm0ds_logic.v(15854)
  not u19305 (Kc7pw6, n5498);  // ../RTL/cortexm0ds_logic.v(15854)
  and u19306 (n5499, E8now6, vis_r4_o[1]);  // ../RTL/cortexm0ds_logic.v(15855)
  not u19307 (Dc7pw6, n5499);  // ../RTL/cortexm0ds_logic.v(15855)
  and u19308 (Na7pw6, Rc7pw6, Yc7pw6);  // ../RTL/cortexm0ds_logic.v(15856)
  and u19309 (Yc7pw6, Fd7pw6, Md7pw6);  // ../RTL/cortexm0ds_logic.v(15857)
  not u1931 (Jk2iu6, n213);  // ../RTL/cortexm0ds_logic.v(3781)
  and u19310 (n5500, N9now6, vis_r1_o[1]);  // ../RTL/cortexm0ds_logic.v(15858)
  not u19311 (Md7pw6, n5500);  // ../RTL/cortexm0ds_logic.v(15858)
  and u19312 (n5501, U9now6, vis_r0_o[1]);  // ../RTL/cortexm0ds_logic.v(15859)
  not u19313 (Fd7pw6, n5501);  // ../RTL/cortexm0ds_logic.v(15859)
  and u19314 (Rc7pw6, Td7pw6, Ae7pw6);  // ../RTL/cortexm0ds_logic.v(15860)
  and u19315 (n5502, Panow6, vis_r3_o[1]);  // ../RTL/cortexm0ds_logic.v(15861)
  not u19316 (Ae7pw6, n5502);  // ../RTL/cortexm0ds_logic.v(15861)
  and u19317 (n5503, Wanow6, vis_r7_o[1]);  // ../RTL/cortexm0ds_logic.v(15862)
  not u19318 (Td7pw6, n5503);  // ../RTL/cortexm0ds_logic.v(15862)
  and u19319 (Ga7pw6, He7pw6, Oe7pw6);  // ../RTL/cortexm0ds_logic.v(15863)
  and u1932 (Ck2iu6, Qk2iu6, Xk2iu6);  // ../RTL/cortexm0ds_logic.v(3782)
  and u19320 (n5504, Ds4ju6, vis_r9_o[1]);  // ../RTL/cortexm0ds_logic.v(15864)
  not u19321 (Oe7pw6, n5504);  // ../RTL/cortexm0ds_logic.v(15864)
  and u19322 (n5505, Rs4ju6, vis_r8_o[1]);  // ../RTL/cortexm0ds_logic.v(15865)
  not u19323 (He7pw6, n5505);  // ../RTL/cortexm0ds_logic.v(15865)
  not u19324 (Rjliu6, Fkfpw6[1]);  // ../RTL/cortexm0ds_logic.v(15866)
  and u19325 (H77pw6, Ve7pw6, Cf7pw6);  // ../RTL/cortexm0ds_logic.v(15867)
  and u19326 (n5506, Jf7pw6, Sdaiu6);  // ../RTL/cortexm0ds_logic.v(15868)
  not u19327 (Cf7pw6, n5506);  // ../RTL/cortexm0ds_logic.v(15868)
  or u19328 (n5507, Qf7pw6, Vtzhu6);  // ../RTL/cortexm0ds_logic.v(15869)
  not u19329 (Jf7pw6, n5507);  // ../RTL/cortexm0ds_logic.v(15869)
  and u1933 (n214, Uthpw6[18], Vk1iu6);  // ../RTL/cortexm0ds_logic.v(3783)
  and u19330 (Vtzhu6, Pkciu6, vis_pc_o[0]);  // ../RTL/cortexm0ds_logic.v(15870)
  or u19331 (n5508, Pkciu6, vis_pc_o[0]);  // ../RTL/cortexm0ds_logic.v(15871)
  not u19332 (Qf7pw6, n5508);  // ../RTL/cortexm0ds_logic.v(15871)
  and u19333 (n5509, Eafpw6[1], A3iiu6);  // ../RTL/cortexm0ds_logic.v(15872)
  not u19334 (Ve7pw6, n5509);  // ../RTL/cortexm0ds_logic.v(15872)
  and u19335 (n5510, Xf7pw6, Eg7pw6);  // ../RTL/cortexm0ds_logic.v(15874)
  not u19336 (Kydpw6, n5510);  // ../RTL/cortexm0ds_logic.v(15874)
  or u19337 (Eg7pw6, T2iiu6, Ol0iu6);  // ../RTL/cortexm0ds_logic.v(15875)
  AL_MUX u19338 (
    .i0(W3miu6),
    .i1(Lg7pw6),
    .sel(Mm4ju6),
    .o(Ol0iu6));  // ../RTL/cortexm0ds_logic.v(15876)
  and u19339 (Lg7pw6, Sg7pw6, Zg7pw6);  // ../RTL/cortexm0ds_logic.v(15877)
  not u1934 (Xk2iu6, n214);  // ../RTL/cortexm0ds_logic.v(3783)
  and u19340 (Zg7pw6, Gh7pw6, Nh7pw6);  // ../RTL/cortexm0ds_logic.v(15878)
  and u19341 (Nh7pw6, Uh7pw6, Bi7pw6);  // ../RTL/cortexm0ds_logic.v(15879)
  and u19342 (n5511, Jo4ju6, vis_r14_o[19]);  // ../RTL/cortexm0ds_logic.v(15880)
  not u19343 (Bi7pw6, n5511);  // ../RTL/cortexm0ds_logic.v(15880)
  and u19344 (Uh7pw6, Ii7pw6, Pi7pw6);  // ../RTL/cortexm0ds_logic.v(15881)
  and u19345 (n5512, Ep4ju6, vis_psp_o[17]);  // ../RTL/cortexm0ds_logic.v(15882)
  not u19346 (Pi7pw6, n5512);  // ../RTL/cortexm0ds_logic.v(15882)
  and u19347 (n5513, Lp4ju6, vis_msp_o[17]);  // ../RTL/cortexm0ds_logic.v(15883)
  not u19348 (Ii7pw6, n5513);  // ../RTL/cortexm0ds_logic.v(15883)
  and u19349 (Gh7pw6, Wi7pw6, Dj7pw6);  // ../RTL/cortexm0ds_logic.v(15884)
  and u1935 (n215, Iahpw6[17], Xl1iu6);  // ../RTL/cortexm0ds_logic.v(3784)
  and u19350 (n5514, Gq4ju6, vis_r12_o[19]);  // ../RTL/cortexm0ds_logic.v(15885)
  not u19351 (Dj7pw6, n5514);  // ../RTL/cortexm0ds_logic.v(15885)
  and u19352 (n5515, Nq4ju6, vis_r11_o[19]);  // ../RTL/cortexm0ds_logic.v(15886)
  not u19353 (Wi7pw6, n5515);  // ../RTL/cortexm0ds_logic.v(15886)
  and u19354 (Sg7pw6, Kj7pw6, Rj7pw6);  // ../RTL/cortexm0ds_logic.v(15887)
  and u19355 (Rj7pw6, Yj7pw6, Fk7pw6);  // ../RTL/cortexm0ds_logic.v(15888)
  and u19356 (n5516, Wr4ju6, vis_r10_o[19]);  // ../RTL/cortexm0ds_logic.v(15889)
  not u19357 (Fk7pw6, n5516);  // ../RTL/cortexm0ds_logic.v(15889)
  and u19358 (n5517, Ds4ju6, vis_r9_o[19]);  // ../RTL/cortexm0ds_logic.v(15890)
  not u19359 (Yj7pw6, n5517);  // ../RTL/cortexm0ds_logic.v(15890)
  not u1936 (Qk2iu6, n215);  // ../RTL/cortexm0ds_logic.v(3784)
  and u19360 (Kj7pw6, L90iu6, Mk7pw6);  // ../RTL/cortexm0ds_logic.v(15891)
  and u19361 (n5518, Rs4ju6, vis_r8_o[19]);  // ../RTL/cortexm0ds_logic.v(15892)
  not u19362 (Mk7pw6, n5518);  // ../RTL/cortexm0ds_logic.v(15892)
  and u19363 (L90iu6, Tk7pw6, Al7pw6);  // ../RTL/cortexm0ds_logic.v(15893)
  and u19364 (Al7pw6, Hl7pw6, Ol7pw6);  // ../RTL/cortexm0ds_logic.v(15894)
  and u19365 (Ol7pw6, Vl7pw6, Cm7pw6);  // ../RTL/cortexm0ds_logic.v(15895)
  and u19366 (n5519, V6now6, vis_r2_o[19]);  // ../RTL/cortexm0ds_logic.v(15896)
  not u19367 (Cm7pw6, n5519);  // ../RTL/cortexm0ds_logic.v(15896)
  and u19368 (n5520, C7now6, vis_r6_o[19]);  // ../RTL/cortexm0ds_logic.v(15897)
  not u19369 (Vl7pw6, n5520);  // ../RTL/cortexm0ds_logic.v(15897)
  and u1937 (n216, El2iu6, Ll2iu6);  // ../RTL/cortexm0ds_logic.v(3785)
  and u19370 (Hl7pw6, Jm7pw6, Qm7pw6);  // ../RTL/cortexm0ds_logic.v(15898)
  and u19371 (n5521, X7now6, vis_r5_o[19]);  // ../RTL/cortexm0ds_logic.v(15899)
  not u19372 (Qm7pw6, n5521);  // ../RTL/cortexm0ds_logic.v(15899)
  and u19373 (n5522, E8now6, vis_r4_o[19]);  // ../RTL/cortexm0ds_logic.v(15900)
  not u19374 (Jm7pw6, n5522);  // ../RTL/cortexm0ds_logic.v(15900)
  and u19375 (Tk7pw6, Xm7pw6, En7pw6);  // ../RTL/cortexm0ds_logic.v(15901)
  and u19376 (En7pw6, Ln7pw6, Sn7pw6);  // ../RTL/cortexm0ds_logic.v(15902)
  and u19377 (n5523, N9now6, vis_r1_o[19]);  // ../RTL/cortexm0ds_logic.v(15903)
  not u19378 (Sn7pw6, n5523);  // ../RTL/cortexm0ds_logic.v(15903)
  and u19379 (n5524, U9now6, vis_r0_o[19]);  // ../RTL/cortexm0ds_logic.v(15904)
  not u1938 (Gyxhu6, n216);  // ../RTL/cortexm0ds_logic.v(3785)
  not u19380 (Ln7pw6, n5524);  // ../RTL/cortexm0ds_logic.v(15904)
  and u19381 (Xm7pw6, Zn7pw6, Go7pw6);  // ../RTL/cortexm0ds_logic.v(15905)
  and u19382 (n5525, Panow6, vis_r3_o[19]);  // ../RTL/cortexm0ds_logic.v(15906)
  not u19383 (Go7pw6, n5525);  // ../RTL/cortexm0ds_logic.v(15906)
  and u19384 (n5526, Wanow6, vis_r7_o[19]);  // ../RTL/cortexm0ds_logic.v(15907)
  not u19385 (Zn7pw6, n5526);  // ../RTL/cortexm0ds_logic.v(15907)
  not u19386 (W3miu6, Fkfpw6[19]);  // ../RTL/cortexm0ds_logic.v(15908)
  and u19387 (Xf7pw6, No7pw6, Uo7pw6);  // ../RTL/cortexm0ds_logic.v(15909)
  and u19388 (n5527, N5fpw6[18], Sdaiu6);  // ../RTL/cortexm0ds_logic.v(15910)
  not u19389 (Uo7pw6, n5527);  // ../RTL/cortexm0ds_logic.v(15910)
  and u1939 (n217, Iahpw6[17], Z4yhu6);  // ../RTL/cortexm0ds_logic.v(3786)
  and u19390 (n5528, Eafpw6[19], A3iiu6);  // ../RTL/cortexm0ds_logic.v(15911)
  not u19391 (No7pw6, n5528);  // ../RTL/cortexm0ds_logic.v(15911)
  and u19392 (n5529, Bp7pw6, Ip7pw6);  // ../RTL/cortexm0ds_logic.v(15913)
  not u19393 (Dydpw6, n5529);  // ../RTL/cortexm0ds_logic.v(15913)
  or u19394 (Ip7pw6, T2iiu6, Vl0iu6);  // ../RTL/cortexm0ds_logic.v(15914)
  AL_MUX u19395 (
    .i0(V6miu6),
    .i1(Pp7pw6),
    .sel(Mm4ju6),
    .o(Vl0iu6));  // ../RTL/cortexm0ds_logic.v(15915)
  and u19396 (Pp7pw6, Wp7pw6, Dq7pw6);  // ../RTL/cortexm0ds_logic.v(15916)
  and u19397 (Dq7pw6, Kq7pw6, Rq7pw6);  // ../RTL/cortexm0ds_logic.v(15917)
  and u19398 (Rq7pw6, Yq7pw6, Fr7pw6);  // ../RTL/cortexm0ds_logic.v(15918)
  and u19399 (n5530, Jo4ju6, vis_r14_o[18]);  // ../RTL/cortexm0ds_logic.v(15919)
  buf u194 (vis_r8_o[11], Ca7bx6);  // ../RTL/cortexm0ds_logic.v(2579)
  not u1940 (Ll2iu6, n217);  // ../RTL/cortexm0ds_logic.v(3786)
  not u19400 (Fr7pw6, n5530);  // ../RTL/cortexm0ds_logic.v(15919)
  and u19401 (Yq7pw6, Mr7pw6, Tr7pw6);  // ../RTL/cortexm0ds_logic.v(15920)
  and u19402 (n5531, Ep4ju6, vis_psp_o[16]);  // ../RTL/cortexm0ds_logic.v(15921)
  not u19403 (Tr7pw6, n5531);  // ../RTL/cortexm0ds_logic.v(15921)
  and u19404 (n5532, Lp4ju6, vis_msp_o[16]);  // ../RTL/cortexm0ds_logic.v(15922)
  not u19405 (Mr7pw6, n5532);  // ../RTL/cortexm0ds_logic.v(15922)
  and u19406 (Kq7pw6, As7pw6, Hs7pw6);  // ../RTL/cortexm0ds_logic.v(15923)
  and u19407 (n5533, Gq4ju6, vis_r12_o[18]);  // ../RTL/cortexm0ds_logic.v(15924)
  not u19408 (Hs7pw6, n5533);  // ../RTL/cortexm0ds_logic.v(15924)
  and u19409 (n5534, Nq4ju6, vis_r11_o[18]);  // ../RTL/cortexm0ds_logic.v(15925)
  and u1941 (El2iu6, Sl2iu6, Zl2iu6);  // ../RTL/cortexm0ds_logic.v(3787)
  not u19410 (As7pw6, n5534);  // ../RTL/cortexm0ds_logic.v(15925)
  and u19411 (Wp7pw6, Os7pw6, Vs7pw6);  // ../RTL/cortexm0ds_logic.v(15926)
  and u19412 (Vs7pw6, Ct7pw6, Jt7pw6);  // ../RTL/cortexm0ds_logic.v(15927)
  and u19413 (n5535, Wr4ju6, vis_r10_o[18]);  // ../RTL/cortexm0ds_logic.v(15928)
  not u19414 (Jt7pw6, n5535);  // ../RTL/cortexm0ds_logic.v(15928)
  and u19415 (n5536, Ds4ju6, vis_r9_o[18]);  // ../RTL/cortexm0ds_logic.v(15929)
  not u19416 (Ct7pw6, n5536);  // ../RTL/cortexm0ds_logic.v(15929)
  and u19417 (Os7pw6, S90iu6, Qt7pw6);  // ../RTL/cortexm0ds_logic.v(15930)
  and u19418 (n5537, Rs4ju6, vis_r8_o[18]);  // ../RTL/cortexm0ds_logic.v(15931)
  not u19419 (Qt7pw6, n5537);  // ../RTL/cortexm0ds_logic.v(15931)
  and u1942 (n218, Uthpw6[17], Vk1iu6);  // ../RTL/cortexm0ds_logic.v(3788)
  and u19420 (S90iu6, Xt7pw6, Eu7pw6);  // ../RTL/cortexm0ds_logic.v(15932)
  and u19421 (Eu7pw6, Lu7pw6, Su7pw6);  // ../RTL/cortexm0ds_logic.v(15933)
  and u19422 (Su7pw6, Zu7pw6, Gv7pw6);  // ../RTL/cortexm0ds_logic.v(15934)
  and u19423 (n5538, V6now6, vis_r2_o[18]);  // ../RTL/cortexm0ds_logic.v(15935)
  not u19424 (Gv7pw6, n5538);  // ../RTL/cortexm0ds_logic.v(15935)
  and u19425 (n5539, C7now6, vis_r6_o[18]);  // ../RTL/cortexm0ds_logic.v(15936)
  not u19426 (Zu7pw6, n5539);  // ../RTL/cortexm0ds_logic.v(15936)
  and u19427 (Lu7pw6, Nv7pw6, Uv7pw6);  // ../RTL/cortexm0ds_logic.v(15937)
  and u19428 (n5540, X7now6, vis_r5_o[18]);  // ../RTL/cortexm0ds_logic.v(15938)
  not u19429 (Uv7pw6, n5540);  // ../RTL/cortexm0ds_logic.v(15938)
  not u1943 (Zl2iu6, n218);  // ../RTL/cortexm0ds_logic.v(3788)
  and u19430 (n5541, E8now6, vis_r4_o[18]);  // ../RTL/cortexm0ds_logic.v(15939)
  not u19431 (Nv7pw6, n5541);  // ../RTL/cortexm0ds_logic.v(15939)
  and u19432 (Xt7pw6, Bw7pw6, Iw7pw6);  // ../RTL/cortexm0ds_logic.v(15940)
  and u19433 (Iw7pw6, Pw7pw6, Ww7pw6);  // ../RTL/cortexm0ds_logic.v(15941)
  and u19434 (n5542, N9now6, vis_r1_o[18]);  // ../RTL/cortexm0ds_logic.v(15942)
  not u19435 (Ww7pw6, n5542);  // ../RTL/cortexm0ds_logic.v(15942)
  and u19436 (n5543, U9now6, vis_r0_o[18]);  // ../RTL/cortexm0ds_logic.v(15943)
  not u19437 (Pw7pw6, n5543);  // ../RTL/cortexm0ds_logic.v(15943)
  and u19438 (Bw7pw6, Dx7pw6, Kx7pw6);  // ../RTL/cortexm0ds_logic.v(15944)
  and u19439 (n5544, Panow6, vis_r3_o[18]);  // ../RTL/cortexm0ds_logic.v(15945)
  and u1944 (n219, Iahpw6[16], Xl1iu6);  // ../RTL/cortexm0ds_logic.v(3789)
  not u19440 (Kx7pw6, n5544);  // ../RTL/cortexm0ds_logic.v(15945)
  and u19441 (n5545, Wanow6, vis_r7_o[18]);  // ../RTL/cortexm0ds_logic.v(15946)
  not u19442 (Dx7pw6, n5545);  // ../RTL/cortexm0ds_logic.v(15946)
  not u19443 (V6miu6, Fkfpw6[18]);  // ../RTL/cortexm0ds_logic.v(15947)
  and u19444 (Bp7pw6, Rx7pw6, Yx7pw6);  // ../RTL/cortexm0ds_logic.v(15948)
  and u19445 (n5546, N5fpw6[17], Sdaiu6);  // ../RTL/cortexm0ds_logic.v(15949)
  not u19446 (Yx7pw6, n5546);  // ../RTL/cortexm0ds_logic.v(15949)
  and u19447 (n5547, Eafpw6[18], A3iiu6);  // ../RTL/cortexm0ds_logic.v(15950)
  not u19448 (Rx7pw6, n5547);  // ../RTL/cortexm0ds_logic.v(15950)
  and u19449 (n5548, Fy7pw6, My7pw6);  // ../RTL/cortexm0ds_logic.v(15952)
  not u1945 (Sl2iu6, n219);  // ../RTL/cortexm0ds_logic.v(3789)
  not u19450 (Wxdpw6, n5548);  // ../RTL/cortexm0ds_logic.v(15952)
  or u19451 (My7pw6, T2iiu6, Cm0iu6);  // ../RTL/cortexm0ds_logic.v(15953)
  AL_MUX u19452 (
    .i0(U9miu6),
    .i1(Ty7pw6),
    .sel(Mm4ju6),
    .o(Cm0iu6));  // ../RTL/cortexm0ds_logic.v(15954)
  and u19453 (Ty7pw6, Az7pw6, Hz7pw6);  // ../RTL/cortexm0ds_logic.v(15955)
  and u19454 (Hz7pw6, Oz7pw6, Vz7pw6);  // ../RTL/cortexm0ds_logic.v(15956)
  and u19455 (Vz7pw6, C08pw6, J08pw6);  // ../RTL/cortexm0ds_logic.v(15957)
  and u19456 (n5549, Jo4ju6, vis_r14_o[17]);  // ../RTL/cortexm0ds_logic.v(15958)
  not u19457 (J08pw6, n5549);  // ../RTL/cortexm0ds_logic.v(15958)
  and u19458 (C08pw6, Q08pw6, X08pw6);  // ../RTL/cortexm0ds_logic.v(15959)
  and u19459 (n5550, Ep4ju6, vis_psp_o[15]);  // ../RTL/cortexm0ds_logic.v(15960)
  and u1946 (n220, Gm2iu6, Nm2iu6);  // ../RTL/cortexm0ds_logic.v(3790)
  not u19460 (X08pw6, n5550);  // ../RTL/cortexm0ds_logic.v(15960)
  and u19461 (n5551, Lp4ju6, vis_msp_o[15]);  // ../RTL/cortexm0ds_logic.v(15961)
  not u19462 (Q08pw6, n5551);  // ../RTL/cortexm0ds_logic.v(15961)
  and u19463 (Oz7pw6, E18pw6, L18pw6);  // ../RTL/cortexm0ds_logic.v(15962)
  and u19464 (n5552, Gq4ju6, vis_r12_o[17]);  // ../RTL/cortexm0ds_logic.v(15963)
  not u19465 (L18pw6, n5552);  // ../RTL/cortexm0ds_logic.v(15963)
  and u19466 (n5553, Nq4ju6, vis_r11_o[17]);  // ../RTL/cortexm0ds_logic.v(15964)
  not u19467 (E18pw6, n5553);  // ../RTL/cortexm0ds_logic.v(15964)
  and u19468 (Az7pw6, S18pw6, Z18pw6);  // ../RTL/cortexm0ds_logic.v(15965)
  and u19469 (Z18pw6, G28pw6, N28pw6);  // ../RTL/cortexm0ds_logic.v(15966)
  not u1947 (Zxxhu6, n220);  // ../RTL/cortexm0ds_logic.v(3790)
  and u19470 (n5554, Wr4ju6, vis_r10_o[17]);  // ../RTL/cortexm0ds_logic.v(15967)
  not u19471 (N28pw6, n5554);  // ../RTL/cortexm0ds_logic.v(15967)
  and u19472 (n5555, Ds4ju6, vis_r9_o[17]);  // ../RTL/cortexm0ds_logic.v(15968)
  not u19473 (G28pw6, n5555);  // ../RTL/cortexm0ds_logic.v(15968)
  and u19474 (S18pw6, Z90iu6, U28pw6);  // ../RTL/cortexm0ds_logic.v(15969)
  and u19475 (n5556, Rs4ju6, vis_r8_o[17]);  // ../RTL/cortexm0ds_logic.v(15970)
  not u19476 (U28pw6, n5556);  // ../RTL/cortexm0ds_logic.v(15970)
  and u19477 (Z90iu6, B38pw6, I38pw6);  // ../RTL/cortexm0ds_logic.v(15971)
  and u19478 (I38pw6, P38pw6, W38pw6);  // ../RTL/cortexm0ds_logic.v(15972)
  and u19479 (W38pw6, D48pw6, K48pw6);  // ../RTL/cortexm0ds_logic.v(15973)
  and u1948 (Nm2iu6, Um2iu6, L72iu6);  // ../RTL/cortexm0ds_logic.v(3791)
  and u19480 (n5557, V6now6, vis_r2_o[17]);  // ../RTL/cortexm0ds_logic.v(15974)
  not u19481 (K48pw6, n5557);  // ../RTL/cortexm0ds_logic.v(15974)
  and u19482 (n5558, C7now6, vis_r6_o[17]);  // ../RTL/cortexm0ds_logic.v(15975)
  not u19483 (D48pw6, n5558);  // ../RTL/cortexm0ds_logic.v(15975)
  and u19484 (P38pw6, R48pw6, Y48pw6);  // ../RTL/cortexm0ds_logic.v(15976)
  and u19485 (n5559, X7now6, vis_r5_o[17]);  // ../RTL/cortexm0ds_logic.v(15977)
  not u19486 (Y48pw6, n5559);  // ../RTL/cortexm0ds_logic.v(15977)
  and u19487 (n5560, E8now6, vis_r4_o[17]);  // ../RTL/cortexm0ds_logic.v(15978)
  not u19488 (R48pw6, n5560);  // ../RTL/cortexm0ds_logic.v(15978)
  and u19489 (B38pw6, F58pw6, M58pw6);  // ../RTL/cortexm0ds_logic.v(15979)
  and u1949 (n221, Uthpw6[16], Vk1iu6);  // ../RTL/cortexm0ds_logic.v(3792)
  and u19490 (M58pw6, T58pw6, A68pw6);  // ../RTL/cortexm0ds_logic.v(15980)
  and u19491 (n5561, N9now6, vis_r1_o[17]);  // ../RTL/cortexm0ds_logic.v(15981)
  not u19492 (A68pw6, n5561);  // ../RTL/cortexm0ds_logic.v(15981)
  and u19493 (n5562, U9now6, vis_r0_o[17]);  // ../RTL/cortexm0ds_logic.v(15982)
  not u19494 (T58pw6, n5562);  // ../RTL/cortexm0ds_logic.v(15982)
  and u19495 (F58pw6, H68pw6, O68pw6);  // ../RTL/cortexm0ds_logic.v(15983)
  and u19496 (n5563, Panow6, vis_r3_o[17]);  // ../RTL/cortexm0ds_logic.v(15984)
  not u19497 (O68pw6, n5563);  // ../RTL/cortexm0ds_logic.v(15984)
  and u19498 (n5564, Wanow6, vis_r7_o[17]);  // ../RTL/cortexm0ds_logic.v(15985)
  not u19499 (H68pw6, n5564);  // ../RTL/cortexm0ds_logic.v(15985)
  buf u195 (Uthpw6[2], Hg7ax6);  // ../RTL/cortexm0ds_logic.v(1882)
  not u1950 (Um2iu6, n221);  // ../RTL/cortexm0ds_logic.v(3792)
  not u19500 (U9miu6, Fkfpw6[17]);  // ../RTL/cortexm0ds_logic.v(15986)
  and u19501 (Fy7pw6, V68pw6, C78pw6);  // ../RTL/cortexm0ds_logic.v(15987)
  and u19502 (n5565, N5fpw6[16], Sdaiu6);  // ../RTL/cortexm0ds_logic.v(15988)
  not u19503 (C78pw6, n5565);  // ../RTL/cortexm0ds_logic.v(15988)
  and u19504 (n5566, Eafpw6[17], A3iiu6);  // ../RTL/cortexm0ds_logic.v(15989)
  not u19505 (V68pw6, n5566);  // ../RTL/cortexm0ds_logic.v(15989)
  and u19506 (n5567, J78pw6, Q78pw6);  // ../RTL/cortexm0ds_logic.v(15991)
  not u19507 (Pxdpw6, n5567);  // ../RTL/cortexm0ds_logic.v(15991)
  or u19508 (Q78pw6, T2iiu6, Jm0iu6);  // ../RTL/cortexm0ds_logic.v(15992)
  AL_MUX u19509 (
    .i0(Tcmiu6),
    .i1(X78pw6),
    .sel(Mm4ju6),
    .o(Jm0iu6));  // ../RTL/cortexm0ds_logic.v(15993)
  and u1951 (Gm2iu6, Bn2iu6, In2iu6);  // ../RTL/cortexm0ds_logic.v(3793)
  and u19510 (X78pw6, E88pw6, L88pw6);  // ../RTL/cortexm0ds_logic.v(15994)
  and u19511 (L88pw6, S88pw6, Z88pw6);  // ../RTL/cortexm0ds_logic.v(15995)
  and u19512 (Z88pw6, G98pw6, N98pw6);  // ../RTL/cortexm0ds_logic.v(15996)
  and u19513 (n5568, Jo4ju6, vis_r14_o[16]);  // ../RTL/cortexm0ds_logic.v(15997)
  not u19514 (N98pw6, n5568);  // ../RTL/cortexm0ds_logic.v(15997)
  and u19515 (G98pw6, U98pw6, Ba8pw6);  // ../RTL/cortexm0ds_logic.v(15998)
  and u19516 (n5569, Ep4ju6, vis_psp_o[14]);  // ../RTL/cortexm0ds_logic.v(15999)
  not u19517 (Ba8pw6, n5569);  // ../RTL/cortexm0ds_logic.v(15999)
  and u19518 (n5570, Lp4ju6, vis_msp_o[14]);  // ../RTL/cortexm0ds_logic.v(16000)
  not u19519 (U98pw6, n5570);  // ../RTL/cortexm0ds_logic.v(16000)
  and u1952 (n222, Iahpw6[15], Xl1iu6);  // ../RTL/cortexm0ds_logic.v(3794)
  and u19520 (S88pw6, Ia8pw6, Pa8pw6);  // ../RTL/cortexm0ds_logic.v(16001)
  and u19521 (n5571, Gq4ju6, vis_r12_o[16]);  // ../RTL/cortexm0ds_logic.v(16002)
  not u19522 (Pa8pw6, n5571);  // ../RTL/cortexm0ds_logic.v(16002)
  and u19523 (n5572, Nq4ju6, vis_r11_o[16]);  // ../RTL/cortexm0ds_logic.v(16003)
  not u19524 (Ia8pw6, n5572);  // ../RTL/cortexm0ds_logic.v(16003)
  and u19525 (E88pw6, Wa8pw6, Db8pw6);  // ../RTL/cortexm0ds_logic.v(16004)
  and u19526 (Db8pw6, Kb8pw6, Rb8pw6);  // ../RTL/cortexm0ds_logic.v(16005)
  and u19527 (n5573, Wr4ju6, vis_r10_o[16]);  // ../RTL/cortexm0ds_logic.v(16006)
  not u19528 (Rb8pw6, n5573);  // ../RTL/cortexm0ds_logic.v(16006)
  and u19529 (n5574, Ds4ju6, vis_r9_o[16]);  // ../RTL/cortexm0ds_logic.v(16007)
  not u1953 (In2iu6, n222);  // ../RTL/cortexm0ds_logic.v(3794)
  not u19530 (Kb8pw6, n5574);  // ../RTL/cortexm0ds_logic.v(16007)
  and u19531 (Wa8pw6, Ga0iu6, Yb8pw6);  // ../RTL/cortexm0ds_logic.v(16008)
  and u19532 (n5575, Rs4ju6, vis_r8_o[16]);  // ../RTL/cortexm0ds_logic.v(16009)
  not u19533 (Yb8pw6, n5575);  // ../RTL/cortexm0ds_logic.v(16009)
  and u19534 (Ga0iu6, Fc8pw6, Mc8pw6);  // ../RTL/cortexm0ds_logic.v(16010)
  and u19535 (Mc8pw6, Tc8pw6, Ad8pw6);  // ../RTL/cortexm0ds_logic.v(16011)
  and u19536 (Ad8pw6, Hd8pw6, Od8pw6);  // ../RTL/cortexm0ds_logic.v(16012)
  and u19537 (n5576, V6now6, vis_r2_o[16]);  // ../RTL/cortexm0ds_logic.v(16013)
  not u19538 (Od8pw6, n5576);  // ../RTL/cortexm0ds_logic.v(16013)
  and u19539 (n5577, C7now6, vis_r6_o[16]);  // ../RTL/cortexm0ds_logic.v(16014)
  and u1954 (n223, Iahpw6[16], Z4yhu6);  // ../RTL/cortexm0ds_logic.v(3795)
  not u19540 (Hd8pw6, n5577);  // ../RTL/cortexm0ds_logic.v(16014)
  and u19541 (Tc8pw6, Vd8pw6, Ce8pw6);  // ../RTL/cortexm0ds_logic.v(16015)
  and u19542 (n5578, X7now6, vis_r5_o[16]);  // ../RTL/cortexm0ds_logic.v(16016)
  not u19543 (Ce8pw6, n5578);  // ../RTL/cortexm0ds_logic.v(16016)
  and u19544 (n5579, E8now6, vis_r4_o[16]);  // ../RTL/cortexm0ds_logic.v(16017)
  not u19545 (Vd8pw6, n5579);  // ../RTL/cortexm0ds_logic.v(16017)
  and u19546 (Fc8pw6, Je8pw6, Qe8pw6);  // ../RTL/cortexm0ds_logic.v(16018)
  and u19547 (Qe8pw6, Xe8pw6, Ef8pw6);  // ../RTL/cortexm0ds_logic.v(16019)
  and u19548 (n5580, N9now6, vis_r1_o[16]);  // ../RTL/cortexm0ds_logic.v(16020)
  not u19549 (Ef8pw6, n5580);  // ../RTL/cortexm0ds_logic.v(16020)
  not u1955 (Bn2iu6, n223);  // ../RTL/cortexm0ds_logic.v(3795)
  and u19550 (n5581, U9now6, vis_r0_o[16]);  // ../RTL/cortexm0ds_logic.v(16021)
  not u19551 (Xe8pw6, n5581);  // ../RTL/cortexm0ds_logic.v(16021)
  and u19552 (Je8pw6, Lf8pw6, Sf8pw6);  // ../RTL/cortexm0ds_logic.v(16022)
  and u19553 (n5582, Panow6, vis_r3_o[16]);  // ../RTL/cortexm0ds_logic.v(16023)
  not u19554 (Sf8pw6, n5582);  // ../RTL/cortexm0ds_logic.v(16023)
  and u19555 (n5583, Wanow6, vis_r7_o[16]);  // ../RTL/cortexm0ds_logic.v(16024)
  not u19556 (Lf8pw6, n5583);  // ../RTL/cortexm0ds_logic.v(16024)
  not u19557 (Tcmiu6, Fkfpw6[16]);  // ../RTL/cortexm0ds_logic.v(16025)
  and u19558 (J78pw6, Zf8pw6, Gg8pw6);  // ../RTL/cortexm0ds_logic.v(16026)
  and u19559 (n5584, N5fpw6[15], Sdaiu6);  // ../RTL/cortexm0ds_logic.v(16027)
  and u1956 (n224, Pn2iu6, Wn2iu6);  // ../RTL/cortexm0ds_logic.v(3796)
  not u19560 (Gg8pw6, n5584);  // ../RTL/cortexm0ds_logic.v(16027)
  and u19561 (n5585, Eafpw6[16], A3iiu6);  // ../RTL/cortexm0ds_logic.v(16028)
  not u19562 (Zf8pw6, n5585);  // ../RTL/cortexm0ds_logic.v(16028)
  and u19563 (n5488[0], Fi9pw6, Mi9pw6);  // ../RTL/cortexm0ds_logic.v(15829)
  buf u19564 (Lwgpw6[0], Zx8ax6);  // ../RTL/cortexm0ds_logic.v(2229)
  and u19565 (n5586, N5fpw6[14], Sdaiu6);  // ../RTL/cortexm0ds_logic.v(16031)
  not u19566 (Ug8pw6, n5586);  // ../RTL/cortexm0ds_logic.v(16031)
  and u19567 (Ng8pw6, Bh8pw6, Ih8pw6);  // ../RTL/cortexm0ds_logic.v(16032)
  or u19568 (Ih8pw6, T2iiu6, Qm0iu6);  // ../RTL/cortexm0ds_logic.v(16033)
  AL_MUX u19569 (
    .i0(Sfmiu6),
    .i1(Ph8pw6),
    .sel(Mm4ju6),
    .o(Qm0iu6));  // ../RTL/cortexm0ds_logic.v(16034)
  not u1957 (Sxxhu6, n224);  // ../RTL/cortexm0ds_logic.v(3796)
  and u19570 (Ph8pw6, Wh8pw6, Di8pw6);  // ../RTL/cortexm0ds_logic.v(16035)
  and u19571 (Di8pw6, Ki8pw6, Ri8pw6);  // ../RTL/cortexm0ds_logic.v(16036)
  and u19572 (Ri8pw6, Yi8pw6, Fj8pw6);  // ../RTL/cortexm0ds_logic.v(16037)
  and u19573 (n5587, Jo4ju6, vis_r14_o[15]);  // ../RTL/cortexm0ds_logic.v(16038)
  not u19574 (Fj8pw6, n5587);  // ../RTL/cortexm0ds_logic.v(16038)
  and u19575 (Yi8pw6, Mj8pw6, Tj8pw6);  // ../RTL/cortexm0ds_logic.v(16039)
  and u19576 (n5588, Ep4ju6, vis_psp_o[13]);  // ../RTL/cortexm0ds_logic.v(16040)
  not u19577 (Tj8pw6, n5588);  // ../RTL/cortexm0ds_logic.v(16040)
  and u19578 (n5589, Lp4ju6, vis_msp_o[13]);  // ../RTL/cortexm0ds_logic.v(16041)
  not u19579 (Mj8pw6, n5589);  // ../RTL/cortexm0ds_logic.v(16041)
  and u1958 (n225, Iahpw6[15], Z4yhu6);  // ../RTL/cortexm0ds_logic.v(3797)
  and u19580 (Ki8pw6, Ak8pw6, Hk8pw6);  // ../RTL/cortexm0ds_logic.v(16042)
  and u19581 (n5590, Gq4ju6, vis_r12_o[15]);  // ../RTL/cortexm0ds_logic.v(16043)
  not u19582 (Hk8pw6, n5590);  // ../RTL/cortexm0ds_logic.v(16043)
  and u19583 (n5591, Nq4ju6, vis_r11_o[15]);  // ../RTL/cortexm0ds_logic.v(16044)
  not u19584 (Ak8pw6, n5591);  // ../RTL/cortexm0ds_logic.v(16044)
  and u19585 (Wh8pw6, Ok8pw6, Vk8pw6);  // ../RTL/cortexm0ds_logic.v(16045)
  and u19586 (Vk8pw6, Cl8pw6, Jl8pw6);  // ../RTL/cortexm0ds_logic.v(16046)
  and u19587 (n5592, Wr4ju6, vis_r10_o[15]);  // ../RTL/cortexm0ds_logic.v(16047)
  not u19588 (Jl8pw6, n5592);  // ../RTL/cortexm0ds_logic.v(16047)
  and u19589 (n5593, Ds4ju6, vis_r9_o[15]);  // ../RTL/cortexm0ds_logic.v(16048)
  not u1959 (Wn2iu6, n225);  // ../RTL/cortexm0ds_logic.v(3797)
  not u19590 (Cl8pw6, n5593);  // ../RTL/cortexm0ds_logic.v(16048)
  and u19591 (Ok8pw6, Na0iu6, Ql8pw6);  // ../RTL/cortexm0ds_logic.v(16049)
  and u19592 (n5594, Rs4ju6, vis_r8_o[15]);  // ../RTL/cortexm0ds_logic.v(16050)
  not u19593 (Ql8pw6, n5594);  // ../RTL/cortexm0ds_logic.v(16050)
  and u19594 (Na0iu6, Xl8pw6, Em8pw6);  // ../RTL/cortexm0ds_logic.v(16051)
  and u19595 (Em8pw6, Lm8pw6, Sm8pw6);  // ../RTL/cortexm0ds_logic.v(16052)
  and u19596 (Sm8pw6, Zm8pw6, Gn8pw6);  // ../RTL/cortexm0ds_logic.v(16053)
  and u19597 (n5595, V6now6, vis_r2_o[15]);  // ../RTL/cortexm0ds_logic.v(16054)
  not u19598 (Gn8pw6, n5595);  // ../RTL/cortexm0ds_logic.v(16054)
  and u19599 (n5596, C7now6, vis_r6_o[15]);  // ../RTL/cortexm0ds_logic.v(16055)
  buf u196 (Jshpw6[26], Nlcbx6);  // ../RTL/cortexm0ds_logic.v(2372)
  and u1960 (Pn2iu6, Do2iu6, Ko2iu6);  // ../RTL/cortexm0ds_logic.v(3798)
  not u19600 (Zm8pw6, n5596);  // ../RTL/cortexm0ds_logic.v(16055)
  and u19601 (Lm8pw6, Nn8pw6, Un8pw6);  // ../RTL/cortexm0ds_logic.v(16056)
  and u19602 (n5597, X7now6, vis_r5_o[15]);  // ../RTL/cortexm0ds_logic.v(16057)
  not u19603 (Un8pw6, n5597);  // ../RTL/cortexm0ds_logic.v(16057)
  and u19604 (n5598, E8now6, vis_r4_o[15]);  // ../RTL/cortexm0ds_logic.v(16058)
  not u19605 (Nn8pw6, n5598);  // ../RTL/cortexm0ds_logic.v(16058)
  and u19606 (Xl8pw6, Bo8pw6, Io8pw6);  // ../RTL/cortexm0ds_logic.v(16059)
  and u19607 (Io8pw6, Po8pw6, Wo8pw6);  // ../RTL/cortexm0ds_logic.v(16060)
  and u19608 (n5599, N9now6, vis_r1_o[15]);  // ../RTL/cortexm0ds_logic.v(16061)
  not u19609 (Wo8pw6, n5599);  // ../RTL/cortexm0ds_logic.v(16061)
  and u1961 (n226, Uthpw6[15], Vk1iu6);  // ../RTL/cortexm0ds_logic.v(3799)
  and u19610 (n5600, U9now6, vis_r0_o[15]);  // ../RTL/cortexm0ds_logic.v(16062)
  not u19611 (Po8pw6, n5600);  // ../RTL/cortexm0ds_logic.v(16062)
  and u19612 (Bo8pw6, Dp8pw6, Kp8pw6);  // ../RTL/cortexm0ds_logic.v(16063)
  and u19613 (n5601, Panow6, vis_r3_o[15]);  // ../RTL/cortexm0ds_logic.v(16064)
  not u19614 (Kp8pw6, n5601);  // ../RTL/cortexm0ds_logic.v(16064)
  and u19615 (n5602, Wanow6, vis_r7_o[15]);  // ../RTL/cortexm0ds_logic.v(16065)
  not u19616 (Dp8pw6, n5602);  // ../RTL/cortexm0ds_logic.v(16065)
  not u19617 (Sfmiu6, Fkfpw6[15]);  // ../RTL/cortexm0ds_logic.v(16066)
  and u19618 (n5603, Eafpw6[15], A3iiu6);  // ../RTL/cortexm0ds_logic.v(16067)
  not u19619 (Bh8pw6, n5603);  // ../RTL/cortexm0ds_logic.v(16067)
  not u1962 (Ko2iu6, n226);  // ../RTL/cortexm0ds_logic.v(3799)
  buf u19620 (vis_r7_o[5], Pxvax6);  // ../RTL/cortexm0ds_logic.v(2654)
  buf u19621 (vis_r7_o[17], Lnwax6);  // ../RTL/cortexm0ds_logic.v(2654)
  and u19622 (n5604, N5fpw6[13], Sdaiu6);  // ../RTL/cortexm0ds_logic.v(16070)
  not u19623 (Yp8pw6, n5604);  // ../RTL/cortexm0ds_logic.v(16070)
  and u19624 (Rp8pw6, Fq8pw6, Mq8pw6);  // ../RTL/cortexm0ds_logic.v(16071)
  or u19625 (Mq8pw6, T2iiu6, Xm0iu6);  // ../RTL/cortexm0ds_logic.v(16072)
  AL_MUX u19626 (
    .i0(Kimiu6),
    .i1(Tq8pw6),
    .sel(Mm4ju6),
    .o(Xm0iu6));  // ../RTL/cortexm0ds_logic.v(16073)
  and u19627 (Tq8pw6, Ar8pw6, Hr8pw6);  // ../RTL/cortexm0ds_logic.v(16074)
  and u19628 (Hr8pw6, Or8pw6, Vr8pw6);  // ../RTL/cortexm0ds_logic.v(16075)
  and u19629 (Vr8pw6, Cs8pw6, Js8pw6);  // ../RTL/cortexm0ds_logic.v(16076)
  and u1963 (n227, Iahpw6[14], Xl1iu6);  // ../RTL/cortexm0ds_logic.v(3800)
  and u19630 (n5605, Jo4ju6, vis_r14_o[14]);  // ../RTL/cortexm0ds_logic.v(16077)
  not u19631 (Js8pw6, n5605);  // ../RTL/cortexm0ds_logic.v(16077)
  and u19632 (Cs8pw6, Qs8pw6, Xs8pw6);  // ../RTL/cortexm0ds_logic.v(16078)
  and u19633 (n5606, Ep4ju6, vis_psp_o[12]);  // ../RTL/cortexm0ds_logic.v(16079)
  not u19634 (Xs8pw6, n5606);  // ../RTL/cortexm0ds_logic.v(16079)
  and u19635 (n5607, Lp4ju6, vis_msp_o[12]);  // ../RTL/cortexm0ds_logic.v(16080)
  not u19636 (Qs8pw6, n5607);  // ../RTL/cortexm0ds_logic.v(16080)
  and u19637 (Or8pw6, Et8pw6, Lt8pw6);  // ../RTL/cortexm0ds_logic.v(16081)
  and u19638 (n5608, Gq4ju6, vis_r12_o[14]);  // ../RTL/cortexm0ds_logic.v(16082)
  not u19639 (Lt8pw6, n5608);  // ../RTL/cortexm0ds_logic.v(16082)
  not u1964 (Do2iu6, n227);  // ../RTL/cortexm0ds_logic.v(3800)
  and u19640 (n5609, Nq4ju6, vis_r11_o[14]);  // ../RTL/cortexm0ds_logic.v(16083)
  not u19641 (Et8pw6, n5609);  // ../RTL/cortexm0ds_logic.v(16083)
  and u19642 (Ar8pw6, St8pw6, Zt8pw6);  // ../RTL/cortexm0ds_logic.v(16084)
  and u19643 (Zt8pw6, Gu8pw6, Nu8pw6);  // ../RTL/cortexm0ds_logic.v(16085)
  and u19644 (n5610, Wr4ju6, vis_r10_o[14]);  // ../RTL/cortexm0ds_logic.v(16086)
  not u19645 (Nu8pw6, n5610);  // ../RTL/cortexm0ds_logic.v(16086)
  and u19646 (n5611, Ds4ju6, vis_r9_o[14]);  // ../RTL/cortexm0ds_logic.v(16087)
  not u19647 (Gu8pw6, n5611);  // ../RTL/cortexm0ds_logic.v(16087)
  and u19648 (St8pw6, Ua0iu6, Uu8pw6);  // ../RTL/cortexm0ds_logic.v(16088)
  and u19649 (n5612, Rs4ju6, vis_r8_o[14]);  // ../RTL/cortexm0ds_logic.v(16089)
  and u1965 (n228, Ro2iu6, Yo2iu6);  // ../RTL/cortexm0ds_logic.v(3801)
  not u19650 (Uu8pw6, n5612);  // ../RTL/cortexm0ds_logic.v(16089)
  and u19651 (Ua0iu6, Bv8pw6, Iv8pw6);  // ../RTL/cortexm0ds_logic.v(16090)
  and u19652 (Iv8pw6, Pv8pw6, Wv8pw6);  // ../RTL/cortexm0ds_logic.v(16091)
  and u19653 (Wv8pw6, Dw8pw6, Kw8pw6);  // ../RTL/cortexm0ds_logic.v(16092)
  and u19654 (n5613, V6now6, vis_r2_o[14]);  // ../RTL/cortexm0ds_logic.v(16093)
  not u19655 (Kw8pw6, n5613);  // ../RTL/cortexm0ds_logic.v(16093)
  and u19656 (n5614, C7now6, vis_r6_o[14]);  // ../RTL/cortexm0ds_logic.v(16094)
  not u19657 (Dw8pw6, n5614);  // ../RTL/cortexm0ds_logic.v(16094)
  and u19658 (Pv8pw6, Rw8pw6, Yw8pw6);  // ../RTL/cortexm0ds_logic.v(16095)
  and u19659 (n5615, X7now6, vis_r5_o[14]);  // ../RTL/cortexm0ds_logic.v(16096)
  not u1966 (Lxxhu6, n228);  // ../RTL/cortexm0ds_logic.v(3801)
  not u19660 (Yw8pw6, n5615);  // ../RTL/cortexm0ds_logic.v(16096)
  and u19661 (n5616, E8now6, vis_r4_o[14]);  // ../RTL/cortexm0ds_logic.v(16097)
  not u19662 (Rw8pw6, n5616);  // ../RTL/cortexm0ds_logic.v(16097)
  and u19663 (Bv8pw6, Fx8pw6, Mx8pw6);  // ../RTL/cortexm0ds_logic.v(16098)
  and u19664 (Mx8pw6, Tx8pw6, Ay8pw6);  // ../RTL/cortexm0ds_logic.v(16099)
  and u19665 (n5617, N9now6, vis_r1_o[14]);  // ../RTL/cortexm0ds_logic.v(16100)
  not u19666 (Ay8pw6, n5617);  // ../RTL/cortexm0ds_logic.v(16100)
  and u19667 (n5618, U9now6, vis_r0_o[14]);  // ../RTL/cortexm0ds_logic.v(16101)
  not u19668 (Tx8pw6, n5618);  // ../RTL/cortexm0ds_logic.v(16101)
  and u19669 (Fx8pw6, Hy8pw6, Oy8pw6);  // ../RTL/cortexm0ds_logic.v(16102)
  and u1967 (n229, Iahpw6[14], Z4yhu6);  // ../RTL/cortexm0ds_logic.v(3802)
  and u19670 (n5619, Panow6, vis_r3_o[14]);  // ../RTL/cortexm0ds_logic.v(16103)
  not u19671 (Oy8pw6, n5619);  // ../RTL/cortexm0ds_logic.v(16103)
  and u19672 (n5620, Wanow6, vis_r7_o[14]);  // ../RTL/cortexm0ds_logic.v(16104)
  not u19673 (Hy8pw6, n5620);  // ../RTL/cortexm0ds_logic.v(16104)
  not u19674 (Kimiu6, Fkfpw6[14]);  // ../RTL/cortexm0ds_logic.v(16105)
  and u19675 (n5621, Eafpw6[14], A3iiu6);  // ../RTL/cortexm0ds_logic.v(16106)
  not u19676 (Fq8pw6, n5621);  // ../RTL/cortexm0ds_logic.v(16106)
  buf u19677 (vis_r7_o[6], Ozvax6);  // ../RTL/cortexm0ds_logic.v(2654)
  buf u19678 (vis_r7_o[18], Llwax6);  // ../RTL/cortexm0ds_logic.v(2654)
  and u19679 (n5622, N5fpw6[12], Sdaiu6);  // ../RTL/cortexm0ds_logic.v(16109)
  not u1968 (Yo2iu6, n229);  // ../RTL/cortexm0ds_logic.v(3802)
  not u19680 (Cz8pw6, n5622);  // ../RTL/cortexm0ds_logic.v(16109)
  and u19681 (Vy8pw6, Jz8pw6, Qz8pw6);  // ../RTL/cortexm0ds_logic.v(16110)
  or u19682 (Qz8pw6, T2iiu6, En0iu6);  // ../RTL/cortexm0ds_logic.v(16111)
  AL_MUX u19683 (
    .i0(Clmiu6),
    .i1(Xz8pw6),
    .sel(Mm4ju6),
    .o(En0iu6));  // ../RTL/cortexm0ds_logic.v(16112)
  and u19684 (Xz8pw6, E09pw6, L09pw6);  // ../RTL/cortexm0ds_logic.v(16113)
  and u19685 (L09pw6, S09pw6, Z09pw6);  // ../RTL/cortexm0ds_logic.v(16114)
  and u19686 (Z09pw6, G19pw6, N19pw6);  // ../RTL/cortexm0ds_logic.v(16115)
  and u19687 (n5623, Jo4ju6, vis_r14_o[13]);  // ../RTL/cortexm0ds_logic.v(16116)
  not u19688 (N19pw6, n5623);  // ../RTL/cortexm0ds_logic.v(16116)
  and u19689 (G19pw6, U19pw6, B29pw6);  // ../RTL/cortexm0ds_logic.v(16117)
  and u1969 (Ro2iu6, Fp2iu6, Mp2iu6);  // ../RTL/cortexm0ds_logic.v(3803)
  and u19690 (n5624, Ep4ju6, vis_psp_o[11]);  // ../RTL/cortexm0ds_logic.v(16118)
  not u19691 (B29pw6, n5624);  // ../RTL/cortexm0ds_logic.v(16118)
  and u19692 (n5625, Lp4ju6, vis_msp_o[11]);  // ../RTL/cortexm0ds_logic.v(16119)
  not u19693 (U19pw6, n5625);  // ../RTL/cortexm0ds_logic.v(16119)
  and u19694 (S09pw6, I29pw6, P29pw6);  // ../RTL/cortexm0ds_logic.v(16120)
  and u19695 (n5626, Gq4ju6, vis_r12_o[13]);  // ../RTL/cortexm0ds_logic.v(16121)
  not u19696 (P29pw6, n5626);  // ../RTL/cortexm0ds_logic.v(16121)
  and u19697 (n5627, Nq4ju6, vis_r11_o[13]);  // ../RTL/cortexm0ds_logic.v(16122)
  not u19698 (I29pw6, n5627);  // ../RTL/cortexm0ds_logic.v(16122)
  and u19699 (E09pw6, W29pw6, D39pw6);  // ../RTL/cortexm0ds_logic.v(16123)
  buf u197 (vis_r12_o[25], Ectax6);  // ../RTL/cortexm0ds_logic.v(2599)
  and u1970 (n230, Uthpw6[14], Vk1iu6);  // ../RTL/cortexm0ds_logic.v(3804)
  and u19700 (D39pw6, K39pw6, R39pw6);  // ../RTL/cortexm0ds_logic.v(16124)
  and u19701 (n5628, Wr4ju6, vis_r10_o[13]);  // ../RTL/cortexm0ds_logic.v(16125)
  not u19702 (R39pw6, n5628);  // ../RTL/cortexm0ds_logic.v(16125)
  and u19703 (n5629, Ds4ju6, vis_r9_o[13]);  // ../RTL/cortexm0ds_logic.v(16126)
  not u19704 (K39pw6, n5629);  // ../RTL/cortexm0ds_logic.v(16126)
  and u19705 (W29pw6, Bb0iu6, Y39pw6);  // ../RTL/cortexm0ds_logic.v(16127)
  and u19706 (n5630, Rs4ju6, vis_r8_o[13]);  // ../RTL/cortexm0ds_logic.v(16128)
  not u19707 (Y39pw6, n5630);  // ../RTL/cortexm0ds_logic.v(16128)
  and u19708 (Bb0iu6, F49pw6, M49pw6);  // ../RTL/cortexm0ds_logic.v(16129)
  and u19709 (M49pw6, T49pw6, A59pw6);  // ../RTL/cortexm0ds_logic.v(16130)
  not u1971 (Mp2iu6, n230);  // ../RTL/cortexm0ds_logic.v(3804)
  and u19710 (A59pw6, H59pw6, O59pw6);  // ../RTL/cortexm0ds_logic.v(16131)
  and u19711 (n5631, V6now6, vis_r2_o[13]);  // ../RTL/cortexm0ds_logic.v(16132)
  not u19712 (O59pw6, n5631);  // ../RTL/cortexm0ds_logic.v(16132)
  and u19713 (n5632, C7now6, vis_r6_o[13]);  // ../RTL/cortexm0ds_logic.v(16133)
  not u19714 (H59pw6, n5632);  // ../RTL/cortexm0ds_logic.v(16133)
  and u19715 (T49pw6, V59pw6, C69pw6);  // ../RTL/cortexm0ds_logic.v(16134)
  and u19716 (n5633, X7now6, vis_r5_o[13]);  // ../RTL/cortexm0ds_logic.v(16135)
  not u19717 (C69pw6, n5633);  // ../RTL/cortexm0ds_logic.v(16135)
  and u19718 (n5634, E8now6, vis_r4_o[13]);  // ../RTL/cortexm0ds_logic.v(16136)
  not u19719 (V59pw6, n5634);  // ../RTL/cortexm0ds_logic.v(16136)
  and u1972 (n231, Iahpw6[13], Xl1iu6);  // ../RTL/cortexm0ds_logic.v(3805)
  and u19720 (F49pw6, J69pw6, Q69pw6);  // ../RTL/cortexm0ds_logic.v(16137)
  and u19721 (Q69pw6, X69pw6, E79pw6);  // ../RTL/cortexm0ds_logic.v(16138)
  and u19722 (n5635, N9now6, vis_r1_o[13]);  // ../RTL/cortexm0ds_logic.v(16139)
  not u19723 (E79pw6, n5635);  // ../RTL/cortexm0ds_logic.v(16139)
  and u19724 (n5636, U9now6, vis_r0_o[13]);  // ../RTL/cortexm0ds_logic.v(16140)
  not u19725 (X69pw6, n5636);  // ../RTL/cortexm0ds_logic.v(16140)
  and u19726 (J69pw6, L79pw6, S79pw6);  // ../RTL/cortexm0ds_logic.v(16141)
  and u19727 (n5637, Panow6, vis_r3_o[13]);  // ../RTL/cortexm0ds_logic.v(16142)
  not u19728 (S79pw6, n5637);  // ../RTL/cortexm0ds_logic.v(16142)
  and u19729 (n5638, Wanow6, vis_r7_o[13]);  // ../RTL/cortexm0ds_logic.v(16143)
  not u1973 (Fp2iu6, n231);  // ../RTL/cortexm0ds_logic.v(3805)
  not u19730 (L79pw6, n5638);  // ../RTL/cortexm0ds_logic.v(16143)
  not u19731 (Clmiu6, Fkfpw6[13]);  // ../RTL/cortexm0ds_logic.v(16144)
  and u19732 (n5639, Eafpw6[13], A3iiu6);  // ../RTL/cortexm0ds_logic.v(16145)
  not u19733 (Jz8pw6, n5639);  // ../RTL/cortexm0ds_logic.v(16145)
  and u19734 (n5640, Z79pw6, G89pw6);  // ../RTL/cortexm0ds_logic.v(16147)
  not u19735 (Ixdpw6, n5640);  // ../RTL/cortexm0ds_logic.v(16147)
  or u19736 (G89pw6, T2iiu6, Ln0iu6);  // ../RTL/cortexm0ds_logic.v(16148)
  AL_MUX u19737 (
    .i0(N89pw6),
    .i1(Unmiu6),
    .sel(Cn5ju6),
    .o(Ln0iu6));  // ../RTL/cortexm0ds_logic.v(16149)
  not u19738 (Cn5ju6, Mm4ju6);  // ../RTL/cortexm0ds_logic.v(16150)
  not u19739 (Unmiu6, Fkfpw6[12]);  // ../RTL/cortexm0ds_logic.v(16151)
  and u1974 (n232, Tp2iu6, Aq2iu6);  // ../RTL/cortexm0ds_logic.v(3806)
  and u19740 (N89pw6, U89pw6, B99pw6);  // ../RTL/cortexm0ds_logic.v(16152)
  and u19741 (B99pw6, I99pw6, P99pw6);  // ../RTL/cortexm0ds_logic.v(16153)
  and u19742 (P99pw6, W99pw6, Da9pw6);  // ../RTL/cortexm0ds_logic.v(16154)
  and u19743 (n5641, Jo4ju6, vis_r14_o[12]);  // ../RTL/cortexm0ds_logic.v(16155)
  not u19744 (Da9pw6, n5641);  // ../RTL/cortexm0ds_logic.v(16155)
  and u19745 (W99pw6, Ka9pw6, Ra9pw6);  // ../RTL/cortexm0ds_logic.v(16156)
  and u19746 (n5642, Ep4ju6, vis_psp_o[10]);  // ../RTL/cortexm0ds_logic.v(16157)
  not u19747 (Ra9pw6, n5642);  // ../RTL/cortexm0ds_logic.v(16157)
  and u19748 (Ep4ju6, Ya9pw6, Fb9pw6);  // ../RTL/cortexm0ds_logic.v(16158)
  or u19749 (n5643, Mb9pw6, Vq2pw6);  // ../RTL/cortexm0ds_logic.v(16159)
  not u1975 (Exxhu6, n232);  // ../RTL/cortexm0ds_logic.v(3806)
  not u19750 (Ya9pw6, n5643);  // ../RTL/cortexm0ds_logic.v(16159)
  not u19751 (Vq2pw6, Vrfhu6);  // ../RTL/cortexm0ds_logic.v(16160)
  and u19752 (n5644, Lp4ju6, vis_msp_o[10]);  // ../RTL/cortexm0ds_logic.v(16161)
  not u19753 (Ka9pw6, n5644);  // ../RTL/cortexm0ds_logic.v(16161)
  and u19754 (Lp4ju6, Tb9pw6, Fb9pw6);  // ../RTL/cortexm0ds_logic.v(16162)
  or u19755 (n5645, Mb9pw6, Vrfhu6);  // ../RTL/cortexm0ds_logic.v(16163)
  not u19756 (Tb9pw6, n5645);  // ../RTL/cortexm0ds_logic.v(16163)
  and u19757 (I99pw6, Ac9pw6, Hc9pw6);  // ../RTL/cortexm0ds_logic.v(16164)
  and u19758 (n5646, Gq4ju6, vis_r12_o[12]);  // ../RTL/cortexm0ds_logic.v(16165)
  not u19759 (Hc9pw6, n5646);  // ../RTL/cortexm0ds_logic.v(16165)
  and u1976 (n233, Iahpw6[13], Z4yhu6);  // ../RTL/cortexm0ds_logic.v(3807)
  and u19760 (n5647, Nq4ju6, vis_r11_o[12]);  // ../RTL/cortexm0ds_logic.v(16166)
  not u19761 (Ac9pw6, n5647);  // ../RTL/cortexm0ds_logic.v(16166)
  and u19762 (U89pw6, Oc9pw6, Vc9pw6);  // ../RTL/cortexm0ds_logic.v(16167)
  and u19763 (Vc9pw6, Cd9pw6, Jd9pw6);  // ../RTL/cortexm0ds_logic.v(16168)
  and u19764 (n5648, Wr4ju6, vis_r10_o[12]);  // ../RTL/cortexm0ds_logic.v(16169)
  not u19765 (Jd9pw6, n5648);  // ../RTL/cortexm0ds_logic.v(16169)
  and u19766 (n5649, Ds4ju6, vis_r9_o[12]);  // ../RTL/cortexm0ds_logic.v(16170)
  not u19767 (Cd9pw6, n5649);  // ../RTL/cortexm0ds_logic.v(16170)
  and u19768 (Oc9pw6, Ib0iu6, Qd9pw6);  // ../RTL/cortexm0ds_logic.v(16171)
  and u19769 (n5650, Rs4ju6, vis_r8_o[12]);  // ../RTL/cortexm0ds_logic.v(16172)
  not u1977 (Aq2iu6, n233);  // ../RTL/cortexm0ds_logic.v(3807)
  not u19770 (Qd9pw6, n5650);  // ../RTL/cortexm0ds_logic.v(16172)
  and u19771 (Ib0iu6, Xd9pw6, Ee9pw6);  // ../RTL/cortexm0ds_logic.v(16173)
  and u19772 (Ee9pw6, Le9pw6, Se9pw6);  // ../RTL/cortexm0ds_logic.v(16174)
  and u19773 (Se9pw6, Ze9pw6, Gf9pw6);  // ../RTL/cortexm0ds_logic.v(16175)
  and u19774 (n5651, V6now6, vis_r2_o[12]);  // ../RTL/cortexm0ds_logic.v(16176)
  not u19775 (Gf9pw6, n5651);  // ../RTL/cortexm0ds_logic.v(16176)
  and u19776 (n5652, C7now6, vis_r6_o[12]);  // ../RTL/cortexm0ds_logic.v(16177)
  not u19777 (Ze9pw6, n5652);  // ../RTL/cortexm0ds_logic.v(16177)
  and u19778 (Le9pw6, Nf9pw6, Uf9pw6);  // ../RTL/cortexm0ds_logic.v(16178)
  and u19779 (n5653, X7now6, vis_r5_o[12]);  // ../RTL/cortexm0ds_logic.v(16179)
  and u1978 (Tp2iu6, Hq2iu6, Oq2iu6);  // ../RTL/cortexm0ds_logic.v(3808)
  not u19780 (Uf9pw6, n5653);  // ../RTL/cortexm0ds_logic.v(16179)
  and u19781 (n5654, E8now6, vis_r4_o[12]);  // ../RTL/cortexm0ds_logic.v(16180)
  not u19782 (Nf9pw6, n5654);  // ../RTL/cortexm0ds_logic.v(16180)
  and u19783 (Xd9pw6, Bg9pw6, Ig9pw6);  // ../RTL/cortexm0ds_logic.v(16181)
  and u19784 (Ig9pw6, Pg9pw6, Wg9pw6);  // ../RTL/cortexm0ds_logic.v(16182)
  and u19785 (n5655, N9now6, vis_r1_o[12]);  // ../RTL/cortexm0ds_logic.v(16183)
  not u19786 (Wg9pw6, n5655);  // ../RTL/cortexm0ds_logic.v(16183)
  and u19787 (n5656, U9now6, vis_r0_o[12]);  // ../RTL/cortexm0ds_logic.v(16184)
  not u19788 (Pg9pw6, n5656);  // ../RTL/cortexm0ds_logic.v(16184)
  and u19789 (Bg9pw6, Dh9pw6, Kh9pw6);  // ../RTL/cortexm0ds_logic.v(16185)
  and u1979 (n234, Uthpw6[13], Vk1iu6);  // ../RTL/cortexm0ds_logic.v(3809)
  and u19790 (n5657, Panow6, vis_r3_o[12]);  // ../RTL/cortexm0ds_logic.v(16186)
  not u19791 (Kh9pw6, n5657);  // ../RTL/cortexm0ds_logic.v(16186)
  and u19792 (n5658, Wanow6, vis_r7_o[12]);  // ../RTL/cortexm0ds_logic.v(16187)
  not u19793 (Dh9pw6, n5658);  // ../RTL/cortexm0ds_logic.v(16187)
  not u19794 (T2iiu6, B7iiu6);  // ../RTL/cortexm0ds_logic.v(16188)
  and u19795 (Z79pw6, Rh9pw6, Yh9pw6);  // ../RTL/cortexm0ds_logic.v(16189)
  and u19796 (n5659, N5fpw6[11], Sdaiu6);  // ../RTL/cortexm0ds_logic.v(16190)
  not u19797 (Yh9pw6, n5659);  // ../RTL/cortexm0ds_logic.v(16190)
  and u19798 (n5660, Eafpw6[12], A3iiu6);  // ../RTL/cortexm0ds_logic.v(16191)
  not u19799 (Rh9pw6, n5660);  // ../RTL/cortexm0ds_logic.v(16191)
  buf u198 (Aghhu6, Pexpw6);  // ../RTL/cortexm0ds_logic.v(2058)
  not u1980 (Oq2iu6, n234);  // ../RTL/cortexm0ds_logic.v(3809)
  and u19800 (n5661, Ti9pw6, E4yhu6);  // ../RTL/cortexm0ds_logic.v(16193)
  not u19801 (Mi9pw6, n5661);  // ../RTL/cortexm0ds_logic.v(16193)
  or u19802 (n5662, Aphpw6[1], Aphpw6[2]);  // ../RTL/cortexm0ds_logic.v(16194)
  not u19803 (E4yhu6, n5662);  // ../RTL/cortexm0ds_logic.v(16194)
  and u19804 (Ti9pw6, Ne3pw6, Tnhpw6[0]);  // ../RTL/cortexm0ds_logic.v(16195)
  or u19805 (n5663, Ze9iu6, Wqzhu6);  // ../RTL/cortexm0ds_logic.v(16196)
  not u19806 (Ne3pw6, n5663);  // ../RTL/cortexm0ds_logic.v(16196)
  and u19807 (Wqzhu6, Ho4iu6, H9xiu6);  // ../RTL/cortexm0ds_logic.v(16197)
  not u19808 (H9xiu6, Eq4iu6);  // ../RTL/cortexm0ds_logic.v(16198)
  and u19809 (Eq4iu6, Cjhpw6[3], Iqzhu6);  // ../RTL/cortexm0ds_logic.v(16199)
  and u1981 (n235, Iahpw6[12], Xl1iu6);  // ../RTL/cortexm0ds_logic.v(3810)
  and u19810 (Ho4iu6, Cjhpw6[2], Iqzhu6);  // ../RTL/cortexm0ds_logic.v(16200)
  xor u19811 (Iqzhu6, Lznhu6, Dtnhu6);  // ../RTL/cortexm0ds_logic.v(16201)
  and u19812 (n5664, My0iu6, Ze9iu6);  // ../RTL/cortexm0ds_logic.v(16202)
  not u19813 (Fi9pw6, n5664);  // ../RTL/cortexm0ds_logic.v(16202)
  and u19814 (Xg6iu6, Aj9pw6, Krzhu6);  // ../RTL/cortexm0ds_logic.v(16203)
  not u19815 (Ze9iu6, Xg6iu6);  // ../RTL/cortexm0ds_logic.v(16203)
  or u19816 (n5665, Gpzhu6, Sqhpw6[1]);  // ../RTL/cortexm0ds_logic.v(16204)
  not u19817 (Krzhu6, n5665);  // ../RTL/cortexm0ds_logic.v(16204)
  not u19818 (Gpzhu6, Sqhpw6[0]);  // ../RTL/cortexm0ds_logic.v(16205)
  and u19819 (n7[4], Wkyhu6, Dlyhu6);  // ../RTL/cortexm0ds_logic.v(3185)
  not u1982 (Hq2iu6, n235);  // ../RTL/cortexm0ds_logic.v(3810)
  not u19820 (Ebxiu6, Jzmhu6);  // ../RTL/cortexm0ds_logic.v(16207)
  or u19821 (n5666, Ympiu6, S18iu6);  // ../RTL/cortexm0ds_logic.v(16208)
  not u19822 (HMASTER, n5666);  // ../RTL/cortexm0ds_logic.v(16208)
  and u19823 (S18iu6, Hj9pw6, Oj9pw6);  // ../RTL/cortexm0ds_logic.v(16209)
  or u19824 (n5667, Sdaiu6, Vj9pw6);  // ../RTL/cortexm0ds_logic.v(16210)
  not u19825 (Oj9pw6, n5667);  // ../RTL/cortexm0ds_logic.v(16210)
  buf u19826 (Bhmhu6, Nvkbx6[4]);  // ../RTL/cortexm0ds_logic.v(3137)
  and u19827 (Hj9pw6, Lrhiu6, I1aiu6);  // ../RTL/cortexm0ds_logic.v(16212)
  and u19828 (My0iu6, Jk9pw6, J71iu6);  // ../RTL/cortexm0ds_logic.v(16213)
  or u19829 (n5668, X71iu6, Mnxow6);  // ../RTL/cortexm0ds_logic.v(16214)
  and u1983 (n236, Vq2iu6, Cr2iu6);  // ../RTL/cortexm0ds_logic.v(3811)
  not u19830 (J71iu6, n5668);  // ../RTL/cortexm0ds_logic.v(16214)
  and u19831 (Mnxow6, Ed3pw6, Qk9pw6);  // ../RTL/cortexm0ds_logic.v(16215)
  and u19832 (n5669, Xk9pw6, El9pw6);  // ../RTL/cortexm0ds_logic.v(16216)
  not u19833 (Qk9pw6, n5669);  // ../RTL/cortexm0ds_logic.v(16216)
  and u19834 (n5670, Frziu6, Xe8iu6);  // ../RTL/cortexm0ds_logic.v(16217)
  not u19835 (El9pw6, n5670);  // ../RTL/cortexm0ds_logic.v(16217)
  or u19836 (n5671, Es1ju6, Vjhow6);  // ../RTL/cortexm0ds_logic.v(16218)
  not u19837 (Xk9pw6, n5671);  // ../RTL/cortexm0ds_logic.v(16218)
  buf u19838 (Iimhu6, Nvkbx6[3]);  // ../RTL/cortexm0ds_logic.v(3137)
  and u19839 (Ed3pw6, Ll9pw6, Sl9pw6);  // ../RTL/cortexm0ds_logic.v(16220)
  not u1984 (Xwxhu6, n236);  // ../RTL/cortexm0ds_logic.v(3811)
  not u19840 (X71iu6, Ed3pw6);  // ../RTL/cortexm0ds_logic.v(16220)
  and u19841 (Sl9pw6, Zl9pw6, Gm9pw6);  // ../RTL/cortexm0ds_logic.v(16221)
  or u19842 (Zl9pw6, Mzlow6, Nlaiu6);  // ../RTL/cortexm0ds_logic.v(16222)
  or u19843 (Mzlow6, Ey2ju6, Tfjiu6);  // ../RTL/cortexm0ds_logic.v(16223)
  not u19844 (Ey2ju6, Fd0iu6);  // ../RTL/cortexm0ds_logic.v(16224)
  and u19845 (Ll9pw6, Nm9pw6, He6ju6);  // ../RTL/cortexm0ds_logic.v(16225)
  not u19846 (He6ju6, Ww8ow6);  // ../RTL/cortexm0ds_logic.v(16226)
  and u19847 (Ww8ow6, Tr0iu6, Nlaiu6);  // ../RTL/cortexm0ds_logic.v(16227)
  and u19848 (n5672, H3aju6, Sq3ju6);  // ../RTL/cortexm0ds_logic.v(16228)
  not u19849 (Nm9pw6, n5672);  // ../RTL/cortexm0ds_logic.v(16228)
  and u1985 (Cr2iu6, Jr2iu6, L72iu6);  // ../RTL/cortexm0ds_logic.v(3812)
  or u19850 (n5673, Ympiu6, Ta3pw6);  // ../RTL/cortexm0ds_logic.v(16229)
  not u19851 (Jk9pw6, n5673);  // ../RTL/cortexm0ds_logic.v(16229)
  buf u19852 (Pjmhu6, Nvkbx6[2]);  // ../RTL/cortexm0ds_logic.v(3137)
  and u19853 (Ta3pw6, Um9pw6, Bn9pw6);  // ../RTL/cortexm0ds_logic.v(16231)
  not u19854 (Ay8iu6, Ta3pw6);  // ../RTL/cortexm0ds_logic.v(16231)
  and u19855 (n5674, B7iiu6, Go0iu6);  // ../RTL/cortexm0ds_logic.v(16232)
  not u19856 (Bn9pw6, n5674);  // ../RTL/cortexm0ds_logic.v(16232)
  AL_MUX u19857 (
    .i0(Fkfpw6[0]),
    .i1(In9pw6),
    .sel(Mm4ju6),
    .o(Go0iu6));  // ../RTL/cortexm0ds_logic.v(16233)
  and u19858 (Mm4ju6, Pn9pw6, Wn9pw6);  // ../RTL/cortexm0ds_logic.v(16234)
  and u19859 (Wn9pw6, Do9pw6, Ko9pw6);  // ../RTL/cortexm0ds_logic.v(16235)
  and u1986 (n237, Uthpw6[12], Vk1iu6);  // ../RTL/cortexm0ds_logic.v(3813)
  and u19860 (Ko9pw6, Ro9pw6, Kgaiu6);  // ../RTL/cortexm0ds_logic.v(16236)
  or u19861 (Ro9pw6, Yo9pw6, Fp9pw6);  // ../RTL/cortexm0ds_logic.v(16237)
  and u19862 (Do9pw6, Mp9pw6, Ty8ow6);  // ../RTL/cortexm0ds_logic.v(16238)
  or u19863 (Ty8ow6, Qxaiu6, K9aiu6);  // ../RTL/cortexm0ds_logic.v(16239)
  and u19864 (n5675, Tp9pw6, Toaiu6);  // ../RTL/cortexm0ds_logic.v(16240)
  not u19865 (Mp9pw6, n5675);  // ../RTL/cortexm0ds_logic.v(16240)
  and u19866 (Toaiu6, Pugiu6, Ii0iu6);  // ../RTL/cortexm0ds_logic.v(16241)
  or u19867 (n5676, Nlaiu6, Cyfpw6[4]);  // ../RTL/cortexm0ds_logic.v(16242)
  not u19868 (Tp9pw6, n5676);  // ../RTL/cortexm0ds_logic.v(16242)
  and u19869 (Pn9pw6, Aq9pw6, Hq9pw6);  // ../RTL/cortexm0ds_logic.v(16243)
  not u1987 (Jr2iu6, n237);  // ../RTL/cortexm0ds_logic.v(3813)
  and u19870 (n5677, Tr0iu6, Oq9pw6);  // ../RTL/cortexm0ds_logic.v(16244)
  not u19871 (Hq9pw6, n5677);  // ../RTL/cortexm0ds_logic.v(16244)
  or u19872 (Oq9pw6, W8aiu6, Oiaiu6);  // ../RTL/cortexm0ds_logic.v(16245)
  and u19873 (Aq9pw6, Vq9pw6, Cr9pw6);  // ../RTL/cortexm0ds_logic.v(16246)
  and u19874 (n5678, Jr9pw6, Frziu6);  // ../RTL/cortexm0ds_logic.v(16247)
  not u19875 (Cr9pw6, n5678);  // ../RTL/cortexm0ds_logic.v(16247)
  or u19876 (n5679, Lkaiu6, C0ehu6);  // ../RTL/cortexm0ds_logic.v(16248)
  not u19877 (Jr9pw6, n5679);  // ../RTL/cortexm0ds_logic.v(16248)
  and u19878 (n5680, Qr9pw6, Fhaiu6);  // ../RTL/cortexm0ds_logic.v(16249)
  not u19879 (Vq9pw6, n5680);  // ../RTL/cortexm0ds_logic.v(16249)
  and u1988 (Vq2iu6, Qr2iu6, Xr2iu6);  // ../RTL/cortexm0ds_logic.v(3814)
  and u19880 (Fhaiu6, Nlaiu6, Mr0iu6);  // ../RTL/cortexm0ds_logic.v(16250)
  or u19881 (n5681, As0iu6, Cyfpw6[3]);  // ../RTL/cortexm0ds_logic.v(16251)
  not u19882 (Qr9pw6, n5681);  // ../RTL/cortexm0ds_logic.v(16251)
  and u19883 (n5682, Xr9pw6, Es9pw6);  // ../RTL/cortexm0ds_logic.v(16252)
  not u19884 (In9pw6, n5682);  // ../RTL/cortexm0ds_logic.v(16252)
  and u19885 (Es9pw6, Ls9pw6, Ss9pw6);  // ../RTL/cortexm0ds_logic.v(16253)
  and u19886 (Ss9pw6, Zs9pw6, Gt9pw6);  // ../RTL/cortexm0ds_logic.v(16254)
  and u19887 (n5683, Jo4ju6, vis_r14_o[0]);  // ../RTL/cortexm0ds_logic.v(16255)
  not u19888 (Gt9pw6, n5683);  // ../RTL/cortexm0ds_logic.v(16255)
  or u19889 (n5684, Yo9pw6, Nt9pw6);  // ../RTL/cortexm0ds_logic.v(16256)
  and u1989 (n238, Iahpw6[11], Xl1iu6);  // ../RTL/cortexm0ds_logic.v(3815)
  not u19890 (Jo4ju6, n5684);  // ../RTL/cortexm0ds_logic.v(16256)
  and u19891 (n5685, Gq4ju6, vis_r12_o[0]);  // ../RTL/cortexm0ds_logic.v(16257)
  not u19892 (Zs9pw6, n5685);  // ../RTL/cortexm0ds_logic.v(16257)
  or u19893 (n5686, Yo9pw6, Ut9pw6);  // ../RTL/cortexm0ds_logic.v(16258)
  not u19894 (Gq4ju6, n5686);  // ../RTL/cortexm0ds_logic.v(16258)
  buf u19895 (Wkmhu6, Nvkbx6[1]);  // ../RTL/cortexm0ds_logic.v(3137)
  or u19896 (Yo9pw6, Ssniu6, Fpniu6);  // ../RTL/cortexm0ds_logic.v(16260)
  not u19897 (Fb9pw6, Yo9pw6);  // ../RTL/cortexm0ds_logic.v(16260)
  and u19898 (Ls9pw6, Bu9pw6, Iu9pw6);  // ../RTL/cortexm0ds_logic.v(16261)
  and u19899 (n5687, Nq4ju6, vis_r11_o[0]);  // ../RTL/cortexm0ds_logic.v(16262)
  buf u199 (vis_r2_o[26], Vgqax6);  // ../RTL/cortexm0ds_logic.v(2551)
  not u1990 (Xr2iu6, n238);  // ../RTL/cortexm0ds_logic.v(3815)
  not u19900 (Iu9pw6, n5687);  // ../RTL/cortexm0ds_logic.v(16262)
  or u19901 (n5688, Pu9pw6, Fp9pw6);  // ../RTL/cortexm0ds_logic.v(16263)
  not u19902 (Nq4ju6, n5688);  // ../RTL/cortexm0ds_logic.v(16263)
  and u19903 (n5689, Wr4ju6, vis_r10_o[0]);  // ../RTL/cortexm0ds_logic.v(16264)
  not u19904 (Bu9pw6, n5689);  // ../RTL/cortexm0ds_logic.v(16264)
  or u19905 (n5690, Pu9pw6, Nt9pw6);  // ../RTL/cortexm0ds_logic.v(16265)
  not u19906 (Wr4ju6, n5690);  // ../RTL/cortexm0ds_logic.v(16265)
  and u19907 (Xr9pw6, Wu9pw6, Dc0iu6);  // ../RTL/cortexm0ds_logic.v(16266)
  and u19908 (Dc0iu6, Dv9pw6, Kv9pw6);  // ../RTL/cortexm0ds_logic.v(16267)
  and u19909 (Kv9pw6, Rv9pw6, Yv9pw6);  // ../RTL/cortexm0ds_logic.v(16268)
  and u1991 (n239, Iahpw6[12], Z4yhu6);  // ../RTL/cortexm0ds_logic.v(3816)
  and u19910 (Yv9pw6, Fw9pw6, Mw9pw6);  // ../RTL/cortexm0ds_logic.v(16269)
  and u19911 (n5691, V6now6, vis_r2_o[0]);  // ../RTL/cortexm0ds_logic.v(16270)
  not u19912 (Mw9pw6, n5691);  // ../RTL/cortexm0ds_logic.v(16270)
  or u19913 (n5692, Tw9pw6, Nt9pw6);  // ../RTL/cortexm0ds_logic.v(16271)
  not u19914 (V6now6, n5692);  // ../RTL/cortexm0ds_logic.v(16271)
  and u19915 (n5693, C7now6, vis_r6_o[0]);  // ../RTL/cortexm0ds_logic.v(16272)
  not u19916 (Fw9pw6, n5693);  // ../RTL/cortexm0ds_logic.v(16272)
  or u19917 (n5694, Ax9pw6, Nt9pw6);  // ../RTL/cortexm0ds_logic.v(16273)
  not u19918 (C7now6, n5694);  // ../RTL/cortexm0ds_logic.v(16273)
  or u19919 (Nt9pw6, Mxuow6, H2fpw6[0]);  // ../RTL/cortexm0ds_logic.v(16274)
  not u1992 (Qr2iu6, n239);  // ../RTL/cortexm0ds_logic.v(3816)
  and u19920 (Rv9pw6, Hx9pw6, Ox9pw6);  // ../RTL/cortexm0ds_logic.v(16275)
  and u19921 (n5695, X7now6, vis_r5_o[0]);  // ../RTL/cortexm0ds_logic.v(16276)
  not u19922 (Ox9pw6, n5695);  // ../RTL/cortexm0ds_logic.v(16276)
  or u19923 (n5696, Mb9pw6, Ax9pw6);  // ../RTL/cortexm0ds_logic.v(16277)
  not u19924 (X7now6, n5696);  // ../RTL/cortexm0ds_logic.v(16277)
  and u19925 (n5697, E8now6, vis_r4_o[0]);  // ../RTL/cortexm0ds_logic.v(16278)
  not u19926 (Hx9pw6, n5697);  // ../RTL/cortexm0ds_logic.v(16278)
  or u19927 (n5698, Ut9pw6, Ax9pw6);  // ../RTL/cortexm0ds_logic.v(16279)
  not u19928 (E8now6, n5698);  // ../RTL/cortexm0ds_logic.v(16279)
  and u19929 (Dv9pw6, Vx9pw6, Cy9pw6);  // ../RTL/cortexm0ds_logic.v(16280)
  and u1993 (n240, Es2iu6, Ls2iu6);  // ../RTL/cortexm0ds_logic.v(3817)
  and u19930 (Cy9pw6, Jy9pw6, Qy9pw6);  // ../RTL/cortexm0ds_logic.v(16281)
  and u19931 (n5699, N9now6, vis_r1_o[0]);  // ../RTL/cortexm0ds_logic.v(16282)
  not u19932 (Qy9pw6, n5699);  // ../RTL/cortexm0ds_logic.v(16282)
  or u19933 (n5700, Mb9pw6, Tw9pw6);  // ../RTL/cortexm0ds_logic.v(16283)
  not u19934 (N9now6, n5700);  // ../RTL/cortexm0ds_logic.v(16283)
  and u19935 (n5701, U9now6, vis_r0_o[0]);  // ../RTL/cortexm0ds_logic.v(16284)
  not u19936 (Jy9pw6, n5701);  // ../RTL/cortexm0ds_logic.v(16284)
  or u19937 (n5702, Ut9pw6, Tw9pw6);  // ../RTL/cortexm0ds_logic.v(16285)
  not u19938 (U9now6, n5702);  // ../RTL/cortexm0ds_logic.v(16285)
  and u19939 (Vx9pw6, Xy9pw6, Ez9pw6);  // ../RTL/cortexm0ds_logic.v(16286)
  not u1994 (Qwxhu6, n240);  // ../RTL/cortexm0ds_logic.v(3817)
  and u19940 (n5703, Panow6, vis_r3_o[0]);  // ../RTL/cortexm0ds_logic.v(16287)
  not u19941 (Ez9pw6, n5703);  // ../RTL/cortexm0ds_logic.v(16287)
  or u19942 (n5704, Fp9pw6, Tw9pw6);  // ../RTL/cortexm0ds_logic.v(16288)
  not u19943 (Panow6, n5704);  // ../RTL/cortexm0ds_logic.v(16288)
  or u19944 (Tw9pw6, H2fpw6[2], H2fpw6[3]);  // ../RTL/cortexm0ds_logic.v(16289)
  and u19945 (n5705, Wanow6, vis_r7_o[0]);  // ../RTL/cortexm0ds_logic.v(16290)
  not u19946 (Xy9pw6, n5705);  // ../RTL/cortexm0ds_logic.v(16290)
  or u19947 (n5706, Fp9pw6, Ax9pw6);  // ../RTL/cortexm0ds_logic.v(16291)
  not u19948 (Wanow6, n5706);  // ../RTL/cortexm0ds_logic.v(16291)
  or u19949 (Ax9pw6, Fpniu6, H2fpw6[3]);  // ../RTL/cortexm0ds_logic.v(16292)
  and u1995 (n241, Iahpw6[11], Z4yhu6);  // ../RTL/cortexm0ds_logic.v(3818)
  not u19950 (Fpniu6, H2fpw6[2]);  // ../RTL/cortexm0ds_logic.v(16293)
  or u19951 (Fp9pw6, Vqniu6, Mxuow6);  // ../RTL/cortexm0ds_logic.v(16294)
  not u19952 (Mxuow6, H2fpw6[1]);  // ../RTL/cortexm0ds_logic.v(16295)
  and u19953 (Wu9pw6, Lz9pw6, Sz9pw6);  // ../RTL/cortexm0ds_logic.v(16296)
  and u19954 (n5707, Ds4ju6, vis_r9_o[0]);  // ../RTL/cortexm0ds_logic.v(16297)
  not u19955 (Sz9pw6, n5707);  // ../RTL/cortexm0ds_logic.v(16297)
  or u19956 (n5708, Pu9pw6, Mb9pw6);  // ../RTL/cortexm0ds_logic.v(16298)
  not u19957 (Ds4ju6, n5708);  // ../RTL/cortexm0ds_logic.v(16298)
  or u19958 (Mb9pw6, Vqniu6, H2fpw6[1]);  // ../RTL/cortexm0ds_logic.v(16299)
  not u19959 (Vqniu6, H2fpw6[0]);  // ../RTL/cortexm0ds_logic.v(16300)
  not u1996 (Ls2iu6, n241);  // ../RTL/cortexm0ds_logic.v(3818)
  and u19960 (n5709, Rs4ju6, vis_r8_o[0]);  // ../RTL/cortexm0ds_logic.v(16301)
  not u19961 (Lz9pw6, n5709);  // ../RTL/cortexm0ds_logic.v(16301)
  or u19962 (n5710, Pu9pw6, Ut9pw6);  // ../RTL/cortexm0ds_logic.v(16302)
  not u19963 (Rs4ju6, n5710);  // ../RTL/cortexm0ds_logic.v(16302)
  or u19964 (Ut9pw6, H2fpw6[0], H2fpw6[1]);  // ../RTL/cortexm0ds_logic.v(16303)
  or u19965 (Pu9pw6, Ssniu6, H2fpw6[2]);  // ../RTL/cortexm0ds_logic.v(16304)
  not u19966 (Ssniu6, H2fpw6[3]);  // ../RTL/cortexm0ds_logic.v(16305)
  and u19967 (B7iiu6, Zz9pw6, Ck9pw6);  // ../RTL/cortexm0ds_logic.v(16306)
  and u19968 (n5711, G0apw6, N0apw6);  // ../RTL/cortexm0ds_logic.v(16307)
  not u19969 (Zz9pw6, n5711);  // ../RTL/cortexm0ds_logic.v(16307)
  and u1997 (Es2iu6, Ss2iu6, Zs2iu6);  // ../RTL/cortexm0ds_logic.v(3819)
  and u19970 (N0apw6, U0apw6, B1apw6);  // ../RTL/cortexm0ds_logic.v(16308)
  and u19971 (n5712, Vxniu6, Cyfpw6[0]);  // ../RTL/cortexm0ds_logic.v(16309)
  not u19972 (B1apw6, n5712);  // ../RTL/cortexm0ds_logic.v(16309)
  or u19973 (n5713, Mjfiu6, Tr0iu6);  // ../RTL/cortexm0ds_logic.v(16310)
  not u19974 (Vxniu6, n5713);  // ../RTL/cortexm0ds_logic.v(16310)
  and u19975 (U0apw6, I1apw6, P1apw6);  // ../RTL/cortexm0ds_logic.v(16311)
  and u19976 (n5714, W1apw6, Fq8iu6);  // ../RTL/cortexm0ds_logic.v(16312)
  not u19977 (P1apw6, n5714);  // ../RTL/cortexm0ds_logic.v(16312)
  and u19978 (Fq8iu6, H4ghu6, Nlaiu6);  // ../RTL/cortexm0ds_logic.v(16313)
  and u19979 (n7[3], Spyhu6, Zpyhu6);  // ../RTL/cortexm0ds_logic.v(3185)
  and u1998 (n242, Uthpw6[11], Vk1iu6);  // ../RTL/cortexm0ds_logic.v(3820)
  not u19980 (W1apw6, Mq8iu6);  // ../RTL/cortexm0ds_logic.v(16314)
  and u19981 (n5715, F9aju6, Kr7ow6);  // ../RTL/cortexm0ds_logic.v(16315)
  not u19982 (I1apw6, n5715);  // ../RTL/cortexm0ds_logic.v(16315)
  and u19983 (F9aju6, Cyfpw6[1], Ii0iu6);  // ../RTL/cortexm0ds_logic.v(16316)
  and u19984 (G0apw6, D2apw6, K2apw6);  // ../RTL/cortexm0ds_logic.v(16317)
  or u19985 (K2apw6, Uvziu6, Cyfpw6[5]);  // ../RTL/cortexm0ds_logic.v(16318)
  and u19986 (D2apw6, R2apw6, Y2apw6);  // ../RTL/cortexm0ds_logic.v(16319)
  and u19987 (n5716, Z6aiu6, Y2oiu6);  // ../RTL/cortexm0ds_logic.v(16320)
  not u19988 (Y2apw6, n5716);  // ../RTL/cortexm0ds_logic.v(16320)
  and u19989 (n5717, F3aiu6, Tr0iu6);  // ../RTL/cortexm0ds_logic.v(16321)
  not u1999 (Zs2iu6, n242);  // ../RTL/cortexm0ds_logic.v(3820)
  not u19990 (R2apw6, n5717);  // ../RTL/cortexm0ds_logic.v(16321)
  and u19991 (n5718, Eafpw6[0], A3iiu6);  // ../RTL/cortexm0ds_logic.v(16322)
  not u19992 (Um9pw6, n5718);  // ../RTL/cortexm0ds_logic.v(16322)
  and u19993 (A3iiu6, F3apw6, Ck9pw6);  // ../RTL/cortexm0ds_logic.v(16323)
  and u19994 (Sdaiu6, M3apw6, T3apw6);  // ../RTL/cortexm0ds_logic.v(16324)
  not u19995 (Ck9pw6, Sdaiu6);  // ../RTL/cortexm0ds_logic.v(16324)
  and u19996 (T3apw6, A4apw6, H4apw6);  // ../RTL/cortexm0ds_logic.v(16325)
  and u19997 (H4apw6, O4apw6, V4apw6);  // ../RTL/cortexm0ds_logic.v(16326)
  and u19998 (n5719, C5apw6, Mfjiu6);  // ../RTL/cortexm0ds_logic.v(16327)
  not u19999 (V4apw6, n5719);  // ../RTL/cortexm0ds_logic.v(16327)
  buf u2 (R4gpw6[36], Nhgbx6);  // ../RTL/cortexm0ds_logic.v(2815)
  buf u20 (vis_r14_o[19], Ntnax6);  // ../RTL/cortexm0ds_logic.v(2497)
  buf u200 (vis_r1_o[1], Sfypw6);  // ../RTL/cortexm0ds_logic.v(1876)
  and u2000 (n243, Iahpw6[10], Xl1iu6);  // ../RTL/cortexm0ds_logic.v(3821)
  or u20000 (n5720, Sbghu6, Cyfpw6[6]);  // ../RTL/cortexm0ds_logic.v(16328)
  not u20001 (C5apw6, n5720);  // ../RTL/cortexm0ds_logic.v(16328)
  and u20002 (O4apw6, J5apw6, Td0iu6);  // ../RTL/cortexm0ds_logic.v(16329)
  and u20003 (n5721, Cyfpw6[7], Q5apw6);  // ../RTL/cortexm0ds_logic.v(16330)
  not u20004 (J5apw6, n5721);  // ../RTL/cortexm0ds_logic.v(16330)
  or u20005 (Q5apw6, X5apw6, I82ju6);  // ../RTL/cortexm0ds_logic.v(16331)
  and u20006 (I82ju6, Apaiu6, L45iu6);  // ../RTL/cortexm0ds_logic.v(16332)
  AL_MUX u20007 (
    .i0(N1aow6),
    .i1(Z6aiu6),
    .sel(Cyfpw6[4]),
    .o(X5apw6));  // ../RTL/cortexm0ds_logic.v(16333)
  and u20008 (N1aow6, Wwziu6, Sijiu6);  // ../RTL/cortexm0ds_logic.v(16334)
  not u20009 (Sijiu6, N2ghu6);  // ../RTL/cortexm0ds_logic.v(16335)
  not u2001 (Ss2iu6, n243);  // ../RTL/cortexm0ds_logic.v(3821)
  and u20010 (A4apw6, E6apw6, L6apw6);  // ../RTL/cortexm0ds_logic.v(16336)
  and u20011 (n5722, S6apw6, Gwyiu6);  // ../RTL/cortexm0ds_logic.v(16337)
  not u20012 (L6apw6, n5722);  // ../RTL/cortexm0ds_logic.v(16337)
  or u20013 (n5723, Kq0iu6, Ae0iu6);  // ../RTL/cortexm0ds_logic.v(16338)
  not u20014 (S6apw6, n5723);  // ../RTL/cortexm0ds_logic.v(16338)
  and u20015 (E6apw6, Z6apw6, G7apw6);  // ../RTL/cortexm0ds_logic.v(16339)
  and u20016 (n5724, N7apw6, Hzziu6);  // ../RTL/cortexm0ds_logic.v(16340)
  not u20017 (G7apw6, n5724);  // ../RTL/cortexm0ds_logic.v(16340)
  or u20018 (n5725, Tr0iu6, H4ghu6);  // ../RTL/cortexm0ds_logic.v(16341)
  not u20019 (N7apw6, n5725);  // ../RTL/cortexm0ds_logic.v(16341)
  and u2002 (n244, Gt2iu6, Nt2iu6);  // ../RTL/cortexm0ds_logic.v(3822)
  and u20020 (n5726, U7apw6, B8apw6);  // ../RTL/cortexm0ds_logic.v(16342)
  not u20021 (Z6apw6, n5726);  // ../RTL/cortexm0ds_logic.v(16342)
  or u20022 (n5727, Nloiu6, Cyfpw6[4]);  // ../RTL/cortexm0ds_logic.v(16343)
  not u20023 (U7apw6, n5727);  // ../RTL/cortexm0ds_logic.v(16343)
  and u20024 (M3apw6, I8apw6, P8apw6);  // ../RTL/cortexm0ds_logic.v(16344)
  and u20025 (P8apw6, W8apw6, Cq3pw6);  // ../RTL/cortexm0ds_logic.v(16345)
  or u20026 (Cq3pw6, Mjfiu6, Mr0iu6);  // ../RTL/cortexm0ds_logic.v(16346)
  not u20027 (Mjfiu6, Xzmiu6);  // ../RTL/cortexm0ds_logic.v(16347)
  and u20028 (Xzmiu6, Ii0iu6, Tfjiu6);  // ../RTL/cortexm0ds_logic.v(16348)
  and u20029 (W8apw6, D9apw6, Oq1ju6);  // ../RTL/cortexm0ds_logic.v(16349)
  not u2003 (Jwxhu6, n244);  // ../RTL/cortexm0ds_logic.v(3822)
  and u20030 (n5728, Qe8iu6, G47ow6);  // ../RTL/cortexm0ds_logic.v(16350)
  not u20031 (Oq1ju6, n5728);  // ../RTL/cortexm0ds_logic.v(16350)
  and u20032 (G47ow6, Xe8iu6, Tfjiu6);  // ../RTL/cortexm0ds_logic.v(16351)
  or u20033 (n5729, P1bow6, C0ehu6);  // ../RTL/cortexm0ds_logic.v(16352)
  not u20034 (Qe8iu6, n5729);  // ../RTL/cortexm0ds_logic.v(16352)
  and u20035 (n5730, K9apw6, R9apw6);  // ../RTL/cortexm0ds_logic.v(16353)
  not u20036 (D9apw6, n5730);  // ../RTL/cortexm0ds_logic.v(16353)
  or u20037 (n5731, Qxaiu6, Cyfpw6[5]);  // ../RTL/cortexm0ds_logic.v(16354)
  not u20038 (R9apw6, n5731);  // ../RTL/cortexm0ds_logic.v(16354)
  and u20039 (K9apw6, Yljiu6, Qyniu6);  // ../RTL/cortexm0ds_logic.v(16355)
  and u2004 (Nt2iu6, Ut2iu6, L72iu6);  // ../RTL/cortexm0ds_logic.v(3823)
  and u20040 (I8apw6, Y9apw6, Rcziu6);  // ../RTL/cortexm0ds_logic.v(16356)
  and u20041 (Rcziu6, Faapw6, Oe8ow6);  // ../RTL/cortexm0ds_logic.v(16357)
  or u20042 (Oe8ow6, K9aiu6, Tr0iu6);  // ../RTL/cortexm0ds_logic.v(16358)
  and u20043 (n5732, Gwyiu6, Maapw6);  // ../RTL/cortexm0ds_logic.v(16359)
  not u20044 (Faapw6, n5732);  // ../RTL/cortexm0ds_logic.v(16359)
  or u20045 (Maapw6, Vbiow6, Y0jiu6);  // ../RTL/cortexm0ds_logic.v(16360)
  and u20046 (Y0jiu6, H4ghu6, It2ju6);  // ../RTL/cortexm0ds_logic.v(16361)
  or u20047 (n5733, Xojiu6, Kq0iu6);  // ../RTL/cortexm0ds_logic.v(16362)
  not u20048 (Vbiow6, n5733);  // ../RTL/cortexm0ds_logic.v(16362)
  and u20049 (Y9apw6, Taapw6, Abapw6);  // ../RTL/cortexm0ds_logic.v(16363)
  and u2005 (n245, Uthpw6[10], Vk1iu6);  // ../RTL/cortexm0ds_logic.v(3824)
  and u20050 (n5734, Hbapw6, Hiaiu6);  // ../RTL/cortexm0ds_logic.v(16364)
  not u20051 (Abapw6, n5734);  // ../RTL/cortexm0ds_logic.v(16364)
  or u20052 (n5735, Iuniu6, Nlaiu6);  // ../RTL/cortexm0ds_logic.v(16365)
  not u20053 (Hbapw6, n5735);  // ../RTL/cortexm0ds_logic.v(16365)
  and u20054 (n5736, Ls1ju6, Md0iu6);  // ../RTL/cortexm0ds_logic.v(16366)
  not u20055 (Taapw6, n5736);  // ../RTL/cortexm0ds_logic.v(16366)
  or u20056 (n5737, Cyfpw6[0], Cyfpw6[4]);  // ../RTL/cortexm0ds_logic.v(16367)
  not u20057 (Md0iu6, n5737);  // ../RTL/cortexm0ds_logic.v(16367)
  and u20058 (Ls1ju6, Apaiu6, Jjhiu6);  // ../RTL/cortexm0ds_logic.v(16368)
  or u20059 (n5738, Jcaiu6, Sbghu6);  // ../RTL/cortexm0ds_logic.v(16369)
  not u2006 (Ut2iu6, n245);  // ../RTL/cortexm0ds_logic.v(3824)
  not u20060 (Apaiu6, n5738);  // ../RTL/cortexm0ds_logic.v(16369)
  and u20061 (n5739, Obapw6, Vbapw6);  // ../RTL/cortexm0ds_logic.v(16370)
  not u20062 (F3apw6, n5739);  // ../RTL/cortexm0ds_logic.v(16370)
  and u20063 (Vbapw6, Ccapw6, Jcapw6);  // ../RTL/cortexm0ds_logic.v(16371)
  or u20064 (n5740, Jf6ju6, Pthiu6);  // ../RTL/cortexm0ds_logic.v(16372)
  not u20065 (Jcapw6, n5740);  // ../RTL/cortexm0ds_logic.v(16372)
  and u20066 (Jf6ju6, Tr0iu6, Ii0iu6);  // ../RTL/cortexm0ds_logic.v(16373)
  and u20067 (Ccapw6, Qcapw6, Xcapw6);  // ../RTL/cortexm0ds_logic.v(16374)
  and u20068 (n5741, Edapw6, Owoiu6);  // ../RTL/cortexm0ds_logic.v(16375)
  not u20069 (Xcapw6, n5741);  // ../RTL/cortexm0ds_logic.v(16375)
  and u2007 (Gt2iu6, Bu2iu6, Iu2iu6);  // ../RTL/cortexm0ds_logic.v(3825)
  and u20070 (Owoiu6, Cyfpw6[3], Xe8iu6);  // ../RTL/cortexm0ds_logic.v(16376)
  and u20071 (n7[2], Auyhu6, Huyhu6);  // ../RTL/cortexm0ds_logic.v(3185)
  not u20072 (Edapw6, E0vow6);  // ../RTL/cortexm0ds_logic.v(16377)
  and u20073 (n5742, H4ghu6, Ldapw6);  // ../RTL/cortexm0ds_logic.v(16378)
  not u20074 (Qcapw6, n5742);  // ../RTL/cortexm0ds_logic.v(16378)
  or u20075 (Ldapw6, Cyfpw6[4], A3aju6);  // ../RTL/cortexm0ds_logic.v(16379)
  and u20076 (A3aju6, Cyfpw6[0], Cyfpw6[1]);  // ../RTL/cortexm0ds_logic.v(16380)
  and u20077 (Obapw6, Sdapw6, Zdapw6);  // ../RTL/cortexm0ds_logic.v(16381)
  and u20078 (Zdapw6, Geapw6, Wh7ju6);  // ../RTL/cortexm0ds_logic.v(16382)
  or u20079 (Wh7ju6, O60ju6, Cyfpw6[0]);  // ../RTL/cortexm0ds_logic.v(16383)
  and u2008 (n246, Iahpw6[9], Xl1iu6);  // ../RTL/cortexm0ds_logic.v(3826)
  not u20080 (O60ju6, Vjhow6);  // ../RTL/cortexm0ds_logic.v(16384)
  and u20081 (Vjhow6, H4ghu6, Cyfpw6[5]);  // ../RTL/cortexm0ds_logic.v(16385)
  or u20082 (Geapw6, Tfjiu6, Lkaiu6);  // ../RTL/cortexm0ds_logic.v(16386)
  and u20083 (Sdapw6, Cyfpw6[7], Neapw6);  // ../RTL/cortexm0ds_logic.v(16387)
  or u20084 (Neapw6, Qxaiu6, Tr0iu6);  // ../RTL/cortexm0ds_logic.v(16388)
  buf u20085 (Caehu6, Nxkbx6[33]);  // ../RTL/cortexm0ds_logic.v(3167)
  and u20086 (Ympiu6, Ueapw6, Bfapw6);  // ../RTL/cortexm0ds_logic.v(16390)
  not u20087 (Ob3pw6, Ympiu6);  // ../RTL/cortexm0ds_logic.v(16390)
  and u20088 (Bfapw6, Aphiu6, Ifapw6);  // ../RTL/cortexm0ds_logic.v(16391)
  and u20089 (n5743, Pfapw6, Srhiu6);  // ../RTL/cortexm0ds_logic.v(16392)
  not u2009 (Iu2iu6, n246);  // ../RTL/cortexm0ds_logic.v(3826)
  not u20090 (Ifapw6, n5743);  // ../RTL/cortexm0ds_logic.v(16392)
  and u20091 (Spcpw6, B7qow6, Et8iu6);  // ../RTL/cortexm0ds_logic.v(16393)
  not u20092 (Srhiu6, Spcpw6);  // ../RTL/cortexm0ds_logic.v(16393)
  AL_MUX u20093 (
    .i0(Wfapw6),
    .i1(Dgapw6),
    .sel(vis_pc_o[0]),
    .o(Pfapw6));  // ../RTL/cortexm0ds_logic.v(16394)
  and u20094 (Dgapw6, Kgapw6, Rgapw6);  // ../RTL/cortexm0ds_logic.v(16395)
  and u20095 (n5744, Juzhu6, Ophiu6);  // ../RTL/cortexm0ds_logic.v(16396)
  not u20096 (Rgapw6, n5744);  // ../RTL/cortexm0ds_logic.v(16396)
  and u20097 (n5745, Sufpw6[1], Ygapw6);  // ../RTL/cortexm0ds_logic.v(16397)
  not u20098 (Juzhu6, n5745);  // ../RTL/cortexm0ds_logic.v(16397)
  or u20099 (Kgapw6, Jjhiu6, Dxfhu6);  // ../RTL/cortexm0ds_logic.v(16398)
  buf u201 (Shhpw6[2], Bk7ax6);  // ../RTL/cortexm0ds_logic.v(1941)
  and u2010 (n247, Iahpw6[10], Z4yhu6);  // ../RTL/cortexm0ds_logic.v(3827)
  and u20100 (n5746, Ophiu6, N6piu6);  // ../RTL/cortexm0ds_logic.v(16399)
  not u20101 (Wfapw6, n5746);  // ../RTL/cortexm0ds_logic.v(16399)
  not u20102 (N6piu6, Pkciu6);  // ../RTL/cortexm0ds_logic.v(16400)
  and u20103 (Pkciu6, Sufpw6[0], Ygapw6);  // ../RTL/cortexm0ds_logic.v(16401)
  and u20104 (n5747, B7qow6, U6qow6);  // ../RTL/cortexm0ds_logic.v(16402)
  not u20105 (Ophiu6, n5747);  // ../RTL/cortexm0ds_logic.v(16402)
  not u20106 (U6qow6, Gu8iu6);  // ../RTL/cortexm0ds_logic.v(16403)
  and u20107 (Gu8iu6, Kgaiu6, Fhapw6);  // ../RTL/cortexm0ds_logic.v(16404)
  and u20108 (n5748, Yp8iu6, Hzziu6);  // ../RTL/cortexm0ds_logic.v(16405)
  not u20109 (Fhapw6, n5748);  // ../RTL/cortexm0ds_logic.v(16405)
  not u2011 (Bu2iu6, n247);  // ../RTL/cortexm0ds_logic.v(3827)
  and u20110 (Yp8iu6, Cyfpw6[5], Nlaiu6);  // ../RTL/cortexm0ds_logic.v(16406)
  not u20111 (Kgaiu6, Uoziu6);  // ../RTL/cortexm0ds_logic.v(16407)
  and u20112 (Uoziu6, L78ju6, Y7ghu6);  // ../RTL/cortexm0ds_logic.v(16408)
  and u20113 (Aphiu6, I1aiu6, Dp8iu6);  // ../RTL/cortexm0ds_logic.v(16409)
  buf u20114 (Eafpw6[31], Nxkbx6[32]);  // ../RTL/cortexm0ds_logic.v(3167)
  and u20115 (Dp8iu6, Mhapw6, Thapw6);  // ../RTL/cortexm0ds_logic.v(16411)
  not u20116 (LOCKUP, Dp8iu6);  // ../RTL/cortexm0ds_logic.v(16411)
  and u20117 (n5749, Aiapw6, H3aju6);  // ../RTL/cortexm0ds_logic.v(16412)
  not u20118 (Thapw6, n5749);  // ../RTL/cortexm0ds_logic.v(16412)
  and u20119 (Aiapw6, Mfjiu6, Sbghu6);  // ../RTL/cortexm0ds_logic.v(16413)
  and u2012 (n248, Pu2iu6, Wu2iu6);  // ../RTL/cortexm0ds_logic.v(3828)
  and u20120 (Mhapw6, Hiapw6, Oiapw6);  // ../RTL/cortexm0ds_logic.v(16414)
  and u20121 (n5750, Omyiu6, Viapw6);  // ../RTL/cortexm0ds_logic.v(16415)
  not u20122 (Oiapw6, n5750);  // ../RTL/cortexm0ds_logic.v(16415)
  and u20123 (n5751, Cjapw6, Jjapw6);  // ../RTL/cortexm0ds_logic.v(16416)
  not u20124 (Viapw6, n5751);  // ../RTL/cortexm0ds_logic.v(16416)
  and u20125 (n5752, Qjapw6, Xjapw6);  // ../RTL/cortexm0ds_logic.v(16417)
  not u20126 (Jjapw6, n5752);  // ../RTL/cortexm0ds_logic.v(16417)
  and u20127 (Xjapw6, Kxziu6, Kr7ow6);  // ../RTL/cortexm0ds_logic.v(16418)
  or u20128 (n5753, Vwaiu6, H4ghu6);  // ../RTL/cortexm0ds_logic.v(16419)
  not u20129 (Kr7ow6, n5753);  // ../RTL/cortexm0ds_logic.v(16419)
  not u2013 (Cwxhu6, n248);  // ../RTL/cortexm0ds_logic.v(3828)
  or u20130 (n5754, Ruaiu6, Wfoiu6);  // ../RTL/cortexm0ds_logic.v(16420)
  not u20131 (Qjapw6, n5754);  // ../RTL/cortexm0ds_logic.v(16420)
  not u20132 (Ruaiu6, V9ghu6);  // ../RTL/cortexm0ds_logic.v(16421)
  and u20133 (n5755, Ekapw6, Lkapw6);  // ../RTL/cortexm0ds_logic.v(16422)
  not u20134 (Cjapw6, n5755);  // ../RTL/cortexm0ds_logic.v(16422)
  or u20135 (n5756, Y7ghu6, H4ghu6);  // ../RTL/cortexm0ds_logic.v(16423)
  not u20136 (Lkapw6, n5756);  // ../RTL/cortexm0ds_logic.v(16423)
  or u20137 (n5757, Qjaiu6, Cyfpw6[5]);  // ../RTL/cortexm0ds_logic.v(16424)
  not u20138 (Ekapw6, n5757);  // ../RTL/cortexm0ds_logic.v(16424)
  and u20139 (n5758, V9ghu6, Skapw6);  // ../RTL/cortexm0ds_logic.v(16425)
  and u2014 (n249, Iahpw6[9], Z4yhu6);  // ../RTL/cortexm0ds_logic.v(3829)
  not u20140 (Hiapw6, n5758);  // ../RTL/cortexm0ds_logic.v(16425)
  and u20141 (n5759, Xxaiu6, Zkapw6);  // ../RTL/cortexm0ds_logic.v(16426)
  not u20142 (Skapw6, n5759);  // ../RTL/cortexm0ds_logic.v(16426)
  and u20143 (Xxaiu6, Glapw6, Nlapw6);  // ../RTL/cortexm0ds_logic.v(16427)
  and u20144 (Nlapw6, Ulapw6, Bmapw6);  // ../RTL/cortexm0ds_logic.v(16428)
  and u20145 (n5760, Imapw6, Buaow6);  // ../RTL/cortexm0ds_logic.v(16429)
  not u20146 (Bmapw6, n5760);  // ../RTL/cortexm0ds_logic.v(16429)
  or u20147 (n5761, Ntgiu6, P0biu6);  // ../RTL/cortexm0ds_logic.v(16430)
  not u20148 (Imapw6, n5761);  // ../RTL/cortexm0ds_logic.v(16430)
  and u20149 (P0biu6, Pmapw6, Wmapw6);  // ../RTL/cortexm0ds_logic.v(16431)
  not u2015 (Wu2iu6, n249);  // ../RTL/cortexm0ds_logic.v(3829)
  and u20150 (n5762, Dnapw6, Knapw6);  // ../RTL/cortexm0ds_logic.v(16432)
  not u20151 (Wmapw6, n5762);  // ../RTL/cortexm0ds_logic.v(16432)
  or u20152 (Knapw6, Sbrow6, B3gpw6[1]);  // ../RTL/cortexm0ds_logic.v(16433)
  and u20153 (Dnapw6, Rnapw6, Gcrow6);  // ../RTL/cortexm0ds_logic.v(16434)
  and u20154 (n5763, Ynapw6, Foapw6);  // ../RTL/cortexm0ds_logic.v(16435)
  not u20155 (Gcrow6, n5763);  // ../RTL/cortexm0ds_logic.v(16435)
  and u20156 (Foapw6, Moapw6, Toapw6);  // ../RTL/cortexm0ds_logic.v(16436)
  and u20157 (Toapw6, Apapw6, Hpapw6);  // ../RTL/cortexm0ds_logic.v(16437)
  and u20158 (Hpapw6, Opapw6, Vpapw6);  // ../RTL/cortexm0ds_logic.v(16438)
  and u20159 (Vpapw6, Cqapw6, Oyfiu6);  // ../RTL/cortexm0ds_logic.v(16439)
  and u2016 (Pu2iu6, Dv2iu6, Kv2iu6);  // ../RTL/cortexm0ds_logic.v(3830)
  or u20160 (n5764, Arfiu6, Ahbiu6);  // ../RTL/cortexm0ds_logic.v(16440)
  not u20161 (Cqapw6, n5764);  // ../RTL/cortexm0ds_logic.v(16440)
  or u20162 (n5765, Lhdiu6, Nbdiu6);  // ../RTL/cortexm0ds_logic.v(16441)
  not u20163 (Opapw6, n5765);  // ../RTL/cortexm0ds_logic.v(16441)
  and u20164 (Apapw6, Jqapw6, Qqapw6);  // ../RTL/cortexm0ds_logic.v(16442)
  or u20165 (n5766, Jndiu6, Kkdiu6);  // ../RTL/cortexm0ds_logic.v(16443)
  not u20166 (Qqapw6, n5766);  // ../RTL/cortexm0ds_logic.v(16443)
  or u20167 (n5767, V5giu6, Iqdiu6);  // ../RTL/cortexm0ds_logic.v(16444)
  not u20168 (Jqapw6, n5767);  // ../RTL/cortexm0ds_logic.v(16444)
  and u20169 (Moapw6, Xqapw6, Erapw6);  // ../RTL/cortexm0ds_logic.v(16445)
  and u2017 (n250, Uthpw6[9], Vk1iu6);  // ../RTL/cortexm0ds_logic.v(3831)
  and u20170 (Erapw6, Lrapw6, Srapw6);  // ../RTL/cortexm0ds_logic.v(16446)
  and u20171 (Srapw6, Zrapw6, Coxiu6);  // ../RTL/cortexm0ds_logic.v(16447)
  or u20172 (n5768, Bggiu6, Z7giu6);  // ../RTL/cortexm0ds_logic.v(16448)
  not u20173 (Zrapw6, n5768);  // ../RTL/cortexm0ds_logic.v(16448)
  or u20174 (n5769, Umgiu6, Odfiu6);  // ../RTL/cortexm0ds_logic.v(16449)
  not u20175 (Lrapw6, n5769);  // ../RTL/cortexm0ds_logic.v(16449)
  and u20176 (Xqapw6, Gsapw6, Nsapw6);  // ../RTL/cortexm0ds_logic.v(16450)
  or u20177 (n5770, Hl7iu6, Yogiu6);  // ../RTL/cortexm0ds_logic.v(16451)
  not u20178 (Nsapw6, n5770);  // ../RTL/cortexm0ds_logic.v(16451)
  or u20179 (n5771, Ajgiu6, Qrgiu6);  // ../RTL/cortexm0ds_logic.v(16452)
  not u2018 (Kv2iu6, n250);  // ../RTL/cortexm0ds_logic.v(3831)
  not u20180 (Gsapw6, n5771);  // ../RTL/cortexm0ds_logic.v(16452)
  and u20181 (Ynapw6, Usapw6, Btapw6);  // ../RTL/cortexm0ds_logic.v(16453)
  and u20182 (Btapw6, Itapw6, Ptapw6);  // ../RTL/cortexm0ds_logic.v(16454)
  and u20183 (Ptapw6, Wtapw6, Duapw6);  // ../RTL/cortexm0ds_logic.v(16455)
  and u20184 (Duapw6, Kuapw6, Giyiu6);  // ../RTL/cortexm0ds_logic.v(16456)
  or u20185 (n5772, Webiu6, Rhgiu6);  // ../RTL/cortexm0ds_logic.v(16457)
  not u20186 (Kuapw6, n5772);  // ../RTL/cortexm0ds_logic.v(16457)
  or u20187 (n5773, Ivfiu6, Etfiu6);  // ../RTL/cortexm0ds_logic.v(16458)
  not u20188 (Wtapw6, n5773);  // ../RTL/cortexm0ds_logic.v(16458)
  not u20189 (Ivfiu6, Ubyiu6);  // ../RTL/cortexm0ds_logic.v(16459)
  and u2019 (n251, Iahpw6[8], Xl1iu6);  // ../RTL/cortexm0ds_logic.v(3832)
  and u20190 (Itapw6, Ruapw6, Yuapw6);  // ../RTL/cortexm0ds_logic.v(16460)
  or u20191 (n5774, O8diu6, Mxfiu6);  // ../RTL/cortexm0ds_logic.v(16461)
  not u20192 (Yuapw6, n5774);  // ../RTL/cortexm0ds_logic.v(16461)
  or u20193 (n5775, N1giu6, Mediu6);  // ../RTL/cortexm0ds_logic.v(16462)
  not u20194 (Ruapw6, n5775);  // ../RTL/cortexm0ds_logic.v(16462)
  and u20195 (Usapw6, Fvapw6, Mvapw6);  // ../RTL/cortexm0ds_logic.v(16463)
  and u20196 (Mvapw6, Tvapw6, Awapw6);  // ../RTL/cortexm0ds_logic.v(16464)
  or u20197 (n5776, R3giu6, Hwhiu6);  // ../RTL/cortexm0ds_logic.v(16465)
  not u20198 (Awapw6, n5776);  // ../RTL/cortexm0ds_logic.v(16465)
  or u20199 (n5777, Hcgiu6, Dagiu6);  // ../RTL/cortexm0ds_logic.v(16466)
  buf u202 (vis_psp_o[7], O1jbx6);  // ../RTL/cortexm0ds_logic.v(2085)
  not u2020 (Dv2iu6, n251);  // ../RTL/cortexm0ds_logic.v(3832)
  not u20200 (Tvapw6, n5777);  // ../RTL/cortexm0ds_logic.v(16466)
  not u20201 (Hcgiu6, Spxiu6);  // ../RTL/cortexm0ds_logic.v(16467)
  and u20202 (Fvapw6, Hwapw6, Owapw6);  // ../RTL/cortexm0ds_logic.v(16468)
  or u20203 (n5778, G9fiu6, Eegiu6);  // ../RTL/cortexm0ds_logic.v(16469)
  not u20204 (Owapw6, n5778);  // ../RTL/cortexm0ds_logic.v(16469)
  or u20205 (n5779, Sffiu6, Kbfiu6);  // ../RTL/cortexm0ds_logic.v(16470)
  not u20206 (Hwapw6, n5779);  // ../RTL/cortexm0ds_logic.v(16470)
  and u20207 (n5780, Vwapw6, Cxapw6);  // ../RTL/cortexm0ds_logic.v(16471)
  not u20208 (Rnapw6, n5780);  // ../RTL/cortexm0ds_logic.v(16471)
  and u20209 (n5781, Sbrow6, B3gpw6[1]);  // ../RTL/cortexm0ds_logic.v(16472)
  and u2021 (n252, Rv2iu6, Yv2iu6);  // ../RTL/cortexm0ds_logic.v(3833)
  not u20210 (Cxapw6, n5781);  // ../RTL/cortexm0ds_logic.v(16472)
  and u20211 (Sbrow6, Jxapw6, Qxapw6);  // ../RTL/cortexm0ds_logic.v(16473)
  and u20212 (Qxapw6, Xxapw6, Eyapw6);  // ../RTL/cortexm0ds_logic.v(16474)
  and u20213 (Eyapw6, Lyapw6, Syapw6);  // ../RTL/cortexm0ds_logic.v(16475)
  and u20214 (Syapw6, Zyapw6, Gzapw6);  // ../RTL/cortexm0ds_logic.v(16476)
  and u20215 (Gzapw6, Nzapw6, Uzapw6);  // ../RTL/cortexm0ds_logic.v(16477)
  and u20216 (n5782, B3gpw6[1], Qrgiu6);  // ../RTL/cortexm0ds_logic.v(16478)
  not u20217 (Uzapw6, n5782);  // ../RTL/cortexm0ds_logic.v(16478)
  and u20218 (Nzapw6, B0bpw6, I0bpw6);  // ../RTL/cortexm0ds_logic.v(16479)
  and u20219 (n5783, L1gpw6[1], Rhgiu6);  // ../RTL/cortexm0ds_logic.v(16480)
  not u2022 (Vvxhu6, n252);  // ../RTL/cortexm0ds_logic.v(3833)
  not u20220 (I0bpw6, n5783);  // ../RTL/cortexm0ds_logic.v(16480)
  and u20221 (n5784, H8gpw6[1], Ajgiu6);  // ../RTL/cortexm0ds_logic.v(16481)
  not u20222 (B0bpw6, n5784);  // ../RTL/cortexm0ds_logic.v(16481)
  and u20223 (Zyapw6, P0bpw6, W0bpw6);  // ../RTL/cortexm0ds_logic.v(16482)
  or u20224 (W0bpw6, U2uow6, Ucxiu6);  // ../RTL/cortexm0ds_logic.v(16483)
  not u20225 (U2uow6, R4gpw6[1]);  // ../RTL/cortexm0ds_logic.v(16484)
  and u20226 (n5785, R4gpw6[3], Yogiu6);  // ../RTL/cortexm0ds_logic.v(16485)
  not u20227 (P0bpw6, n5785);  // ../RTL/cortexm0ds_logic.v(16485)
  and u20228 (Lyapw6, D1bpw6, K1bpw6);  // ../RTL/cortexm0ds_logic.v(16486)
  and u20229 (K1bpw6, R1bpw6, Y1bpw6);  // ../RTL/cortexm0ds_logic.v(16487)
  and u2023 (n253, Iahpw6[8], Z4yhu6);  // ../RTL/cortexm0ds_logic.v(3834)
  or u20230 (Y1bpw6, Fytow6, Agxiu6);  // ../RTL/cortexm0ds_logic.v(16488)
  not u20231 (Fytow6, R4gpw6[5]);  // ../RTL/cortexm0ds_logic.v(16489)
  or u20232 (R1bpw6, Yxtow6, Qhxiu6);  // ../RTL/cortexm0ds_logic.v(16490)
  not u20233 (Qhxiu6, Sffiu6);  // ../RTL/cortexm0ds_logic.v(16491)
  not u20234 (Yxtow6, R4gpw6[7]);  // ../RTL/cortexm0ds_logic.v(16492)
  and u20235 (D1bpw6, F2bpw6, M2bpw6);  // ../RTL/cortexm0ds_logic.v(16493)
  and u20236 (n5786, R4gpw6[9], Odfiu6);  // ../RTL/cortexm0ds_logic.v(16494)
  not u20237 (M2bpw6, n5786);  // ../RTL/cortexm0ds_logic.v(16494)
  or u20238 (F2bpw6, Yqtow6, Wkxiu6);  // ../RTL/cortexm0ds_logic.v(16495)
  not u20239 (Wkxiu6, Kbfiu6);  // ../RTL/cortexm0ds_logic.v(16496)
  not u2024 (Yv2iu6, n253);  // ../RTL/cortexm0ds_logic.v(3834)
  not u20240 (Yqtow6, R4gpw6[11]);  // ../RTL/cortexm0ds_logic.v(16497)
  and u20241 (Xxapw6, T2bpw6, A3bpw6);  // ../RTL/cortexm0ds_logic.v(16498)
  and u20242 (A3bpw6, H3bpw6, O3bpw6);  // ../RTL/cortexm0ds_logic.v(16499)
  and u20243 (O3bpw6, V3bpw6, C4bpw6);  // ../RTL/cortexm0ds_logic.v(16500)
  or u20244 (C4bpw6, Mrtow6, Mmxiu6);  // ../RTL/cortexm0ds_logic.v(16501)
  buf u20245 (Eafpw6[30], Nxkbx6[31]);  // ../RTL/cortexm0ds_logic.v(3167)
  not u20246 (Mrtow6, R4gpw6[13]);  // ../RTL/cortexm0ds_logic.v(16503)
  and u20247 (V3bpw6, J4bpw6, Q4bpw6);  // ../RTL/cortexm0ds_logic.v(16504)
  or u20248 (Q4bpw6, Frtow6, Coxiu6);  // ../RTL/cortexm0ds_logic.v(16505)
  not u20249 (Frtow6, R4gpw6[15]);  // ../RTL/cortexm0ds_logic.v(16506)
  and u2025 (Rv2iu6, Fw2iu6, Mw2iu6);  // ../RTL/cortexm0ds_logic.v(3835)
  or u20250 (J4bpw6, Xluow6, Gfgiu6);  // ../RTL/cortexm0ds_logic.v(16507)
  not u20251 (Xluow6, R4gpw6[17]);  // ../RTL/cortexm0ds_logic.v(16508)
  and u20252 (H3bpw6, X4bpw6, E5bpw6);  // ../RTL/cortexm0ds_logic.v(16509)
  or u20253 (E5bpw6, Qluow6, Jdgiu6);  // ../RTL/cortexm0ds_logic.v(16510)
  not u20254 (Qluow6, R4gpw6[19]);  // ../RTL/cortexm0ds_logic.v(16511)
  or u20255 (X4bpw6, Pouow6, Spxiu6);  // ../RTL/cortexm0ds_logic.v(16512)
  not u20256 (Pouow6, R4gpw6[21]);  // ../RTL/cortexm0ds_logic.v(16513)
  and u20257 (T2bpw6, L5bpw6, S5bpw6);  // ../RTL/cortexm0ds_logic.v(16514)
  and u20258 (S5bpw6, Z5bpw6, G6bpw6);  // ../RTL/cortexm0ds_logic.v(16515)
  or u20259 (G6bpw6, Wouow6, Irxiu6);  // ../RTL/cortexm0ds_logic.v(16516)
  and u2026 (n254, Uthpw6[8], Vk1iu6);  // ../RTL/cortexm0ds_logic.v(3836)
  not u20260 (Wouow6, R4gpw6[23]);  // ../RTL/cortexm0ds_logic.v(16517)
  and u20261 (n5787, R4gpw6[25], Z7giu6);  // ../RTL/cortexm0ds_logic.v(16518)
  not u20262 (Z5bpw6, n5787);  // ../RTL/cortexm0ds_logic.v(16518)
  and u20263 (L5bpw6, N6bpw6, U6bpw6);  // ../RTL/cortexm0ds_logic.v(16519)
  or u20264 (U6bpw6, Ihuow6, Ouxiu6);  // ../RTL/cortexm0ds_logic.v(16520)
  not u20265 (Ihuow6, R4gpw6[27]);  // ../RTL/cortexm0ds_logic.v(16521)
  and u20266 (n5788, R4gpw6[29], R3giu6);  // ../RTL/cortexm0ds_logic.v(16522)
  not u20267 (N6bpw6, n5788);  // ../RTL/cortexm0ds_logic.v(16522)
  and u20268 (Jxapw6, B7bpw6, I7bpw6);  // ../RTL/cortexm0ds_logic.v(16523)
  and u20269 (I7bpw6, P7bpw6, W7bpw6);  // ../RTL/cortexm0ds_logic.v(16524)
  not u2027 (Mw2iu6, n254);  // ../RTL/cortexm0ds_logic.v(3836)
  and u20270 (W7bpw6, D8bpw6, K8bpw6);  // ../RTL/cortexm0ds_logic.v(16525)
  and u20271 (K8bpw6, R8bpw6, Y8bpw6);  // ../RTL/cortexm0ds_logic.v(16526)
  or u20272 (Y8bpw6, Mcuow6, Nxxiu6);  // ../RTL/cortexm0ds_logic.v(16527)
  not u20273 (Mcuow6, R4gpw6[31]);  // ../RTL/cortexm0ds_logic.v(16528)
  and u20274 (R8bpw6, F9bpw6, M9bpw6);  // ../RTL/cortexm0ds_logic.v(16529)
  and u20275 (n5789, R4gpw6[33], Hwhiu6);  // ../RTL/cortexm0ds_logic.v(16530)
  not u20276 (M9bpw6, n5789);  // ../RTL/cortexm0ds_logic.v(16530)
  or u20277 (F9bpw6, Dksow6, M0yiu6);  // ../RTL/cortexm0ds_logic.v(16531)
  not u20278 (M0yiu6, Iqdiu6);  // ../RTL/cortexm0ds_logic.v(16532)
  not u20279 (Dksow6, R4gpw6[35]);  // ../RTL/cortexm0ds_logic.v(16533)
  and u2028 (n255, Iahpw6[7], Xl1iu6);  // ../RTL/cortexm0ds_logic.v(3837)
  and u20280 (D8bpw6, T9bpw6, Aabpw6);  // ../RTL/cortexm0ds_logic.v(16534)
  or u20281 (Aabpw6, Ehsow6, C2yiu6);  // ../RTL/cortexm0ds_logic.v(16535)
  not u20282 (C2yiu6, Jndiu6);  // ../RTL/cortexm0ds_logic.v(16536)
  not u20283 (Ehsow6, R4gpw6[37]);  // ../RTL/cortexm0ds_logic.v(16537)
  and u20284 (n5790, R4gpw6[39], Kkdiu6);  // ../RTL/cortexm0ds_logic.v(16538)
  not u20285 (T9bpw6, n5790);  // ../RTL/cortexm0ds_logic.v(16538)
  and u20286 (P7bpw6, Habpw6, Oabpw6);  // ../RTL/cortexm0ds_logic.v(16539)
  and u20287 (Oabpw6, Vabpw6, Cbbpw6);  // ../RTL/cortexm0ds_logic.v(16540)
  and u20288 (n5791, R4gpw6[41], Lhdiu6);  // ../RTL/cortexm0ds_logic.v(16541)
  not u20289 (Cbbpw6, n5791);  // ../RTL/cortexm0ds_logic.v(16541)
  not u2029 (Fw2iu6, n255);  // ../RTL/cortexm0ds_logic.v(3837)
  or u20290 (Vabpw6, Q9sow6, Y6yiu6);  // ../RTL/cortexm0ds_logic.v(16542)
  not u20291 (Y6yiu6, Mediu6);  // ../RTL/cortexm0ds_logic.v(16543)
  not u20292 (Q9sow6, R4gpw6[43]);  // ../RTL/cortexm0ds_logic.v(16544)
  and u20293 (Habpw6, Jbbpw6, Qbbpw6);  // ../RTL/cortexm0ds_logic.v(16545)
  or u20294 (Qbbpw6, Ubsow6, O8yiu6);  // ../RTL/cortexm0ds_logic.v(16546)
  buf u20295 (Eafpw6[29], Nxkbx6[30]);  // ../RTL/cortexm0ds_logic.v(3167)
  not u20296 (Ubsow6, R4gpw6[45]);  // ../RTL/cortexm0ds_logic.v(16548)
  and u20297 (n5792, R4gpw6[47], O8diu6);  // ../RTL/cortexm0ds_logic.v(16549)
  not u20298 (Jbbpw6, n5792);  // ../RTL/cortexm0ds_logic.v(16549)
  and u20299 (B7bpw6, Xbbpw6, Ecbpw6);  // ../RTL/cortexm0ds_logic.v(16550)
  buf u203 (vis_r4_o[13], V9vax6);  // ../RTL/cortexm0ds_logic.v(2626)
  AL_MUX u2030 (
    .i0(SWDITMS),
    .i1(Mdhpw6[3]),
    .sel(Tw2iu6),
    .o(Ovxhu6));  // ../RTL/cortexm0ds_logic.v(3838)
  and u20300 (Ecbpw6, Lcbpw6, Scbpw6);  // ../RTL/cortexm0ds_logic.v(16551)
  and u20301 (Scbpw6, Zcbpw6, Gdbpw6);  // ../RTL/cortexm0ds_logic.v(16552)
  or u20302 (Gdbpw6, Otsow6, Oyfiu6);  // ../RTL/cortexm0ds_logic.v(16553)
  not u20303 (Otsow6, R4gpw6[49]);  // ../RTL/cortexm0ds_logic.v(16554)
  or u20304 (Zcbpw6, Htsow6, Rwfiu6);  // ../RTL/cortexm0ds_logic.v(16555)
  not u20305 (Htsow6, R4gpw6[51]);  // ../RTL/cortexm0ds_logic.v(16556)
  and u20306 (Lcbpw6, Ndbpw6, Udbpw6);  // ../RTL/cortexm0ds_logic.v(16557)
  or u20307 (Udbpw6, Vtsow6, Ubyiu6);  // ../RTL/cortexm0ds_logic.v(16558)
  not u20308 (Vtsow6, R4gpw6[53]);  // ../RTL/cortexm0ds_logic.v(16559)
  or u20309 (Ndbpw6, Cusow6, Kdyiu6);  // ../RTL/cortexm0ds_logic.v(16560)
  and u2031 (Tw2iu6, Ax2iu6, Hx2iu6);  // ../RTL/cortexm0ds_logic.v(3839)
  not u20310 (Cusow6, R4gpw6[55]);  // ../RTL/cortexm0ds_logic.v(16561)
  and u20311 (Xbbpw6, Bebpw6, Iebpw6);  // ../RTL/cortexm0ds_logic.v(16562)
  and u20312 (Iebpw6, Pebpw6, Webpw6);  // ../RTL/cortexm0ds_logic.v(16563)
  and u20313 (n5793, R4gpw6[57], Arfiu6);  // ../RTL/cortexm0ds_logic.v(16564)
  not u20314 (Webpw6, n5793);  // ../RTL/cortexm0ds_logic.v(16564)
  or u20315 (Pebpw6, V7tow6, Qgyiu6);  // ../RTL/cortexm0ds_logic.v(16565)
  not u20316 (V7tow6, R4gpw6[59]);  // ../RTL/cortexm0ds_logic.v(16566)
  and u20317 (Bebpw6, Dfbpw6, Kfbpw6);  // ../RTL/cortexm0ds_logic.v(16567)
  or u20318 (Kfbpw6, E2tow6, Giyiu6);  // ../RTL/cortexm0ds_logic.v(16568)
  not u20319 (Giyiu6, Lyhiu6);  // ../RTL/cortexm0ds_logic.v(16569)
  and u2032 (Hx2iu6, Ox2iu6, Vx2iu6);  // ../RTL/cortexm0ds_logic.v(3840)
  not u20320 (E2tow6, R4gpw6[61]);  // ../RTL/cortexm0ds_logic.v(16570)
  and u20321 (n5794, R4gpw6[63], Webiu6);  // ../RTL/cortexm0ds_logic.v(16571)
  not u20322 (Dfbpw6, n5794);  // ../RTL/cortexm0ds_logic.v(16571)
  and u20323 (Vwapw6, Idrow6, Xglow6);  // ../RTL/cortexm0ds_logic.v(16572)
  not u20324 (Xglow6, B3gpw6[0]);  // ../RTL/cortexm0ds_logic.v(16573)
  and u20325 (n5795, Rfbpw6, Yfbpw6);  // ../RTL/cortexm0ds_logic.v(16574)
  not u20326 (Idrow6, n5795);  // ../RTL/cortexm0ds_logic.v(16574)
  and u20327 (Yfbpw6, Fgbpw6, Mgbpw6);  // ../RTL/cortexm0ds_logic.v(16575)
  and u20328 (Mgbpw6, Tgbpw6, Ahbpw6);  // ../RTL/cortexm0ds_logic.v(16576)
  and u20329 (Ahbpw6, Hhbpw6, Ohbpw6);  // ../RTL/cortexm0ds_logic.v(16577)
  and u2033 (n256, Cy2iu6, Ujyhu6);  // ../RTL/cortexm0ds_logic.v(3841)
  and u20330 (Ohbpw6, Vhbpw6, Cibpw6);  // ../RTL/cortexm0ds_logic.v(16578)
  and u20331 (n5796, B3gpw6[0], Qrgiu6);  // ../RTL/cortexm0ds_logic.v(16579)
  not u20332 (Cibpw6, n5796);  // ../RTL/cortexm0ds_logic.v(16579)
  and u20333 (Qrgiu6, F8row6, Jibpw6);  // ../RTL/cortexm0ds_logic.v(16580)
  and u20334 (Vhbpw6, Qibpw6, Xibpw6);  // ../RTL/cortexm0ds_logic.v(16581)
  and u20335 (n5797, L1gpw6[0], Rhgiu6);  // ../RTL/cortexm0ds_logic.v(16582)
  not u20336 (Xibpw6, n5797);  // ../RTL/cortexm0ds_logic.v(16582)
  and u20337 (Rhgiu6, Ejbpw6, A9row6);  // ../RTL/cortexm0ds_logic.v(16583)
  and u20338 (Ejbpw6, Ljbpw6, H9row6);  // ../RTL/cortexm0ds_logic.v(16584)
  and u20339 (n5798, H8gpw6[0], Ajgiu6);  // ../RTL/cortexm0ds_logic.v(16585)
  not u2034 (Ox2iu6, n256);  // ../RTL/cortexm0ds_logic.v(3841)
  not u20340 (Qibpw6, n5798);  // ../RTL/cortexm0ds_logic.v(16585)
  and u20341 (Ajgiu6, F8row6, Ljbpw6);  // ../RTL/cortexm0ds_logic.v(16586)
  and u20342 (F8row6, Sjbpw6, H9row6);  // ../RTL/cortexm0ds_logic.v(16587)
  and u20343 (Hhbpw6, Zjbpw6, Gkbpw6);  // ../RTL/cortexm0ds_logic.v(16588)
  or u20344 (Gkbpw6, B3uow6, Ucxiu6);  // ../RTL/cortexm0ds_logic.v(16589)
  not u20345 (Ucxiu6, Hl7iu6);  // ../RTL/cortexm0ds_logic.v(16590)
  and u20346 (Hl7iu6, Nkbpw6, Ukbpw6);  // ../RTL/cortexm0ds_logic.v(16591)
  not u20347 (B3uow6, R4gpw6[0]);  // ../RTL/cortexm0ds_logic.v(16592)
  and u20348 (n5799, R4gpw6[2], Yogiu6);  // ../RTL/cortexm0ds_logic.v(16593)
  not u20349 (Zjbpw6, n5799);  // ../RTL/cortexm0ds_logic.v(16593)
  or u2035 (Cy2iu6, Jy2iu6, Qy2iu6);  // ../RTL/cortexm0ds_logic.v(3842)
  or u20350 (Kexiu6, Blbpw6, Ilbpw6);  // ../RTL/cortexm0ds_logic.v(16594)
  not u20351 (Yogiu6, Kexiu6);  // ../RTL/cortexm0ds_logic.v(16594)
  and u20352 (Tgbpw6, Plbpw6, Wlbpw6);  // ../RTL/cortexm0ds_logic.v(16595)
  and u20353 (Wlbpw6, Dmbpw6, Kmbpw6);  // ../RTL/cortexm0ds_logic.v(16596)
  or u20354 (Kmbpw6, J0uow6, Agxiu6);  // ../RTL/cortexm0ds_logic.v(16597)
  not u20355 (Agxiu6, Umgiu6);  // ../RTL/cortexm0ds_logic.v(16598)
  and u20356 (Umgiu6, Nkbpw6, A9row6);  // ../RTL/cortexm0ds_logic.v(16599)
  not u20357 (J0uow6, R4gpw6[4]);  // ../RTL/cortexm0ds_logic.v(16600)
  and u20358 (n5800, R4gpw6[6], Sffiu6);  // ../RTL/cortexm0ds_logic.v(16601)
  not u20359 (Dmbpw6, n5800);  // ../RTL/cortexm0ds_logic.v(16601)
  AL_MUX u2036 (
    .i0(Xy2iu6),
    .i1(Iyyhu6),
    .sel(Ighpw6[1]),
    .o(Qy2iu6));  // ../RTL/cortexm0ds_logic.v(3843)
  and u20360 (Sffiu6, Nkbpw6, Sjbpw6);  // ../RTL/cortexm0ds_logic.v(16602)
  buf u20361 (Eafpw6[28], Nxkbx6[29]);  // ../RTL/cortexm0ds_logic.v(3167)
  and u20362 (Nkbpw6, Rmbpw6, M8row6);  // ../RTL/cortexm0ds_logic.v(16604)
  not u20363 (Blbpw6, Nkbpw6);  // ../RTL/cortexm0ds_logic.v(16604)
  and u20364 (Plbpw6, Ymbpw6, Fnbpw6);  // ../RTL/cortexm0ds_logic.v(16605)
  and u20365 (n5801, R4gpw6[8], Odfiu6);  // ../RTL/cortexm0ds_logic.v(16606)
  not u20366 (Fnbpw6, n5801);  // ../RTL/cortexm0ds_logic.v(16606)
  or u20367 (Gjxiu6, Mnbpw6, Tnbpw6);  // ../RTL/cortexm0ds_logic.v(16607)
  not u20368 (Odfiu6, Gjxiu6);  // ../RTL/cortexm0ds_logic.v(16607)
  and u20369 (n5802, R4gpw6[10], Kbfiu6);  // ../RTL/cortexm0ds_logic.v(16608)
  and u2037 (Xy2iu6, Ez2iu6, Lz2iu6);  // ../RTL/cortexm0ds_logic.v(3844)
  not u20370 (Ymbpw6, n5802);  // ../RTL/cortexm0ds_logic.v(16608)
  and u20371 (Kbfiu6, Aobpw6, Hobpw6);  // ../RTL/cortexm0ds_logic.v(16609)
  and u20372 (Fgbpw6, Oobpw6, Vobpw6);  // ../RTL/cortexm0ds_logic.v(16610)
  and u20373 (Vobpw6, Cpbpw6, Jpbpw6);  // ../RTL/cortexm0ds_logic.v(16611)
  and u20374 (Jpbpw6, Qpbpw6, Xpbpw6);  // ../RTL/cortexm0ds_logic.v(16612)
  and u20375 (n5803, R4gpw6[12], G9fiu6);  // ../RTL/cortexm0ds_logic.v(16613)
  not u20376 (Xpbpw6, n5803);  // ../RTL/cortexm0ds_logic.v(16613)
  or u20377 (Mmxiu6, Mnbpw6, Eqbpw6);  // ../RTL/cortexm0ds_logic.v(16614)
  not u20378 (G9fiu6, Mmxiu6);  // ../RTL/cortexm0ds_logic.v(16614)
  not u20379 (Mnbpw6, Aobpw6);  // ../RTL/cortexm0ds_logic.v(16615)
  and u2038 (n257, Wdyhu6, Sz2iu6);  // ../RTL/cortexm0ds_logic.v(3845)
  and u20380 (Qpbpw6, Lqbpw6, Sqbpw6);  // ../RTL/cortexm0ds_logic.v(16616)
  or u20381 (Sqbpw6, Qttow6, Coxiu6);  // ../RTL/cortexm0ds_logic.v(16617)
  not u20382 (Coxiu6, C7fiu6);  // ../RTL/cortexm0ds_logic.v(16618)
  and u20383 (C7fiu6, Aobpw6, Sjbpw6);  // ../RTL/cortexm0ds_logic.v(16619)
  and u20384 (Aobpw6, Zqbpw6, Rmbpw6);  // ../RTL/cortexm0ds_logic.v(16620)
  not u20385 (Qttow6, R4gpw6[14]);  // ../RTL/cortexm0ds_logic.v(16621)
  or u20386 (Lqbpw6, Iouow6, Gfgiu6);  // ../RTL/cortexm0ds_logic.v(16622)
  buf u20387 (Eafpw6[27], Nxkbx6[28]);  // ../RTL/cortexm0ds_logic.v(3167)
  or u20388 (Gfgiu6, Grbpw6, Tnbpw6);  // ../RTL/cortexm0ds_logic.v(16624)
  not u20389 (Bggiu6, Gfgiu6);  // ../RTL/cortexm0ds_logic.v(16624)
  not u2039 (Lz2iu6, n257);  // ../RTL/cortexm0ds_logic.v(3845)
  not u20390 (Iouow6, R4gpw6[16]);  // ../RTL/cortexm0ds_logic.v(16625)
  and u20391 (Cpbpw6, Nrbpw6, Urbpw6);  // ../RTL/cortexm0ds_logic.v(16626)
  and u20392 (n5804, R4gpw6[18], Eegiu6);  // ../RTL/cortexm0ds_logic.v(16627)
  not u20393 (Urbpw6, n5804);  // ../RTL/cortexm0ds_logic.v(16627)
  not u20394 (Eegiu6, Jdgiu6);  // ../RTL/cortexm0ds_logic.v(16628)
  or u20395 (Jdgiu6, Grbpw6, Ilbpw6);  // ../RTL/cortexm0ds_logic.v(16629)
  or u20396 (Nrbpw6, Aruow6, Spxiu6);  // ../RTL/cortexm0ds_logic.v(16630)
  or u20397 (Spxiu6, Grbpw6, Eqbpw6);  // ../RTL/cortexm0ds_logic.v(16631)
  not u20398 (Aruow6, R4gpw6[20]);  // ../RTL/cortexm0ds_logic.v(16632)
  and u20399 (Oobpw6, Bsbpw6, Isbpw6);  // ../RTL/cortexm0ds_logic.v(16633)
  buf u204 (vis_r14_o[10], N7oax6);  // ../RTL/cortexm0ds_logic.v(2497)
  or u2040 (Sz2iu6, Mdhpw6[0], Ighpw6[0]);  // ../RTL/cortexm0ds_logic.v(3846)
  and u20400 (Isbpw6, Psbpw6, Wsbpw6);  // ../RTL/cortexm0ds_logic.v(16634)
  and u20401 (n5805, R4gpw6[22], Dagiu6);  // ../RTL/cortexm0ds_logic.v(16635)
  not u20402 (Wsbpw6, n5805);  // ../RTL/cortexm0ds_logic.v(16635)
  not u20403 (Dagiu6, Irxiu6);  // ../RTL/cortexm0ds_logic.v(16636)
  or u20404 (Irxiu6, Grbpw6, Dtbpw6);  // ../RTL/cortexm0ds_logic.v(16637)
  and u20405 (n5806, Rmbpw6, Jibpw6);  // ../RTL/cortexm0ds_logic.v(16638)
  not u20406 (Grbpw6, n5806);  // ../RTL/cortexm0ds_logic.v(16638)
  and u20407 (n5807, R4gpw6[24], Z7giu6);  // ../RTL/cortexm0ds_logic.v(16639)
  not u20408 (Psbpw6, n5807);  // ../RTL/cortexm0ds_logic.v(16639)
  buf u20409 (Eafpw6[26], Nxkbx6[27]);  // ../RTL/cortexm0ds_logic.v(3167)
  and u2041 (n258, Zz2iu6, G03iu6);  // ../RTL/cortexm0ds_logic.v(3847)
  and u20410 (Z7giu6, Ktbpw6, Rmbpw6);  // ../RTL/cortexm0ds_logic.v(16641)
  not u20411 (Ysxiu6, Z7giu6);  // ../RTL/cortexm0ds_logic.v(16641)
  and u20412 (Ktbpw6, Ljbpw6, Ukbpw6);  // ../RTL/cortexm0ds_logic.v(16642)
  and u20413 (Bsbpw6, Rtbpw6, Ytbpw6);  // ../RTL/cortexm0ds_logic.v(16643)
  and u20414 (n5808, R4gpw6[26], V5giu6);  // ../RTL/cortexm0ds_logic.v(16644)
  not u20415 (Ytbpw6, n5808);  // ../RTL/cortexm0ds_logic.v(16644)
  buf u20416 (Eafpw6[25], Nxkbx6[26]);  // ../RTL/cortexm0ds_logic.v(3167)
  and u20417 (V5giu6, Fubpw6, Rmbpw6);  // ../RTL/cortexm0ds_logic.v(16646)
  not u20418 (Ouxiu6, V5giu6);  // ../RTL/cortexm0ds_logic.v(16646)
  and u20419 (Fubpw6, Ljbpw6, Hobpw6);  // ../RTL/cortexm0ds_logic.v(16647)
  not u2042 (Jy2iu6, n258);  // ../RTL/cortexm0ds_logic.v(3847)
  and u20420 (n5809, R4gpw6[28], R3giu6);  // ../RTL/cortexm0ds_logic.v(16648)
  not u20421 (Rtbpw6, n5809);  // ../RTL/cortexm0ds_logic.v(16648)
  and u20422 (R3giu6, Mubpw6, Rmbpw6);  // ../RTL/cortexm0ds_logic.v(16649)
  and u20423 (Mubpw6, A9row6, Ljbpw6);  // ../RTL/cortexm0ds_logic.v(16650)
  and u20424 (Rfbpw6, Tubpw6, Avbpw6);  // ../RTL/cortexm0ds_logic.v(16651)
  and u20425 (Avbpw6, Hvbpw6, Ovbpw6);  // ../RTL/cortexm0ds_logic.v(16652)
  and u20426 (Ovbpw6, Vvbpw6, Cwbpw6);  // ../RTL/cortexm0ds_logic.v(16653)
  and u20427 (Cwbpw6, Jwbpw6, Qwbpw6);  // ../RTL/cortexm0ds_logic.v(16654)
  and u20428 (n5810, R4gpw6[30], N1giu6);  // ../RTL/cortexm0ds_logic.v(16655)
  not u20429 (Qwbpw6, n5810);  // ../RTL/cortexm0ds_logic.v(16655)
  and u2043 (n259, N03iu6, Ighpw6[2]);  // ../RTL/cortexm0ds_logic.v(3848)
  buf u20430 (Eafpw6[24], Nxkbx6[25]);  // ../RTL/cortexm0ds_logic.v(3167)
  and u20431 (N1giu6, Xwbpw6, Rmbpw6);  // ../RTL/cortexm0ds_logic.v(16657)
  not u20432 (Nxxiu6, N1giu6);  // ../RTL/cortexm0ds_logic.v(16657)
  and u20433 (Rmbpw6, vis_ipsr_o[4], Vhbiu6);  // ../RTL/cortexm0ds_logic.v(16658)
  and u20434 (Xwbpw6, Sjbpw6, Ljbpw6);  // ../RTL/cortexm0ds_logic.v(16659)
  and u20435 (Jwbpw6, Exbpw6, Lxbpw6);  // ../RTL/cortexm0ds_logic.v(16660)
  and u20436 (n5811, R4gpw6[32], Hwhiu6);  // ../RTL/cortexm0ds_logic.v(16661)
  not u20437 (Lxbpw6, n5811);  // ../RTL/cortexm0ds_logic.v(16661)
  or u20438 (n5812, Sxbpw6, Tnbpw6);  // ../RTL/cortexm0ds_logic.v(16662)
  not u20439 (Hwhiu6, n5812);  // ../RTL/cortexm0ds_logic.v(16662)
  not u2044 (G03iu6, n259);  // ../RTL/cortexm0ds_logic.v(3848)
  and u20440 (n5813, R4gpw6[34], Iqdiu6);  // ../RTL/cortexm0ds_logic.v(16663)
  not u20441 (Exbpw6, n5813);  // ../RTL/cortexm0ds_logic.v(16663)
  and u20442 (Iqdiu6, Zxbpw6, Hobpw6);  // ../RTL/cortexm0ds_logic.v(16664)
  and u20443 (Vvbpw6, Gybpw6, Nybpw6);  // ../RTL/cortexm0ds_logic.v(16665)
  and u20444 (n5814, R4gpw6[36], Jndiu6);  // ../RTL/cortexm0ds_logic.v(16666)
  not u20445 (Nybpw6, n5814);  // ../RTL/cortexm0ds_logic.v(16666)
  and u20446 (Jndiu6, Zxbpw6, A9row6);  // ../RTL/cortexm0ds_logic.v(16667)
  or u20447 (Gybpw6, Lhsow6, S3yiu6);  // ../RTL/cortexm0ds_logic.v(16668)
  not u20448 (S3yiu6, Kkdiu6);  // ../RTL/cortexm0ds_logic.v(16669)
  and u20449 (Kkdiu6, Sjbpw6, Zxbpw6);  // ../RTL/cortexm0ds_logic.v(16670)
  and u2045 (N03iu6, Gjyhu6, Eiyhu6);  // ../RTL/cortexm0ds_logic.v(3849)
  buf u20450 (Eafpw6[23], Nxkbx6[24]);  // ../RTL/cortexm0ds_logic.v(3167)
  and u20451 (Zxbpw6, Uybpw6, M8row6);  // ../RTL/cortexm0ds_logic.v(16672)
  not u20452 (Sxbpw6, Zxbpw6);  // ../RTL/cortexm0ds_logic.v(16672)
  not u20453 (Lhsow6, R4gpw6[38]);  // ../RTL/cortexm0ds_logic.v(16673)
  and u20454 (Hvbpw6, Bzbpw6, Izbpw6);  // ../RTL/cortexm0ds_logic.v(16674)
  and u20455 (Izbpw6, Pzbpw6, Wzbpw6);  // ../RTL/cortexm0ds_logic.v(16675)
  and u20456 (n5815, R4gpw6[40], Lhdiu6);  // ../RTL/cortexm0ds_logic.v(16676)
  not u20457 (Wzbpw6, n5815);  // ../RTL/cortexm0ds_logic.v(16676)
  or u20458 (I5yiu6, D0cpw6, Tnbpw6);  // ../RTL/cortexm0ds_logic.v(16677)
  not u20459 (Lhdiu6, I5yiu6);  // ../RTL/cortexm0ds_logic.v(16677)
  or u2046 (Zz2iu6, Deyhu6, Ighpw6[3]);  // ../RTL/cortexm0ds_logic.v(3850)
  and u20460 (n5816, R4gpw6[42], Mediu6);  // ../RTL/cortexm0ds_logic.v(16678)
  not u20461 (Pzbpw6, n5816);  // ../RTL/cortexm0ds_logic.v(16678)
  and u20462 (Mediu6, K0cpw6, Hobpw6);  // ../RTL/cortexm0ds_logic.v(16679)
  and u20463 (Bzbpw6, R0cpw6, Y0cpw6);  // ../RTL/cortexm0ds_logic.v(16680)
  and u20464 (n5817, R4gpw6[44], Nbdiu6);  // ../RTL/cortexm0ds_logic.v(16681)
  not u20465 (Y0cpw6, n5817);  // ../RTL/cortexm0ds_logic.v(16681)
  or u20466 (O8yiu6, Eqbpw6, D0cpw6);  // ../RTL/cortexm0ds_logic.v(16682)
  not u20467 (Nbdiu6, O8yiu6);  // ../RTL/cortexm0ds_logic.v(16682)
  not u20468 (D0cpw6, K0cpw6);  // ../RTL/cortexm0ds_logic.v(16683)
  or u20469 (R0cpw6, Bcsow6, Eayiu6);  // ../RTL/cortexm0ds_logic.v(16684)
  and u2047 (Ax2iu6, U03iu6, B13iu6);  // ../RTL/cortexm0ds_logic.v(3851)
  not u20470 (Eayiu6, O8diu6);  // ../RTL/cortexm0ds_logic.v(16685)
  and u20471 (O8diu6, Sjbpw6, K0cpw6);  // ../RTL/cortexm0ds_logic.v(16686)
  and u20472 (K0cpw6, Zqbpw6, Uybpw6);  // ../RTL/cortexm0ds_logic.v(16687)
  or u20473 (n5818, Tfciu6, vis_ipsr_o[3]);  // ../RTL/cortexm0ds_logic.v(16688)
  not u20474 (Zqbpw6, n5818);  // ../RTL/cortexm0ds_logic.v(16688)
  not u20475 (Bcsow6, R4gpw6[46]);  // ../RTL/cortexm0ds_logic.v(16689)
  and u20476 (Tubpw6, F1cpw6, M1cpw6);  // ../RTL/cortexm0ds_logic.v(16690)
  and u20477 (M1cpw6, T1cpw6, A2cpw6);  // ../RTL/cortexm0ds_logic.v(16691)
  and u20478 (A2cpw6, H2cpw6, O2cpw6);  // ../RTL/cortexm0ds_logic.v(16692)
  or u20479 (O2cpw6, Yysow6, Oyfiu6);  // ../RTL/cortexm0ds_logic.v(16693)
  or u2048 (B13iu6, L02iu6, Mdhpw6[0]);  // ../RTL/cortexm0ds_logic.v(3852)
  buf u20480 (Eafpw6[22], Nxkbx6[23]);  // ../RTL/cortexm0ds_logic.v(3167)
  or u20481 (Oyfiu6, V2cpw6, Tnbpw6);  // ../RTL/cortexm0ds_logic.v(16695)
  not u20482 (Jzfiu6, Oyfiu6);  // ../RTL/cortexm0ds_logic.v(16695)
  buf u20483 (Eafpw6[21], Nxkbx6[22]);  // ../RTL/cortexm0ds_logic.v(3167)
  not u20484 (Yysow6, R4gpw6[48]);  // ../RTL/cortexm0ds_logic.v(16697)
  and u20485 (n5819, R4gpw6[50], Mxfiu6);  // ../RTL/cortexm0ds_logic.v(16698)
  not u20486 (H2cpw6, n5819);  // ../RTL/cortexm0ds_logic.v(16698)
  not u20487 (Mxfiu6, Rwfiu6);  // ../RTL/cortexm0ds_logic.v(16699)
  or u20488 (Rwfiu6, V2cpw6, Ilbpw6);  // ../RTL/cortexm0ds_logic.v(16700)
  and u20489 (T1cpw6, C3cpw6, J3cpw6);  // ../RTL/cortexm0ds_logic.v(16701)
  AL_MUX u2049 (
    .i0(I13iu6),
    .i1(P13iu6),
    .sel(W13iu6),
    .o(Hvxhu6));  // ../RTL/cortexm0ds_logic.v(3853)
  or u20490 (J3cpw6, Uwsow6, Ubyiu6);  // ../RTL/cortexm0ds_logic.v(16702)
  or u20491 (Ubyiu6, Eqbpw6, V2cpw6);  // ../RTL/cortexm0ds_logic.v(16703)
  buf u20492 (Eafpw6[20], Nxkbx6[21]);  // ../RTL/cortexm0ds_logic.v(3167)
  not u20493 (Uwsow6, R4gpw6[52]);  // ../RTL/cortexm0ds_logic.v(16705)
  and u20494 (n5820, R4gpw6[54], Etfiu6);  // ../RTL/cortexm0ds_logic.v(16706)
  not u20495 (C3cpw6, n5820);  // ../RTL/cortexm0ds_logic.v(16706)
  not u20496 (Etfiu6, Kdyiu6);  // ../RTL/cortexm0ds_logic.v(16707)
  or u20497 (Kdyiu6, Dtbpw6, V2cpw6);  // ../RTL/cortexm0ds_logic.v(16708)
  and u20498 (n5821, Jibpw6, Uybpw6);  // ../RTL/cortexm0ds_logic.v(16709)
  not u20499 (V2cpw6, n5821);  // ../RTL/cortexm0ds_logic.v(16709)
  buf u205 (vis_r8_o[19], Oyrax6);  // ../RTL/cortexm0ds_logic.v(2579)
  and u2050 (I13iu6, D23iu6, K23iu6);  // ../RTL/cortexm0ds_logic.v(3854)
  or u20500 (n5822, Ngfiu6, vis_ipsr_o[2]);  // ../RTL/cortexm0ds_logic.v(16710)
  not u20501 (Jibpw6, n5822);  // ../RTL/cortexm0ds_logic.v(16710)
  not u20502 (Dtbpw6, Sjbpw6);  // ../RTL/cortexm0ds_logic.v(16711)
  and u20503 (F1cpw6, Q3cpw6, X3cpw6);  // ../RTL/cortexm0ds_logic.v(16712)
  and u20504 (X3cpw6, E4cpw6, L4cpw6);  // ../RTL/cortexm0ds_logic.v(16713)
  and u20505 (n5823, R4gpw6[56], Arfiu6);  // ../RTL/cortexm0ds_logic.v(16714)
  not u20506 (L4cpw6, n5823);  // ../RTL/cortexm0ds_logic.v(16714)
  buf u20507 (Eafpw6[19], Nxkbx6[20]);  // ../RTL/cortexm0ds_logic.v(3167)
  and u20508 (Arfiu6, S4cpw6, Ljbpw6);  // ../RTL/cortexm0ds_logic.v(16716)
  not u20509 (Afyiu6, Arfiu6);  // ../RTL/cortexm0ds_logic.v(16716)
  and u2051 (K23iu6, R23iu6, Y23iu6);  // ../RTL/cortexm0ds_logic.v(3855)
  and u20510 (S4cpw6, Uybpw6, Ukbpw6);  // ../RTL/cortexm0ds_logic.v(16717)
  and u20511 (n5824, R4gpw6[58], Ahbiu6);  // ../RTL/cortexm0ds_logic.v(16718)
  not u20512 (E4cpw6, n5824);  // ../RTL/cortexm0ds_logic.v(16718)
  buf u20513 (Eafpw6[18], Nxkbx6[19]);  // ../RTL/cortexm0ds_logic.v(3167)
  and u20514 (Ahbiu6, Z4cpw6, Ljbpw6);  // ../RTL/cortexm0ds_logic.v(16720)
  not u20515 (Qgyiu6, Ahbiu6);  // ../RTL/cortexm0ds_logic.v(16720)
  and u20516 (Z4cpw6, Uybpw6, Hobpw6);  // ../RTL/cortexm0ds_logic.v(16721)
  buf u20517 (Eafpw6[17], Nxkbx6[18]);  // ../RTL/cortexm0ds_logic.v(3167)
  and u20518 (Hobpw6, vis_ipsr_o[0], Siciu6);  // ../RTL/cortexm0ds_logic.v(16723)
  not u20519 (Ilbpw6, Hobpw6);  // ../RTL/cortexm0ds_logic.v(16723)
  or u2052 (n260, Iahpw6[29], Iahpw6[30]);  // ../RTL/cortexm0ds_logic.v(3856)
  and u20520 (Q3cpw6, G5cpw6, N5cpw6);  // ../RTL/cortexm0ds_logic.v(16724)
  and u20521 (n5825, R4gpw6[60], Lyhiu6);  // ../RTL/cortexm0ds_logic.v(16725)
  not u20522 (N5cpw6, n5825);  // ../RTL/cortexm0ds_logic.v(16725)
  and u20523 (Lyhiu6, U5cpw6, A9row6);  // ../RTL/cortexm0ds_logic.v(16726)
  and u20524 (n5826, R4gpw6[62], Webiu6);  // ../RTL/cortexm0ds_logic.v(16727)
  not u20525 (G5cpw6, n5826);  // ../RTL/cortexm0ds_logic.v(16727)
  and u20526 (Webiu6, U5cpw6, Sjbpw6);  // ../RTL/cortexm0ds_logic.v(16728)
  and u20527 (U5cpw6, Ljbpw6, Uybpw6);  // ../RTL/cortexm0ds_logic.v(16729)
  or u20528 (n5827, Vhbiu6, vis_ipsr_o[4]);  // ../RTL/cortexm0ds_logic.v(16730)
  not u20529 (Uybpw6, n5827);  // ../RTL/cortexm0ds_logic.v(16730)
  not u2053 (Y23iu6, n260);  // ../RTL/cortexm0ds_logic.v(3856)
  not u20530 (Vhbiu6, vis_ipsr_o[5]);  // ../RTL/cortexm0ds_logic.v(16731)
  or u20531 (n5828, Ngfiu6, Tfciu6);  // ../RTL/cortexm0ds_logic.v(16732)
  not u20532 (Ljbpw6, n5828);  // ../RTL/cortexm0ds_logic.v(16732)
  not u20533 (Tfciu6, vis_ipsr_o[2]);  // ../RTL/cortexm0ds_logic.v(16733)
  not u20534 (Ngfiu6, vis_ipsr_o[3]);  // ../RTL/cortexm0ds_logic.v(16734)
  or u20535 (n5829, B6cpw6, vis_primask_o);  // ../RTL/cortexm0ds_logic.v(16735)
  not u20536 (Pmapw6, n5829);  // ../RTL/cortexm0ds_logic.v(16735)
  and u20537 (B6cpw6, I6cpw6, H9row6);  // ../RTL/cortexm0ds_logic.v(16736)
  and u20538 (I6cpw6, M8row6, P6cpw6);  // ../RTL/cortexm0ds_logic.v(16737)
  or u20539 (P6cpw6, A9row6, Sjbpw6);  // ../RTL/cortexm0ds_logic.v(16738)
  or u2054 (n261, Iahpw6[27], Iahpw6[28]);  // ../RTL/cortexm0ds_logic.v(3857)
  and u20540 (Sjbpw6, vis_ipsr_o[1], vis_ipsr_o[0]);  // ../RTL/cortexm0ds_logic.v(16739)
  or u20541 (Eqbpw6, Siciu6, vis_ipsr_o[0]);  // ../RTL/cortexm0ds_logic.v(16740)
  not u20542 (A9row6, Eqbpw6);  // ../RTL/cortexm0ds_logic.v(16740)
  not u20543 (Siciu6, vis_ipsr_o[1]);  // ../RTL/cortexm0ds_logic.v(16741)
  and u20544 (n5830, W6cpw6, D7cpw6);  // ../RTL/cortexm0ds_logic.v(16742)
  not u20545 (Ulapw6, n5830);  // ../RTL/cortexm0ds_logic.v(16742)
  and u20546 (D7cpw6, K7cpw6, Kxziu6);  // ../RTL/cortexm0ds_logic.v(16743)
  or u20547 (n5831, R75iu6, Hbbow6);  // ../RTL/cortexm0ds_logic.v(16744)
  not u20548 (K7cpw6, n5831);  // ../RTL/cortexm0ds_logic.v(16744)
  not u20549 (R75iu6, Omyiu6);  // ../RTL/cortexm0ds_logic.v(16745)
  not u2055 (R23iu6, n261);  // ../RTL/cortexm0ds_logic.v(3857)
  and u20550 (W6cpw6, L78ju6, Frziu6);  // ../RTL/cortexm0ds_logic.v(16746)
  and u20551 (Glapw6, Erhiu6, R7cpw6);  // ../RTL/cortexm0ds_logic.v(16747)
  and u20552 (n5832, Jxaiu6, Y7cpw6);  // ../RTL/cortexm0ds_logic.v(16748)
  not u20553 (R7cpw6, n5832);  // ../RTL/cortexm0ds_logic.v(16748)
  and u20554 (n5833, F8cpw6, M8cpw6);  // ../RTL/cortexm0ds_logic.v(16749)
  not u20555 (Y7cpw6, n5833);  // ../RTL/cortexm0ds_logic.v(16749)
  and u20556 (n5834, T8cpw6, A9cpw6);  // ../RTL/cortexm0ds_logic.v(16750)
  not u20557 (M8cpw6, n5834);  // ../RTL/cortexm0ds_logic.v(16750)
  or u20558 (A9cpw6, Ftjiu6, D7fpw6[14]);  // ../RTL/cortexm0ds_logic.v(16751)
  or u20559 (n5835, Xjbow6, D7fpw6[12]);  // ../RTL/cortexm0ds_logic.v(16752)
  and u2056 (D23iu6, F33iu6, M33iu6);  // ../RTL/cortexm0ds_logic.v(3858)
  not u20560 (T8cpw6, n5835);  // ../RTL/cortexm0ds_logic.v(16752)
  and u20561 (Xjbow6, D7fpw6[14], S1ehu6);  // ../RTL/cortexm0ds_logic.v(16753)
  or u20562 (n5836, Y40ju6, Jiiiu6);  // ../RTL/cortexm0ds_logic.v(16754)
  not u20563 (F8cpw6, n5836);  // ../RTL/cortexm0ds_logic.v(16754)
  and u20564 (Jxaiu6, H9cpw6, O9cpw6);  // ../RTL/cortexm0ds_logic.v(16755)
  or u20565 (n5837, Y2oiu6, Jcaiu6);  // ../RTL/cortexm0ds_logic.v(16756)
  not u20566 (O9cpw6, n5837);  // ../RTL/cortexm0ds_logic.v(16756)
  or u20567 (n5838, Wfoiu6, Ccoiu6);  // ../RTL/cortexm0ds_logic.v(16757)
  not u20568 (H9cpw6, n5838);  // ../RTL/cortexm0ds_logic.v(16757)
  and u20569 (n5839, Pu1ju6, B8apw6);  // ../RTL/cortexm0ds_logic.v(16758)
  or u2057 (n262, Iahpw6[25], Iahpw6[26]);  // ../RTL/cortexm0ds_logic.v(3859)
  not u20570 (I1aiu6, n5839);  // ../RTL/cortexm0ds_logic.v(16758)
  and u20571 (Ueapw6, Erhiu6, Lrhiu6);  // ../RTL/cortexm0ds_logic.v(16759)
  and u20572 (Lrhiu6, V9cpw6, Cacpw6);  // ../RTL/cortexm0ds_logic.v(16760)
  and u20573 (Cacpw6, Jacpw6, Qacpw6);  // ../RTL/cortexm0ds_logic.v(16761)
  and u20574 (Qacpw6, Xacpw6, Uloiu6);  // ../RTL/cortexm0ds_logic.v(16762)
  and u20575 (n5840, Ebcpw6, N2ghu6);  // ../RTL/cortexm0ds_logic.v(16763)
  not u20576 (Uloiu6, n5840);  // ../RTL/cortexm0ds_logic.v(16763)
  and u20577 (Ebcpw6, Whfiu6, D6kiu6);  // ../RTL/cortexm0ds_logic.v(16764)
  and u20578 (Whfiu6, Cyfpw6[3], Cyfpw6[5]);  // ../RTL/cortexm0ds_logic.v(16765)
  and u20579 (Xacpw6, Kz6ow6, Td0iu6);  // ../RTL/cortexm0ds_logic.v(16766)
  not u2058 (M33iu6, n262);  // ../RTL/cortexm0ds_logic.v(3859)
  and u20580 (n5841, Omyiu6, Pfiow6);  // ../RTL/cortexm0ds_logic.v(16767)
  not u20581 (Td0iu6, n5841);  // ../RTL/cortexm0ds_logic.v(16767)
  and u20582 (Pfiow6, Lbcpw6, Oiaiu6);  // ../RTL/cortexm0ds_logic.v(16768)
  and u20583 (Lbcpw6, Sq3ju6, Cyfpw6[5]);  // ../RTL/cortexm0ds_logic.v(16769)
  and u20584 (n5842, Sbcpw6, Pthiu6);  // ../RTL/cortexm0ds_logic.v(16770)
  not u20585 (Kz6ow6, n5842);  // ../RTL/cortexm0ds_logic.v(16770)
  and u20586 (n7[1], H1zhu6, O1zhu6);  // ../RTL/cortexm0ds_logic.v(3185)
  not u20587 (Sbcpw6, Bwziu6);  // ../RTL/cortexm0ds_logic.v(16771)
  buf u20588 (Eafpw6[16], Nxkbx6[17]);  // ../RTL/cortexm0ds_logic.v(3167)
  or u20589 (Jojiu6, Mr0iu6, K9aiu6);  // ../RTL/cortexm0ds_logic.v(16773)
  or u2059 (n263, Iahpw6[23], Iahpw6[24]);  // ../RTL/cortexm0ds_logic.v(3860)
  not u20590 (Pu1ju6, Jojiu6);  // ../RTL/cortexm0ds_logic.v(16773)
  or u20591 (n5843, Zbcpw6, Iepiu6);  // ../RTL/cortexm0ds_logic.v(16774)
  not u20592 (Jacpw6, n5843);  // ../RTL/cortexm0ds_logic.v(16774)
  and u20593 (Iepiu6, W8aiu6, Ldoiu6);  // ../RTL/cortexm0ds_logic.v(16775)
  and u20594 (Zbcpw6, Wp0iu6, D6kiu6);  // ../RTL/cortexm0ds_logic.v(16776)
  and u20595 (V9cpw6, Gccpw6, Nccpw6);  // ../RTL/cortexm0ds_logic.v(16777)
  and u20596 (Nccpw6, Zkapw6, Uccpw6);  // ../RTL/cortexm0ds_logic.v(16778)
  and u20597 (n5844, Ae0iu6, Bdcpw6);  // ../RTL/cortexm0ds_logic.v(16779)
  not u20598 (Uccpw6, n5844);  // ../RTL/cortexm0ds_logic.v(16779)
  and u20599 (n5845, Idcpw6, Pdcpw6);  // ../RTL/cortexm0ds_logic.v(16780)
  buf u206 (Vbgpw6[13], Fb0bx6);  // ../RTL/cortexm0ds_logic.v(3092)
  not u2060 (F33iu6, n263);  // ../RTL/cortexm0ds_logic.v(3860)
  not u20600 (Bdcpw6, n5845);  // ../RTL/cortexm0ds_logic.v(16780)
  and u20601 (Pdcpw6, Wdcpw6, Decpw6);  // ../RTL/cortexm0ds_logic.v(16781)
  and u20602 (n5846, N3ziu6, Kecpw6);  // ../RTL/cortexm0ds_logic.v(16782)
  not u20603 (Decpw6, n5846);  // ../RTL/cortexm0ds_logic.v(16782)
  or u20604 (Kecpw6, Y2oiu6, X97ow6);  // ../RTL/cortexm0ds_logic.v(16783)
  and u20605 (N3ziu6, Yljiu6, Nlaiu6);  // ../RTL/cortexm0ds_logic.v(16784)
  and u20606 (Wdcpw6, Recpw6, Iw8ow6);  // ../RTL/cortexm0ds_logic.v(16785)
  and u20607 (n5847, Yecpw6, Wwziu6);  // ../RTL/cortexm0ds_logic.v(16786)
  not u20608 (Iw8ow6, n5847);  // ../RTL/cortexm0ds_logic.v(16786)
  buf u20609 (Eafpw6[15], Nxkbx6[16]);  // ../RTL/cortexm0ds_logic.v(3167)
  AL_MUX u2061 (
    .i0(T33iu6),
    .i1(Pifax6),
    .sel(W13iu6),
    .o(Avxhu6));  // ../RTL/cortexm0ds_logic.v(3861)
  and u20610 (Wwziu6, D6kiu6, H4ghu6);  // ../RTL/cortexm0ds_logic.v(16788)
  not u20611 (Nloiu6, Wwziu6);  // ../RTL/cortexm0ds_logic.v(16788)
  or u20612 (n5848, Y2oiu6, Xe8iu6);  // ../RTL/cortexm0ds_logic.v(16789)
  not u20613 (Yecpw6, n5848);  // ../RTL/cortexm0ds_logic.v(16789)
  and u20614 (n5849, Ffcpw6, Pt2ju6);  // ../RTL/cortexm0ds_logic.v(16790)
  not u20615 (Recpw6, n5849);  // ../RTL/cortexm0ds_logic.v(16790)
  or u20616 (n5850, C0ehu6, Cyfpw6[6]);  // ../RTL/cortexm0ds_logic.v(16791)
  not u20617 (Ffcpw6, n5850);  // ../RTL/cortexm0ds_logic.v(16791)
  and u20618 (Idcpw6, Mfcpw6, Tfcpw6);  // ../RTL/cortexm0ds_logic.v(16792)
  or u20619 (Tfcpw6, Qjaiu6, Kw0ju6);  // ../RTL/cortexm0ds_logic.v(16793)
  AL_MUX u2062 (
    .i0(n6026),
    .i1(1'b0),
    .sel(Romhu6),
    .o(n6023));  // ../RTL/cortexm0ds_logic.v(3132)
  and u20620 (Mfcpw6, Agcpw6, Hgcpw6);  // ../RTL/cortexm0ds_logic.v(16794)
  and u20621 (n5851, S6aiu6, Ogcpw6);  // ../RTL/cortexm0ds_logic.v(16795)
  not u20622 (Hgcpw6, n5851);  // ../RTL/cortexm0ds_logic.v(16795)
  and u20623 (n5852, Owaiu6, Vgcpw6);  // ../RTL/cortexm0ds_logic.v(16796)
  not u20624 (Ogcpw6, n5852);  // ../RTL/cortexm0ds_logic.v(16796)
  or u20625 (Vgcpw6, Xmliu6, Cyfpw6[0]);  // ../RTL/cortexm0ds_logic.v(16797)
  not u20626 (Owaiu6, Cp3ju6);  // ../RTL/cortexm0ds_logic.v(16798)
  and u20627 (n5853, Chcpw6, K9aiu6);  // ../RTL/cortexm0ds_logic.v(16799)
  not u20628 (Agcpw6, n5853);  // ../RTL/cortexm0ds_logic.v(16799)
  and u20629 (n5854, Jhcpw6, Qhcpw6);  // ../RTL/cortexm0ds_logic.v(16800)
  AL_MUX u2063 (
    .i0(Cjhpw6[3]),
    .i1(H43iu6),
    .sel(Em1iu6),
    .o(Tuxhu6));  // ../RTL/cortexm0ds_logic.v(3863)
  not u20630 (Chcpw6, n5854);  // ../RTL/cortexm0ds_logic.v(16800)
  buf u20631 (Tnhpw6[3], P23qw6);  // ../RTL/cortexm0ds_logic.v(2163)
  not u20632 (Qhcpw6, Qkaow6);  // ../RTL/cortexm0ds_logic.v(16801)
  or u20633 (n5855, Gm9pw6, Cyfpw6[4]);  // ../RTL/cortexm0ds_logic.v(16802)
  not u20634 (L45iu6, n5855);  // ../RTL/cortexm0ds_logic.v(16802)
  or u20635 (Gm9pw6, Cyfpw6[3], C0ehu6);  // ../RTL/cortexm0ds_logic.v(16803)
  buf u20636 (Tnhpw6[2], Xn7ax6);  // ../RTL/cortexm0ds_logic.v(2163)
  and u20637 (n5856, Xhcpw6, Eicpw6);  // ../RTL/cortexm0ds_logic.v(16805)
  not u20638 (Zkapw6, n5856);  // ../RTL/cortexm0ds_logic.v(16805)
  or u20639 (n5857, Knaiu6, Cyfpw6[5]);  // ../RTL/cortexm0ds_logic.v(16806)
  and u2064 (n264, Omdpw6, O43iu6);  // ../RTL/cortexm0ds_logic.v(3864)
  not u20640 (Eicpw6, n5857);  // ../RTL/cortexm0ds_logic.v(16806)
  or u20641 (n5858, As0iu6, Qxaiu6);  // ../RTL/cortexm0ds_logic.v(16807)
  not u20642 (Xhcpw6, n5858);  // ../RTL/cortexm0ds_logic.v(16807)
  and u20643 (Gccpw6, Licpw6, Sicpw6);  // ../RTL/cortexm0ds_logic.v(16808)
  and u20644 (n5859, Zicpw6, Mmjiu6);  // ../RTL/cortexm0ds_logic.v(16809)
  not u20645 (Sicpw6, n5859);  // ../RTL/cortexm0ds_logic.v(16809)
  not u20646 (Mmjiu6, Qu7ow6);  // ../RTL/cortexm0ds_logic.v(16810)
  or u20647 (Qu7ow6, Nsaiu6, Pxyiu6);  // ../RTL/cortexm0ds_logic.v(16811)
  and u20648 (n5860, Gjcpw6, vis_pc_o[2]);  // ../RTL/cortexm0ds_logic.v(16812)
  not u20649 (Pxyiu6, n5860);  // ../RTL/cortexm0ds_logic.v(16812)
  not u2065 (H43iu6, n264);  // ../RTL/cortexm0ds_logic.v(3864)
  and u20650 (Gjcpw6, Qqdhu6, El1ju6);  // ../RTL/cortexm0ds_logic.v(16813)
  and u20651 (L62ju6, Njcpw6, Q5aiu6);  // ../RTL/cortexm0ds_logic.v(16814)
  not u20652 (Nsaiu6, L62ju6);  // ../RTL/cortexm0ds_logic.v(16814)
  or u20653 (Njcpw6, El1ju6, E6phu6);  // ../RTL/cortexm0ds_logic.v(16815)
  not u20654 (El1ju6, Stdhu6);  // ../RTL/cortexm0ds_logic.v(16816)
  buf u20655 (Tnhpw6[1], Vj3qw6);  // ../RTL/cortexm0ds_logic.v(2163)
  not u20656 (Zicpw6, Tfcpw6);  // ../RTL/cortexm0ds_logic.v(16817)
  and u20657 (n5861, I30ju6, Ii0iu6);  // ../RTL/cortexm0ds_logic.v(16818)
  not u20658 (Kw0ju6, n5861);  // ../RTL/cortexm0ds_logic.v(16818)
  or u20659 (n5862, R2aiu6, Dxziu6);  // ../RTL/cortexm0ds_logic.v(16819)
  AL_MUX u2066 (
    .i0(Lznhu6),
    .i1(Dtnhu6),
    .sel(n265),
    .o(Muxhu6));  // ../RTL/cortexm0ds_logic.v(3865)
  not u20660 (I30ju6, n5862);  // ../RTL/cortexm0ds_logic.v(16819)
  buf u20661 (Eafpw6[14], Nxkbx6[15]);  // ../RTL/cortexm0ds_logic.v(3167)
  and u20662 (Dxziu6, Ujcpw6, Bkcpw6);  // ../RTL/cortexm0ds_logic.v(16821)
  not u20663 (Xojiu6, Dxziu6);  // ../RTL/cortexm0ds_logic.v(16821)
  and u20664 (Bkcpw6, Ikcpw6, Pkcpw6);  // ../RTL/cortexm0ds_logic.v(16822)
  or u20665 (n5863, Xkhow6, Qbiiu6);  // ../RTL/cortexm0ds_logic.v(16823)
  not u20666 (Pkcpw6, n5863);  // ../RTL/cortexm0ds_logic.v(16823)
  and u20667 (Qbiiu6, S8fpw6[9], S8fpw6[8]);  // ../RTL/cortexm0ds_logic.v(16824)
  and u20668 (Xkhow6, S8fpw6[7], L28ow6);  // ../RTL/cortexm0ds_logic.v(16825)
  or u20669 (L28ow6, G55iu6, S8fpw6[6]);  // ../RTL/cortexm0ds_logic.v(16826)
  or u2067 (n265, Npzhu6, Gpzhu6);  // ../RTL/cortexm0ds_logic.v(3866)
  and u20670 (Ikcpw6, Wj7ow6, G7iow6);  // ../RTL/cortexm0ds_logic.v(16827)
  and u20671 (n5864, S8fpw6[6], G55iu6);  // ../RTL/cortexm0ds_logic.v(16828)
  not u20672 (G7iow6, n5864);  // ../RTL/cortexm0ds_logic.v(16828)
  or u20673 (G55iu6, Wkcpw6, S8fpw6[5]);  // ../RTL/cortexm0ds_logic.v(16829)
  and u20674 (n5865, S8fpw6[5], Wkcpw6);  // ../RTL/cortexm0ds_logic.v(16830)
  not u20675 (Wj7ow6, n5865);  // ../RTL/cortexm0ds_logic.v(16830)
  not u20676 (Wkcpw6, Zoyiu6);  // ../RTL/cortexm0ds_logic.v(16831)
  and u20677 (Zoyiu6, N55iu6, Qjoiu6);  // ../RTL/cortexm0ds_logic.v(16832)
  and u20678 (Ujcpw6, Dlcpw6, Klcpw6);  // ../RTL/cortexm0ds_logic.v(16833)
  and u20679 (n5866, S8fpw6[10], Weiiu6);  // ../RTL/cortexm0ds_logic.v(16834)
  buf u2068 (Eafpw6[5], Nxkbx6[6]);  // ../RTL/cortexm0ds_logic.v(3167)
  not u20680 (Klcpw6, n5866);  // ../RTL/cortexm0ds_logic.v(16834)
  and u20681 (Dlcpw6, Voiiu6, Btbow6);  // ../RTL/cortexm0ds_logic.v(16835)
  or u20682 (Btbow6, Qjoiu6, N55iu6);  // ../RTL/cortexm0ds_logic.v(16836)
  or u20683 (n5867, B65iu6, S8fpw6[11]);  // ../RTL/cortexm0ds_logic.v(16837)
  not u20684 (N55iu6, n5867);  // ../RTL/cortexm0ds_logic.v(16837)
  not u20685 (Qjoiu6, S8fpw6[4]);  // ../RTL/cortexm0ds_logic.v(16838)
  and u20686 (n5868, S8fpw6[11], B65iu6);  // ../RTL/cortexm0ds_logic.v(16839)
  not u20687 (Voiiu6, n5868);  // ../RTL/cortexm0ds_logic.v(16839)
  or u20688 (B65iu6, Weiiu6, S8fpw6[10]);  // ../RTL/cortexm0ds_logic.v(16840)
  or u20689 (Weiiu6, S8fpw6[8], S8fpw6[9]);  // ../RTL/cortexm0ds_logic.v(16841)
  xor u2069 (n266, C53iu6, G2ohu6);  // ../RTL/cortexm0ds_logic.v(3867)
  AL_MUX u20690 (
    .i0(Rlcpw6),
    .i1(Ylcpw6),
    .sel(Cyfpw6[4]),
    .o(Licpw6));  // ../RTL/cortexm0ds_logic.v(16842)
  or u20691 (Ylcpw6, Ccoiu6, Geaiu6);  // ../RTL/cortexm0ds_logic.v(16843)
  and u20692 (Rlcpw6, Fmcpw6, Mmcpw6);  // ../RTL/cortexm0ds_logic.v(16844)
  and u20693 (n5869, Z6aiu6, Oiaiu6);  // ../RTL/cortexm0ds_logic.v(16845)
  not u20694 (Mmcpw6, n5869);  // ../RTL/cortexm0ds_logic.v(16845)
  and u20695 (Fmcpw6, Tmcpw6, Ancpw6);  // ../RTL/cortexm0ds_logic.v(16846)
  and u20696 (n5870, Hncpw6, K2aiu6);  // ../RTL/cortexm0ds_logic.v(16847)
  not u20697 (Ancpw6, n5870);  // ../RTL/cortexm0ds_logic.v(16847)
  and u20698 (Hncpw6, N2ghu6, D6kiu6);  // ../RTL/cortexm0ds_logic.v(16848)
  or u20699 (Tmcpw6, Jc2ju6, R2aiu6);  // ../RTL/cortexm0ds_logic.v(16849)
  buf u207 (Gqgpw6[25], Tkdax6);  // ../RTL/cortexm0ds_logic.v(2377)
  not u2070 (Fuxhu6, n266);  // ../RTL/cortexm0ds_logic.v(3867)
  not u20700 (R2aiu6, W8aiu6);  // ../RTL/cortexm0ds_logic.v(16850)
  not u20701 (Jc2ju6, Es1ju6);  // ../RTL/cortexm0ds_logic.v(16851)
  and u20702 (Es1ju6, Nlaiu6, Xe8iu6);  // ../RTL/cortexm0ds_logic.v(16852)
  or u20703 (n5871, CDBGPWRUPACK, Oncpw6);  // ../RTL/cortexm0ds_logic.v(16853)
  not u20704 (GATEHCLK, n5871);  // ../RTL/cortexm0ds_logic.v(16853)
  or u20705 (n5872, E6phu6, SLEEPING);  // ../RTL/cortexm0ds_logic.v(16854)
  not u20706 (Oncpw6, n5872);  // ../RTL/cortexm0ds_logic.v(16854)
  and u20707 (SLEEPING, Qnghu6, Vncpw6);  // ../RTL/cortexm0ds_logic.v(16855)
  and u20708 (n5873, Cocpw6, Jocpw6);  // ../RTL/cortexm0ds_logic.v(16856)
  not u20709 (CODENSEQ, n5873);  // ../RTL/cortexm0ds_logic.v(16856)
  AL_MUX u2071 (
    .i0(Punhu6),
    .i1(Xkqpw6),
    .sel(n267),
    .o(Ytxhu6));  // ../RTL/cortexm0ds_logic.v(3868)
  and u20710 (Jocpw6, Qocpw6, Uriiu6);  // ../RTL/cortexm0ds_logic.v(16857)
  or u20711 (n5874, Hrfpw6[16], Yyfhu6);  // ../RTL/cortexm0ds_logic.v(16858)
  not u20712 (Qocpw6, n5874);  // ../RTL/cortexm0ds_logic.v(16858)
  and u20713 (Cocpw6, Xocpw6, Epcpw6);  // ../RTL/cortexm0ds_logic.v(16859)
  and u20714 (n5875, Ppfpw6[16], Ntfhu6);  // ../RTL/cortexm0ds_logic.v(16860)
  not u20715 (Epcpw6, n5875);  // ../RTL/cortexm0ds_logic.v(16860)
  and u20716 (Xocpw6, Lpcpw6, Ygapw6);  // ../RTL/cortexm0ds_logic.v(16861)
  and u20717 (n5876, Spcpw6, Gc5iu6);  // ../RTL/cortexm0ds_logic.v(16862)
  not u20718 (Ygapw6, n5876);  // ../RTL/cortexm0ds_logic.v(16862)
  buf u20719 (Eafpw6[13], Nxkbx6[14]);  // ../RTL/cortexm0ds_logic.v(3167)
  or u2072 (n267, Rrnhu6, G2ohu6);  // ../RTL/cortexm0ds_logic.v(3869)
  and u20720 (Gc5iu6, L6aiu6, Zpcpw6);  // ../RTL/cortexm0ds_logic.v(16864)
  not u20721 (Wofiu6, Gc5iu6);  // ../RTL/cortexm0ds_logic.v(16864)
  and u20722 (n5877, B8apw6, D6kiu6);  // ../RTL/cortexm0ds_logic.v(16865)
  not u20723 (Zpcpw6, n5877);  // ../RTL/cortexm0ds_logic.v(16865)
  or u20724 (n5878, Ccoiu6, Ii0iu6);  // ../RTL/cortexm0ds_logic.v(16866)
  not u20725 (B8apw6, n5878);  // ../RTL/cortexm0ds_logic.v(16866)
  not u20726 (Ccoiu6, H3aju6);  // ../RTL/cortexm0ds_logic.v(16867)
  and u20727 (H3aju6, Cyfpw6[7], Xe8iu6);  // ../RTL/cortexm0ds_logic.v(16868)
  and u20728 (n5879, Wp0iu6, Mfjiu6);  // ../RTL/cortexm0ds_logic.v(16869)
  not u20729 (L6aiu6, n5879);  // ../RTL/cortexm0ds_logic.v(16869)
  buf u2073 (Eafpw6[4], Nxkbx6[5]);  // ../RTL/cortexm0ds_logic.v(3167)
  and u20730 (Mfjiu6, Cyfpw6[4], Y7ghu6);  // ../RTL/cortexm0ds_logic.v(16870)
  and u20731 (n101[1], Lozhu6, Sozhu6);  // ../RTL/cortexm0ds_logic.v(3356)
  or u20732 (Et8iu6, U0aiu6, Gqcpw6);  // ../RTL/cortexm0ds_logic.v(16872)
  and u20733 (Gqcpw6, D1piu6, Tr0iu6);  // ../RTL/cortexm0ds_logic.v(16873)
  and u20734 (U0aiu6, Hzziu6, Cyfpw6[0]);  // ../RTL/cortexm0ds_logic.v(16874)
  and u20735 (n5880, Nqcpw6, Uqcpw6);  // ../RTL/cortexm0ds_logic.v(16875)
  not u20736 (B7qow6, n5880);  // ../RTL/cortexm0ds_logic.v(16875)
  and u20737 (Uqcpw6, Brcpw6, Ircpw6);  // ../RTL/cortexm0ds_logic.v(16876)
  or u20738 (n5881, Prcpw6, Nz2ju6);  // ../RTL/cortexm0ds_logic.v(16877)
  not u20739 (Ircpw6, n5881);  // ../RTL/cortexm0ds_logic.v(16877)
  and u2074 (n268, X53iu6, E63iu6);  // ../RTL/cortexm0ds_logic.v(3871)
  and u20740 (Nz2ju6, F23ju6, D31ju6);  // ../RTL/cortexm0ds_logic.v(16878)
  and u20741 (D31ju6, Cyfpw6[5], Tfjiu6);  // ../RTL/cortexm0ds_logic.v(16879)
  and u20742 (F23ju6, Cyfpw6[0], Hs0iu6);  // ../RTL/cortexm0ds_logic.v(16880)
  and u20743 (Prcpw6, Wrcpw6, Obbow6);  // ../RTL/cortexm0ds_logic.v(16881)
  or u20744 (n5882, Jcaiu6, Mr0iu6);  // ../RTL/cortexm0ds_logic.v(16882)
  not u20745 (Obbow6, n5882);  // ../RTL/cortexm0ds_logic.v(16882)
  and u20746 (Wrcpw6, Dscpw6, Lkaiu6);  // ../RTL/cortexm0ds_logic.v(16883)
  not u20747 (Lkaiu6, Gwyiu6);  // ../RTL/cortexm0ds_logic.v(16884)
  and u20748 (Gwyiu6, Cyfpw6[5], Ii0iu6);  // ../RTL/cortexm0ds_logic.v(16885)
  or u20749 (Dscpw6, U4kiu6, Buaow6);  // ../RTL/cortexm0ds_logic.v(16886)
  not u2075 (Rtxhu6, n268);  // ../RTL/cortexm0ds_logic.v(3871)
  and u20750 (Buaow6, Tr0iu6, Xe8iu6);  // ../RTL/cortexm0ds_logic.v(16887)
  and u20751 (Brcpw6, Kscpw6, Rscpw6);  // ../RTL/cortexm0ds_logic.v(16888)
  and u20752 (n5883, Yscpw6, W2aow6);  // ../RTL/cortexm0ds_logic.v(16889)
  not u20753 (Rscpw6, n5883);  // ../RTL/cortexm0ds_logic.v(16889)
  and u20754 (W2aow6, Cyfpw6[5], Hs0iu6);  // ../RTL/cortexm0ds_logic.v(16890)
  or u20755 (n5884, Mr0iu6, Y7ghu6);  // ../RTL/cortexm0ds_logic.v(16891)
  not u20756 (Yscpw6, n5884);  // ../RTL/cortexm0ds_logic.v(16891)
  and u20757 (n5885, Imaiu6, Ftcpw6);  // ../RTL/cortexm0ds_logic.v(16892)
  not u20758 (Kscpw6, n5885);  // ../RTL/cortexm0ds_logic.v(16892)
  and u20759 (n5886, Mtcpw6, Ttcpw6);  // ../RTL/cortexm0ds_logic.v(16893)
  and u2076 (n269, Rgnhu6, L63iu6);  // ../RTL/cortexm0ds_logic.v(3872)
  not u20760 (Ftcpw6, n5886);  // ../RTL/cortexm0ds_logic.v(16893)
  or u20761 (n5887, Wp0iu6, Cyfpw6[7]);  // ../RTL/cortexm0ds_logic.v(16894)
  not u20762 (Ttcpw6, n5887);  // ../RTL/cortexm0ds_logic.v(16894)
  or u20763 (n5888, Cp3ju6, Sq3ju6);  // ../RTL/cortexm0ds_logic.v(16895)
  not u20764 (Mtcpw6, n5888);  // ../RTL/cortexm0ds_logic.v(16895)
  and u20765 (Sq3ju6, Cyfpw6[6], Nlaiu6);  // ../RTL/cortexm0ds_logic.v(16896)
  and u20766 (Cp3ju6, Cyfpw6[1], Y2oiu6);  // ../RTL/cortexm0ds_logic.v(16897)
  and u20767 (Nqcpw6, Aucpw6, Hucpw6);  // ../RTL/cortexm0ds_logic.v(16898)
  and u20768 (Hucpw6, Oucpw6, Vucpw6);  // ../RTL/cortexm0ds_logic.v(16899)
  and u20769 (n5889, Ae0iu6, Cvcpw6);  // ../RTL/cortexm0ds_logic.v(16900)
  not u2077 (E63iu6, n269);  // ../RTL/cortexm0ds_logic.v(3872)
  not u20770 (Vucpw6, n5889);  // ../RTL/cortexm0ds_logic.v(16900)
  and u20771 (n5890, Jvcpw6, Qvcpw6);  // ../RTL/cortexm0ds_logic.v(16901)
  not u20772 (Cvcpw6, n5890);  // ../RTL/cortexm0ds_logic.v(16901)
  and u20773 (n5891, Xvcpw6, Pfoiu6);  // ../RTL/cortexm0ds_logic.v(16902)
  not u20774 (Qvcpw6, n5891);  // ../RTL/cortexm0ds_logic.v(16902)
  and u20775 (Pfoiu6, Xe8iu6, Hs0iu6);  // ../RTL/cortexm0ds_logic.v(16903)
  not u20776 (Hs0iu6, Cyfpw6[7]);  // ../RTL/cortexm0ds_logic.v(16904)
  and u20777 (Xvcpw6, Frziu6, Cyfpw6[0]);  // ../RTL/cortexm0ds_logic.v(16905)
  or u20778 (n5892, Tfjiu6, H4ghu6);  // ../RTL/cortexm0ds_logic.v(16906)
  not u20779 (Frziu6, n5892);  // ../RTL/cortexm0ds_logic.v(16906)
  and u2078 (n270, S63iu6, Fmyhu6);  // ../RTL/cortexm0ds_logic.v(3873)
  and u20780 (n5893, Ewcpw6, Fd0iu6);  // ../RTL/cortexm0ds_logic.v(16907)
  not u20781 (Jvcpw6, n5893);  // ../RTL/cortexm0ds_logic.v(16907)
  and u20782 (Fd0iu6, Cyfpw6[5], Cyfpw6[1]);  // ../RTL/cortexm0ds_logic.v(16908)
  and u20783 (Ewcpw6, F3aiu6, Tfjiu6);  // ../RTL/cortexm0ds_logic.v(16909)
  and u20784 (n5894, V9ghu6, Lwcpw6);  // ../RTL/cortexm0ds_logic.v(16910)
  not u20785 (Oucpw6, n5894);  // ../RTL/cortexm0ds_logic.v(16910)
  and u20786 (n5895, Erhiu6, Swcpw6);  // ../RTL/cortexm0ds_logic.v(16911)
  not u20787 (Lwcpw6, n5895);  // ../RTL/cortexm0ds_logic.v(16911)
  and u20788 (n5896, Zwcpw6, Pt2ju6);  // ../RTL/cortexm0ds_logic.v(16912)
  not u20789 (Swcpw6, n5896);  // ../RTL/cortexm0ds_logic.v(16912)
  not u2079 (L63iu6, n270);  // ../RTL/cortexm0ds_logic.v(3873)
  and u20790 (Pt2ju6, Cyfpw6[1], Xe8iu6);  // ../RTL/cortexm0ds_logic.v(16913)
  or u20791 (n5897, Qxaiu6, Knaiu6);  // ../RTL/cortexm0ds_logic.v(16914)
  not u20792 (Zwcpw6, n5897);  // ../RTL/cortexm0ds_logic.v(16914)
  buf u20793 (Eafpw6[12], Nxkbx6[13]);  // ../RTL/cortexm0ds_logic.v(3167)
  and u20794 (Erhiu6, Tq9ow6, Gxcpw6);  // ../RTL/cortexm0ds_logic.v(16916)
  and u20795 (n5898, Y8aju6, Vj9pw6);  // ../RTL/cortexm0ds_logic.v(16917)
  not u20796 (Gxcpw6, n5898);  // ../RTL/cortexm0ds_logic.v(16917)
  buf u20797 (Ppfpw6[16], L4lax6);  // ../RTL/cortexm0ds_logic.v(2461)
  not u20798 (Y8aju6, G1vow6);  // ../RTL/cortexm0ds_logic.v(16918)
  or u20799 (Tq9ow6, W8oiu6, Knaiu6);  // ../RTL/cortexm0ds_logic.v(16919)
  buf u208 (Ntfhu6, X7ypw6);  // ../RTL/cortexm0ds_logic.v(2073)
  or u2080 (n271, Z63iu6, G73iu6);  // ../RTL/cortexm0ds_logic.v(3874)
  not u20800 (W8oiu6, Vj9pw6);  // ../RTL/cortexm0ds_logic.v(16920)
  and u20801 (Vj9pw6, Sbghu6, K9aiu6);  // ../RTL/cortexm0ds_logic.v(16921)
  and u20802 (Aucpw6, Nxcpw6, Uxcpw6);  // ../RTL/cortexm0ds_logic.v(16922)
  and u20803 (n5899, J4aju6, Qyniu6);  // ../RTL/cortexm0ds_logic.v(16923)
  not u20804 (Uxcpw6, n5899);  // ../RTL/cortexm0ds_logic.v(16923)
  or u20805 (n5900, Cyfpw6[1], Cyfpw6[6]);  // ../RTL/cortexm0ds_logic.v(16924)
  not u20806 (Qyniu6, n5900);  // ../RTL/cortexm0ds_logic.v(16924)
  and u20807 (J4aju6, Bycpw6, Omyiu6);  // ../RTL/cortexm0ds_logic.v(16925)
  and u20808 (Omyiu6, Cyfpw6[3], Jjhiu6);  // ../RTL/cortexm0ds_logic.v(16926)
  or u20809 (n5901, Cyfpw6[5], Y7ghu6);  // ../RTL/cortexm0ds_logic.v(16927)
  not u2081 (S63iu6, n271);  // ../RTL/cortexm0ds_logic.v(3874)
  not u20810 (Bycpw6, n5901);  // ../RTL/cortexm0ds_logic.v(16927)
  and u20811 (n5902, Cyfpw6[4], Iycpw6);  // ../RTL/cortexm0ds_logic.v(16928)
  not u20812 (Nxcpw6, n5902);  // ../RTL/cortexm0ds_logic.v(16928)
  and u20813 (n5903, Pycpw6, Wycpw6);  // ../RTL/cortexm0ds_logic.v(16929)
  not u20814 (Iycpw6, n5903);  // ../RTL/cortexm0ds_logic.v(16929)
  and u20815 (Wycpw6, Dzcpw6, Kzcpw6);  // ../RTL/cortexm0ds_logic.v(16930)
  or u20816 (n5904, Z6aiu6, N20ju6);  // ../RTL/cortexm0ds_logic.v(16931)
  not u20817 (Kzcpw6, n5904);  // ../RTL/cortexm0ds_logic.v(16931)
  and u20818 (N20ju6, W8aiu6, Cyfpw6[6]);  // ../RTL/cortexm0ds_logic.v(16932)
  and u20819 (Z6aiu6, Vo3ju6, Pugiu6);  // ../RTL/cortexm0ds_logic.v(16933)
  or u2082 (n272, N73iu6, R7yhu6);  // ../RTL/cortexm0ds_logic.v(3875)
  and u20820 (Pugiu6, Cyfpw6[5], Tr0iu6);  // ../RTL/cortexm0ds_logic.v(16934)
  and u20821 (Dzcpw6, Rzcpw6, Yzcpw6);  // ../RTL/cortexm0ds_logic.v(16935)
  and u20822 (n5905, V9ghu6, F0dpw6);  // ../RTL/cortexm0ds_logic.v(16936)
  not u20823 (Yzcpw6, n5905);  // ../RTL/cortexm0ds_logic.v(16936)
  and u20824 (n5906, M0dpw6, T0dpw6);  // ../RTL/cortexm0ds_logic.v(16937)
  not u20825 (F0dpw6, n5906);  // ../RTL/cortexm0ds_logic.v(16937)
  and u20826 (n5907, A1dpw6, Vo3ju6);  // ../RTL/cortexm0ds_logic.v(16938)
  not u20827 (T0dpw6, n5907);  // ../RTL/cortexm0ds_logic.v(16938)
  or u20828 (n5908, Jcaiu6, D7fpw6[14]);  // ../RTL/cortexm0ds_logic.v(16939)
  not u20829 (A1dpw6, n5908);  // ../RTL/cortexm0ds_logic.v(16939)
  not u2083 (G73iu6, n272);  // ../RTL/cortexm0ds_logic.v(3875)
  buf u20830 (Eafpw6[11], Nxkbx6[12]);  // ../RTL/cortexm0ds_logic.v(3167)
  and u20831 (n5909, H1dpw6, Mr0iu6);  // ../RTL/cortexm0ds_logic.v(16941)
  not u20832 (M0dpw6, n5909);  // ../RTL/cortexm0ds_logic.v(16941)
  and u20833 (n5910, O1dpw6, V1dpw6);  // ../RTL/cortexm0ds_logic.v(16942)
  not u20834 (H1dpw6, n5910);  // ../RTL/cortexm0ds_logic.v(16942)
  and u20835 (n5911, C2dpw6, Kxziu6);  // ../RTL/cortexm0ds_logic.v(16943)
  not u20836 (V1dpw6, n5911);  // ../RTL/cortexm0ds_logic.v(16943)
  or u20837 (Qpaju6, Ae0iu6, D7fpw6[14]);  // ../RTL/cortexm0ds_logic.v(16944)
  not u20838 (Kxziu6, Qpaju6);  // ../RTL/cortexm0ds_logic.v(16944)
  or u20839 (n5912, Ii0iu6, Hbbow6);  // ../RTL/cortexm0ds_logic.v(16945)
  AL_MUX u2084 (
    .i0(Ubnhu6),
    .i1(Mmyhu6),
    .sel(U73iu6),
    .o(Ktxhu6));  // ../RTL/cortexm0ds_logic.v(3876)
  not u20840 (C2dpw6, n5912);  // ../RTL/cortexm0ds_logic.v(16945)
  and u20841 (Hbbow6, Dcziu6, J2dpw6);  // ../RTL/cortexm0ds_logic.v(16946)
  or u20842 (J2dpw6, Dzjiu6, A1kiu6);  // ../RTL/cortexm0ds_logic.v(16947)
  not u20843 (A1kiu6, D7fpw6[4]);  // ../RTL/cortexm0ds_logic.v(16948)
  not u20844 (Dzjiu6, D7fpw6[5]);  // ../RTL/cortexm0ds_logic.v(16949)
  and u20845 (n5913, Llaow6, Q2dpw6);  // ../RTL/cortexm0ds_logic.v(16950)
  not u20846 (O1dpw6, n5913);  // ../RTL/cortexm0ds_logic.v(16950)
  and u20847 (n5914, X2dpw6, Mpaow6);  // ../RTL/cortexm0ds_logic.v(16951)
  not u20848 (Q2dpw6, n5914);  // ../RTL/cortexm0ds_logic.v(16951)
  or u20849 (n5915, Y40ju6, Vk9ow6);  // ../RTL/cortexm0ds_logic.v(16952)
  and u2085 (U73iu6, B83iu6, Mdhpw6[0]);  // ../RTL/cortexm0ds_logic.v(3877)
  not u20850 (Mpaow6, n5915);  // ../RTL/cortexm0ds_logic.v(16952)
  and u20851 (Vk9ow6, X1ziu6, Ftjiu6);  // ../RTL/cortexm0ds_logic.v(16953)
  and u20852 (Y40ju6, D7fpw6[12], X1ziu6);  // ../RTL/cortexm0ds_logic.v(16954)
  or u20853 (n5916, E3dpw6, Jiiiu6);  // ../RTL/cortexm0ds_logic.v(16955)
  not u20854 (X2dpw6, n5916);  // ../RTL/cortexm0ds_logic.v(16955)
  and u20855 (Jiiiu6, Uriiu6, Ftjiu6);  // ../RTL/cortexm0ds_logic.v(16956)
  and u20856 (E3dpw6, Ya1ju6, D7fpw6[14]);  // ../RTL/cortexm0ds_logic.v(16957)
  or u20857 (n5917, Ftjiu6, D7fpw6[12]);  // ../RTL/cortexm0ds_logic.v(16958)
  not u20858 (Ya1ju6, n5917);  // ../RTL/cortexm0ds_logic.v(16958)
  or u20859 (Jcaiu6, Ae0iu6, Y7ghu6);  // ../RTL/cortexm0ds_logic.v(16959)
  or u2086 (n273, N5yhu6, I83iu6);  // ../RTL/cortexm0ds_logic.v(3878)
  not u20860 (Llaow6, Jcaiu6);  // ../RTL/cortexm0ds_logic.v(16959)
  and u20861 (n5918, K2aiu6, D6kiu6);  // ../RTL/cortexm0ds_logic.v(16960)
  not u20862 (Rzcpw6, n5918);  // ../RTL/cortexm0ds_logic.v(16960)
  or u20863 (n5919, Tfjiu6, K9aiu6);  // ../RTL/cortexm0ds_logic.v(16961)
  not u20864 (D6kiu6, n5919);  // ../RTL/cortexm0ds_logic.v(16961)
  and u20865 (K2aiu6, Ii0iu6, Xe8iu6);  // ../RTL/cortexm0ds_logic.v(16962)
  or u20866 (n5920, L3dpw6, S3dpw6);  // ../RTL/cortexm0ds_logic.v(16963)
  not u20867 (Pycpw6, n5920);  // ../RTL/cortexm0ds_logic.v(16963)
  AL_MUX u20868 (
    .i0(Z3dpw6),
    .i1(W8aiu6),
    .sel(Sbghu6),
    .o(S3dpw6));  // ../RTL/cortexm0ds_logic.v(16964)
  or u20869 (n5921, Knaiu6, Tr0iu6);  // ../RTL/cortexm0ds_logic.v(16965)
  not u2087 (B83iu6, n273);  // ../RTL/cortexm0ds_logic.v(3878)
  not u20870 (Z3dpw6, n5921);  // ../RTL/cortexm0ds_logic.v(16965)
  and u20871 (n5922, G4dpw6, N4dpw6);  // ../RTL/cortexm0ds_logic.v(16966)
  not u20872 (L3dpw6, n5922);  // ../RTL/cortexm0ds_logic.v(16966)
  or u20873 (N4dpw6, K9bow6, Xkaow6);  // ../RTL/cortexm0ds_logic.v(16967)
  not u20874 (Xkaow6, Hiaiu6);  // ../RTL/cortexm0ds_logic.v(16968)
  and u20875 (Hiaiu6, Zraiu6, Geaiu6);  // ../RTL/cortexm0ds_logic.v(16969)
  not u20876 (K9bow6, X97ow6);  // ../RTL/cortexm0ds_logic.v(16970)
  and u20877 (X97ow6, Cyfpw6[5], Mr0iu6);  // ../RTL/cortexm0ds_logic.v(16971)
  or u20878 (G4dpw6, P1bow6, Nlaiu6);  // ../RTL/cortexm0ds_logic.v(16972)
  not u20879 (P1bow6, Neoiu6);  // ../RTL/cortexm0ds_logic.v(16973)
  and u2088 (n274, P83iu6, W83iu6);  // ../RTL/cortexm0ds_logic.v(3879)
  and u20880 (Neoiu6, Cyfpw6[1], Zraiu6);  // ../RTL/cortexm0ds_logic.v(16974)
  buf u20881 (Eafpw6[10], Nxkbx6[11]);  // ../RTL/cortexm0ds_logic.v(3167)
  or u20882 (Lpcpw6, Sufpw6[0], Sufpw6[1]);  // ../RTL/cortexm0ds_logic.v(16976)
  and u20883 (n5923, U4dpw6, B5dpw6);  // ../RTL/cortexm0ds_logic.v(16977)
  and u20884 (n1272[0], S5iiu6, Z5iiu6);  // ../RTL/cortexm0ds_logic.v(16030)
  and u20885 (B5dpw6, I5dpw6, P5dpw6);  // ../RTL/cortexm0ds_logic.v(16978)
  or u20886 (n5924, W5dpw6, Nriiu6);  // ../RTL/cortexm0ds_logic.v(16979)
  not u20887 (P5dpw6, n5924);  // ../RTL/cortexm0ds_logic.v(16979)
  and u20888 (Nriiu6, D6dpw6, Vboiu6);  // ../RTL/cortexm0ds_logic.v(16980)
  or u20889 (n5925, E4jiu6, Cyfpw6[5]);  // ../RTL/cortexm0ds_logic.v(16981)
  not u2089 (Dtxhu6, n274);  // ../RTL/cortexm0ds_logic.v(3879)
  not u20890 (D6dpw6, n5925);  // ../RTL/cortexm0ds_logic.v(16981)
  not u20891 (E4jiu6, Hzziu6);  // ../RTL/cortexm0ds_logic.v(16982)
  and u20892 (Hzziu6, Cyfpw6[4], Jjhiu6);  // ../RTL/cortexm0ds_logic.v(16983)
  and u20893 (W5dpw6, K6dpw6, De6ow6);  // ../RTL/cortexm0ds_logic.v(16984)
  or u20894 (n5926, Vwaiu6, C0ehu6);  // ../RTL/cortexm0ds_logic.v(16985)
  not u20895 (De6ow6, n5926);  // ../RTL/cortexm0ds_logic.v(16985)
  not u20896 (Vwaiu6, Wp0iu6);  // ../RTL/cortexm0ds_logic.v(16986)
  and u20897 (Wp0iu6, Cyfpw6[0], Xe8iu6);  // ../RTL/cortexm0ds_logic.v(16987)
  not u20898 (Xe8iu6, Cyfpw6[5]);  // ../RTL/cortexm0ds_logic.v(16988)
  or u20899 (n5927, As0iu6, Knaiu6);  // ../RTL/cortexm0ds_logic.v(16989)
  buf u209 (Iahpw6[0], W6ipw6);  // ../RTL/cortexm0ds_logic.v(1883)
  and u2090 (W83iu6, D93iu6, K93iu6);  // ../RTL/cortexm0ds_logic.v(3880)
  not u20900 (K6dpw6, n5927);  // ../RTL/cortexm0ds_logic.v(16989)
  buf u20901 (Eafpw6[9], Nxkbx6[10]);  // ../RTL/cortexm0ds_logic.v(3167)
  or u20902 (As0iu6, Tfjiu6, Cyfpw6[4]);  // ../RTL/cortexm0ds_logic.v(16991)
  not u20903 (Ldoiu6, As0iu6);  // ../RTL/cortexm0ds_logic.v(16991)
  and u20904 (I5dpw6, R6dpw6, Y6dpw6);  // ../RTL/cortexm0ds_logic.v(16992)
  and u20905 (n5928, F7dpw6, F3aiu6);  // ../RTL/cortexm0ds_logic.v(16993)
  not u20906 (Y6dpw6, n5928);  // ../RTL/cortexm0ds_logic.v(16993)
  and u20907 (F3aiu6, Vo3ju6, Mr0iu6);  // ../RTL/cortexm0ds_logic.v(16994)
  or u20908 (Qxaiu6, Nlaiu6, Ii0iu6);  // ../RTL/cortexm0ds_logic.v(16995)
  not u20909 (Vo3ju6, Qxaiu6);  // ../RTL/cortexm0ds_logic.v(16995)
  and u2091 (n275, Uthpw6[6], Vk1iu6);  // ../RTL/cortexm0ds_logic.v(3881)
  or u20910 (n5929, Qjaiu6, C0ehu6);  // ../RTL/cortexm0ds_logic.v(16996)
  not u20911 (F7dpw6, n5929);  // ../RTL/cortexm0ds_logic.v(16996)
  not u20912 (Qjaiu6, U4kiu6);  // ../RTL/cortexm0ds_logic.v(16997)
  and u20913 (U4kiu6, Tr0iu6, Y2oiu6);  // ../RTL/cortexm0ds_logic.v(16998)
  and u20914 (n5930, Cyfpw6[7], M7dpw6);  // ../RTL/cortexm0ds_logic.v(16999)
  not u20915 (R6dpw6, n5930);  // ../RTL/cortexm0ds_logic.v(16999)
  and u20916 (n5931, Fmjiu6, T7dpw6);  // ../RTL/cortexm0ds_logic.v(17000)
  not u20917 (M7dpw6, n5931);  // ../RTL/cortexm0ds_logic.v(17000)
  or u20918 (T7dpw6, Uvziu6, Cyfpw6[0]);  // ../RTL/cortexm0ds_logic.v(17001)
  not u20919 (Uvziu6, Gsbow6);  // ../RTL/cortexm0ds_logic.v(17002)
  not u2092 (K93iu6, n275);  // ../RTL/cortexm0ds_logic.v(3881)
  and u20920 (Gsbow6, Cyfpw6[3], Y7ghu6);  // ../RTL/cortexm0ds_logic.v(17003)
  and u20921 (n5932, Pthiu6, Y7ghu6);  // ../RTL/cortexm0ds_logic.v(17004)
  not u20922 (Fmjiu6, n5932);  // ../RTL/cortexm0ds_logic.v(17004)
  and u20923 (U4dpw6, A8dpw6, H8dpw6);  // ../RTL/cortexm0ds_logic.v(17005)
  and u20924 (H8dpw6, O8dpw6, V8dpw6);  // ../RTL/cortexm0ds_logic.v(17006)
  and u20925 (n5933, C9dpw6, Ii0iu6);  // ../RTL/cortexm0ds_logic.v(17007)
  not u20926 (V8dpw6, n5933);  // ../RTL/cortexm0ds_logic.v(17007)
  not u20927 (Ii0iu6, Cyfpw6[3]);  // ../RTL/cortexm0ds_logic.v(17008)
  and u20928 (n5934, J9dpw6, Q9dpw6);  // ../RTL/cortexm0ds_logic.v(17009)
  not u20929 (C9dpw6, n5934);  // ../RTL/cortexm0ds_logic.v(17009)
  and u2093 (D93iu6, R93iu6, L72iu6);  // ../RTL/cortexm0ds_logic.v(3882)
  or u20930 (n5935, W8aiu6, Ae0iu6);  // ../RTL/cortexm0ds_logic.v(17010)
  not u20931 (Q9dpw6, n5935);  // ../RTL/cortexm0ds_logic.v(17010)
  and u20932 (W8aiu6, Y7ghu6, Mr0iu6);  // ../RTL/cortexm0ds_logic.v(17011)
  and u20933 (J9dpw6, X9dpw6, Kq0iu6);  // ../RTL/cortexm0ds_logic.v(17012)
  not u20934 (Kq0iu6, It2ju6);  // ../RTL/cortexm0ds_logic.v(17013)
  and u20935 (It2ju6, Y7ghu6, Y2oiu6);  // ../RTL/cortexm0ds_logic.v(17014)
  not u20936 (Y2oiu6, Cyfpw6[4]);  // ../RTL/cortexm0ds_logic.v(17015)
  or u20937 (X9dpw6, Pd6ow6, Sbghu6);  // ../RTL/cortexm0ds_logic.v(17016)
  and u20938 (n5936, Eadpw6, D1piu6);  // ../RTL/cortexm0ds_logic.v(17017)
  not u20939 (Pd6ow6, n5936);  // ../RTL/cortexm0ds_logic.v(17017)
  and u2094 (n276, Y93iu6, Pinhu6);  // ../RTL/cortexm0ds_logic.v(3883)
  or u20940 (n5937, Nlaiu6, C0ehu6);  // ../RTL/cortexm0ds_logic.v(17018)
  not u20941 (D1piu6, n5937);  // ../RTL/cortexm0ds_logic.v(17018)
  or u20942 (n5938, Wfoiu6, Knaiu6);  // ../RTL/cortexm0ds_logic.v(17019)
  not u20943 (Eadpw6, n5938);  // ../RTL/cortexm0ds_logic.v(17019)
  not u20944 (Knaiu6, Oiaiu6);  // ../RTL/cortexm0ds_logic.v(17020)
  and u20945 (Oiaiu6, Cyfpw6[7], Mr0iu6);  // ../RTL/cortexm0ds_logic.v(17021)
  not u20946 (Mr0iu6, H4ghu6);  // ../RTL/cortexm0ds_logic.v(17022)
  not u20947 (Wfoiu6, Vboiu6);  // ../RTL/cortexm0ds_logic.v(17023)
  and u20948 (Vboiu6, Cyfpw6[6], Tr0iu6);  // ../RTL/cortexm0ds_logic.v(17024)
  not u20949 (Tr0iu6, Cyfpw6[1]);  // ../RTL/cortexm0ds_logic.v(17025)
  not u2095 (R93iu6, n276);  // ../RTL/cortexm0ds_logic.v(3883)
  or u20950 (O8dpw6, S5qow6, Y31ju6);  // ../RTL/cortexm0ds_logic.v(17026)
  and u20951 (Y31ju6, Q5aiu6, Uriiu6);  // ../RTL/cortexm0ds_logic.v(17027)
  not u20952 (Uriiu6, S1ehu6);  // ../RTL/cortexm0ds_logic.v(17028)
  not u20953 (S5qow6, Imaiu6);  // ../RTL/cortexm0ds_logic.v(17029)
  and u20954 (Imaiu6, C0ehu6, Geaiu6);  // ../RTL/cortexm0ds_logic.v(17030)
  and u20955 (A8dpw6, Pmbow6, Ladpw6);  // ../RTL/cortexm0ds_logic.v(17031)
  and u20956 (n5939, Sadpw6, Geaiu6);  // ../RTL/cortexm0ds_logic.v(17032)
  not u20957 (Ladpw6, n5939);  // ../RTL/cortexm0ds_logic.v(17032)
  and u20958 (n5940, Zadpw6, Gbdpw6);  // ../RTL/cortexm0ds_logic.v(17033)
  not u20959 (Sadpw6, n5940);  // ../RTL/cortexm0ds_logic.v(17033)
  and u2096 (P83iu6, Fa3iu6, Ma3iu6);  // ../RTL/cortexm0ds_logic.v(3884)
  and u20960 (Gbdpw6, Nbdpw6, Ubdpw6);  // ../RTL/cortexm0ds_logic.v(17034)
  and u20961 (n5941, Bcdpw6, J5iow6);  // ../RTL/cortexm0ds_logic.v(17035)
  not u20962 (Ubdpw6, n5941);  // ../RTL/cortexm0ds_logic.v(17035)
  and u20963 (J5iow6, Icdpw6, D7fpw6[14]);  // ../RTL/cortexm0ds_logic.v(17036)
  or u20964 (n5942, D7fpw6[13], D7fpw6[15]);  // ../RTL/cortexm0ds_logic.v(17037)
  not u20965 (Icdpw6, n5942);  // ../RTL/cortexm0ds_logic.v(17037)
  and u20966 (Bcdpw6, P0piu6, Pcdpw6);  // ../RTL/cortexm0ds_logic.v(17038)
  and u20967 (n5943, Qjiow6, Wcdpw6);  // ../RTL/cortexm0ds_logic.v(17039)
  not u20968 (Pcdpw6, n5943);  // ../RTL/cortexm0ds_logic.v(17039)
  or u20969 (Wcdpw6, L7aow6, I6jiu6);  // ../RTL/cortexm0ds_logic.v(17040)
  and u2097 (n277, Iahpw6[6], Z4yhu6);  // ../RTL/cortexm0ds_logic.v(3885)
  not u20970 (I6jiu6, D7fpw6[10]);  // ../RTL/cortexm0ds_logic.v(17041)
  or u20971 (L7aow6, Rg2ju6, D7fpw6[8]);  // ../RTL/cortexm0ds_logic.v(17042)
  and u20972 (Qe0ju6, Dddpw6, Kddpw6);  // ../RTL/cortexm0ds_logic.v(17043)
  not u20973 (Rg2ju6, Qe0ju6);  // ../RTL/cortexm0ds_logic.v(17043)
  or u20974 (n5944, Ccaiu6, Prjiu6);  // ../RTL/cortexm0ds_logic.v(17044)
  not u20975 (Kddpw6, n5944);  // ../RTL/cortexm0ds_logic.v(17044)
  not u20976 (Prjiu6, D7fpw6[2]);  // ../RTL/cortexm0ds_logic.v(17045)
  or u20977 (n5945, O95iu6, Rb8iu6);  // ../RTL/cortexm0ds_logic.v(17046)
  not u20978 (Dddpw6, n5945);  // ../RTL/cortexm0ds_logic.v(17046)
  not u20979 (Qjiow6, Q6aow6);  // ../RTL/cortexm0ds_logic.v(17047)
  not u2098 (Ma3iu6, n277);  // ../RTL/cortexm0ds_logic.v(3885)
  and u20980 (Q6aow6, Qxoiu6, D7fpw6[8]);  // ../RTL/cortexm0ds_logic.v(17048)
  and u20981 (P0piu6, Mtjiu6, Oviiu6);  // ../RTL/cortexm0ds_logic.v(17049)
  and u20982 (Mtjiu6, C0ehu6, Gkiiu6);  // ../RTL/cortexm0ds_logic.v(17050)
  not u20983 (Gkiiu6, D7fpw6[12]);  // ../RTL/cortexm0ds_logic.v(17051)
  and u20984 (n5946, Rddpw6, A95iu6);  // ../RTL/cortexm0ds_logic.v(17052)
  not u20985 (Nbdpw6, n5946);  // ../RTL/cortexm0ds_logic.v(17052)
  or u20986 (n5947, N38ow6, D7fpw6[10]);  // ../RTL/cortexm0ds_logic.v(17053)
  not u20987 (A95iu6, n5947);  // ../RTL/cortexm0ds_logic.v(17053)
  not u20988 (N38ow6, Xiiiu6);  // ../RTL/cortexm0ds_logic.v(17054)
  and u20989 (Xiiiu6, D7fpw6[13], C0ehu6);  // ../RTL/cortexm0ds_logic.v(17055)
  and u2099 (Fa3iu6, Ta3iu6, Ab3iu6);  // ../RTL/cortexm0ds_logic.v(3886)
  and u20990 (Rddpw6, Aujiu6, Yddpw6);  // ../RTL/cortexm0ds_logic.v(17056)
  and u20991 (n5948, Fedpw6, Medpw6);  // ../RTL/cortexm0ds_logic.v(17057)
  not u20992 (Yddpw6, n5948);  // ../RTL/cortexm0ds_logic.v(17057)
  or u20993 (Medpw6, Kcziu6, Oviiu6);  // ../RTL/cortexm0ds_logic.v(17058)
  not u20994 (Kcziu6, L01ju6);  // ../RTL/cortexm0ds_logic.v(17059)
  and u20995 (L01ju6, D7fpw6[7], Ad8iu6);  // ../RTL/cortexm0ds_logic.v(17060)
  not u20996 (Ad8iu6, D7fpw6[6]);  // ../RTL/cortexm0ds_logic.v(17061)
  or u20997 (n5949, Il3ju6, D7fpw6[8]);  // ../RTL/cortexm0ds_logic.v(17062)
  not u20998 (Fedpw6, n5949);  // ../RTL/cortexm0ds_logic.v(17062)
  and u20999 (Aujiu6, D7fpw6[15], D7fpw6[12]);  // ../RTL/cortexm0ds_logic.v(17063)
  buf u21 (vis_r8_o[28], Rbibx6);  // ../RTL/cortexm0ds_logic.v(2579)
  buf u210 (vis_r2_o[11], C67bx6);  // ../RTL/cortexm0ds_logic.v(2551)
  and u2100 (n278, Ubnhu6, Cl1iu6);  // ../RTL/cortexm0ds_logic.v(3887)
  and u21000 (Zadpw6, Tedpw6, Afdpw6);  // ../RTL/cortexm0ds_logic.v(17064)
  and u21001 (n5950, J9kiu6, Hfdpw6);  // ../RTL/cortexm0ds_logic.v(17065)
  not u21002 (Afdpw6, n5950);  // ../RTL/cortexm0ds_logic.v(17065)
  and u21003 (n5951, Co6ow6, Ofdpw6);  // ../RTL/cortexm0ds_logic.v(17066)
  not u21004 (Hfdpw6, n5951);  // ../RTL/cortexm0ds_logic.v(17066)
  and u21005 (n5952, D7fpw6[12], Vfdpw6);  // ../RTL/cortexm0ds_logic.v(17067)
  not u21006 (Ofdpw6, n5952);  // ../RTL/cortexm0ds_logic.v(17067)
  and u21007 (n5953, Cgdpw6, Jgdpw6);  // ../RTL/cortexm0ds_logic.v(17068)
  not u21008 (Vfdpw6, n5953);  // ../RTL/cortexm0ds_logic.v(17068)
  and u21009 (n5954, D7fpw6[13], Qgdpw6);  // ../RTL/cortexm0ds_logic.v(17069)
  not u2101 (Ab3iu6, n278);  // ../RTL/cortexm0ds_logic.v(3887)
  not u21010 (Jgdpw6, n5954);  // ../RTL/cortexm0ds_logic.v(17069)
  or u21011 (Qgdpw6, Xgdpw6, Ehdpw6);  // ../RTL/cortexm0ds_logic.v(17070)
  and u21012 (Ehdpw6, Lhdpw6, Qxoiu6);  // ../RTL/cortexm0ds_logic.v(17071)
  or u21013 (n5955, Cwiiu6, D7fpw6[11]);  // ../RTL/cortexm0ds_logic.v(17072)
  not u21014 (Lhdpw6, n5955);  // ../RTL/cortexm0ds_logic.v(17072)
  and u21015 (Cwiiu6, Dcziu6, D7fpw6[5]);  // ../RTL/cortexm0ds_logic.v(17073)
  and u21016 (Dcziu6, D7fpw6[6], O95iu6);  // ../RTL/cortexm0ds_logic.v(17074)
  AL_MUX u21017 (
    .i0(F6ziu6),
    .i1(Shdpw6),
    .sel(D7fpw6[8]),
    .o(Xgdpw6));  // ../RTL/cortexm0ds_logic.v(17075)
  and u21018 (n5956, Zhdpw6, Gidpw6);  // ../RTL/cortexm0ds_logic.v(17076)
  not u21019 (Shdpw6, n5956);  // ../RTL/cortexm0ds_logic.v(17076)
  and u2102 (n279, Iahpw6[5], Xl1iu6);  // ../RTL/cortexm0ds_logic.v(3888)
  or u21020 (Gidpw6, Oviiu6, Wh0ju6);  // ../RTL/cortexm0ds_logic.v(17077)
  and u21021 (Wh0ju6, Nidpw6, R9aiu6);  // ../RTL/cortexm0ds_logic.v(17078)
  and u21022 (R9aiu6, Rb8iu6, Ccaiu6);  // ../RTL/cortexm0ds_logic.v(17079)
  not u21023 (Ccaiu6, D7fpw6[1]);  // ../RTL/cortexm0ds_logic.v(17080)
  not u21024 (Rb8iu6, D7fpw6[0]);  // ../RTL/cortexm0ds_logic.v(17081)
  or u21025 (n5957, D7fpw6[2], D7fpw6[3]);  // ../RTL/cortexm0ds_logic.v(17082)
  not u21026 (Nidpw6, n5957);  // ../RTL/cortexm0ds_logic.v(17082)
  buf u21027 (Ppfpw6[15], W8hbx6);  // ../RTL/cortexm0ds_logic.v(2461)
  not u21028 (Zhdpw6, Bl3ju6);  // ../RTL/cortexm0ds_logic.v(17083)
  and u21029 (Il3ju6, D7fpw6[11], Tniiu6);  // ../RTL/cortexm0ds_logic.v(17084)
  not u2103 (Ta3iu6, n279);  // ../RTL/cortexm0ds_logic.v(3888)
  not u21030 (Tniiu6, D7fpw6[9]);  // ../RTL/cortexm0ds_logic.v(17085)
  and u21031 (Zroiu6, D7fpw6[9], Oviiu6);  // ../RTL/cortexm0ds_logic.v(17086)
  and u21032 (n5958, F6ziu6, D7fpw6[14]);  // ../RTL/cortexm0ds_logic.v(17087)
  not u21033 (Cgdpw6, n5958);  // ../RTL/cortexm0ds_logic.v(17087)
  and u21034 (F6ziu6, Qxoiu6, D7fpw6[11]);  // ../RTL/cortexm0ds_logic.v(17088)
  not u21035 (Co6ow6, Hl8ow6);  // ../RTL/cortexm0ds_logic.v(17089)
  and u21036 (Hl8ow6, D7fpw6[13], D7fpw6[14]);  // ../RTL/cortexm0ds_logic.v(17090)
  or u21037 (n5959, Jjhiu6, Ftjiu6);  // ../RTL/cortexm0ds_logic.v(17091)
  not u21038 (J9kiu6, n5959);  // ../RTL/cortexm0ds_logic.v(17091)
  not u21039 (Ftjiu6, D7fpw6[15]);  // ../RTL/cortexm0ds_logic.v(17092)
  and u2104 (n280, Hb3iu6, Ob3iu6);  // ../RTL/cortexm0ds_logic.v(3889)
  or u21040 (Tedpw6, Ntgiu6, Cyfpw6[1]);  // ../RTL/cortexm0ds_logic.v(17093)
  and u21041 (n5960, Pthiu6, Yljiu6);  // ../RTL/cortexm0ds_logic.v(17094)
  not u21042 (Ntgiu6, n5960);  // ../RTL/cortexm0ds_logic.v(17094)
  and u21043 (Pthiu6, Nlaiu6, Tfjiu6);  // ../RTL/cortexm0ds_logic.v(17095)
  not u21044 (Tfjiu6, Cyfpw6[6]);  // ../RTL/cortexm0ds_logic.v(17096)
  and u21045 (Pmbow6, Faaiu6, Uidpw6);  // ../RTL/cortexm0ds_logic.v(17097)
  and u21046 (n5961, Xmliu6, Bjdpw6);  // ../RTL/cortexm0ds_logic.v(17098)
  not u21047 (Uidpw6, n5961);  // ../RTL/cortexm0ds_logic.v(17098)
  and u21048 (n5962, Ijdpw6, Pjdpw6);  // ../RTL/cortexm0ds_logic.v(17099)
  not u21049 (Bjdpw6, n5962);  // ../RTL/cortexm0ds_logic.v(17099)
  not u2105 (Wsxhu6, n280);  // ../RTL/cortexm0ds_logic.v(3889)
  and u21050 (n5963, Wjdpw6, Yljiu6);  // ../RTL/cortexm0ds_logic.v(17100)
  not u21051 (Pjdpw6, n5963);  // ../RTL/cortexm0ds_logic.v(17100)
  or u21052 (n5964, Cyfpw6[1], Cyfpw6[7]);  // ../RTL/cortexm0ds_logic.v(17101)
  not u21053 (Wjdpw6, n5964);  // ../RTL/cortexm0ds_logic.v(17101)
  or u21054 (Ijdpw6, G7oiu6, Iuniu6);  // ../RTL/cortexm0ds_logic.v(17102)
  not u21055 (Iuniu6, S6aiu6);  // ../RTL/cortexm0ds_logic.v(17103)
  and u21056 (S6aiu6, Yljiu6, H4ghu6);  // ../RTL/cortexm0ds_logic.v(17104)
  and u21057 (Yljiu6, Jjhiu6, K9aiu6);  // ../RTL/cortexm0ds_logic.v(17105)
  not u21058 (G7oiu6, L78ju6);  // ../RTL/cortexm0ds_logic.v(17106)
  and u21059 (L78ju6, Cyfpw6[4], Nlaiu6);  // ../RTL/cortexm0ds_logic.v(17107)
  and u2106 (Ob3iu6, Vb3iu6, Cc3iu6);  // ../RTL/cortexm0ds_logic.v(3890)
  not u21060 (Nlaiu6, Cyfpw6[0]);  // ../RTL/cortexm0ds_logic.v(17108)
  buf u21061 (Eafpw6[8], Nxkbx6[9]);  // ../RTL/cortexm0ds_logic.v(3167)
  and u21062 (Xmliu6, Dkdpw6, Kkdpw6);  // ../RTL/cortexm0ds_logic.v(17110)
  not u21063 (Taaiu6, Xmliu6);  // ../RTL/cortexm0ds_logic.v(17110)
  and u21064 (Kkdpw6, Rkdpw6, vis_pc_o[27]);  // ../RTL/cortexm0ds_logic.v(17111)
  or u21065 (n5965, Noliu6, Hlliu6);  // ../RTL/cortexm0ds_logic.v(17112)
  not u21066 (Rkdpw6, n5965);  // ../RTL/cortexm0ds_logic.v(17112)
  and u21067 (Hlliu6, Ykdpw6, H9row6);  // ../RTL/cortexm0ds_logic.v(17113)
  or u21068 (n5966, vis_ipsr_o[4], vis_ipsr_o[5]);  // ../RTL/cortexm0ds_logic.v(17114)
  not u21069 (H9row6, n5966);  // ../RTL/cortexm0ds_logic.v(17114)
  and u2107 (n281, Cl1iu6, Fanhu6);  // ../RTL/cortexm0ds_logic.v(3891)
  and u21070 (Ykdpw6, Ukbpw6, M8row6);  // ../RTL/cortexm0ds_logic.v(17115)
  or u21071 (n5967, vis_ipsr_o[2], vis_ipsr_o[3]);  // ../RTL/cortexm0ds_logic.v(17116)
  not u21072 (M8row6, n5967);  // ../RTL/cortexm0ds_logic.v(17116)
  or u21073 (Tnbpw6, vis_ipsr_o[0], vis_ipsr_o[1]);  // ../RTL/cortexm0ds_logic.v(17117)
  not u21074 (Ukbpw6, Tnbpw6);  // ../RTL/cortexm0ds_logic.v(17117)
  not u21075 (Noliu6, T6ehu6);  // ../RTL/cortexm0ds_logic.v(17118)
  and u21076 (Dkdpw6, Fldpw6, vis_pc_o[30]);  // ../RTL/cortexm0ds_logic.v(17119)
  and u21077 (Fldpw6, vis_pc_o[29], vis_pc_o[28]);  // ../RTL/cortexm0ds_logic.v(17120)
  not u21078 (Faaiu6, O4oiu6);  // ../RTL/cortexm0ds_logic.v(17121)
  and u21079 (O4oiu6, Ae0iu6, K9aiu6);  // ../RTL/cortexm0ds_logic.v(17122)
  not u2108 (Cc3iu6, n281);  // ../RTL/cortexm0ds_logic.v(3891)
  not u21080 (K9aiu6, Y7ghu6);  // ../RTL/cortexm0ds_logic.v(17123)
  or u21081 (n5968[0], Oi2ju6, D7fpw6[7]);  // ../RTL/cortexm0ds_logic.v(17124)
  not u21082 (O95iu6, D7fpw6[7]);  // ../RTL/cortexm0ds_logic.v(17125)
  not u21083 (Oi2ju6, Wf2ju6);  // ../RTL/cortexm0ds_logic.v(17127)
  and u21084 (Wf2ju6, Mldpw6, Tldpw6);  // ../RTL/cortexm0ds_logic.v(17128)
  and u21085 (Tldpw6, Amdpw6, Geaiu6);  // ../RTL/cortexm0ds_logic.v(17129)
  not u21086 (Geaiu6, Sbghu6);  // ../RTL/cortexm0ds_logic.v(17130)
  or u21087 (Amdpw6, Uyiiu6, Hmdpw6);  // ../RTL/cortexm0ds_logic.v(17131)
  or u21088 (n5969, Lraiu6, Qxoiu6);  // ../RTL/cortexm0ds_logic.v(17132)
  not u21089 (Hmdpw6, n5969);  // ../RTL/cortexm0ds_logic.v(17132)
  and u2109 (Vb3iu6, Jc3iu6, L72iu6);  // ../RTL/cortexm0ds_logic.v(3892)
  and u21090 (Qxoiu6, D7fpw6[10], D7fpw6[9]);  // ../RTL/cortexm0ds_logic.v(17133)
  and u21091 (Uyiiu6, Q5aiu6, Oviiu6);  // ../RTL/cortexm0ds_logic.v(17134)
  not u21092 (Oviiu6, D7fpw6[11]);  // ../RTL/cortexm0ds_logic.v(17135)
  not u21093 (Q5aiu6, Lraiu6);  // ../RTL/cortexm0ds_logic.v(17136)
  and u21094 (Lraiu6, Pzwiu6, Xbopw6);  // ../RTL/cortexm0ds_logic.v(17137)
  buf u21095 (Eafpw6[7], Nxkbx6[8]);  // ../RTL/cortexm0ds_logic.v(3167)
  and u21096 (Pzwiu6, Vchhu6, Jehhu6);  // ../RTL/cortexm0ds_logic.v(17139)
  and u21097 (Mldpw6, R7jiu6, Ia8iu6);  // ../RTL/cortexm0ds_logic.v(17140)
  or u21098 (n5970, X1ziu6, Ae0iu6);  // ../RTL/cortexm0ds_logic.v(17141)
  not u21099 (Ia8iu6, n5970);  // ../RTL/cortexm0ds_logic.v(17141)
  buf u211 (D7fpw6[6], W4jax6);  // ../RTL/cortexm0ds_logic.v(2074)
  and u2110 (n282, Uthpw6[5], Vk1iu6);  // ../RTL/cortexm0ds_logic.v(3893)
  or u21100 (Zraiu6, Vncpw6, E6phu6);  // ../RTL/cortexm0ds_logic.v(17142)
  not u21101 (Ae0iu6, Zraiu6);  // ../RTL/cortexm0ds_logic.v(17142)
  not u21102 (Vncpw6, Fvdhu6);  // ../RTL/cortexm0ds_logic.v(17143)
  not u21103 (X1ziu6, D7fpw6[14]);  // ../RTL/cortexm0ds_logic.v(17144)
  and u21104 (R7jiu6, Ozziu6, D7fpw6[15]);  // ../RTL/cortexm0ds_logic.v(17145)
  and u21105 (Ozziu6, Nbkiu6, D7fpw6[12]);  // ../RTL/cortexm0ds_logic.v(17146)
  or u21106 (Yb9ow6, Jjhiu6, D7fpw6[13]);  // ../RTL/cortexm0ds_logic.v(17147)
  not u21107 (Nbkiu6, Yb9ow6);  // ../RTL/cortexm0ds_logic.v(17147)
  not u21108 (Jjhiu6, C0ehu6);  // ../RTL/cortexm0ds_logic.v(17148)
  buf u21109 (R4gpw6[31], Oa5bx6);  // ../RTL/cortexm0ds_logic.v(2815)
  not u2111 (Jc3iu6, n282);  // ../RTL/cortexm0ds_logic.v(3893)
  not u21110 (n5971, PORESETn);  // ../RTL/cortexm0ds_logic.v(17151)
  buf u21111 (R4gpw6[30], M85bx6);  // ../RTL/cortexm0ds_logic.v(2815)
  buf u21112 (Ppfpw6[14], E6iax6);  // ../RTL/cortexm0ds_logic.v(2461)
  buf u21113 (R4gpw6[29], K65bx6);  // ../RTL/cortexm0ds_logic.v(2815)
  buf u21114 (Ppfpw6[13], W2jax6);  // ../RTL/cortexm0ds_logic.v(2461)
  buf u21115 (R4gpw6[28], Pjgbx6);  // ../RTL/cortexm0ds_logic.v(2815)
  not u21116 (n5972, Fmdhu6);  // ../RTL/cortexm0ds_logic.v(17169)
  buf u21117 (R4gpw6[27], I45bx6);  // ../RTL/cortexm0ds_logic.v(2815)
  buf u21118 (Ppfpw6[12], W0jax6);  // ../RTL/cortexm0ds_logic.v(2461)
  buf u21119 (R4gpw6[26], G25bx6);  // ../RTL/cortexm0ds_logic.v(2815)
  and u2112 (Hb3iu6, Qc3iu6, Xc3iu6);  // ../RTL/cortexm0ds_logic.v(3894)
  buf u21120 (Ppfpw6[11], Wyiax6);  // ../RTL/cortexm0ds_logic.v(2461)
  buf u21121 (R4gpw6[25], E05bx6);  // ../RTL/cortexm0ds_logic.v(2815)
  not u21122 (n5973, HRESETn);  // ../RTL/cortexm0ds_logic.v(17190)
  buf u21123 (R4gpw6[24], X7abx6);  // ../RTL/cortexm0ds_logic.v(2815)
  buf u21124 (Ppfpw6[10], Wwiax6);  // ../RTL/cortexm0ds_logic.v(2461)
  buf u21125 (R4gpw6[23], Sh4bx6);  // ../RTL/cortexm0ds_logic.v(2815)
  buf u21126 (Ppfpw6[9], Xuiax6);  // ../RTL/cortexm0ds_logic.v(2461)
  buf u21127 (Ppfpw6[8], Ysiax6);  // ../RTL/cortexm0ds_logic.v(2461)
  buf u21128 (R4gpw6[22], Qf4bx6);  // ../RTL/cortexm0ds_logic.v(2815)
  buf u21129 (Ppfpw6[7], Zqiax6);  // ../RTL/cortexm0ds_logic.v(2461)
  and u2113 (n283, Iahpw6[4], Xl1iu6);  // ../RTL/cortexm0ds_logic.v(3895)
  buf u21130 (R4gpw6[21], Od4bx6);  // ../RTL/cortexm0ds_logic.v(2815)
  buf u21131 (Ppfpw6[6], E8iax6);  // ../RTL/cortexm0ds_logic.v(2461)
  buf u21132 (R4gpw6[20], Rlgbx6);  // ../RTL/cortexm0ds_logic.v(2815)
  buf u21133 (Ppfpw6[5], F4iax6);  // ../RTL/cortexm0ds_logic.v(2461)
  buf u21134 (R4gpw6[19], Mb4bx6);  // ../RTL/cortexm0ds_logic.v(2815)
  buf u21135 (Ppfpw6[4], G2iax6);  // ../RTL/cortexm0ds_logic.v(2461)
  buf u21136 (R4gpw6[18], K94bx6);  // ../RTL/cortexm0ds_logic.v(2815)
  buf u21137 (Ppfpw6[3], Xiipw6);  // ../RTL/cortexm0ds_logic.v(2461)
  buf u21138 (R4gpw6[17], I74bx6);  // ../RTL/cortexm0ds_logic.v(2815)
  buf u21139 (Ppfpw6[2], Jpmpw6);  // ../RTL/cortexm0ds_logic.v(2461)
  not u2114 (Xc3iu6, n283);  // ../RTL/cortexm0ds_logic.v(3895)
  buf u21140 (R4gpw6[16], Z9abx6);  // ../RTL/cortexm0ds_logic.v(2815)
  not u21141 (n5974, DBGRESETn);  // ../RTL/cortexm0ds_logic.v(17262)
  buf u21142 (R4gpw6[15], Eyyax6);  // ../RTL/cortexm0ds_logic.v(2815)
  buf u21143 (Ppfpw6[1], T5mpw6);  // ../RTL/cortexm0ds_logic.v(2461)
  buf u21144 (R4gpw6[14], Cwyax6);  // ../RTL/cortexm0ds_logic.v(2815)
  not u21145 (Mifpw6[31], n112[31]);  // ../RTL/cortexm0ds_logic.v(3417)
  buf u21146 (R4gpw6[13], Auyax6);  // ../RTL/cortexm0ds_logic.v(2815)
  not u21147 (Mifpw6[30], n112[30]);  // ../RTL/cortexm0ds_logic.v(3417)
  buf u21148 (R4gpw6[12], Tngbx6);  // ../RTL/cortexm0ds_logic.v(2815)
  not u21149 (Mifpw6[29], n112[29]);  // ../RTL/cortexm0ds_logic.v(3417)
  and u2115 (n284, Iahpw6[5], Z4yhu6);  // ../RTL/cortexm0ds_logic.v(3896)
  buf u21150 (R4gpw6[11], Yryax6);  // ../RTL/cortexm0ds_logic.v(2815)
  not u21151 (Mifpw6[28], n112[28]);  // ../RTL/cortexm0ds_logic.v(3417)
  buf u21152 (R4gpw6[10], Vbspw6);  // ../RTL/cortexm0ds_logic.v(2815)
  not u21153 (Mifpw6[27], n112[27]);  // ../RTL/cortexm0ds_logic.v(3417)
  buf u21154 (R4gpw6[9], S3mpw6);  // ../RTL/cortexm0ds_logic.v(2815)
  not u21155 (Mifpw6[26], n112[26]);  // ../RTL/cortexm0ds_logic.v(3417)
  buf u21156 (R4gpw6[8], Bcabx6);  // ../RTL/cortexm0ds_logic.v(2815)
  not u21157 (Mifpw6[25], n112[25]);  // ../RTL/cortexm0ds_logic.v(3417)
  buf u21158 (R4gpw6[7], Tgzax6);  // ../RTL/cortexm0ds_logic.v(2815)
  not u21159 (Mifpw6[24], n112[24]);  // ../RTL/cortexm0ds_logic.v(3417)
  not u2116 (Qc3iu6, n284);  // ../RTL/cortexm0ds_logic.v(3896)
  buf u21160 (R4gpw6[6], Uizax6);  // ../RTL/cortexm0ds_logic.v(2815)
  not u21161 (Mifpw6[23], n112[23]);  // ../RTL/cortexm0ds_logic.v(3417)
  buf u21162 (R4gpw6[5], Vkzax6);  // ../RTL/cortexm0ds_logic.v(2815)
  not u21163 (Mifpw6[22], n112[22]);  // ../RTL/cortexm0ds_logic.v(3417)
  buf u21164 (R4gpw6[4], C5gbx6);  // ../RTL/cortexm0ds_logic.v(2815)
  not u21165 (Mifpw6[21], n112[21]);  // ../RTL/cortexm0ds_logic.v(3417)
  buf u21166 (R4gpw6[3], Wmzax6);  // ../RTL/cortexm0ds_logic.v(2815)
  not u21167 (Mifpw6[20], n112[20]);  // ../RTL/cortexm0ds_logic.v(3417)
  buf u21168 (R4gpw6[2], Xozax6);  // ../RTL/cortexm0ds_logic.v(2815)
  not u21169 (Mifpw6[19], n112[19]);  // ../RTL/cortexm0ds_logic.v(3417)
  and u2117 (n285, Ed3iu6, Ld3iu6);  // ../RTL/cortexm0ds_logic.v(3897)
  buf u21170 (R4gpw6[1], Yqzax6);  // ../RTL/cortexm0ds_logic.v(2815)
  not u21171 (Mifpw6[18], n112[18]);  // ../RTL/cortexm0ds_logic.v(3417)
  buf u21172 (H8gpw6[1], Elnpw6);  // ../RTL/cortexm0ds_logic.v(1877)
  not u21173 (Mifpw6[17], n112[17]);  // ../RTL/cortexm0ds_logic.v(3417)
  buf u21174 (Cyfpw6[7], Yvjpw6);  // ../RTL/cortexm0ds_logic.v(1807)
  not u21175 (Mifpw6[16], n112[16]);  // ../RTL/cortexm0ds_logic.v(3417)
  buf u21176 (Cyfpw6[6], Aujpw6);  // ../RTL/cortexm0ds_logic.v(1807)
  not u21177 (Mifpw6[15], n112[15]);  // ../RTL/cortexm0ds_logic.v(3417)
  buf u21178 (Cyfpw6[5], R3vpw6);  // ../RTL/cortexm0ds_logic.v(1807)
  not u21179 (Mifpw6[14], n112[14]);  // ../RTL/cortexm0ds_logic.v(3417)
  not u2118 (Psxhu6, n285);  // ../RTL/cortexm0ds_logic.v(3897)
  buf u21180 (Cyfpw6[4], T1vpw6);  // ../RTL/cortexm0ds_logic.v(1807)
  not u21181 (Mifpw6[13], n112[13]);  // ../RTL/cortexm0ds_logic.v(3417)
  buf u21182 (Cyfpw6[3], Ufopw6);  // ../RTL/cortexm0ds_logic.v(1807)
  not u21183 (Mifpw6[12], n112[12]);  // ../RTL/cortexm0ds_logic.v(3417)
  buf u21184 (Cyfpw6[1], Xxupw6);  // ../RTL/cortexm0ds_logic.v(1807)
  not u21185 (Mifpw6[11], n112[11]);  // ../RTL/cortexm0ds_logic.v(3417)
  buf u21186 (Odgpw6[31], Hg3bx6);  // ../RTL/cortexm0ds_logic.v(2789)
  not u21187 (Mifpw6[10], n112[10]);  // ../RTL/cortexm0ds_logic.v(3417)
  buf u21188 (Odgpw6[30], Tcipw6);  // ../RTL/cortexm0ds_logic.v(2789)
  not u21189 (Mifpw6[9], n112[9]);  // ../RTL/cortexm0ds_logic.v(3417)
  and u2119 (Ld3iu6, Sd3iu6, L72iu6);  // ../RTL/cortexm0ds_logic.v(3898)
  buf u21190 (Odgpw6[29], Bc3bx6);  // ../RTL/cortexm0ds_logic.v(2789)
  not u21191 (Mifpw6[8], n112[8]);  // ../RTL/cortexm0ds_logic.v(3417)
  buf u21192 (Odgpw6[28], V73bx6);  // ../RTL/cortexm0ds_logic.v(2789)
  not u21193 (Mifpw6[7], n112[7]);  // ../RTL/cortexm0ds_logic.v(3417)
  buf u21194 (Odgpw6[27], P33bx6);  // ../RTL/cortexm0ds_logic.v(2789)
  not u21195 (Mifpw6[6], n112[6]);  // ../RTL/cortexm0ds_logic.v(3417)
  buf u21196 (Odgpw6[26], Jz2bx6);  // ../RTL/cortexm0ds_logic.v(2789)
  not u21197 (Mifpw6[5], n112[5]);  // ../RTL/cortexm0ds_logic.v(3417)
  buf u21198 (Odgpw6[25], Rm2bx6);  // ../RTL/cortexm0ds_logic.v(2789)
  not u21199 (Mifpw6[4], n112[4]);  // ../RTL/cortexm0ds_logic.v(3417)
  buf u212 (vis_control_o, Npypw6);  // ../RTL/cortexm0ds_logic.v(2082)
  and u2120 (n286, Uthpw6[4], Vk1iu6);  // ../RTL/cortexm0ds_logic.v(3899)
  buf u21200 (Odgpw6[24], Dv2bx6);  // ../RTL/cortexm0ds_logic.v(2789)
  not u21201 (Mifpw6[3], n112[3]);  // ../RTL/cortexm0ds_logic.v(3417)
  buf u21202 (Odgpw6[23], Xq2bx6);  // ../RTL/cortexm0ds_logic.v(2789)
  not u21203 (Mifpw6[2], n112[2]);  // ../RTL/cortexm0ds_logic.v(3417)
  buf u21204 (Odgpw6[22], Y0gbx6);  // ../RTL/cortexm0ds_logic.v(2789)
  not u21205 (Mifpw6[1], n112[1]);  // ../RTL/cortexm0ds_logic.v(3417)
  buf u21206 (Odgpw6[21], Li2bx6);  // ../RTL/cortexm0ds_logic.v(2789)
  or u21207 (n111[31], Xuzhu6, Bxzhu6);  // ../RTL/cortexm0ds_logic.v(3385)
  buf u21208 (Odgpw6[20], Fe2bx6);  // ../RTL/cortexm0ds_logic.v(2789)
  or u21209 (n111[30], Xuzhu6, Ixzhu6);  // ../RTL/cortexm0ds_logic.v(3385)
  not u2121 (Sd3iu6, n286);  // ../RTL/cortexm0ds_logic.v(3899)
  buf u21210 (Odgpw6[19], V52bx6);  // ../RTL/cortexm0ds_logic.v(2789)
  or u21211 (n111[29], Xuzhu6, Wxzhu6);  // ../RTL/cortexm0ds_logic.v(3385)
  buf u21212 (Odgpw6[18], P12bx6);  // ../RTL/cortexm0ds_logic.v(2789)
  or u21213 (n111[28], Xuzhu6, Dyzhu6);  // ../RTL/cortexm0ds_logic.v(3385)
  buf u21214 (Odgpw6[17], Dt1bx6);  // ../RTL/cortexm0ds_logic.v(2789)
  or u21215 (n111[27], Kyzhu6, Xuzhu6);  // ../RTL/cortexm0ds_logic.v(3385)
  buf u21216 (Odgpw6[16], Jx1bx6);  // ../RTL/cortexm0ds_logic.v(2789)
  or u21217 (n111[26], Ryzhu6, Xuzhu6);  // ../RTL/cortexm0ds_logic.v(3385)
  buf u21218 (Odgpw6[15], Yxrpw6);  // ../RTL/cortexm0ds_logic.v(2789)
  or u21219 (n111[25], Yyzhu6, Xuzhu6);  // ../RTL/cortexm0ds_logic.v(3385)
  and u2122 (Ed3iu6, Zd3iu6, Ge3iu6);  // ../RTL/cortexm0ds_logic.v(3900)
  buf u21220 (Odgpw6[14], Xo1bx6);  // ../RTL/cortexm0ds_logic.v(2789)
  or u21221 (n111[24], Fzzhu6, Xuzhu6);  // ../RTL/cortexm0ds_logic.v(3385)
  buf u21222 (Odgpw6[13], Rk1bx6);  // ../RTL/cortexm0ds_logic.v(2789)
  or u21223 (n111[23], Mzzhu6, Xuzhu6);  // ../RTL/cortexm0ds_logic.v(3385)
  buf u21224 (Odgpw6[12], Z71bx6);  // ../RTL/cortexm0ds_logic.v(2789)
  or u21225 (n111[22], Tzzhu6, Xuzhu6);  // ../RTL/cortexm0ds_logic.v(3385)
  buf u21226 (Odgpw6[11], Lg1bx6);  // ../RTL/cortexm0ds_logic.v(2789)
  or u21227 (n111[21], A00iu6, Xuzhu6);  // ../RTL/cortexm0ds_logic.v(3385)
  buf u21228 (Odgpw6[10], Fc1bx6);  // ../RTL/cortexm0ds_logic.v(2789)
  or u21229 (n111[20], H00iu6, Xuzhu6);  // ../RTL/cortexm0ds_logic.v(3385)
  and u2123 (n287, Iahpw6[3], Xl1iu6);  // ../RTL/cortexm0ds_logic.v(3901)
  buf u21230 (Odgpw6[9], Rijbx6);  // ../RTL/cortexm0ds_logic.v(2789)
  or u21231 (n111[19], V00iu6, Xuzhu6);  // ../RTL/cortexm0ds_logic.v(3385)
  buf u21232 (Odgpw6[8], Us3bx6);  // ../RTL/cortexm0ds_logic.v(2789)
  or u21233 (n111[18], C10iu6, Xuzhu6);  // ../RTL/cortexm0ds_logic.v(3385)
  buf u21234 (Odgpw6[7], Qo3bx6);  // ../RTL/cortexm0ds_logic.v(2789)
  or u21235 (n111[17], J10iu6, Xuzhu6);  // ../RTL/cortexm0ds_logic.v(3385)
  buf u21236 (Odgpw6[6], Lr9bx6);  // ../RTL/cortexm0ds_logic.v(2789)
  or u21237 (n111[16], Q10iu6, Xuzhu6);  // ../RTL/cortexm0ds_logic.v(3385)
  buf u21238 (Odgpw6[5], Mk3bx6);  // ../RTL/cortexm0ds_logic.v(2789)
  or u21239 (n111[15], X10iu6, Xuzhu6);  // ../RTL/cortexm0ds_logic.v(3385)
  not u2124 (Ge3iu6, n287);  // ../RTL/cortexm0ds_logic.v(3901)
  buf u21240 (Odgpw6[4], Gihbx6);  // ../RTL/cortexm0ds_logic.v(2789)
  or u21241 (n111[14], Xuzhu6, E20iu6);  // ../RTL/cortexm0ds_logic.v(3385)
  buf u21242 (Odgpw6[3], Muhbx6);  // ../RTL/cortexm0ds_logic.v(2789)
  or u21243 (n111[13], L20iu6, Xuzhu6);  // ../RTL/cortexm0ds_logic.v(3385)
  buf u21244 (Odgpw6[2], N5bbx6);  // ../RTL/cortexm0ds_logic.v(2789)
  or u21245 (n111[12], Xuzhu6, S20iu6);  // ../RTL/cortexm0ds_logic.v(3385)
  buf u21246 (Odgpw6[1], Aa2bx6);  // ../RTL/cortexm0ds_logic.v(2789)
  or u21247 (n111[11], Xuzhu6, Z20iu6);  // ../RTL/cortexm0ds_logic.v(3385)
  buf u21248 (Gmhpw6[9], Vrkbx6[10]);  // ../RTL/cortexm0ds_logic.v(3109)
  or u21249 (n111[10], Xuzhu6, G30iu6);  // ../RTL/cortexm0ds_logic.v(3385)
  and u2125 (n288, Iahpw6[4], Z4yhu6);  // ../RTL/cortexm0ds_logic.v(3902)
  buf u21250 (Gmhpw6[8], Vrkbx6[9]);  // ../RTL/cortexm0ds_logic.v(3109)
  or u21251 (n111[9], Xuzhu6, Evzhu6);  // ../RTL/cortexm0ds_logic.v(3385)
  buf u21252 (Gmhpw6[7], Vrkbx6[8]);  // ../RTL/cortexm0ds_logic.v(3109)
  or u21253 (n111[8], Xuzhu6, Lvzhu6);  // ../RTL/cortexm0ds_logic.v(3385)
  buf u21254 (Gmhpw6[6], Vrkbx6[7]);  // ../RTL/cortexm0ds_logic.v(3109)
  or u21255 (n111[7], Xuzhu6, Svzhu6);  // ../RTL/cortexm0ds_logic.v(3385)
  buf u21256 (Gmhpw6[5], Vrkbx6[6]);  // ../RTL/cortexm0ds_logic.v(3109)
  or u21257 (n111[6], Xuzhu6, Zvzhu6);  // ../RTL/cortexm0ds_logic.v(3385)
  buf u21258 (Gmhpw6[4], Vrkbx6[5]);  // ../RTL/cortexm0ds_logic.v(3109)
  or u21259 (n111[5], Xuzhu6, Gwzhu6);  // ../RTL/cortexm0ds_logic.v(3385)
  not u2126 (Zd3iu6, n288);  // ../RTL/cortexm0ds_logic.v(3902)
  buf u21260 (Gmhpw6[3], Vrkbx6[4]);  // ../RTL/cortexm0ds_logic.v(3109)
  or u21261 (n111[4], Xuzhu6, Nwzhu6);  // ../RTL/cortexm0ds_logic.v(3385)
  buf u21262 (Gmhpw6[2], Vrkbx6[3]);  // ../RTL/cortexm0ds_logic.v(3109)
  or u21263 (n111[3], Xuzhu6, Uwzhu6);  // ../RTL/cortexm0ds_logic.v(3385)
  buf u21264 (Gmhpw6[1], Vrkbx6[2]);  // ../RTL/cortexm0ds_logic.v(3109)
  or u21265 (n111[2], Xuzhu6, Pxzhu6);  // ../RTL/cortexm0ds_logic.v(3385)
  AL_MUX u21266 (
    .i0(n5975),
    .i1(1'b0),
    .sel(Oakhu6),
    .o(Ntkbx6[0]));  // ../RTL/cortexm0ds_logic.v(3118)
  or u21267 (n111[1], Xuzhu6, O00iu6);  // ../RTL/cortexm0ds_logic.v(3385)
  AL_MUX u21268 (
    .i0(n5976),
    .i1(1'b0),
    .sel(Oakhu6),
    .o(Ntkbx6[1]));  // ../RTL/cortexm0ds_logic.v(3118)
  buf u21269 (Fkfpw6[31], Usnpw6);  // ../RTL/cortexm0ds_logic.v(1881)
  AL_MUX u2127 (
    .i0(Ne3iu6),
    .i1(N3nhu6),
    .sel(W13iu6),
    .o(Isxhu6));  // ../RTL/cortexm0ds_logic.v(3903)
  AL_MUX u21270 (
    .i0(n5977),
    .i1(1'b0),
    .sel(Oakhu6),
    .o(Ntkbx6[2]));  // ../RTL/cortexm0ds_logic.v(3118)
  buf u21271 (Fkfpw6[30], F6dbx6);  // ../RTL/cortexm0ds_logic.v(1881)
  AL_MUX u21272 (
    .i0(n5978),
    .i1(1'b0),
    .sel(Oakhu6),
    .o(Ntkbx6[3]));  // ../RTL/cortexm0ds_logic.v(3118)
  buf u21273 (Fkfpw6[29], Sx3qw6);  // ../RTL/cortexm0ds_logic.v(1881)
  AL_MUX u21274 (
    .i0(n5979),
    .i1(1'b0),
    .sel(Oakhu6),
    .o(Ntkbx6[4]));  // ../RTL/cortexm0ds_logic.v(3118)
  buf u21275 (Fkfpw6[28], Ibqpw6);  // ../RTL/cortexm0ds_logic.v(1881)
  AL_MUX u21276 (
    .i0(n5980),
    .i1(1'b0),
    .sel(Oakhu6),
    .o(Ntkbx6[5]));  // ../RTL/cortexm0ds_logic.v(3118)
  buf u21277 (Fkfpw6[27], Nybbx6);  // ../RTL/cortexm0ds_logic.v(1881)
  AL_MUX u21278 (
    .i0(n5981),
    .i1(1'b0),
    .sel(Oakhu6),
    .o(Ntkbx6[6]));  // ../RTL/cortexm0ds_logic.v(3118)
  buf u21279 (Fkfpw6[26], F8cbx6);  // ../RTL/cortexm0ds_logic.v(1881)
  and u2128 (Ne3iu6, Iahpw6[3], Ue3iu6);  // ../RTL/cortexm0ds_logic.v(3904)
  AL_MUX u21280 (
    .i0(n5982),
    .i1(1'b0),
    .sel(Oakhu6),
    .o(Ntkbx6[7]));  // ../RTL/cortexm0ds_logic.v(3118)
  buf u21281 (Fkfpw6[25], Nwbbx6);  // ../RTL/cortexm0ds_logic.v(1881)
  AL_MUX u21282 (
    .i0(n5983),
    .i1(1'b0),
    .sel(Oakhu6),
    .o(Ntkbx6[8]));  // ../RTL/cortexm0ds_logic.v(3118)
  buf u21283 (Fkfpw6[24], Tgkbx6);  // ../RTL/cortexm0ds_logic.v(1881)
  AL_MUX u21284 (
    .i0(n5984),
    .i1(1'b0),
    .sel(Oakhu6),
    .o(Ntkbx6[9]));  // ../RTL/cortexm0ds_logic.v(3118)
  buf u21285 (Fkfpw6[23], Ztgbx6);  // ../RTL/cortexm0ds_logic.v(1881)
  AL_MUX u21286 (
    .i0(n5985),
    .i1(1'b0),
    .sel(Oakhu6),
    .o(Ntkbx6[10]));  // ../RTL/cortexm0ds_logic.v(3118)
  buf u21287 (Fkfpw6[22], Tlebx6);  // ../RTL/cortexm0ds_logic.v(1881)
  AL_MUX u21288 (
    .i0(n5986),
    .i1(1'b0),
    .sel(Oakhu6),
    .o(Ntkbx6[11]));  // ../RTL/cortexm0ds_logic.v(3118)
  buf u21289 (Fkfpw6[21], M2ebx6);  // ../RTL/cortexm0ds_logic.v(1881)
  and u2129 (n289, T33iu6, Bf3iu6);  // ../RTL/cortexm0ds_logic.v(3905)
  AL_MUX u21290 (
    .i0(n5987),
    .i1(1'b0),
    .sel(Oakhu6),
    .o(Ntkbx6[12]));  // ../RTL/cortexm0ds_logic.v(3118)
  buf u21291 (Fkfpw6[20], Fjdbx6);  // ../RTL/cortexm0ds_logic.v(1881)
  AL_MUX u21292 (
    .i0(n5988),
    .i1(1'b0),
    .sel(Oakhu6),
    .o(Ntkbx6[13]));  // ../RTL/cortexm0ds_logic.v(3118)
  buf u21293 (Fkfpw6[19], T6kbx6);  // ../RTL/cortexm0ds_logic.v(1881)
  AL_MUX u21294 (
    .i0(n5989),
    .i1(1'b0),
    .sel(Oakhu6),
    .o(Ntkbx6[14]));  // ../RTL/cortexm0ds_logic.v(3118)
  buf u21295 (Fkfpw6[18], Syjbx6);  // ../RTL/cortexm0ds_logic.v(1881)
  buf u21296 (Fkfpw6[17], Pbbbx6);  // ../RTL/cortexm0ds_logic.v(1881)
  AL_MUX u21297 (
    .i0(1'b1),
    .i1(n5975),
    .sel(Oakhu6),
    .o(Ntkbx6[16]));  // ../RTL/cortexm0ds_logic.v(3118)
  buf u21298 (Fkfpw6[16], Chwpw6);  // ../RTL/cortexm0ds_logic.v(1881)
  AL_MUX u21299 (
    .i0(1'b1),
    .i1(n5976),
    .sel(Oakhu6),
    .o(Ntkbx6[17]));  // ../RTL/cortexm0ds_logic.v(3118)
  buf u213 (Vrfhu6, Jrypw6);  // ../RTL/cortexm0ds_logic.v(2083)
  not u2130 (Ue3iu6, n289);  // ../RTL/cortexm0ds_logic.v(3905)
  buf u21300 (Fkfpw6[15], Z47ax6);  // ../RTL/cortexm0ds_logic.v(1881)
  AL_MUX u21301 (
    .i0(1'b1),
    .i1(n5977),
    .sel(Oakhu6),
    .o(Ntkbx6[18]));  // ../RTL/cortexm0ds_logic.v(3118)
  buf u21302 (Fkfpw6[14], Sb8ax6);  // ../RTL/cortexm0ds_logic.v(1881)
  AL_MUX u21303 (
    .i0(1'b1),
    .i1(n5978),
    .sel(Oakhu6),
    .o(Ntkbx6[19]));  // ../RTL/cortexm0ds_logic.v(3118)
  buf u21304 (Fkfpw6[13], Xpxax6);  // ../RTL/cortexm0ds_logic.v(1881)
  AL_MUX u21305 (
    .i0(1'b1),
    .i1(n5979),
    .sel(Oakhu6),
    .o(Ntkbx6[20]));  // ../RTL/cortexm0ds_logic.v(3118)
  buf u21306 (Fkfpw6[12], Dm6bx6);  // ../RTL/cortexm0ds_logic.v(1881)
  AL_MUX u21307 (
    .i0(1'b1),
    .i1(n5980),
    .sel(Oakhu6),
    .o(Ntkbx6[21]));  // ../RTL/cortexm0ds_logic.v(3118)
  buf u21308 (Fkfpw6[11], C07bx6);  // ../RTL/cortexm0ds_logic.v(1881)
  AL_MUX u21309 (
    .i0(1'b1),
    .i1(n5981),
    .sel(Oakhu6),
    .o(Ntkbx6[22]));  // ../RTL/cortexm0ds_logic.v(3118)
  and u2131 (n290, If3iu6, Iahpw6[4]);  // ../RTL/cortexm0ds_logic.v(3906)
  buf u21310 (Fkfpw6[10], Gwxpw6);  // ../RTL/cortexm0ds_logic.v(1881)
  AL_MUX u21311 (
    .i0(1'b1),
    .i1(n5982),
    .sel(Oakhu6),
    .o(Ntkbx6[23]));  // ../RTL/cortexm0ds_logic.v(3118)
  buf u21312 (Fkfpw6[9], Kn1qw6);  // ../RTL/cortexm0ds_logic.v(1881)
  AL_MUX u21313 (
    .i0(1'b1),
    .i1(n5983),
    .sel(Oakhu6),
    .o(Ntkbx6[24]));  // ../RTL/cortexm0ds_logic.v(3118)
  buf u21314 (Fkfpw6[8], N61qw6);  // ../RTL/cortexm0ds_logic.v(1881)
  AL_MUX u21315 (
    .i0(1'b1),
    .i1(n5984),
    .sel(Oakhu6),
    .o(Ntkbx6[25]));  // ../RTL/cortexm0ds_logic.v(3118)
  buf u21316 (Fkfpw6[7], Asupw6);  // ../RTL/cortexm0ds_logic.v(1881)
  AL_MUX u21317 (
    .i0(1'b1),
    .i1(n5985),
    .sel(Oakhu6),
    .o(Ntkbx6[26]));  // ../RTL/cortexm0ds_logic.v(3118)
  buf u21318 (Fkfpw6[6], Ua9bx6);  // ../RTL/cortexm0ds_logic.v(1881)
  AL_MUX u21319 (
    .i0(1'b1),
    .i1(n5986),
    .sel(Oakhu6),
    .o(Ntkbx6[27]));  // ../RTL/cortexm0ds_logic.v(3118)
  not u2132 (Bf3iu6, n290);  // ../RTL/cortexm0ds_logic.v(3906)
  buf u21320 (Fkfpw6[5], Qc5bx6);  // ../RTL/cortexm0ds_logic.v(1881)
  AL_MUX u21321 (
    .i0(1'b1),
    .i1(n5987),
    .sel(Oakhu6),
    .o(Ntkbx6[28]));  // ../RTL/cortexm0ds_logic.v(3118)
  buf u21322 (Fkfpw6[4], Wtxax6);  // ../RTL/cortexm0ds_logic.v(1881)
  AL_MUX u21323 (
    .i0(1'b1),
    .i1(n5988),
    .sel(Oakhu6),
    .o(Ntkbx6[29]));  // ../RTL/cortexm0ds_logic.v(3118)
  buf u21324 (Fkfpw6[3], T5yax6);  // ../RTL/cortexm0ds_logic.v(1881)
  AL_MUX u21325 (
    .i0(1'b1),
    .i1(n5989),
    .sel(Oakhu6),
    .o(Ntkbx6[30]));  // ../RTL/cortexm0ds_logic.v(3118)
  buf u21326 (Fkfpw6[2], Xrxax6);  // ../RTL/cortexm0ds_logic.v(1881)
  not u21327 (Ntkbx6[15], Oakhu6);  // ../RTL/cortexm0ds_logic.v(3118)
  buf u21328 (Fkfpw6[1], Nu5bx6);  // ../RTL/cortexm0ds_logic.v(1881)
  AL_MUX u21329 (
    .i0(n5990),
    .i1(1'b0),
    .sel(G9khu6),
    .o(n5975));  // ../RTL/cortexm0ds_logic.v(3118)
  and u2133 (If3iu6, Iahpw6[5], Iahpw6[6]);  // ../RTL/cortexm0ds_logic.v(3907)
  or u21330 (n112[31], Xuzhu6, R50iu6);  // ../RTL/cortexm0ds_logic.v(3417)
  AL_MUX u21331 (
    .i0(n5991),
    .i1(1'b0),
    .sel(G9khu6),
    .o(n5976));  // ../RTL/cortexm0ds_logic.v(3118)
  or u21332 (n112[30], Xuzhu6, Y50iu6);  // ../RTL/cortexm0ds_logic.v(3417)
  AL_MUX u21333 (
    .i0(n5992),
    .i1(1'b0),
    .sel(G9khu6),
    .o(n5977));  // ../RTL/cortexm0ds_logic.v(3118)
  or u21334 (n112[29], Xuzhu6, M60iu6);  // ../RTL/cortexm0ds_logic.v(3417)
  AL_MUX u21335 (
    .i0(n5993),
    .i1(1'b0),
    .sel(G9khu6),
    .o(n5978));  // ../RTL/cortexm0ds_logic.v(3118)
  or u21336 (n112[28], Xuzhu6, T60iu6);  // ../RTL/cortexm0ds_logic.v(3417)
  AL_MUX u21337 (
    .i0(n5994),
    .i1(1'b0),
    .sel(G9khu6),
    .o(n5979));  // ../RTL/cortexm0ds_logic.v(3118)
  or u21338 (n112[27], Xuzhu6, A70iu6);  // ../RTL/cortexm0ds_logic.v(3417)
  AL_MUX u21339 (
    .i0(n5995),
    .i1(1'b0),
    .sel(G9khu6),
    .o(n5980));  // ../RTL/cortexm0ds_logic.v(3118)
  or u2134 (T33iu6, Pf3iu6, Iahpw6[4]);  // ../RTL/cortexm0ds_logic.v(3908)
  or u21340 (n112[26], Xuzhu6, H70iu6);  // ../RTL/cortexm0ds_logic.v(3417)
  AL_MUX u21341 (
    .i0(n5996),
    .i1(1'b0),
    .sel(G9khu6),
    .o(n5981));  // ../RTL/cortexm0ds_logic.v(3118)
  or u21342 (n112[25], Xuzhu6, O70iu6);  // ../RTL/cortexm0ds_logic.v(3417)
  or u21343 (n112[24], Xuzhu6, V70iu6);  // ../RTL/cortexm0ds_logic.v(3417)
  AL_MUX u21344 (
    .i0(1'b1),
    .i1(n5990),
    .sel(G9khu6),
    .o(n5983));  // ../RTL/cortexm0ds_logic.v(3118)
  or u21345 (n112[23], Xuzhu6, C80iu6);  // ../RTL/cortexm0ds_logic.v(3417)
  AL_MUX u21346 (
    .i0(1'b1),
    .i1(n5991),
    .sel(G9khu6),
    .o(n5984));  // ../RTL/cortexm0ds_logic.v(3118)
  or u21347 (n112[22], Xuzhu6, J80iu6);  // ../RTL/cortexm0ds_logic.v(3417)
  AL_MUX u21348 (
    .i0(1'b1),
    .i1(n5992),
    .sel(G9khu6),
    .o(n5985));  // ../RTL/cortexm0ds_logic.v(3118)
  or u21349 (n112[21], Xuzhu6, Q80iu6);  // ../RTL/cortexm0ds_logic.v(3417)
  or u2135 (Pf3iu6, Iahpw6[5], Iahpw6[6]);  // ../RTL/cortexm0ds_logic.v(3909)
  AL_MUX u21350 (
    .i0(1'b1),
    .i1(n5993),
    .sel(G9khu6),
    .o(n5986));  // ../RTL/cortexm0ds_logic.v(3118)
  or u21351 (n112[20], Xuzhu6, X80iu6);  // ../RTL/cortexm0ds_logic.v(3417)
  AL_MUX u21352 (
    .i0(1'b1),
    .i1(n5994),
    .sel(G9khu6),
    .o(n5987));  // ../RTL/cortexm0ds_logic.v(3118)
  or u21353 (n112[19], Xuzhu6, L90iu6);  // ../RTL/cortexm0ds_logic.v(3417)
  AL_MUX u21354 (
    .i0(1'b1),
    .i1(n5995),
    .sel(G9khu6),
    .o(n5988));  // ../RTL/cortexm0ds_logic.v(3118)
  or u21355 (n112[18], Xuzhu6, S90iu6);  // ../RTL/cortexm0ds_logic.v(3417)
  AL_MUX u21356 (
    .i0(1'b1),
    .i1(n5996),
    .sel(G9khu6),
    .o(n5989));  // ../RTL/cortexm0ds_logic.v(3118)
  or u21357 (n112[17], Xuzhu6, Z90iu6);  // ../RTL/cortexm0ds_logic.v(3417)
  not u21358 (n5982, G9khu6);  // ../RTL/cortexm0ds_logic.v(3118)
  or u21359 (n112[16], Xuzhu6, Ga0iu6);  // ../RTL/cortexm0ds_logic.v(3417)
  and u2136 (n291, Wf3iu6, Dg3iu6);  // ../RTL/cortexm0ds_logic.v(3910)
  or u21360 (n112[15], Xuzhu6, Na0iu6);  // ../RTL/cortexm0ds_logic.v(3417)
  or u21361 (n112[14], Xuzhu6, Ua0iu6);  // ../RTL/cortexm0ds_logic.v(3417)
  or u21362 (n112[13], Xuzhu6, Bb0iu6);  // ../RTL/cortexm0ds_logic.v(3417)
  or u21363 (n112[12], Xuzhu6, Ib0iu6);  // ../RTL/cortexm0ds_logic.v(3417)
  or u21364 (n112[11], Xuzhu6, Pb0iu6);  // ../RTL/cortexm0ds_logic.v(3417)
  or u21365 (n112[10], Xuzhu6, Wb0iu6);  // ../RTL/cortexm0ds_logic.v(3417)
  or u21366 (n112[9], Xuzhu6, U30iu6);  // ../RTL/cortexm0ds_logic.v(3417)
  or u21367 (n112[8], Xuzhu6, B40iu6);  // ../RTL/cortexm0ds_logic.v(3417)
  or u21368 (n112[7], Xuzhu6, I40iu6);  // ../RTL/cortexm0ds_logic.v(3417)
  or u21369 (n112[6], Xuzhu6, P40iu6);  // ../RTL/cortexm0ds_logic.v(3417)
  not u2137 (Bsxhu6, n291);  // ../RTL/cortexm0ds_logic.v(3910)
  or u21370 (n112[5], Xuzhu6, W40iu6);  // ../RTL/cortexm0ds_logic.v(3417)
  or u21371 (n112[4], Xuzhu6, D50iu6);  // ../RTL/cortexm0ds_logic.v(3417)
  or u21372 (n112[3], Xuzhu6, K50iu6);  // ../RTL/cortexm0ds_logic.v(3417)
  or u21373 (n112[2], Xuzhu6, F60iu6);  // ../RTL/cortexm0ds_logic.v(3417)
  or u21374 (n112[1], Xuzhu6, E90iu6);  // ../RTL/cortexm0ds_logic.v(3417)
  not u21375 (Tgfpw6[31], n111[31]);  // ../RTL/cortexm0ds_logic.v(3385)
  AL_MUX u21376 (
    .i0(n5997),
    .i1(1'b0),
    .sel(Y7khu6),
    .o(n5990));  // ../RTL/cortexm0ds_logic.v(3118)
  not u21377 (Tgfpw6[30], n111[30]);  // ../RTL/cortexm0ds_logic.v(3385)
  AL_MUX u21378 (
    .i0(n5998),
    .i1(1'b0),
    .sel(Y7khu6),
    .o(n5991));  // ../RTL/cortexm0ds_logic.v(3118)
  not u21379 (Tgfpw6[29], n111[29]);  // ../RTL/cortexm0ds_logic.v(3385)
  and u2138 (n292, Iahpw6[3], Z4yhu6);  // ../RTL/cortexm0ds_logic.v(3911)
  AL_MUX u21380 (
    .i0(n5999),
    .i1(1'b0),
    .sel(Y7khu6),
    .o(n5992));  // ../RTL/cortexm0ds_logic.v(3118)
  not u21381 (Tgfpw6[28], n111[28]);  // ../RTL/cortexm0ds_logic.v(3385)
  not u21382 (Tgfpw6[27], n111[27]);  // ../RTL/cortexm0ds_logic.v(3385)
  AL_MUX u21383 (
    .i0(1'b1),
    .i1(n5997),
    .sel(Y7khu6),
    .o(n5994));  // ../RTL/cortexm0ds_logic.v(3118)
  not u21384 (Tgfpw6[26], n111[26]);  // ../RTL/cortexm0ds_logic.v(3385)
  AL_MUX u21385 (
    .i0(1'b1),
    .i1(n5998),
    .sel(Y7khu6),
    .o(n5995));  // ../RTL/cortexm0ds_logic.v(3118)
  not u21386 (Tgfpw6[25], n111[25]);  // ../RTL/cortexm0ds_logic.v(3385)
  AL_MUX u21387 (
    .i0(1'b1),
    .i1(n5999),
    .sel(Y7khu6),
    .o(n5996));  // ../RTL/cortexm0ds_logic.v(3118)
  not u21388 (Tgfpw6[24], n111[24]);  // ../RTL/cortexm0ds_logic.v(3385)
  not u21389 (n5993, Y7khu6);  // ../RTL/cortexm0ds_logic.v(3118)
  not u2139 (Dg3iu6, n292);  // ../RTL/cortexm0ds_logic.v(3911)
  not u21390 (Tgfpw6[23], n111[23]);  // ../RTL/cortexm0ds_logic.v(3385)
  not u21391 (Tgfpw6[22], n111[22]);  // ../RTL/cortexm0ds_logic.v(3385)
  not u21392 (Tgfpw6[21], n111[21]);  // ../RTL/cortexm0ds_logic.v(3385)
  not u21393 (Tgfpw6[20], n111[20]);  // ../RTL/cortexm0ds_logic.v(3385)
  not u21394 (Tgfpw6[19], n111[19]);  // ../RTL/cortexm0ds_logic.v(3385)
  not u21395 (Tgfpw6[18], n111[18]);  // ../RTL/cortexm0ds_logic.v(3385)
  not u21396 (Tgfpw6[17], n111[17]);  // ../RTL/cortexm0ds_logic.v(3385)
  not u21397 (Tgfpw6[16], n111[16]);  // ../RTL/cortexm0ds_logic.v(3385)
  not u21398 (Tgfpw6[15], n111[15]);  // ../RTL/cortexm0ds_logic.v(3385)
  not u21399 (Tgfpw6[14], n111[14]);  // ../RTL/cortexm0ds_logic.v(3385)
  buf u214 (Shhpw6[10], C2ypw6);  // ../RTL/cortexm0ds_logic.v(1941)
  and u2140 (Wf3iu6, Kg3iu6, Rg3iu6);  // ../RTL/cortexm0ds_logic.v(3912)
  not u21400 (Tgfpw6[13], n111[13]);  // ../RTL/cortexm0ds_logic.v(3385)
  not u21401 (Tgfpw6[12], n111[12]);  // ../RTL/cortexm0ds_logic.v(3385)
  not u21402 (Tgfpw6[11], n111[11]);  // ../RTL/cortexm0ds_logic.v(3385)
  not u21403 (Tgfpw6[10], n111[10]);  // ../RTL/cortexm0ds_logic.v(3385)
  not u21404 (Tgfpw6[9], n111[9]);  // ../RTL/cortexm0ds_logic.v(3385)
  not u21405 (Tgfpw6[8], n111[8]);  // ../RTL/cortexm0ds_logic.v(3385)
  not u21406 (Tgfpw6[7], n111[7]);  // ../RTL/cortexm0ds_logic.v(3385)
  not u21407 (Tgfpw6[6], n111[6]);  // ../RTL/cortexm0ds_logic.v(3385)
  not u21408 (Tgfpw6[5], n111[5]);  // ../RTL/cortexm0ds_logic.v(3385)
  not u21409 (Tgfpw6[4], n111[4]);  // ../RTL/cortexm0ds_logic.v(3385)
  and u2141 (n293, Uthpw6[3], Vk1iu6);  // ../RTL/cortexm0ds_logic.v(3913)
  not u21410 (Tgfpw6[3], n111[3]);  // ../RTL/cortexm0ds_logic.v(3385)
  not u21411 (Tgfpw6[2], n111[2]);  // ../RTL/cortexm0ds_logic.v(3385)
  not u21412 (Tgfpw6[1], n111[1]);  // ../RTL/cortexm0ds_logic.v(3385)
  or u21413 (n114[23], Sg0iu6, Cf0iu6);  // ../RTL/cortexm0ds_logic.v(3453)
  or u21414 (n114[22], Pi0iu6, Cf0iu6);  // ../RTL/cortexm0ds_logic.v(3453)
  AL_MUX u21415 (
    .i0(n6000),
    .i1(1'b0),
    .sel(Q6khu6),
    .o(n5997));  // ../RTL/cortexm0ds_logic.v(3118)
  or u21416 (n114[21], Wi0iu6, Cf0iu6);  // ../RTL/cortexm0ds_logic.v(3453)
  or u21417 (n114[20], Yj0iu6, Cf0iu6);  // ../RTL/cortexm0ds_logic.v(3453)
  AL_MUX u21418 (
    .i0(1'b1),
    .i1(n6000),
    .sel(Q6khu6),
    .o(n5999));  // ../RTL/cortexm0ds_logic.v(3118)
  or u21419 (n114[19], Fk0iu6, Cf0iu6);  // ../RTL/cortexm0ds_logic.v(3453)
  not u2142 (Rg3iu6, n293);  // ../RTL/cortexm0ds_logic.v(3913)
  not u21420 (n5998, Q6khu6);  // ../RTL/cortexm0ds_logic.v(3118)
  or u21421 (n114[18], Mk0iu6, Cf0iu6);  // ../RTL/cortexm0ds_logic.v(3453)
  or u21422 (n114[17], Tk0iu6, Cf0iu6);  // ../RTL/cortexm0ds_logic.v(3453)
  or u21423 (n114[16], Al0iu6, Cf0iu6);  // ../RTL/cortexm0ds_logic.v(3453)
  or u21424 (n114[15], Ol0iu6, Cf0iu6);  // ../RTL/cortexm0ds_logic.v(3453)
  or u21425 (n114[14], Vl0iu6, Cf0iu6);  // ../RTL/cortexm0ds_logic.v(3453)
  or u21426 (n114[13], Cm0iu6, Cf0iu6);  // ../RTL/cortexm0ds_logic.v(3453)
  or u21427 (n114[12], Jm0iu6, Cf0iu6);  // ../RTL/cortexm0ds_logic.v(3453)
  or u21428 (n114[11], Qm0iu6, Cf0iu6);  // ../RTL/cortexm0ds_logic.v(3453)
  or u21429 (n114[10], Xm0iu6, Cf0iu6);  // ../RTL/cortexm0ds_logic.v(3453)
  and u2143 (n294, Xl1iu6, Iahpw6[2]);  // ../RTL/cortexm0ds_logic.v(3914)
  or u21430 (n114[9], En0iu6, Cf0iu6);  // ../RTL/cortexm0ds_logic.v(3453)
  or u21431 (n114[8], Ln0iu6, Cf0iu6);  // ../RTL/cortexm0ds_logic.v(3453)
  or u21432 (n114[7], Sn0iu6, Cf0iu6);  // ../RTL/cortexm0ds_logic.v(3453)
  or u21433 (n114[6], Zn0iu6, Cf0iu6);  // ../RTL/cortexm0ds_logic.v(3453)
  or u21434 (n114[5], Ve0iu6, Cf0iu6);  // ../RTL/cortexm0ds_logic.v(3453)
  or u21435 (n114[4], Jf0iu6, Cf0iu6);  // ../RTL/cortexm0ds_logic.v(3453)
  or u21436 (n114[3], Xf0iu6, Cf0iu6);  // ../RTL/cortexm0ds_logic.v(3453)
  or u21437 (n114[2], Eg0iu6, Cf0iu6);  // ../RTL/cortexm0ds_logic.v(3453)
  or u21438 (n114[1], Lg0iu6, Cf0iu6);  // ../RTL/cortexm0ds_logic.v(3453)
  not u21439 (Idfpw6[30], n114[23]);  // ../RTL/cortexm0ds_logic.v(3453)
  not u2144 (Kg3iu6, n294);  // ../RTL/cortexm0ds_logic.v(3914)
  not u21440 (Idfpw6[29], n114[22]);  // ../RTL/cortexm0ds_logic.v(3453)
  not u21441 (Idfpw6[28], n114[21]);  // ../RTL/cortexm0ds_logic.v(3453)
  not u21442 (Idfpw6[24], n114[20]);  // ../RTL/cortexm0ds_logic.v(3453)
  not u21443 (Idfpw6[23], n114[19]);  // ../RTL/cortexm0ds_logic.v(3453)
  not u21444 (Idfpw6[22], n114[18]);  // ../RTL/cortexm0ds_logic.v(3453)
  not u21445 (Idfpw6[21], n114[17]);  // ../RTL/cortexm0ds_logic.v(3453)
  not u21446 (Idfpw6[20], n114[16]);  // ../RTL/cortexm0ds_logic.v(3453)
  not u21447 (Idfpw6[19], n114[15]);  // ../RTL/cortexm0ds_logic.v(3453)
  not u21448 (Idfpw6[18], n114[14]);  // ../RTL/cortexm0ds_logic.v(3453)
  not u21449 (Idfpw6[17], n114[13]);  // ../RTL/cortexm0ds_logic.v(3453)
  and u2145 (n295, Yg3iu6, Fh3iu6);  // ../RTL/cortexm0ds_logic.v(3915)
  not u21450 (Idfpw6[16], n114[12]);  // ../RTL/cortexm0ds_logic.v(3453)
  not u21451 (Idfpw6[15], n114[11]);  // ../RTL/cortexm0ds_logic.v(3453)
  not u21452 (Idfpw6[14], n114[10]);  // ../RTL/cortexm0ds_logic.v(3453)
  not u21453 (Idfpw6[13], n114[9]);  // ../RTL/cortexm0ds_logic.v(3453)
  not u21454 (Idfpw6[12], n114[8]);  // ../RTL/cortexm0ds_logic.v(3453)
  not u21455 (Idfpw6[11], n114[7]);  // ../RTL/cortexm0ds_logic.v(3453)
  not u21456 (Idfpw6[10], n114[6]);  // ../RTL/cortexm0ds_logic.v(3453)
  not u21457 (Idfpw6[8], n114[5]);  // ../RTL/cortexm0ds_logic.v(3453)
  not u21458 (Idfpw6[7], n114[4]);  // ../RTL/cortexm0ds_logic.v(3453)
  not u21459 (Idfpw6[5], n114[3]);  // ../RTL/cortexm0ds_logic.v(3453)
  not u2146 (Urxhu6, n295);  // ../RTL/cortexm0ds_logic.v(3915)
  not u21460 (Idfpw6[4], n114[2]);  // ../RTL/cortexm0ds_logic.v(3453)
  not u21461 (Idfpw6[3], n114[1]);  // ../RTL/cortexm0ds_logic.v(3453)
  not u21462 (Qbfpw6[23], n2661[7]);  // ../RTL/cortexm0ds_logic.v(9500)
  not u21463 (Qbfpw6[10], n2661[6]);  // ../RTL/cortexm0ds_logic.v(9500)
  not u21464 (Qbfpw6[5], n2661[5]);  // ../RTL/cortexm0ds_logic.v(9500)
  not u21465 (Qbfpw6[4], n2661[4]);  // ../RTL/cortexm0ds_logic.v(9500)
  not u21466 (Qbfpw6[3], n2661[3]);  // ../RTL/cortexm0ds_logic.v(9500)
  not u21467 (Qbfpw6[2], n2661[2]);  // ../RTL/cortexm0ds_logic.v(9500)
  not u21468 (Qbfpw6[1], n2661[1]);  // ../RTL/cortexm0ds_logic.v(9500)
  and u21469 (Idfpw6[31], To2ju6, Oe0iu6);  // ../RTL/cortexm0ds_logic.v(9222)
  and u2147 (Fh3iu6, Mh3iu6, L72iu6);  // ../RTL/cortexm0ds_logic.v(3916)
  and u21470 (Idfpw6[27], Dj0iu6, Oe0iu6);  // ../RTL/cortexm0ds_logic.v(9222)
  and u21471 (Idfpw6[26], Kj0iu6, Oe0iu6);  // ../RTL/cortexm0ds_logic.v(9222)
  and u21472 (Idfpw6[25], Rj0iu6, Oe0iu6);  // ../RTL/cortexm0ds_logic.v(9222)
  and u21473 (Idfpw6[9], He0iu6, Oe0iu6);  // ../RTL/cortexm0ds_logic.v(9222)
  and u21474 (Idfpw6[6], Qf0iu6, Oe0iu6);  // ../RTL/cortexm0ds_logic.v(9222)
  and u21475 (Idfpw6[2], Zg0iu6, Gh0iu6);  // ../RTL/cortexm0ds_logic.v(9222)
  xor u21476 (n2661[7], Sh5ju6, Hu4ju6);  // ../RTL/cortexm0ds_logic.v(9500)
  xor u21477 (n2661[6], Fb8ju6, Hu4ju6);  // ../RTL/cortexm0ds_logic.v(9500)
  xor u21478 (n2661[5], Ua6ju6, Hu4ju6);  // ../RTL/cortexm0ds_logic.v(9500)
  xor u21479 (n2661[4], Au4ju6, Hu4ju6);  // ../RTL/cortexm0ds_logic.v(9500)
  and u2148 (n296, Uthpw6[2], Vk1iu6);  // ../RTL/cortexm0ds_logic.v(3917)
  xor u21480 (n2661[3], J16ju6, Hu4ju6);  // ../RTL/cortexm0ds_logic.v(9500)
  xor u21481 (n2661[2], Rr5ju6, Hu4ju6);  // ../RTL/cortexm0ds_logic.v(9500)
  buf u21482 (U0jhu6, Ntkbx6[30]);  // ../RTL/cortexm0ds_logic.v(3123)
  xor u21483 (n2661[1], Vd7ju6, Hu4ju6);  // ../RTL/cortexm0ds_logic.v(9500)
  buf u21484 (C2jhu6, Ntkbx6[29]);  // ../RTL/cortexm0ds_logic.v(3123)
  not u21485 (CODEHINTDE[2], n5923);  // ../RTL/cortexm0ds_logic.v(16977)
  buf u21486 (K3jhu6, Ntkbx6[28]);  // ../RTL/cortexm0ds_logic.v(3123)
  not u21487 (CODEHINTDE[1], n5968[1]);  // ../RTL/cortexm0ds_logic.v(16977)
  buf u21488 (S4jhu6, Ntkbx6[27]);  // ../RTL/cortexm0ds_logic.v(3123)
  and u21489 (n4277[31], Dhvow6, Khvow6);  // ../RTL/cortexm0ds_logic.v(14039)
  not u2149 (Mh3iu6, n296);  // ../RTL/cortexm0ds_logic.v(3917)
  buf u21490 (A6jhu6, Ntkbx6[26]);  // ../RTL/cortexm0ds_logic.v(3123)
  and u21491 (n4277[30], Crvow6, Jrvow6);  // ../RTL/cortexm0ds_logic.v(14039)
  buf u21492 (I7jhu6, Ntkbx6[25]);  // ../RTL/cortexm0ds_logic.v(3123)
  and u21493 (n4277[29], Lqqow6, Sqqow6);  // ../RTL/cortexm0ds_logic.v(14039)
  buf u21494 (Q8jhu6, Ntkbx6[24]);  // ../RTL/cortexm0ds_logic.v(3123)
  and u21495 (n4277[28], P1wow6, W1wow6);  // ../RTL/cortexm0ds_logic.v(14039)
  buf u21496 (Y9jhu6, Ntkbx6[23]);  // ../RTL/cortexm0ds_logic.v(3123)
  and u21497 (n4277[27], Obwow6, Vbwow6);  // ../RTL/cortexm0ds_logic.v(14039)
  buf u21498 (Gbjhu6, Ntkbx6[22]);  // ../RTL/cortexm0ds_logic.v(3123)
  and u21499 (n4277[26], Ulwow6, Bmwow6);  // ../RTL/cortexm0ds_logic.v(14039)
  buf u215 (S8fpw6[0], Sqkax6);  // ../RTL/cortexm0ds_logic.v(2451)
  and u2150 (Yg3iu6, Th3iu6, Ai3iu6);  // ../RTL/cortexm0ds_logic.v(3918)
  buf u21500 (Ocjhu6, Ntkbx6[21]);  // ../RTL/cortexm0ds_logic.v(3123)
  and u21501 (n4277[25], Tvwow6, Awwow6);  // ../RTL/cortexm0ds_logic.v(14039)
  buf u21502 (Wdjhu6, Ntkbx6[20]);  // ../RTL/cortexm0ds_logic.v(3123)
  and u21503 (n4277[24], Bexow6, Iexow6);  // ../RTL/cortexm0ds_logic.v(14039)
  buf u21504 (Efjhu6, Ntkbx6[19]);  // ../RTL/cortexm0ds_logic.v(3123)
  and u21505 (n4277[23], Jwxow6, Qwxow6);  // ../RTL/cortexm0ds_logic.v(14039)
  buf u21506 (Mgjhu6, Ntkbx6[18]);  // ../RTL/cortexm0ds_logic.v(3123)
  and u21507 (n4277[22], U5yow6, B6yow6);  // ../RTL/cortexm0ds_logic.v(14039)
  buf u21508 (Uhjhu6, Ntkbx6[17]);  // ../RTL/cortexm0ds_logic.v(3123)
  and u21509 (n4277[21], Ffyow6, Mfyow6);  // ../RTL/cortexm0ds_logic.v(14039)
  and u2151 (n297, Xl1iu6, Iahpw6[1]);  // ../RTL/cortexm0ds_logic.v(3919)
  buf u21510 (Cjjhu6, Ntkbx6[16]);  // ../RTL/cortexm0ds_logic.v(3123)
  and u21511 (n4277[20], Qoyow6, Xoyow6);  // ../RTL/cortexm0ds_logic.v(14039)
  buf u21512 (Kkjhu6, Ntkbx6[15]);  // ../RTL/cortexm0ds_logic.v(3123)
  and u21513 (n4277[19], Pyyow6, Wyyow6);  // ../RTL/cortexm0ds_logic.v(14039)
  buf u21514 (Sljhu6, Ntkbx6[14]);  // ../RTL/cortexm0ds_logic.v(3123)
  and u21515 (n4277[18], A8zow6, H8zow6);  // ../RTL/cortexm0ds_logic.v(14039)
  buf u21516 (Anjhu6, Ntkbx6[13]);  // ../RTL/cortexm0ds_logic.v(3123)
  and u21517 (n4277[17], Lhzow6, Shzow6);  // ../RTL/cortexm0ds_logic.v(14039)
  buf u21518 (Iojhu6, Ntkbx6[12]);  // ../RTL/cortexm0ds_logic.v(3123)
  and u21519 (n4277[16], Xbqow6, Ecqow6);  // ../RTL/cortexm0ds_logic.v(14039)
  not u2152 (Ai3iu6, n297);  // ../RTL/cortexm0ds_logic.v(3919)
  buf u21520 (Qpjhu6, Ntkbx6[11]);  // ../RTL/cortexm0ds_logic.v(3123)
  and u21521 (n4277[15], Kyzow6, Ryzow6);  // ../RTL/cortexm0ds_logic.v(14039)
  buf u21522 (Yqjhu6, Ntkbx6[10]);  // ../RTL/cortexm0ds_logic.v(3123)
  and u21523 (n4277[14], Eg0pw6, Lg0pw6);  // ../RTL/cortexm0ds_logic.v(14039)
  buf u21524 (Gsjhu6, Ntkbx6[9]);  // ../RTL/cortexm0ds_logic.v(3123)
  and u21525 (n4277[13], Rx0pw6, Yx0pw6);  // ../RTL/cortexm0ds_logic.v(14039)
  buf u21526 (Otjhu6, Ntkbx6[8]);  // ../RTL/cortexm0ds_logic.v(3123)
  and u21527 (n4277[12], Ef1pw6, Lf1pw6);  // ../RTL/cortexm0ds_logic.v(14039)
  buf u21528 (Wujhu6, Ntkbx6[7]);  // ../RTL/cortexm0ds_logic.v(3123)
  and u21529 (n4277[11], Rw1pw6, Yw1pw6);  // ../RTL/cortexm0ds_logic.v(14039)
  and u2153 (n298, Iahpw6[2], Z4yhu6);  // ../RTL/cortexm0ds_logic.v(3920)
  buf u21530 (Ewjhu6, Ntkbx6[6]);  // ../RTL/cortexm0ds_logic.v(3123)
  and u21531 (n4277[10], Ee2pw6, Le2pw6);  // ../RTL/cortexm0ds_logic.v(14039)
  buf u21532 (Mxjhu6, Ntkbx6[5]);  // ../RTL/cortexm0ds_logic.v(3123)
  and u21533 (n4277[9], Tbvow6, Acvow6);  // ../RTL/cortexm0ds_logic.v(14039)
  buf u21534 (Uyjhu6, Ntkbx6[4]);  // ../RTL/cortexm0ds_logic.v(3123)
  and u21535 (n4277[8], Cdvow6, Jdvow6);  // ../RTL/cortexm0ds_logic.v(14039)
  buf u21536 (C0khu6, Ntkbx6[3]);  // ../RTL/cortexm0ds_logic.v(3123)
  and u21537 (n4277[7], Eevow6, Levow6);  // ../RTL/cortexm0ds_logic.v(14039)
  buf u21538 (K1khu6, Ntkbx6[2]);  // ../RTL/cortexm0ds_logic.v(3123)
  and u21539 (n4277[6], Zevow6, Gfvow6);  // ../RTL/cortexm0ds_logic.v(14039)
  not u2154 (Th3iu6, n298);  // ../RTL/cortexm0ds_logic.v(3920)
  buf u21540 (S2khu6, Ntkbx6[1]);  // ../RTL/cortexm0ds_logic.v(3123)
  and u21541 (n4277[5], Nfvow6, Ufvow6);  // ../RTL/cortexm0ds_logic.v(14039)
  AL_MUX u21542 (
    .i0(n6001),
    .i1(1'b0),
    .sel(Msmhu6),
    .o(Nvkbx6[0]));  // ../RTL/cortexm0ds_logic.v(3132)
  and u21543 (n4277[4], Bgvow6, Igvow6);  // ../RTL/cortexm0ds_logic.v(14039)
  AL_MUX u21544 (
    .i0(n6002),
    .i1(1'b0),
    .sel(Msmhu6),
    .o(Nvkbx6[1]));  // ../RTL/cortexm0ds_logic.v(3132)
  and u21545 (n4277[3], Pgvow6, Wgvow6);  // ../RTL/cortexm0ds_logic.v(14039)
  AL_MUX u21546 (
    .i0(n6003),
    .i1(1'b0),
    .sel(Msmhu6),
    .o(Nvkbx6[2]));  // ../RTL/cortexm0ds_logic.v(3132)
  and u21547 (n4277[2], B1wow6, I1wow6);  // ../RTL/cortexm0ds_logic.v(14039)
  AL_MUX u21548 (
    .i0(n6004),
    .i1(1'b0),
    .sel(Msmhu6),
    .o(Nvkbx6[3]));  // ../RTL/cortexm0ds_logic.v(3132)
  and u21549 (n4277[1], Byyow6, Iyyow6);  // ../RTL/cortexm0ds_logic.v(14039)
  and u2155 (n299, Hi3iu6, Oi3iu6);  // ../RTL/cortexm0ds_logic.v(3921)
  AL_MUX u21550 (
    .i0(n6005),
    .i1(1'b0),
    .sel(Msmhu6),
    .o(Nvkbx6[4]));  // ../RTL/cortexm0ds_logic.v(3132)
  not u21551 (HWDATA[31], n4277[31]);  // ../RTL/cortexm0ds_logic.v(14039)
  AL_MUX u21552 (
    .i0(n6006),
    .i1(1'b0),
    .sel(Msmhu6),
    .o(Nvkbx6[5]));  // ../RTL/cortexm0ds_logic.v(3132)
  not u21553 (HWDATA[30], n4277[30]);  // ../RTL/cortexm0ds_logic.v(14039)
  AL_MUX u21554 (
    .i0(n6007),
    .i1(1'b0),
    .sel(Msmhu6),
    .o(Nvkbx6[6]));  // ../RTL/cortexm0ds_logic.v(3132)
  not u21555 (HWDATA[29], n4277[29]);  // ../RTL/cortexm0ds_logic.v(14039)
  AL_MUX u21556 (
    .i0(n6008),
    .i1(1'b0),
    .sel(Msmhu6),
    .o(Nvkbx6[7]));  // ../RTL/cortexm0ds_logic.v(3132)
  not u21557 (HWDATA[28], n4277[28]);  // ../RTL/cortexm0ds_logic.v(14039)
  AL_MUX u21558 (
    .i0(n6009),
    .i1(1'b0),
    .sel(Msmhu6),
    .o(Nvkbx6[8]));  // ../RTL/cortexm0ds_logic.v(3132)
  not u21559 (HWDATA[27], n4277[27]);  // ../RTL/cortexm0ds_logic.v(14039)
  not u2156 (Nrxhu6, n299);  // ../RTL/cortexm0ds_logic.v(3921)
  AL_MUX u21560 (
    .i0(n6010),
    .i1(1'b0),
    .sel(Msmhu6),
    .o(Nvkbx6[9]));  // ../RTL/cortexm0ds_logic.v(3132)
  not u21561 (HWDATA[26], n4277[26]);  // ../RTL/cortexm0ds_logic.v(14039)
  AL_MUX u21562 (
    .i0(n6011),
    .i1(1'b0),
    .sel(Msmhu6),
    .o(Nvkbx6[10]));  // ../RTL/cortexm0ds_logic.v(3132)
  not u21563 (HWDATA[25], n4277[25]);  // ../RTL/cortexm0ds_logic.v(14039)
  AL_MUX u21564 (
    .i0(n6012),
    .i1(1'b0),
    .sel(Msmhu6),
    .o(Nvkbx6[11]));  // ../RTL/cortexm0ds_logic.v(3132)
  not u21565 (HWDATA[24], n4277[24]);  // ../RTL/cortexm0ds_logic.v(14039)
  AL_MUX u21566 (
    .i0(n6013),
    .i1(1'b0),
    .sel(Msmhu6),
    .o(Nvkbx6[12]));  // ../RTL/cortexm0ds_logic.v(3132)
  not u21567 (HWDATA[23], n4277[23]);  // ../RTL/cortexm0ds_logic.v(14039)
  AL_MUX u21568 (
    .i0(n6014),
    .i1(1'b0),
    .sel(Msmhu6),
    .o(Nvkbx6[13]));  // ../RTL/cortexm0ds_logic.v(3132)
  not u21569 (HWDATA[22], n4277[22]);  // ../RTL/cortexm0ds_logic.v(14039)
  and u2157 (n300, Vi3iu6, B7nhu6);  // ../RTL/cortexm0ds_logic.v(3922)
  AL_MUX u21570 (
    .i0(n6015),
    .i1(1'b0),
    .sel(Msmhu6),
    .o(Nvkbx6[14]));  // ../RTL/cortexm0ds_logic.v(3132)
  not u21571 (HWDATA[21], n4277[21]);  // ../RTL/cortexm0ds_logic.v(14039)
  not u21572 (HWDATA[20], n4277[20]);  // ../RTL/cortexm0ds_logic.v(14039)
  AL_MUX u21573 (
    .i0(1'b1),
    .i1(n6001),
    .sel(Msmhu6),
    .o(Nvkbx6[16]));  // ../RTL/cortexm0ds_logic.v(3132)
  not u21574 (HWDATA[19], n4277[19]);  // ../RTL/cortexm0ds_logic.v(14039)
  AL_MUX u21575 (
    .i0(1'b1),
    .i1(n6002),
    .sel(Msmhu6),
    .o(Nvkbx6[17]));  // ../RTL/cortexm0ds_logic.v(3132)
  not u21576 (HWDATA[18], n4277[18]);  // ../RTL/cortexm0ds_logic.v(14039)
  AL_MUX u21577 (
    .i0(1'b1),
    .i1(n6003),
    .sel(Msmhu6),
    .o(Nvkbx6[18]));  // ../RTL/cortexm0ds_logic.v(3132)
  not u21578 (HWDATA[17], n4277[17]);  // ../RTL/cortexm0ds_logic.v(14039)
  AL_MUX u21579 (
    .i0(1'b1),
    .i1(n6004),
    .sel(Msmhu6),
    .o(Nvkbx6[19]));  // ../RTL/cortexm0ds_logic.v(3132)
  not u2158 (Oi3iu6, n300);  // ../RTL/cortexm0ds_logic.v(3922)
  not u21580 (HWDATA[16], n4277[16]);  // ../RTL/cortexm0ds_logic.v(14039)
  AL_MUX u21581 (
    .i0(1'b1),
    .i1(n6005),
    .sel(Msmhu6),
    .o(Nvkbx6[20]));  // ../RTL/cortexm0ds_logic.v(3132)
  not u21582 (HWDATA[15], n4277[15]);  // ../RTL/cortexm0ds_logic.v(14039)
  AL_MUX u21583 (
    .i0(1'b1),
    .i1(n6006),
    .sel(Msmhu6),
    .o(Nvkbx6[21]));  // ../RTL/cortexm0ds_logic.v(3132)
  not u21584 (HWDATA[14], n4277[14]);  // ../RTL/cortexm0ds_logic.v(14039)
  AL_MUX u21585 (
    .i0(1'b1),
    .i1(n6007),
    .sel(Msmhu6),
    .o(Nvkbx6[22]));  // ../RTL/cortexm0ds_logic.v(3132)
  not u21586 (HWDATA[13], n4277[13]);  // ../RTL/cortexm0ds_logic.v(14039)
  AL_MUX u21587 (
    .i0(1'b1),
    .i1(n6008),
    .sel(Msmhu6),
    .o(Nvkbx6[23]));  // ../RTL/cortexm0ds_logic.v(3132)
  not u21588 (HWDATA[12], n4277[12]);  // ../RTL/cortexm0ds_logic.v(14039)
  AL_MUX u21589 (
    .i0(1'b1),
    .i1(n6009),
    .sel(Msmhu6),
    .o(Nvkbx6[24]));  // ../RTL/cortexm0ds_logic.v(3132)
  and u2159 (Vi3iu6, Cj3iu6, L02iu6);  // ../RTL/cortexm0ds_logic.v(3923)
  not u21590 (HWDATA[11], n4277[11]);  // ../RTL/cortexm0ds_logic.v(14039)
  AL_MUX u21591 (
    .i0(1'b1),
    .i1(n6010),
    .sel(Msmhu6),
    .o(Nvkbx6[25]));  // ../RTL/cortexm0ds_logic.v(3132)
  not u21592 (HWDATA[10], n4277[10]);  // ../RTL/cortexm0ds_logic.v(14039)
  AL_MUX u21593 (
    .i0(1'b1),
    .i1(n6011),
    .sel(Msmhu6),
    .o(Nvkbx6[26]));  // ../RTL/cortexm0ds_logic.v(3132)
  not u21594 (HWDATA[9], n4277[9]);  // ../RTL/cortexm0ds_logic.v(14039)
  AL_MUX u21595 (
    .i0(1'b1),
    .i1(n6012),
    .sel(Msmhu6),
    .o(Nvkbx6[27]));  // ../RTL/cortexm0ds_logic.v(3132)
  not u21596 (HWDATA[8], n4277[8]);  // ../RTL/cortexm0ds_logic.v(14039)
  AL_MUX u21597 (
    .i0(1'b1),
    .i1(n6013),
    .sel(Msmhu6),
    .o(Nvkbx6[28]));  // ../RTL/cortexm0ds_logic.v(3132)
  not u21598 (HWDATA[7], n4277[7]);  // ../RTL/cortexm0ds_logic.v(14039)
  AL_MUX u21599 (
    .i0(1'b1),
    .i1(n6014),
    .sel(Msmhu6),
    .o(Nvkbx6[29]));  // ../RTL/cortexm0ds_logic.v(3132)
  buf u216 (vis_r12_o[13], Estax6);  // ../RTL/cortexm0ds_logic.v(2599)
  and u2160 (n301, Vx2iu6, Jj3iu6);  // ../RTL/cortexm0ds_logic.v(3924)
  not u21600 (HWDATA[6], n4277[6]);  // ../RTL/cortexm0ds_logic.v(14039)
  AL_MUX u21601 (
    .i0(1'b1),
    .i1(n6015),
    .sel(Msmhu6),
    .o(Nvkbx6[30]));  // ../RTL/cortexm0ds_logic.v(3132)
  not u21602 (HWDATA[5], n4277[5]);  // ../RTL/cortexm0ds_logic.v(14039)
  not u21603 (Nvkbx6[15], Msmhu6);  // ../RTL/cortexm0ds_logic.v(3132)
  not u21604 (HWDATA[4], n4277[4]);  // ../RTL/cortexm0ds_logic.v(14039)
  AL_MUX u21605 (
    .i0(n6016),
    .i1(1'b0),
    .sel(Frmhu6),
    .o(n6001));  // ../RTL/cortexm0ds_logic.v(3132)
  not u21606 (HWDATA[3], n4277[3]);  // ../RTL/cortexm0ds_logic.v(14039)
  AL_MUX u21607 (
    .i0(n6017),
    .i1(1'b0),
    .sel(Frmhu6),
    .o(n6002));  // ../RTL/cortexm0ds_logic.v(3132)
  not u21608 (HWDATA[2], n4277[2]);  // ../RTL/cortexm0ds_logic.v(14039)
  AL_MUX u21609 (
    .i0(n6018),
    .i1(1'b0),
    .sel(Frmhu6),
    .o(n6003));  // ../RTL/cortexm0ds_logic.v(3132)
  not u2161 (Cj3iu6, n301);  // ../RTL/cortexm0ds_logic.v(3924)
  not u21610 (HWDATA[1], n4277[1]);  // ../RTL/cortexm0ds_logic.v(14039)
  AL_MUX u21611 (
    .i0(n6019),
    .i1(1'b0),
    .sel(Frmhu6),
    .o(n6004));  // ../RTL/cortexm0ds_logic.v(3132)
  not u21612 (HSIZE[1], Cc3pw6);  // ../RTL/cortexm0ds_logic.v(15237)
  AL_MUX u21613 (
    .i0(n6020),
    .i1(1'b0),
    .sel(Frmhu6),
    .o(n6005));  // ../RTL/cortexm0ds_logic.v(3132)
  and u21614 (n5200[1], HPROT[2], Ue3pw6);  // ../RTL/cortexm0ds_logic.v(15247)
  AL_MUX u21615 (
    .i0(n6021),
    .i1(1'b0),
    .sel(Frmhu6),
    .o(n6006));  // ../RTL/cortexm0ds_logic.v(3132)
  not u21616 (HADDR[1], n5488[1]);  // ../RTL/cortexm0ds_logic.v(15829)
  AL_MUX u21617 (
    .i0(n6022),
    .i1(1'b0),
    .sel(Frmhu6),
    .o(n6007));  // ../RTL/cortexm0ds_logic.v(3132)
  buf u21618 (HBURST[2], 1'b0);  // ../RTL/cortexm0ds_logic.v(1725)
  buf u21619 (HBURST[1], 1'b0);  // ../RTL/cortexm0ds_logic.v(1725)
  and u2162 (n302, A1zhu6, Qj3iu6);  // ../RTL/cortexm0ds_logic.v(3925)
  AL_MUX u21620 (
    .i0(1'b1),
    .i1(n6016),
    .sel(Frmhu6),
    .o(n6009));  // ../RTL/cortexm0ds_logic.v(3132)
  and u21621 (n5488[1], Y57pw6, F67pw6);  // ../RTL/cortexm0ds_logic.v(15829)
  AL_MUX u21622 (
    .i0(1'b1),
    .i1(n6017),
    .sel(Frmhu6),
    .o(n6010));  // ../RTL/cortexm0ds_logic.v(3132)
  buf u21623 (Lwgpw6[2], Vz8ax6);  // ../RTL/cortexm0ds_logic.v(2229)
  AL_MUX u21624 (
    .i0(1'b1),
    .i1(n6018),
    .sel(Frmhu6),
    .o(n6011));  // ../RTL/cortexm0ds_logic.v(3132)
  buf u21625 (Lwgpw6[1], R19ax6);  // ../RTL/cortexm0ds_logic.v(2229)
  AL_MUX u21626 (
    .i0(1'b1),
    .i1(n6019),
    .sel(Frmhu6),
    .o(n6012));  // ../RTL/cortexm0ds_logic.v(3132)
  and u21627 (n1272[12], Ng8pw6, Ug8pw6);  // ../RTL/cortexm0ds_logic.v(16030)
  AL_MUX u21628 (
    .i0(1'b1),
    .i1(n6020),
    .sel(Frmhu6),
    .o(n6013));  // ../RTL/cortexm0ds_logic.v(3132)
  and u21629 (n1272[11], Rp8pw6, Yp8pw6);  // ../RTL/cortexm0ds_logic.v(16030)
  not u2163 (Jj3iu6, n302);  // ../RTL/cortexm0ds_logic.v(3925)
  AL_MUX u21630 (
    .i0(1'b1),
    .i1(n6021),
    .sel(Frmhu6),
    .o(n6014));  // ../RTL/cortexm0ds_logic.v(3132)
  and u21631 (Iu9iu6, Vy8pw6, Cz8pw6);  // ../RTL/cortexm0ds_logic.v(16030)
  AL_MUX u21632 (
    .i0(1'b1),
    .i1(n6022),
    .sel(Frmhu6),
    .o(n6015));  // ../RTL/cortexm0ds_logic.v(3132)
  and u21633 (n1272[9], Ypmiu6, Fqmiu6);  // ../RTL/cortexm0ds_logic.v(16030)
  not u21634 (n6008, Frmhu6);  // ../RTL/cortexm0ds_logic.v(3132)
  and u21635 (n1272[8], Kwmiu6, Rwmiu6);  // ../RTL/cortexm0ds_logic.v(16030)
  and u21636 (n1272[7], Yu3pw6, Fv3pw6);  // ../RTL/cortexm0ds_logic.v(16030)
  and u21637 (n1272[6], A5niu6, H5niu6);  // ../RTL/cortexm0ds_logic.v(16030)
  and u21638 (n1272[5], Mskiu6, Tskiu6);  // ../RTL/cortexm0ds_logic.v(16030)
  and u21639 (n1272[4], C44pw6, J44pw6);  // ../RTL/cortexm0ds_logic.v(16030)
  or u2164 (Qj3iu6, Hknhu6, K7yhu6);  // ../RTL/cortexm0ds_logic.v(3926)
  and u21640 (n1272[3], Omkiu6, Vmkiu6);  // ../RTL/cortexm0ds_logic.v(16030)
  and u21641 (n1272[2], R1iiu6, Y1iiu6);  // ../RTL/cortexm0ds_logic.v(16030)
  and u21642 (n1272[1], Gikiu6, Nikiu6);  // ../RTL/cortexm0ds_logic.v(16030)
  or u21643 (n5968[1], Oi2ju6, O95iu6);  // ../RTL/cortexm0ds_logic.v(17124)
  buf u21644 (WICSENSE[33], 1'b0);  // ../RTL/cortexm0ds_logic.v(1767)
  buf u21645 (WICSENSE[32], 1'b0);  // ../RTL/cortexm0ds_logic.v(1767)
  buf u21646 (WICSENSE[31], 1'b0);  // ../RTL/cortexm0ds_logic.v(1767)
  buf u21647 (WICSENSE[30], 1'b0);  // ../RTL/cortexm0ds_logic.v(1767)
  buf u21648 (WICSENSE[29], 1'b0);  // ../RTL/cortexm0ds_logic.v(1767)
  buf u21649 (WICSENSE[28], 1'b0);  // ../RTL/cortexm0ds_logic.v(1767)
  AL_MUX u2165 (
    .i0(1'b1),
    .i1(n6026),
    .sel(Romhu6),
    .o(n6025));  // ../RTL/cortexm0ds_logic.v(3132)
  buf u21650 (WICSENSE[27], 1'b0);  // ../RTL/cortexm0ds_logic.v(1767)
  buf u21651 (WICSENSE[26], 1'b0);  // ../RTL/cortexm0ds_logic.v(1767)
  AL_MUX u21652 (
    .i0(n6023),
    .i1(1'b0),
    .sel(Ypmhu6),
    .o(n6016));  // ../RTL/cortexm0ds_logic.v(3132)
  buf u21653 (WICSENSE[25], 1'b0);  // ../RTL/cortexm0ds_logic.v(1767)
  AL_MUX u21654 (
    .i0(n6024),
    .i1(1'b0),
    .sel(Ypmhu6),
    .o(n6017));  // ../RTL/cortexm0ds_logic.v(3132)
  buf u21655 (WICSENSE[24], 1'b0);  // ../RTL/cortexm0ds_logic.v(1767)
  AL_MUX u21656 (
    .i0(n6025),
    .i1(1'b0),
    .sel(Ypmhu6),
    .o(n6018));  // ../RTL/cortexm0ds_logic.v(3132)
  buf u21657 (WICSENSE[23], 1'b0);  // ../RTL/cortexm0ds_logic.v(1767)
  buf u21658 (WICSENSE[22], 1'b0);  // ../RTL/cortexm0ds_logic.v(1767)
  AL_MUX u21659 (
    .i0(1'b1),
    .i1(n6023),
    .sel(Ypmhu6),
    .o(n6020));  // ../RTL/cortexm0ds_logic.v(3132)
  and u2166 (n303, Q8nhu6, Ek3iu6);  // ../RTL/cortexm0ds_logic.v(3928)
  buf u21660 (WICSENSE[21], 1'b0);  // ../RTL/cortexm0ds_logic.v(1767)
  AL_MUX u21661 (
    .i0(1'b1),
    .i1(n6024),
    .sel(Ypmhu6),
    .o(n6021));  // ../RTL/cortexm0ds_logic.v(3132)
  buf u21662 (WICSENSE[20], 1'b0);  // ../RTL/cortexm0ds_logic.v(1767)
  AL_MUX u21663 (
    .i0(1'b1),
    .i1(n6025),
    .sel(Ypmhu6),
    .o(n6022));  // ../RTL/cortexm0ds_logic.v(3132)
  buf u21664 (WICSENSE[19], 1'b0);  // ../RTL/cortexm0ds_logic.v(1767)
  buf u21665 (WICSENSE[18], 1'b0);  // ../RTL/cortexm0ds_logic.v(1767)
  buf u21666 (WICSENSE[17], 1'b0);  // ../RTL/cortexm0ds_logic.v(1767)
  buf u21667 (WICSENSE[16], 1'b0);  // ../RTL/cortexm0ds_logic.v(1767)
  buf u21668 (WICSENSE[15], 1'b0);  // ../RTL/cortexm0ds_logic.v(1767)
  buf u21669 (WICSENSE[14], 1'b0);  // ../RTL/cortexm0ds_logic.v(1767)
  not u2167 (Hi3iu6, n303);  // ../RTL/cortexm0ds_logic.v(3928)
  buf u21670 (WICSENSE[13], 1'b0);  // ../RTL/cortexm0ds_logic.v(1767)
  buf u21671 (WICSENSE[12], 1'b0);  // ../RTL/cortexm0ds_logic.v(1767)
  buf u21672 (WICSENSE[11], 1'b0);  // ../RTL/cortexm0ds_logic.v(1767)
  buf u21673 (WICSENSE[10], 1'b0);  // ../RTL/cortexm0ds_logic.v(1767)
  buf u21674 (WICSENSE[9], 1'b0);  // ../RTL/cortexm0ds_logic.v(1767)
  buf u21675 (WICSENSE[8], 1'b0);  // ../RTL/cortexm0ds_logic.v(1767)
  buf u21676 (WICSENSE[7], 1'b0);  // ../RTL/cortexm0ds_logic.v(1767)
  buf u21677 (WICSENSE[6], 1'b0);  // ../RTL/cortexm0ds_logic.v(1767)
  buf u21678 (WICSENSE[5], 1'b0);  // ../RTL/cortexm0ds_logic.v(1767)
  buf u21679 (WICSENSE[4], 1'b0);  // ../RTL/cortexm0ds_logic.v(1767)
  and u2168 (n304, Iahpw6[3], Di1iu6);  // ../RTL/cortexm0ds_logic.v(3929)
  buf u21680 (WICSENSE[3], 1'b0);  // ../RTL/cortexm0ds_logic.v(1767)
  buf u21681 (WICSENSE[2], 1'b0);  // ../RTL/cortexm0ds_logic.v(1767)
  buf u21682 (WICSENSE[1], 1'b0);  // ../RTL/cortexm0ds_logic.v(1767)
  buf u21683 (WICSENSE[0], 1'b0);  // ../RTL/cortexm0ds_logic.v(1767)
  not u2169 (Ek3iu6, n304);  // ../RTL/cortexm0ds_logic.v(3929)
  buf u217 (Shhpw6[8], Gc1qw6);  // ../RTL/cortexm0ds_logic.v(1941)
  and u2170 (n305, Lk3iu6, Sk3iu6);  // ../RTL/cortexm0ds_logic.v(3930)
  not u2171 (Grxhu6, n305);  // ../RTL/cortexm0ds_logic.v(3930)
  and u2172 (Sk3iu6, Zk3iu6, Gl3iu6);  // ../RTL/cortexm0ds_logic.v(3931)
  and u2173 (n306, Q8nhu6, Cl1iu6);  // ../RTL/cortexm0ds_logic.v(3932)
  not u2174 (Gl3iu6, n306);  // ../RTL/cortexm0ds_logic.v(3932)
  and u2175 (Zk3iu6, Nl3iu6, L72iu6);  // ../RTL/cortexm0ds_logic.v(3933)
  and u2176 (n307, Uthpw6[1], Vk1iu6);  // ../RTL/cortexm0ds_logic.v(3934)
  not u2177 (Nl3iu6, n307);  // ../RTL/cortexm0ds_logic.v(3934)
  and u2178 (Lk3iu6, Ul3iu6, Bm3iu6);  // ../RTL/cortexm0ds_logic.v(3935)
  and u2179 (n308, Iahpw6[0], Xl1iu6);  // ../RTL/cortexm0ds_logic.v(3936)
  buf u218 (Shhpw6[9], Gl1qw6);  // ../RTL/cortexm0ds_logic.v(1941)
  not u2180 (Bm3iu6, n308);  // ../RTL/cortexm0ds_logic.v(3936)
  and u2181 (n309, Iahpw6[1], Z4yhu6);  // ../RTL/cortexm0ds_logic.v(3937)
  not u2182 (Ul3iu6, n309);  // ../RTL/cortexm0ds_logic.v(3937)
  and u2183 (n310, Im3iu6, Pm3iu6);  // ../RTL/cortexm0ds_logic.v(3938)
  not u2184 (Zqxhu6, n310);  // ../RTL/cortexm0ds_logic.v(3938)
  and u2185 (Pm3iu6, Wm3iu6, Dn3iu6);  // ../RTL/cortexm0ds_logic.v(3939)
  and u2186 (n311, B7nhu6, Cl1iu6);  // ../RTL/cortexm0ds_logic.v(3940)
  not u2187 (Dn3iu6, n311);  // ../RTL/cortexm0ds_logic.v(3940)
  and u2188 (Cl1iu6, Kn3iu6, Y93iu6);  // ../RTL/cortexm0ds_logic.v(3941)
  and u2189 (Wm3iu6, Rn3iu6, L72iu6);  // ../RTL/cortexm0ds_logic.v(3942)
  buf u219 (Shhpw6[7], O1mpw6);  // ../RTL/cortexm0ds_logic.v(1941)
  and u2190 (Qz1iu6, Y93iu6, O8zhu6);  // ../RTL/cortexm0ds_logic.v(3943)
  not u2191 (L72iu6, Qz1iu6);  // ../RTL/cortexm0ds_logic.v(3943)
  and u2192 (Y93iu6, Yn3iu6, Fmyhu6);  // ../RTL/cortexm0ds_logic.v(3944)
  and u2193 (n312, Uthpw6[0], Vk1iu6);  // ../RTL/cortexm0ds_logic.v(3945)
  not u2194 (Rn3iu6, n312);  // ../RTL/cortexm0ds_logic.v(3945)
  and u2195 (Vk1iu6, Fo3iu6, Mo3iu6);  // ../RTL/cortexm0ds_logic.v(3946)
  or u2196 (n313, I83iu6, Yenhu6);  // ../RTL/cortexm0ds_logic.v(3947)
  not u2197 (Fo3iu6, n313);  // ../RTL/cortexm0ds_logic.v(3947)
  not u2198 (n6024, Romhu6);  // ../RTL/cortexm0ds_logic.v(3132)
  and u2199 (Im3iu6, To3iu6, Ap3iu6);  // ../RTL/cortexm0ds_logic.v(3949)
  not u22 (Zvdpw6, Qaipw6);  // ../RTL/cortexm0ds_logic.v(1778)
  buf u220 (Shhpw6[6], Q89bx6);  // ../RTL/cortexm0ds_logic.v(1941)
  and u2200 (n314, Tonhu6, Xl1iu6);  // ../RTL/cortexm0ds_logic.v(3950)
  not u2201 (Ap3iu6, n314);  // ../RTL/cortexm0ds_logic.v(3950)
  or u2202 (n315, Z4yhu6, Fmyhu6);  // ../RTL/cortexm0ds_logic.v(3951)
  not u2203 (Xl1iu6, n315);  // ../RTL/cortexm0ds_logic.v(3951)
  and u2204 (n316, Iahpw6[0], Z4yhu6);  // ../RTL/cortexm0ds_logic.v(3952)
  not u2205 (To3iu6, n316);  // ../RTL/cortexm0ds_logic.v(3952)
  AL_MUX u2206 (
    .i0(Tonhu6),
    .i1(Pinhu6),
    .sel(W13iu6),
    .o(Sqxhu6));  // ../RTL/cortexm0ds_logic.v(3953)
  and u2207 (n317, Hp3iu6, Op3iu6);  // ../RTL/cortexm0ds_logic.v(3954)
  not u2208 (W13iu6, n317);  // ../RTL/cortexm0ds_logic.v(3954)
  or u2209 (n318, Vp3iu6, Mdhpw6[1]);  // ../RTL/cortexm0ds_logic.v(3955)
  buf u221 (Shhpw6[5], T3opw6);  // ../RTL/cortexm0ds_logic.v(1941)
  not u2210 (Op3iu6, n318);  // ../RTL/cortexm0ds_logic.v(3955)
  and u2211 (Hp3iu6, Mdhpw6[2], Cq3iu6);  // ../RTL/cortexm0ds_logic.v(3956)
  AL_MUX u2212 (
    .i0(Iahpw6[29]),
    .i1(Zbhpw6[30]),
    .sel(Jq3iu6),
    .o(Lqxhu6));  // ../RTL/cortexm0ds_logic.v(3957)
  AL_MUX u2213 (
    .i0(Cjhpw6[1]),
    .i1(Mdhpw6[2]),
    .sel(Em1iu6),
    .o(Eqxhu6));  // ../RTL/cortexm0ds_logic.v(3958)
  AL_MUX u2214 (
    .i0(Cjhpw6[2]),
    .i1(Qq3iu6),
    .sel(Em1iu6),
    .o(Xpxhu6));  // ../RTL/cortexm0ds_logic.v(3959)
  and u2215 (Qq3iu6, N3nhu6, O43iu6);  // ../RTL/cortexm0ds_logic.v(3960)
  AL_MUX u2216 (
    .i0(Cjhpw6[0]),
    .i1(Mdhpw6[1]),
    .sel(Em1iu6),
    .o(Qpxhu6));  // ../RTL/cortexm0ds_logic.v(3961)
  AL_MUX u2217 (
    .i0(Shhpw6[1]),
    .i1(Iahpw6[0]),
    .sel(Em1iu6),
    .o(Jpxhu6));  // ../RTL/cortexm0ds_logic.v(3962)
  AL_MUX u2218 (
    .i0(Shhpw6[2]),
    .i1(Iahpw6[1]),
    .sel(Em1iu6),
    .o(Cpxhu6));  // ../RTL/cortexm0ds_logic.v(3963)
  AL_MUX u2219 (
    .i0(Shhpw6[3]),
    .i1(Iahpw6[2]),
    .sel(Em1iu6),
    .o(Voxhu6));  // ../RTL/cortexm0ds_logic.v(3964)
  buf u222 (vis_r12_o[19], Eitax6);  // ../RTL/cortexm0ds_logic.v(2599)
  AL_MUX u2220 (
    .i0(Shhpw6[4]),
    .i1(Iahpw6[3]),
    .sel(Em1iu6),
    .o(Ooxhu6));  // ../RTL/cortexm0ds_logic.v(3965)
  AL_MUX u2221 (
    .i0(Shhpw6[5]),
    .i1(Iahpw6[4]),
    .sel(Em1iu6),
    .o(Hoxhu6));  // ../RTL/cortexm0ds_logic.v(3966)
  AL_MUX u2222 (
    .i0(Shhpw6[6]),
    .i1(Iahpw6[5]),
    .sel(Em1iu6),
    .o(Aoxhu6));  // ../RTL/cortexm0ds_logic.v(3967)
  AL_MUX u2223 (
    .i0(Shhpw6[7]),
    .i1(Iahpw6[6]),
    .sel(Em1iu6),
    .o(Tnxhu6));  // ../RTL/cortexm0ds_logic.v(3968)
  AL_MUX u2224 (
    .i0(Shhpw6[8]),
    .i1(Iahpw6[7]),
    .sel(Em1iu6),
    .o(Mnxhu6));  // ../RTL/cortexm0ds_logic.v(3969)
  AL_MUX u2225 (
    .i0(Shhpw6[9]),
    .i1(Iahpw6[8]),
    .sel(Em1iu6),
    .o(Fnxhu6));  // ../RTL/cortexm0ds_logic.v(3970)
  AL_MUX u2226 (
    .i0(Shhpw6[10]),
    .i1(Iahpw6[9]),
    .sel(Em1iu6),
    .o(Ymxhu6));  // ../RTL/cortexm0ds_logic.v(3971)
  AL_MUX u2227 (
    .i0(Shhpw6[11]),
    .i1(Iahpw6[10]),
    .sel(Em1iu6),
    .o(Rmxhu6));  // ../RTL/cortexm0ds_logic.v(3972)
  AL_MUX u2228 (
    .i0(Shhpw6[12]),
    .i1(Iahpw6[11]),
    .sel(Em1iu6),
    .o(Kmxhu6));  // ../RTL/cortexm0ds_logic.v(3973)
  AL_MUX u2229 (
    .i0(Shhpw6[13]),
    .i1(Iahpw6[12]),
    .sel(Em1iu6),
    .o(Dmxhu6));  // ../RTL/cortexm0ds_logic.v(3974)
  buf u223 (vis_r12_o[17], Emtax6);  // ../RTL/cortexm0ds_logic.v(2599)
  AL_MUX u2230 (
    .i0(Shhpw6[14]),
    .i1(Iahpw6[13]),
    .sel(Em1iu6),
    .o(Wlxhu6));  // ../RTL/cortexm0ds_logic.v(3975)
  AL_MUX u2231 (
    .i0(Shhpw6[15]),
    .i1(Iahpw6[14]),
    .sel(Em1iu6),
    .o(Plxhu6));  // ../RTL/cortexm0ds_logic.v(3976)
  AL_MUX u2232 (
    .i0(Shhpw6[16]),
    .i1(Iahpw6[15]),
    .sel(Em1iu6),
    .o(Ilxhu6));  // ../RTL/cortexm0ds_logic.v(3977)
  AL_MUX u2233 (
    .i0(Shhpw6[17]),
    .i1(Iahpw6[16]),
    .sel(Em1iu6),
    .o(Blxhu6));  // ../RTL/cortexm0ds_logic.v(3978)
  AL_MUX u2234 (
    .i0(Shhpw6[18]),
    .i1(Iahpw6[17]),
    .sel(Em1iu6),
    .o(Ukxhu6));  // ../RTL/cortexm0ds_logic.v(3979)
  AL_MUX u2235 (
    .i0(Shhpw6[19]),
    .i1(Iahpw6[18]),
    .sel(Em1iu6),
    .o(Nkxhu6));  // ../RTL/cortexm0ds_logic.v(3980)
  AL_MUX u2236 (
    .i0(Shhpw6[20]),
    .i1(Iahpw6[19]),
    .sel(Em1iu6),
    .o(Gkxhu6));  // ../RTL/cortexm0ds_logic.v(3981)
  AL_MUX u2237 (
    .i0(Shhpw6[21]),
    .i1(Iahpw6[20]),
    .sel(Em1iu6),
    .o(Zjxhu6));  // ../RTL/cortexm0ds_logic.v(3982)
  AL_MUX u2238 (
    .i0(Shhpw6[22]),
    .i1(Iahpw6[21]),
    .sel(Em1iu6),
    .o(Sjxhu6));  // ../RTL/cortexm0ds_logic.v(3983)
  AL_MUX u2239 (
    .i0(Shhpw6[23]),
    .i1(Iahpw6[22]),
    .sel(Em1iu6),
    .o(Ljxhu6));  // ../RTL/cortexm0ds_logic.v(3984)
  buf u224 (vis_r12_o[16], Eotax6);  // ../RTL/cortexm0ds_logic.v(2599)
  AL_MUX u2240 (
    .i0(Shhpw6[24]),
    .i1(Iahpw6[23]),
    .sel(Em1iu6),
    .o(Ejxhu6));  // ../RTL/cortexm0ds_logic.v(3985)
  AL_MUX u2241 (
    .i0(Shhpw6[25]),
    .i1(Iahpw6[24]),
    .sel(Em1iu6),
    .o(Xixhu6));  // ../RTL/cortexm0ds_logic.v(3986)
  AL_MUX u2242 (
    .i0(Shhpw6[26]),
    .i1(Iahpw6[25]),
    .sel(Em1iu6),
    .o(Qixhu6));  // ../RTL/cortexm0ds_logic.v(3987)
  AL_MUX u2243 (
    .i0(Shhpw6[27]),
    .i1(Iahpw6[26]),
    .sel(Em1iu6),
    .o(Jixhu6));  // ../RTL/cortexm0ds_logic.v(3988)
  AL_MUX u2244 (
    .i0(Shhpw6[28]),
    .i1(Iahpw6[27]),
    .sel(Em1iu6),
    .o(Cixhu6));  // ../RTL/cortexm0ds_logic.v(3989)
  AL_MUX u2245 (
    .i0(Shhpw6[29]),
    .i1(Iahpw6[28]),
    .sel(Em1iu6),
    .o(Vhxhu6));  // ../RTL/cortexm0ds_logic.v(3990)
  AL_MUX u2246 (
    .i0(Shhpw6[30]),
    .i1(Iahpw6[29]),
    .sel(Em1iu6),
    .o(Ohxhu6));  // ../RTL/cortexm0ds_logic.v(3991)
  AL_MUX u2247 (
    .i0(Shhpw6[0]),
    .i1(Tonhu6),
    .sel(Em1iu6),
    .o(Hhxhu6));  // ../RTL/cortexm0ds_logic.v(3992)
  AL_MUX u2248 (
    .i0(Iqnhu6),
    .i1(Mdhpw6[0]),
    .sel(Em1iu6),
    .o(Ahxhu6));  // ../RTL/cortexm0ds_logic.v(3993)
  not u2249 (Em1iu6, C53iu6);  // ../RTL/cortexm0ds_logic.v(3994)
  buf u225 (vis_r12_o[14], Eqtax6);  // ../RTL/cortexm0ds_logic.v(2599)
  and u2250 (C53iu6, X53iu6, O43iu6);  // ../RTL/cortexm0ds_logic.v(3995)
  and u2251 (n319, Xq3iu6, G2ohu6);  // ../RTL/cortexm0ds_logic.v(3996)
  not u2252 (O43iu6, n319);  // ../RTL/cortexm0ds_logic.v(3996)
  and u2253 (Xq3iu6, Rrnhu6, A52iu6);  // ../RTL/cortexm0ds_logic.v(3997)
  or u2254 (X53iu6, Bh1iu6, Ng1iu6);  // ../RTL/cortexm0ds_logic.v(3998)
  and u2255 (n320, Er3iu6, Lr3iu6);  // ../RTL/cortexm0ds_logic.v(3999)
  not u2256 (Ng1iu6, n320);  // ../RTL/cortexm0ds_logic.v(3999)
  and u2257 (Lr3iu6, Sr3iu6, P13iu6);  // ../RTL/cortexm0ds_logic.v(4000)
  buf u2258 (Uhehu6, Ozkbx6[29]);  // ../RTL/cortexm0ds_logic.v(3176)
  and u2259 (Er3iu6, Ulnhu6, Fj1iu6);  // ../RTL/cortexm0ds_logic.v(4003)
  buf u226 (H2fpw6[2], Dzvpw6);  // ../RTL/cortexm0ds_logic.v(2444)
  and u2260 (Ug1iu6, Zr3iu6, Gs3iu6);  // ../RTL/cortexm0ds_logic.v(4004)
  not u2261 (Bh1iu6, Ug1iu6);  // ../RTL/cortexm0ds_logic.v(4004)
  buf u2262 (Ijehu6, Ozkbx6[28]);  // ../RTL/cortexm0ds_logic.v(3176)
  not u2263 (Gs3iu6, T42iu6);  // ../RTL/cortexm0ds_logic.v(4005)
  and u2264 (Zr3iu6, Zbhpw6[28], Gwnhu6);  // ../RTL/cortexm0ds_logic.v(4006)
  AL_MUX u2265 (
    .i0(Tonhu6),
    .i1(B7nhu6),
    .sel(Jq3iu6),
    .o(Tgxhu6));  // ../RTL/cortexm0ds_logic.v(4007)
  AL_MUX u2266 (
    .i0(Iahpw6[25]),
    .i1(Zbhpw6[26]),
    .sel(Jq3iu6),
    .o(Mgxhu6));  // ../RTL/cortexm0ds_logic.v(4008)
  AL_MUX u2267 (
    .i0(Iahpw6[27]),
    .i1(Zbhpw6[28]),
    .sel(Jq3iu6),
    .o(Fgxhu6));  // ../RTL/cortexm0ds_logic.v(4009)
  and u2268 (n321, Kn3iu6, Tezhu6);  // ../RTL/cortexm0ds_logic.v(4010)
  not u2269 (Jq3iu6, n321);  // ../RTL/cortexm0ds_logic.v(4010)
  buf u227 (vis_pc_o[0], Lerpw6);  // ../RTL/cortexm0ds_logic.v(2011)
  or u2270 (n322, O8zhu6, Pinhu6);  // ../RTL/cortexm0ds_logic.v(4011)
  not u2271 (Kn3iu6, n322);  // ../RTL/cortexm0ds_logic.v(4011)
  and u2272 (n323, Ns3iu6, Us3iu6);  // ../RTL/cortexm0ds_logic.v(4012)
  not u2273 (Yfxhu6, n323);  // ../RTL/cortexm0ds_logic.v(4012)
  and u2274 (n324, Zbhpw6[28], Bt3iu6);  // ../RTL/cortexm0ds_logic.v(4013)
  not u2275 (Us3iu6, n324);  // ../RTL/cortexm0ds_logic.v(4013)
  and u2276 (n325, Gwnhu6, A52iu6);  // ../RTL/cortexm0ds_logic.v(4014)
  not u2277 (Bt3iu6, n325);  // ../RTL/cortexm0ds_logic.v(4014)
  or u2278 (Ns3iu6, A52iu6, Gwnhu6);  // ../RTL/cortexm0ds_logic.v(4015)
  not u2279 (A52iu6, Punhu6);  // ../RTL/cortexm0ds_logic.v(4016)
  buf u228 (Shhpw6[11], Xx6bx6);  // ../RTL/cortexm0ds_logic.v(1941)
  and u2280 (n326, It3iu6, Pt3iu6);  // ../RTL/cortexm0ds_logic.v(4017)
  not u2281 (Rfxhu6, n326);  // ../RTL/cortexm0ds_logic.v(4017)
  and u2282 (n327, U5yhu6, Wt3iu6);  // ../RTL/cortexm0ds_logic.v(4018)
  not u2283 (Pt3iu6, n327);  // ../RTL/cortexm0ds_logic.v(4018)
  or u2284 (Wt3iu6, Du3iu6, Ku3iu6);  // ../RTL/cortexm0ds_logic.v(4019)
  and u2285 (Ku3iu6, Mmyhu6, Agyhu6);  // ../RTL/cortexm0ds_logic.v(4020)
  and u2286 (Mmyhu6, Ru3iu6, Xj3iu6);  // ../RTL/cortexm0ds_logic.v(4021)
  and u2287 (n328, Yu3iu6, Fv3iu6);  // ../RTL/cortexm0ds_logic.v(4022)
  not u2288 (Ru3iu6, n328);  // ../RTL/cortexm0ds_logic.v(4022)
  and u2289 (Fv3iu6, Mv3iu6, Tv3iu6);  // ../RTL/cortexm0ds_logic.v(4023)
  not u229 (Zehpw6[6], n7[6]);  // ../RTL/cortexm0ds_logic.v(3185)
  or u2290 (Tv3iu6, Aw3iu6, N73iu6);  // ../RTL/cortexm0ds_logic.v(4024)
  and u2291 (I83iu6, Hw3iu6, P5zhu6);  // ../RTL/cortexm0ds_logic.v(4025)
  not u2292 (N73iu6, I83iu6);  // ../RTL/cortexm0ds_logic.v(4025)
  not u2293 (P5zhu6, Ulnhu6);  // ../RTL/cortexm0ds_logic.v(4026)
  and u2294 (n329, Pyyhu6, Mdhpw6[0]);  // ../RTL/cortexm0ds_logic.v(4027)
  not u2295 (Hw3iu6, n329);  // ../RTL/cortexm0ds_logic.v(4027)
  or u2296 (n330, Qgzhu6, O8zhu6);  // ../RTL/cortexm0ds_logic.v(4028)
  not u2297 (Pyyhu6, n330);  // ../RTL/cortexm0ds_logic.v(4028)
  not u2298 (Qgzhu6, Mdhpw6[2]);  // ../RTL/cortexm0ds_logic.v(4029)
  and u2299 (Mv3iu6, Ow3iu6, P13iu6);  // ../RTL/cortexm0ds_logic.v(4030)
  buf u23 (Gqgpw6[28], Bngax6);  // ../RTL/cortexm0ds_logic.v(2377)
  buf u230 (H2fpw6[1], Wxjpw6);  // ../RTL/cortexm0ds_logic.v(2444)
  and u2300 (Yu3iu6, Rgnhu6, Z63iu6);  // ../RTL/cortexm0ds_logic.v(4032)
  AL_MUX u2301 (
    .i0(A1zhu6),
    .i1(Vw3iu6),
    .sel(Xj3iu6),
    .o(Du3iu6));  // ../RTL/cortexm0ds_logic.v(4033)
  and u2302 (Vw3iu6, T0zhu6, Rzyhu6);  // ../RTL/cortexm0ds_logic.v(4034)
  or u2303 (n331, Y7yhu6, Ighpw6[0]);  // ../RTL/cortexm0ds_logic.v(4035)
  not u2304 (A1zhu6, n331);  // ../RTL/cortexm0ds_logic.v(4035)
  AL_MUX u2305 (
    .i0(Cx3iu6),
    .i1(Jx3iu6),
    .sel(Hknhu6),
    .o(It3iu6));  // ../RTL/cortexm0ds_logic.v(4036)
  AL_MUX u2306 (
    .i0(Qx3iu6),
    .i1(Xx3iu6),
    .sel(Ey3iu6),
    .o(Jx3iu6));  // ../RTL/cortexm0ds_logic.v(4037)
  and u2307 (Qx3iu6, U5yhu6, Ly3iu6);  // ../RTL/cortexm0ds_logic.v(4038)
  and u2308 (n332, Sy3iu6, Zy3iu6);  // ../RTL/cortexm0ds_logic.v(4039)
  not u2309 (Ly3iu6, n332);  // ../RTL/cortexm0ds_logic.v(4039)
  not u231 (Zehpw6[5], n7[5]);  // ../RTL/cortexm0ds_logic.v(3185)
  and u2310 (Zy3iu6, Gz3iu6, Y7yhu6);  // ../RTL/cortexm0ds_logic.v(4040)
  and u2311 (n333, Nz3iu6, Ighpw6[2]);  // ../RTL/cortexm0ds_logic.v(4041)
  not u2312 (Y7yhu6, n333);  // ../RTL/cortexm0ds_logic.v(4041)
  or u2313 (n334, Wdyhu6, Ighpw6[1]);  // ../RTL/cortexm0ds_logic.v(4042)
  not u2314 (Nz3iu6, n334);  // ../RTL/cortexm0ds_logic.v(4042)
  or u2315 (n335, T0zhu6, Agyhu6);  // ../RTL/cortexm0ds_logic.v(4043)
  not u2316 (Gz3iu6, n335);  // ../RTL/cortexm0ds_logic.v(4043)
  and u2317 (T0zhu6, Gjyhu6, Vuyhu6);  // ../RTL/cortexm0ds_logic.v(4044)
  and u2318 (Sy3iu6, Uz3iu6, B04iu6);  // ../RTL/cortexm0ds_logic.v(4045)
  or u2319 (B04iu6, C9zhu6, Vmzhu6);  // ../RTL/cortexm0ds_logic.v(4046)
  not u232 (Zehpw6[4], n7[4]);  // ../RTL/cortexm0ds_logic.v(3185)
  and u2320 (Uz3iu6, I04iu6, Joyhu6);  // ../RTL/cortexm0ds_logic.v(4047)
  and u2321 (n336, P04iu6, Epyhu6);  // ../RTL/cortexm0ds_logic.v(4048)
  not u2322 (Joyhu6, n336);  // ../RTL/cortexm0ds_logic.v(4048)
  or u2323 (n337, Deyhu6, Ighpw6[2]);  // ../RTL/cortexm0ds_logic.v(4049)
  not u2324 (P04iu6, n337);  // ../RTL/cortexm0ds_logic.v(4049)
  buf u2325 (Wkehu6, Ozkbx6[27]);  // ../RTL/cortexm0ds_logic.v(3176)
  not u2326 (I04iu6, N03iu6);  // ../RTL/cortexm0ds_logic.v(4050)
  or u2327 (n338, C9zhu6, Wdyhu6);  // ../RTL/cortexm0ds_logic.v(4051)
  not u2328 (Gjyhu6, n338);  // ../RTL/cortexm0ds_logic.v(4051)
  not u2329 (C9zhu6, Cvyhu6);  // ../RTL/cortexm0ds_logic.v(4052)
  not u233 (Zehpw6[3], n7[3]);  // ../RTL/cortexm0ds_logic.v(3185)
  and u2330 (n339, Ey3iu6, Xx3iu6);  // ../RTL/cortexm0ds_logic.v(4053)
  not u2331 (Cx3iu6, n339);  // ../RTL/cortexm0ds_logic.v(4053)
  and u2332 (n340, W04iu6, D14iu6);  // ../RTL/cortexm0ds_logic.v(4054)
  not u2333 (Xx3iu6, n340);  // ../RTL/cortexm0ds_logic.v(4054)
  and u2334 (n341, K14iu6, Z4yhu6);  // ../RTL/cortexm0ds_logic.v(4055)
  not u2335 (D14iu6, n341);  // ../RTL/cortexm0ds_logic.v(4055)
  and u2336 (K14iu6, Mdhpw6[0], SWDO);  // ../RTL/cortexm0ds_logic.v(4056)
  and u2337 (n342, Mdhpw6[3], R14iu6);  // ../RTL/cortexm0ds_logic.v(4057)
  not u2338 (W04iu6, n342);  // ../RTL/cortexm0ds_logic.v(4057)
  or u2339 (R14iu6, L02iu6, R7yhu6);  // ../RTL/cortexm0ds_logic.v(4058)
  buf u234 (Shhpw6[17], Lhbbx6);  // ../RTL/cortexm0ds_logic.v(1941)
  not u2340 (R7yhu6, Mdhpw6[0]);  // ../RTL/cortexm0ds_logic.v(4059)
  not u2341 (L02iu6, Z4yhu6);  // ../RTL/cortexm0ds_logic.v(4060)
  or u2342 (Ey3iu6, Y14iu6, Z4yhu6);  // ../RTL/cortexm0ds_logic.v(4061)
  and u2343 (Z4yhu6, Ighpw6[5], Vx2iu6);  // ../RTL/cortexm0ds_logic.v(4062)
  AL_MUX u2344 (
    .i0(Aphpw6[1]),
    .i1(F24iu6),
    .sel(M24iu6),
    .o(Kfxhu6));  // ../RTL/cortexm0ds_logic.v(4063)
  and u2345 (F24iu6, T24iu6, A34iu6);  // ../RTL/cortexm0ds_logic.v(4064)
  AL_MUX u2346 (
    .i0(Cynhu6),
    .i1(H34iu6),
    .sel(M24iu6),
    .o(Dfxhu6));  // ../RTL/cortexm0ds_logic.v(4065)
  AL_MUX u2347 (
    .i0(Aphpw6[2]),
    .i1(O34iu6),
    .sel(M24iu6),
    .o(Wexhu6));  // ../RTL/cortexm0ds_logic.v(4066)
  and u2348 (M24iu6, V34iu6, C44iu6);  // ../RTL/cortexm0ds_logic.v(4067)
  AL_MUX u2349 (
    .i0(Jshpw6[10]),
    .i1(J44iu6),
    .sel(Sm1iu6),
    .o(Pexhu6));  // ../RTL/cortexm0ds_logic.v(4068)
  buf u235 (Shhpw6[15], Va7ax6);  // ../RTL/cortexm0ds_logic.v(1941)
  AL_MUX u2350 (
    .i0(Jshpw6[11]),
    .i1(Q44iu6),
    .sel(Sm1iu6),
    .o(Iexhu6));  // ../RTL/cortexm0ds_logic.v(4069)
  AL_MUX u2351 (
    .i0(Jshpw6[12]),
    .i1(X44iu6),
    .sel(Sm1iu6),
    .o(Bexhu6));  // ../RTL/cortexm0ds_logic.v(4070)
  AL_MUX u2352 (
    .i0(Jshpw6[13]),
    .i1(E54iu6),
    .sel(Sm1iu6),
    .o(Udxhu6));  // ../RTL/cortexm0ds_logic.v(4071)
  AL_MUX u2353 (
    .i0(Jshpw6[14]),
    .i1(L54iu6),
    .sel(Sm1iu6),
    .o(Ndxhu6));  // ../RTL/cortexm0ds_logic.v(4072)
  AL_MUX u2354 (
    .i0(Jshpw6[15]),
    .i1(S54iu6),
    .sel(Sm1iu6),
    .o(Gdxhu6));  // ../RTL/cortexm0ds_logic.v(4073)
  AL_MUX u2355 (
    .i0(Jshpw6[16]),
    .i1(Z54iu6),
    .sel(Sm1iu6),
    .o(Zcxhu6));  // ../RTL/cortexm0ds_logic.v(4074)
  AL_MUX u2356 (
    .i0(Jshpw6[17]),
    .i1(G64iu6),
    .sel(Sm1iu6),
    .o(Scxhu6));  // ../RTL/cortexm0ds_logic.v(4075)
  AL_MUX u2357 (
    .i0(Jshpw6[18]),
    .i1(N64iu6),
    .sel(Sm1iu6),
    .o(Lcxhu6));  // ../RTL/cortexm0ds_logic.v(4076)
  AL_MUX u2358 (
    .i0(Jshpw6[19]),
    .i1(U64iu6),
    .sel(Sm1iu6),
    .o(Ecxhu6));  // ../RTL/cortexm0ds_logic.v(4077)
  AL_MUX u2359 (
    .i0(Jshpw6[20]),
    .i1(B74iu6),
    .sel(Sm1iu6),
    .o(Xbxhu6));  // ../RTL/cortexm0ds_logic.v(4078)
  buf u236 (Shhpw6[14], Liabx6);  // ../RTL/cortexm0ds_logic.v(1941)
  AL_MUX u2360 (
    .i0(Jshpw6[21]),
    .i1(I74iu6),
    .sel(Sm1iu6),
    .o(Qbxhu6));  // ../RTL/cortexm0ds_logic.v(4079)
  AL_MUX u2361 (
    .i0(Jshpw6[22]),
    .i1(P74iu6),
    .sel(Sm1iu6),
    .o(Jbxhu6));  // ../RTL/cortexm0ds_logic.v(4080)
  AL_MUX u2362 (
    .i0(Jshpw6[23]),
    .i1(W74iu6),
    .sel(Sm1iu6),
    .o(Cbxhu6));  // ../RTL/cortexm0ds_logic.v(4081)
  AL_MUX u2363 (
    .i0(Jshpw6[24]),
    .i1(D84iu6),
    .sel(Sm1iu6),
    .o(Vaxhu6));  // ../RTL/cortexm0ds_logic.v(4082)
  AL_MUX u2364 (
    .i0(Jshpw6[25]),
    .i1(K84iu6),
    .sel(Sm1iu6),
    .o(Oaxhu6));  // ../RTL/cortexm0ds_logic.v(4083)
  AL_MUX u2365 (
    .i0(Jshpw6[26]),
    .i1(R84iu6),
    .sel(Sm1iu6),
    .o(Haxhu6));  // ../RTL/cortexm0ds_logic.v(4084)
  AL_MUX u2366 (
    .i0(Jshpw6[27]),
    .i1(Y84iu6),
    .sel(Sm1iu6),
    .o(Aaxhu6));  // ../RTL/cortexm0ds_logic.v(4085)
  AL_MUX u2367 (
    .i0(Jshpw6[28]),
    .i1(F94iu6),
    .sel(Sm1iu6),
    .o(T9xhu6));  // ../RTL/cortexm0ds_logic.v(4086)
  AL_MUX u2368 (
    .i0(Jshpw6[29]),
    .i1(M94iu6),
    .sel(Sm1iu6),
    .o(M9xhu6));  // ../RTL/cortexm0ds_logic.v(4087)
  AL_MUX u2369 (
    .i0(Jshpw6[30]),
    .i1(T94iu6),
    .sel(Sm1iu6),
    .o(F9xhu6));  // ../RTL/cortexm0ds_logic.v(4088)
  buf u237 (Shhpw6[12], Ns8ax6);  // ../RTL/cortexm0ds_logic.v(1941)
  and u2370 (n343, Aa4iu6, Ha4iu6);  // ../RTL/cortexm0ds_logic.v(4089)
  not u2371 (Y8xhu6, n343);  // ../RTL/cortexm0ds_logic.v(4089)
  and u2372 (n344, Gmhpw6[0], Oa4iu6);  // ../RTL/cortexm0ds_logic.v(4090)
  not u2373 (Ha4iu6, n344);  // ../RTL/cortexm0ds_logic.v(4090)
  and u2374 (Aa4iu6, Va4iu6, Cb4iu6);  // ../RTL/cortexm0ds_logic.v(4091)
  and u2375 (n345, T24iu6, Sm1iu6);  // ../RTL/cortexm0ds_logic.v(4092)
  not u2376 (Cb4iu6, n345);  // ../RTL/cortexm0ds_logic.v(4092)
  and u2377 (n346, Tnhpw6[0], Jb4iu6);  // ../RTL/cortexm0ds_logic.v(4093)
  not u2378 (Va4iu6, n346);  // ../RTL/cortexm0ds_logic.v(4093)
  and u2379 (n347, Qb4iu6, Xb4iu6);  // ../RTL/cortexm0ds_logic.v(4094)
  buf u238 (Shhpw6[16], Ymwpw6);  // ../RTL/cortexm0ds_logic.v(1941)
  not u2380 (R8xhu6, n347);  // ../RTL/cortexm0ds_logic.v(4094)
  and u2381 (n348, Gmhpw6[1], Oa4iu6);  // ../RTL/cortexm0ds_logic.v(4095)
  not u2382 (Xb4iu6, n348);  // ../RTL/cortexm0ds_logic.v(4095)
  and u2383 (Qb4iu6, Ec4iu6, Lc4iu6);  // ../RTL/cortexm0ds_logic.v(4096)
  and u2384 (n349, Sm1iu6, O34iu6);  // ../RTL/cortexm0ds_logic.v(4097)
  not u2385 (Lc4iu6, n349);  // ../RTL/cortexm0ds_logic.v(4097)
  and u2386 (n350, Tnhpw6[1], Jb4iu6);  // ../RTL/cortexm0ds_logic.v(4098)
  not u2387 (Ec4iu6, n350);  // ../RTL/cortexm0ds_logic.v(4098)
  and u2388 (n351, Sc4iu6, Zc4iu6);  // ../RTL/cortexm0ds_logic.v(4099)
  not u2389 (K8xhu6, n351);  // ../RTL/cortexm0ds_logic.v(4099)
  buf u239 (Shhpw6[20], Ahdbx6);  // ../RTL/cortexm0ds_logic.v(1941)
  and u2390 (n352, Gmhpw6[2], Oa4iu6);  // ../RTL/cortexm0ds_logic.v(4100)
  not u2391 (Zc4iu6, n352);  // ../RTL/cortexm0ds_logic.v(4100)
  and u2392 (Sc4iu6, Gd4iu6, Nd4iu6);  // ../RTL/cortexm0ds_logic.v(4101)
  and u2393 (n353, Ud4iu6, Sm1iu6);  // ../RTL/cortexm0ds_logic.v(4102)
  not u2394 (Nd4iu6, n353);  // ../RTL/cortexm0ds_logic.v(4102)
  and u2395 (n354, Tnhpw6[2], Jb4iu6);  // ../RTL/cortexm0ds_logic.v(4103)
  not u2396 (Gd4iu6, n354);  // ../RTL/cortexm0ds_logic.v(4103)
  and u2397 (n355, Be4iu6, Ie4iu6);  // ../RTL/cortexm0ds_logic.v(4104)
  not u2398 (D8xhu6, n355);  // ../RTL/cortexm0ds_logic.v(4104)
  and u2399 (n356, Gmhpw6[3], Oa4iu6);  // ../RTL/cortexm0ds_logic.v(4105)
  buf u24 (Uthpw6[21], Jhebx6);  // ../RTL/cortexm0ds_logic.v(1882)
  buf u240 (Shhpw6[21], H0ebx6);  // ../RTL/cortexm0ds_logic.v(1941)
  not u2400 (Ie4iu6, n356);  // ../RTL/cortexm0ds_logic.v(4105)
  and u2401 (Be4iu6, Pe4iu6, We4iu6);  // ../RTL/cortexm0ds_logic.v(4106)
  and u2402 (n357, Df4iu6, Sm1iu6);  // ../RTL/cortexm0ds_logic.v(4107)
  not u2403 (We4iu6, n357);  // ../RTL/cortexm0ds_logic.v(4107)
  and u2404 (n358, Tnhpw6[3], Jb4iu6);  // ../RTL/cortexm0ds_logic.v(4108)
  not u2405 (Pe4iu6, n358);  // ../RTL/cortexm0ds_logic.v(4108)
  and u2406 (n359, Kf4iu6, Rf4iu6);  // ../RTL/cortexm0ds_logic.v(4109)
  not u2407 (W7xhu6, n359);  // ../RTL/cortexm0ds_logic.v(4109)
  and u2408 (n360, Gmhpw6[4], Oa4iu6);  // ../RTL/cortexm0ds_logic.v(4110)
  not u2409 (Rf4iu6, n360);  // ../RTL/cortexm0ds_logic.v(4110)
  buf u241 (Shhpw6[22], Ojebx6);  // ../RTL/cortexm0ds_logic.v(1941)
  and u2410 (Kf4iu6, Yf4iu6, Fg4iu6);  // ../RTL/cortexm0ds_logic.v(4111)
  and u2411 (n361, H34iu6, Sm1iu6);  // ../RTL/cortexm0ds_logic.v(4112)
  not u2412 (Fg4iu6, n361);  // ../RTL/cortexm0ds_logic.v(4112)
  and u2413 (n362, Jshpw6[4], Jb4iu6);  // ../RTL/cortexm0ds_logic.v(4113)
  not u2414 (Yf4iu6, n362);  // ../RTL/cortexm0ds_logic.v(4113)
  and u2415 (n363, Mg4iu6, Tg4iu6);  // ../RTL/cortexm0ds_logic.v(4114)
  not u2416 (P7xhu6, n363);  // ../RTL/cortexm0ds_logic.v(4114)
  and u2417 (n364, Gmhpw6[5], Oa4iu6);  // ../RTL/cortexm0ds_logic.v(4115)
  not u2418 (Tg4iu6, n364);  // ../RTL/cortexm0ds_logic.v(4115)
  and u2419 (Mg4iu6, Ah4iu6, Hh4iu6);  // ../RTL/cortexm0ds_logic.v(4116)
  buf u242 (Shhpw6[23], Urgbx6);  // ../RTL/cortexm0ds_logic.v(1941)
  and u2420 (n365, Oh4iu6, Sm1iu6);  // ../RTL/cortexm0ds_logic.v(4117)
  not u2421 (Hh4iu6, n365);  // ../RTL/cortexm0ds_logic.v(4117)
  and u2422 (n366, Jshpw6[5], Jb4iu6);  // ../RTL/cortexm0ds_logic.v(4118)
  not u2423 (Ah4iu6, n366);  // ../RTL/cortexm0ds_logic.v(4118)
  and u2424 (n367, Vh4iu6, Ci4iu6);  // ../RTL/cortexm0ds_logic.v(4119)
  not u2425 (I7xhu6, n367);  // ../RTL/cortexm0ds_logic.v(4119)
  and u2426 (n368, Gmhpw6[6], Oa4iu6);  // ../RTL/cortexm0ds_logic.v(4120)
  not u2427 (Ci4iu6, n368);  // ../RTL/cortexm0ds_logic.v(4120)
  and u2428 (Vh4iu6, Ji4iu6, Qi4iu6);  // ../RTL/cortexm0ds_logic.v(4121)
  and u2429 (n369, Xi4iu6, Sm1iu6);  // ../RTL/cortexm0ds_logic.v(4122)
  buf u243 (Shhpw6[24], Jvkpw6);  // ../RTL/cortexm0ds_logic.v(1941)
  not u2430 (Qi4iu6, n369);  // ../RTL/cortexm0ds_logic.v(4122)
  and u2431 (n370, Jshpw6[6], Jb4iu6);  // ../RTL/cortexm0ds_logic.v(4123)
  not u2432 (Ji4iu6, n370);  // ../RTL/cortexm0ds_logic.v(4123)
  and u2433 (n371, Ej4iu6, Lj4iu6);  // ../RTL/cortexm0ds_logic.v(4124)
  not u2434 (B7xhu6, n371);  // ../RTL/cortexm0ds_logic.v(4124)
  and u2435 (n372, Gmhpw6[7], Oa4iu6);  // ../RTL/cortexm0ds_logic.v(4125)
  not u2436 (Lj4iu6, n372);  // ../RTL/cortexm0ds_logic.v(4125)
  and u2437 (Ej4iu6, Sj4iu6, Zj4iu6);  // ../RTL/cortexm0ds_logic.v(4126)
  and u2438 (n373, Gk4iu6, Sm1iu6);  // ../RTL/cortexm0ds_logic.v(4127)
  not u2439 (Zj4iu6, n373);  // ../RTL/cortexm0ds_logic.v(4127)
  buf u244 (Shhpw6[25], Bp2qw6);  // ../RTL/cortexm0ds_logic.v(1941)
  and u2440 (n374, Jshpw6[7], Jb4iu6);  // ../RTL/cortexm0ds_logic.v(4128)
  not u2441 (Sj4iu6, n374);  // ../RTL/cortexm0ds_logic.v(4128)
  and u2442 (n375, Nk4iu6, Uk4iu6);  // ../RTL/cortexm0ds_logic.v(4129)
  not u2443 (U6xhu6, n375);  // ../RTL/cortexm0ds_logic.v(4129)
  and u2444 (n376, Gmhpw6[8], Oa4iu6);  // ../RTL/cortexm0ds_logic.v(4130)
  not u2445 (Uk4iu6, n376);  // ../RTL/cortexm0ds_logic.v(4130)
  and u2446 (Nk4iu6, Bl4iu6, Il4iu6);  // ../RTL/cortexm0ds_logic.v(4131)
  and u2447 (n377, Sm1iu6, Pl4iu6);  // ../RTL/cortexm0ds_logic.v(4132)
  not u2448 (Il4iu6, n377);  // ../RTL/cortexm0ds_logic.v(4132)
  and u2449 (n378, Jshpw6[8], Jb4iu6);  // ../RTL/cortexm0ds_logic.v(4133)
  buf u245 (Shhpw6[28], D2rpw6);  // ../RTL/cortexm0ds_logic.v(1941)
  not u2450 (Bl4iu6, n378);  // ../RTL/cortexm0ds_logic.v(4133)
  and u2451 (n379, Wl4iu6, Dm4iu6);  // ../RTL/cortexm0ds_logic.v(4134)
  not u2452 (N6xhu6, n379);  // ../RTL/cortexm0ds_logic.v(4134)
  and u2453 (n380, Gmhpw6[9], Oa4iu6);  // ../RTL/cortexm0ds_logic.v(4135)
  not u2454 (Dm4iu6, n380);  // ../RTL/cortexm0ds_logic.v(4135)
  and u2455 (Wl4iu6, Km4iu6, Rm4iu6);  // ../RTL/cortexm0ds_logic.v(4136)
  and u2456 (n381, Sm1iu6, Ym4iu6);  // ../RTL/cortexm0ds_logic.v(4137)
  not u2457 (Rm4iu6, n381);  // ../RTL/cortexm0ds_logic.v(4137)
  or u2458 (n382, Jb4iu6, Oa4iu6);  // ../RTL/cortexm0ds_logic.v(4138)
  not u2459 (Sm1iu6, n382);  // ../RTL/cortexm0ds_logic.v(4138)
  buf u246 (Shhpw6[29], Nv3qw6);  // ../RTL/cortexm0ds_logic.v(1941)
  and u2460 (n383, Jshpw6[9], Jb4iu6);  // ../RTL/cortexm0ds_logic.v(4139)
  not u2461 (Km4iu6, n383);  // ../RTL/cortexm0ds_logic.v(4139)
  or u2462 (n384, Fn4iu6, Oa4iu6);  // ../RTL/cortexm0ds_logic.v(4140)
  not u2463 (Jb4iu6, n384);  // ../RTL/cortexm0ds_logic.v(4140)
  and u2464 (Oa4iu6, Mn4iu6, Tn4iu6);  // ../RTL/cortexm0ds_logic.v(4141)
  and u2465 (Tn4iu6, Ao4iu6, Pqzhu6);  // ../RTL/cortexm0ds_logic.v(4142)
  or u2466 (n385, Lf1iu6, Ho4iu6);  // ../RTL/cortexm0ds_logic.v(4143)
  not u2467 (Ao4iu6, n385);  // ../RTL/cortexm0ds_logic.v(4143)
  and u2468 (Lf1iu6, HRESP, R0nhu6);  // ../RTL/cortexm0ds_logic.v(4144)
  and u2469 (Mn4iu6, Cynhu6, Tszhu6);  // ../RTL/cortexm0ds_logic.v(4145)
  buf u247 (Shhpw6[31], Yzqpw6);  // ../RTL/cortexm0ds_logic.v(1941)
  and u2470 (Tszhu6, Oo4iu6, Sqhpw6[1]);  // ../RTL/cortexm0ds_logic.v(4146)
  or u2471 (n386, Fszhu6, Sqhpw6[0]);  // ../RTL/cortexm0ds_logic.v(4147)
  not u2472 (Oo4iu6, n386);  // ../RTL/cortexm0ds_logic.v(4147)
  and u2473 (Fn4iu6, V34iu6, Vo4iu6);  // ../RTL/cortexm0ds_logic.v(4148)
  and u2474 (V34iu6, Cp4iu6, Jp4iu6);  // ../RTL/cortexm0ds_logic.v(4149)
  and u2475 (Jp4iu6, Qp4iu6, Xp4iu6);  // ../RTL/cortexm0ds_logic.v(4150)
  or u2476 (n387, Ho4iu6, Eq4iu6);  // ../RTL/cortexm0ds_logic.v(4151)
  not u2477 (Qp4iu6, n387);  // ../RTL/cortexm0ds_logic.v(4151)
  and u2478 (Cp4iu6, Lq4iu6, Sqhpw6[1]);  // ../RTL/cortexm0ds_logic.v(4152)
  or u2479 (n388, Gpzhu6, Sq4iu6);  // ../RTL/cortexm0ds_logic.v(4153)
  not u248 (Zehpw6[2], n7[2]);  // ../RTL/cortexm0ds_logic.v(3185)
  not u2480 (Lq4iu6, n388);  // ../RTL/cortexm0ds_logic.v(4153)
  not u2481 (G6xhu6, Zq4iu6);  // ../RTL/cortexm0ds_logic.v(4154)
  AL_MUX u2482 (
    .i0(Gr4iu6),
    .i1(Sq4iu6),
    .sel(Nr4iu6),
    .o(Zq4iu6));  // ../RTL/cortexm0ds_logic.v(4155)
  and u2483 (n389, A2nhu6, Ur4iu6);  // ../RTL/cortexm0ds_logic.v(4156)
  not u2484 (Gr4iu6, n389);  // ../RTL/cortexm0ds_logic.v(4156)
  AL_MUX u2485 (
    .i0(T24iu6),
    .i1(Lwgpw6[0]),
    .sel(Bs4iu6),
    .o(Z5xhu6));  // ../RTL/cortexm0ds_logic.v(4157)
  AL_MUX u2486 (
    .i0(Ud4iu6),
    .i1(Lwgpw6[2]),
    .sel(Bs4iu6),
    .o(S5xhu6));  // ../RTL/cortexm0ds_logic.v(4158)
  AL_MUX u2487 (
    .i0(O34iu6),
    .i1(Lwgpw6[1]),
    .sel(Bs4iu6),
    .o(L5xhu6));  // ../RTL/cortexm0ds_logic.v(4159)
  or u2488 (Bs4iu6, Is4iu6, Ps4iu6);  // ../RTL/cortexm0ds_logic.v(4160)
  AL_MUX u2489 (
    .i0(Vchhu6),
    .i1(Dt4iu6),
    .sel(Kt4iu6),
    .o(E5xhu6));  // ../RTL/cortexm0ds_logic.v(4162)
  buf u249 (Uthpw6[12], Ro8ax6);  // ../RTL/cortexm0ds_logic.v(1882)
  and u2490 (Kt4iu6, HREADY, Rt4iu6);  // ../RTL/cortexm0ds_logic.v(4163)
  and u2491 (n390, Yt4iu6, Fu4iu6);  // ../RTL/cortexm0ds_logic.v(4164)
  not u2492 (Rt4iu6, n390);  // ../RTL/cortexm0ds_logic.v(4164)
  or u2493 (n391, Mu4iu6, Tu4iu6);  // ../RTL/cortexm0ds_logic.v(4165)
  not u2494 (Fu4iu6, n391);  // ../RTL/cortexm0ds_logic.v(4165)
  or u2495 (n392, Dt4iu6, Av4iu6);  // ../RTL/cortexm0ds_logic.v(4166)
  not u2496 (Yt4iu6, n392);  // ../RTL/cortexm0ds_logic.v(4166)
  or u2497 (n393, K7vpw6, DBGRESTART);  // ../RTL/cortexm0ds_logic.v(4167)
  not u2498 (Av4iu6, n393);  // ../RTL/cortexm0ds_logic.v(4167)
  and u2499 (n394, Ov4iu6, Vv4iu6);  // ../RTL/cortexm0ds_logic.v(4168)
  buf u25 (K7hpw6[16], Ue9ax6);  // ../RTL/cortexm0ds_logic.v(2366)
  buf u250 (G4hpw6[2], T7bax6);  // ../RTL/cortexm0ds_logic.v(2274)
  not u2500 (Dt4iu6, n394);  // ../RTL/cortexm0ds_logic.v(4168)
  and u2501 (Vv4iu6, Cw4iu6, Jw4iu6);  // ../RTL/cortexm0ds_logic.v(4169)
  and u2502 (Cw4iu6, Qw4iu6, Xw4iu6);  // ../RTL/cortexm0ds_logic.v(4170)
  or u2503 (n395, Ex4iu6, Lx4iu6);  // ../RTL/cortexm0ds_logic.v(4171)
  not u2504 (Ov4iu6, n395);  // ../RTL/cortexm0ds_logic.v(4171)
  and u2505 (n396, Sx4iu6, Zx4iu6);  // ../RTL/cortexm0ds_logic.v(4172)
  not u2506 (X4xhu6, n396);  // ../RTL/cortexm0ds_logic.v(4172)
  and u2507 (Zx4iu6, Gy4iu6, Ny4iu6);  // ../RTL/cortexm0ds_logic.v(4173)
  and u2508 (n397, Hrfpw6[16], Uy4iu6);  // ../RTL/cortexm0ds_logic.v(4174)
  not u2509 (Ny4iu6, n397);  // ../RTL/cortexm0ds_logic.v(4174)
  buf u251 (Shhpw6[4], P93qw6);  // ../RTL/cortexm0ds_logic.v(1941)
  and u2510 (Gy4iu6, Bz4iu6, Iz4iu6);  // ../RTL/cortexm0ds_logic.v(4175)
  and u2511 (n398, Pz4iu6, Wz4iu6);  // ../RTL/cortexm0ds_logic.v(4176)
  not u2512 (Bz4iu6, n398);  // ../RTL/cortexm0ds_logic.v(4176)
  and u2513 (Sx4iu6, D05iu6, K05iu6);  // ../RTL/cortexm0ds_logic.v(4177)
  and u2514 (n399, R05iu6, S1ehu6);  // ../RTL/cortexm0ds_logic.v(4178)
  not u2515 (K05iu6, n399);  // ../RTL/cortexm0ds_logic.v(4178)
  and u2516 (D05iu6, Y05iu6, F15iu6);  // ../RTL/cortexm0ds_logic.v(4179)
  and u2517 (n400, M15iu6, T15iu6);  // ../RTL/cortexm0ds_logic.v(4180)
  not u2518 (F15iu6, n400);  // ../RTL/cortexm0ds_logic.v(4180)
  and u2519 (n401, Ppfpw6[16], A25iu6);  // ../RTL/cortexm0ds_logic.v(4181)
  buf u252 (vis_psp_o[9], Yt8bx6);  // ../RTL/cortexm0ds_logic.v(2085)
  not u2520 (Y05iu6, n401);  // ../RTL/cortexm0ds_logic.v(4181)
  AL_MUX u2521 (
    .i0(H25iu6),
    .i1(X3fpw6[1]),
    .sel(O25iu6),
    .o(Q4xhu6));  // ../RTL/cortexm0ds_logic.v(4182)
  and u2522 (n402, V25iu6, C35iu6);  // ../RTL/cortexm0ds_logic.v(4183)
  not u2523 (H25iu6, n402);  // ../RTL/cortexm0ds_logic.v(4183)
  and u2524 (C35iu6, J35iu6, Q35iu6);  // ../RTL/cortexm0ds_logic.v(4184)
  and u2525 (Q35iu6, X35iu6, E45iu6);  // ../RTL/cortexm0ds_logic.v(4185)
  and u2526 (n403, L45iu6, S45iu6);  // ../RTL/cortexm0ds_logic.v(4186)
  not u2527 (X35iu6, n403);  // ../RTL/cortexm0ds_logic.v(4186)
  and u2528 (n404, Z45iu6, G55iu6);  // ../RTL/cortexm0ds_logic.v(4187)
  not u2529 (S45iu6, n404);  // ../RTL/cortexm0ds_logic.v(4187)
  buf u253 (vis_r4_o[15], Z78bx6);  // ../RTL/cortexm0ds_logic.v(2626)
  AL_MUX u2530 (
    .i0(N55iu6),
    .i1(U55iu6),
    .sel(B65iu6),
    .o(Z45iu6));  // ../RTL/cortexm0ds_logic.v(4188)
  and u2531 (n405, I65iu6, P65iu6);  // ../RTL/cortexm0ds_logic.v(4189)
  not u2532 (U55iu6, n405);  // ../RTL/cortexm0ds_logic.v(4189)
  and u2533 (J35iu6, W65iu6, D75iu6);  // ../RTL/cortexm0ds_logic.v(4190)
  and u2534 (n406, D7fpw6[4], K75iu6);  // ../RTL/cortexm0ds_logic.v(4191)
  not u2535 (D75iu6, n406);  // ../RTL/cortexm0ds_logic.v(4191)
  or u2536 (W65iu6, R75iu6, P65iu6);  // ../RTL/cortexm0ds_logic.v(4192)
  and u2537 (V25iu6, Y75iu6, F85iu6);  // ../RTL/cortexm0ds_logic.v(4193)
  and u2538 (Y75iu6, M85iu6, T85iu6);  // ../RTL/cortexm0ds_logic.v(4194)
  and u2539 (n407, A95iu6, D7fpw6[1]);  // ../RTL/cortexm0ds_logic.v(4195)
  buf u254 (vis_r14_o[12], N5oax6);  // ../RTL/cortexm0ds_logic.v(2497)
  not u2540 (T85iu6, n407);  // ../RTL/cortexm0ds_logic.v(4195)
  or u2541 (M85iu6, H95iu6, O95iu6);  // ../RTL/cortexm0ds_logic.v(4196)
  AL_MUX u2542 (
    .i0(V95iu6),
    .i1(Ca5iu6),
    .sel(Fsdhu6),
    .o(J4xhu6));  // ../RTL/cortexm0ds_logic.v(4197)
  and u2543 (n408, Ja5iu6, Qa5iu6);  // ../RTL/cortexm0ds_logic.v(4198)
  not u2544 (Ca5iu6, n408);  // ../RTL/cortexm0ds_logic.v(4198)
  and u2545 (n409, Xa5iu6, Eb5iu6);  // ../RTL/cortexm0ds_logic.v(4199)
  not u2546 (V95iu6, n409);  // ../RTL/cortexm0ds_logic.v(4199)
  and u2547 (Eb5iu6, Lb5iu6, Sb5iu6);  // ../RTL/cortexm0ds_logic.v(4200)
  or u2548 (n410, RXEV, TXEV);  // ../RTL/cortexm0ds_logic.v(4201)
  not u2549 (Lb5iu6, n410);  // ../RTL/cortexm0ds_logic.v(4201)
  buf u255 (vis_r8_o[21], Ourax6);  // ../RTL/cortexm0ds_logic.v(2579)
  and u2550 (Xa5iu6, Zb5iu6, Gc5iu6);  // ../RTL/cortexm0ds_logic.v(4202)
  and u2551 (Zb5iu6, Nc5iu6, Uc5iu6);  // ../RTL/cortexm0ds_logic.v(4203)
  and u2552 (n411, Gfghu6, Bd5iu6);  // ../RTL/cortexm0ds_logic.v(4204)
  not u2553 (Nc5iu6, n411);  // ../RTL/cortexm0ds_logic.v(4204)
  and u2554 (n412, Id5iu6, Pd5iu6);  // ../RTL/cortexm0ds_logic.v(4205)
  not u2555 (Bd5iu6, n412);  // ../RTL/cortexm0ds_logic.v(4205)
  and u2556 (Pd5iu6, Wd5iu6, De5iu6);  // ../RTL/cortexm0ds_logic.v(4206)
  and u2557 (De5iu6, Ke5iu6, Re5iu6);  // ../RTL/cortexm0ds_logic.v(4207)
  and u2558 (Re5iu6, Ye5iu6, Ff5iu6);  // ../RTL/cortexm0ds_logic.v(4208)
  and u2559 (Ff5iu6, Mf5iu6, Tf5iu6);  // ../RTL/cortexm0ds_logic.v(4209)
  buf u256 (Vbgpw6[15], Hf0bx6);  // ../RTL/cortexm0ds_logic.v(3092)
  or u2560 (Tf5iu6, Ag5iu6, Yyghu6);  // ../RTL/cortexm0ds_logic.v(4210)
  and u2561 (Mf5iu6, Hg5iu6, Og5iu6);  // ../RTL/cortexm0ds_logic.v(4211)
  and u2562 (n413, Vg5iu6, Ch5iu6);  // ../RTL/cortexm0ds_logic.v(4212)
  not u2563 (Og5iu6, n413);  // ../RTL/cortexm0ds_logic.v(4212)
  and u2564 (Vg5iu6, HWDATA[28], Jh5iu6);  // ../RTL/cortexm0ds_logic.v(4213)
  or u2565 (Hg5iu6, Qh5iu6, Zlghu6);  // ../RTL/cortexm0ds_logic.v(4214)
  and u2566 (Ye5iu6, Xh5iu6, Ei5iu6);  // ../RTL/cortexm0ds_logic.v(4215)
  or u2567 (Ei5iu6, Li5iu6, Righu6);  // ../RTL/cortexm0ds_logic.v(4216)
  and u2568 (n414, Cyohu6, Si5iu6);  // ../RTL/cortexm0ds_logic.v(4217)
  not u2569 (Xh5iu6, n414);  // ../RTL/cortexm0ds_logic.v(4217)
  buf u257 (Vbgpw6[14], Gd0bx6);  // ../RTL/cortexm0ds_logic.v(3092)
  not u2570 (Si5iu6, Odgpw6[31]);  // ../RTL/cortexm0ds_logic.v(4218)
  and u2571 (Ke5iu6, Zi5iu6, Gj5iu6);  // ../RTL/cortexm0ds_logic.v(4219)
  and u2572 (Gj5iu6, Nj5iu6, Uj5iu6);  // ../RTL/cortexm0ds_logic.v(4220)
  and u2573 (n415, Xyohu6, Bk5iu6);  // ../RTL/cortexm0ds_logic.v(4221)
  not u2574 (Uj5iu6, n415);  // ../RTL/cortexm0ds_logic.v(4221)
  not u2575 (Bk5iu6, Odgpw6[28]);  // ../RTL/cortexm0ds_logic.v(4222)
  and u2576 (Nj5iu6, Ik5iu6, Pk5iu6);  // ../RTL/cortexm0ds_logic.v(4223)
  and u2577 (n416, Jyohu6, Wk5iu6);  // ../RTL/cortexm0ds_logic.v(4224)
  not u2578 (Pk5iu6, n416);  // ../RTL/cortexm0ds_logic.v(4224)
  not u2579 (Wk5iu6, Odgpw6[30]);  // ../RTL/cortexm0ds_logic.v(4225)
  buf u258 (vis_r4_o[14], V7vax6);  // ../RTL/cortexm0ds_logic.v(2626)
  and u2580 (n417, Qyohu6, Dl5iu6);  // ../RTL/cortexm0ds_logic.v(4226)
  not u2581 (Ik5iu6, n417);  // ../RTL/cortexm0ds_logic.v(4226)
  not u2582 (Dl5iu6, Odgpw6[29]);  // ../RTL/cortexm0ds_logic.v(4227)
  and u2583 (Zi5iu6, Kl5iu6, Rl5iu6);  // ../RTL/cortexm0ds_logic.v(4228)
  and u2584 (n418, Ezohu6, Yl5iu6);  // ../RTL/cortexm0ds_logic.v(4229)
  not u2585 (Rl5iu6, n418);  // ../RTL/cortexm0ds_logic.v(4229)
  not u2586 (Yl5iu6, Odgpw6[27]);  // ../RTL/cortexm0ds_logic.v(4230)
  and u2587 (n419, Lzohu6, Fm5iu6);  // ../RTL/cortexm0ds_logic.v(4231)
  not u2588 (Kl5iu6, n419);  // ../RTL/cortexm0ds_logic.v(4231)
  not u2589 (Fm5iu6, Odgpw6[26]);  // ../RTL/cortexm0ds_logic.v(4232)
  buf u259 (vis_r14_o[11], Zp8bx6);  // ../RTL/cortexm0ds_logic.v(2497)
  and u2590 (Wd5iu6, Mm5iu6, Tm5iu6);  // ../RTL/cortexm0ds_logic.v(4233)
  and u2591 (Tm5iu6, An5iu6, Hn5iu6);  // ../RTL/cortexm0ds_logic.v(4234)
  and u2592 (Hn5iu6, On5iu6, Vn5iu6);  // ../RTL/cortexm0ds_logic.v(4235)
  and u2593 (n420, G0phu6, Co5iu6);  // ../RTL/cortexm0ds_logic.v(4236)
  not u2594 (Vn5iu6, n420);  // ../RTL/cortexm0ds_logic.v(4236)
  not u2595 (Co5iu6, Odgpw6[21]);  // ../RTL/cortexm0ds_logic.v(4237)
  and u2596 (On5iu6, Jo5iu6, Qo5iu6);  // ../RTL/cortexm0ds_logic.v(4238)
  and u2597 (n421, Szohu6, Xo5iu6);  // ../RTL/cortexm0ds_logic.v(4239)
  not u2598 (Qo5iu6, n421);  // ../RTL/cortexm0ds_logic.v(4239)
  not u2599 (Xo5iu6, Odgpw6[23]);  // ../RTL/cortexm0ds_logic.v(4240)
  buf u26 (vis_r2_o[27], Viqax6);  // ../RTL/cortexm0ds_logic.v(2551)
  buf u260 (vis_r8_o[20], Owrax6);  // ../RTL/cortexm0ds_logic.v(2579)
  and u2600 (n422, Zzohu6, Ep5iu6);  // ../RTL/cortexm0ds_logic.v(4241)
  not u2601 (Jo5iu6, n422);  // ../RTL/cortexm0ds_logic.v(4241)
  not u2602 (Ep5iu6, Odgpw6[22]);  // ../RTL/cortexm0ds_logic.v(4242)
  and u2603 (An5iu6, Lp5iu6, Sp5iu6);  // ../RTL/cortexm0ds_logic.v(4243)
  and u2604 (n423, N0phu6, Zp5iu6);  // ../RTL/cortexm0ds_logic.v(4244)
  not u2605 (Sp5iu6, n423);  // ../RTL/cortexm0ds_logic.v(4244)
  not u2606 (Zp5iu6, Odgpw6[20]);  // ../RTL/cortexm0ds_logic.v(4245)
  and u2607 (n424, U0phu6, Gq5iu6);  // ../RTL/cortexm0ds_logic.v(4246)
  not u2608 (Lp5iu6, n424);  // ../RTL/cortexm0ds_logic.v(4246)
  not u2609 (Gq5iu6, Odgpw6[19]);  // ../RTL/cortexm0ds_logic.v(4247)
  buf u261 (vis_psp_o[8], Huxpw6);  // ../RTL/cortexm0ds_logic.v(2085)
  and u2610 (Mm5iu6, Nq5iu6, Uq5iu6);  // ../RTL/cortexm0ds_logic.v(4248)
  and u2611 (Uq5iu6, Br5iu6, Ir5iu6);  // ../RTL/cortexm0ds_logic.v(4249)
  and u2612 (n425, B1phu6, Pr5iu6);  // ../RTL/cortexm0ds_logic.v(4250)
  not u2613 (Ir5iu6, n425);  // ../RTL/cortexm0ds_logic.v(4250)
  not u2614 (Pr5iu6, Odgpw6[18]);  // ../RTL/cortexm0ds_logic.v(4251)
  and u2615 (n426, I1phu6, Wr5iu6);  // ../RTL/cortexm0ds_logic.v(4252)
  not u2616 (Br5iu6, n426);  // ../RTL/cortexm0ds_logic.v(4252)
  not u2617 (Wr5iu6, Odgpw6[17]);  // ../RTL/cortexm0ds_logic.v(4253)
  and u2618 (Nq5iu6, Ds5iu6, Ks5iu6);  // ../RTL/cortexm0ds_logic.v(4254)
  and u2619 (n427, P1phu6, Rs5iu6);  // ../RTL/cortexm0ds_logic.v(4255)
  buf u262 (vis_r1_o[16], C7wpw6);  // ../RTL/cortexm0ds_logic.v(1876)
  not u2620 (Ks5iu6, n427);  // ../RTL/cortexm0ds_logic.v(4255)
  not u2621 (Rs5iu6, Odgpw6[16]);  // ../RTL/cortexm0ds_logic.v(4256)
  and u2622 (n428, W1phu6, Ys5iu6);  // ../RTL/cortexm0ds_logic.v(4257)
  not u2623 (Ds5iu6, n428);  // ../RTL/cortexm0ds_logic.v(4257)
  not u2624 (Ys5iu6, Odgpw6[15]);  // ../RTL/cortexm0ds_logic.v(4258)
  and u2625 (Id5iu6, Ft5iu6, Mt5iu6);  // ../RTL/cortexm0ds_logic.v(4259)
  and u2626 (Mt5iu6, Tt5iu6, Au5iu6);  // ../RTL/cortexm0ds_logic.v(4260)
  and u2627 (Au5iu6, Hu5iu6, Ou5iu6);  // ../RTL/cortexm0ds_logic.v(4261)
  and u2628 (Ou5iu6, Vu5iu6, Cv5iu6);  // ../RTL/cortexm0ds_logic.v(4262)
  and u2629 (n429, R2phu6, Jv5iu6);  // ../RTL/cortexm0ds_logic.v(4263)
  buf u263 (vis_r1_o[14], Sz7ax6);  // ../RTL/cortexm0ds_logic.v(1876)
  not u2630 (Cv5iu6, n429);  // ../RTL/cortexm0ds_logic.v(4263)
  not u2631 (Jv5iu6, Odgpw6[12]);  // ../RTL/cortexm0ds_logic.v(4264)
  and u2632 (Vu5iu6, Qv5iu6, Xv5iu6);  // ../RTL/cortexm0ds_logic.v(4265)
  and u2633 (n430, D2phu6, Ew5iu6);  // ../RTL/cortexm0ds_logic.v(4266)
  not u2634 (Xv5iu6, n430);  // ../RTL/cortexm0ds_logic.v(4266)
  not u2635 (Ew5iu6, Odgpw6[14]);  // ../RTL/cortexm0ds_logic.v(4267)
  and u2636 (n431, K2phu6, Lw5iu6);  // ../RTL/cortexm0ds_logic.v(4268)
  not u2637 (Qv5iu6, n431);  // ../RTL/cortexm0ds_logic.v(4268)
  not u2638 (Lw5iu6, Odgpw6[13]);  // ../RTL/cortexm0ds_logic.v(4269)
  and u2639 (Hu5iu6, Sw5iu6, Zw5iu6);  // ../RTL/cortexm0ds_logic.v(4270)
  buf u264 (R4gpw6[60], Hbgbx6);  // ../RTL/cortexm0ds_logic.v(2815)
  and u2640 (n432, Y2phu6, Gx5iu6);  // ../RTL/cortexm0ds_logic.v(4271)
  not u2641 (Zw5iu6, n432);  // ../RTL/cortexm0ds_logic.v(4271)
  not u2642 (Gx5iu6, Odgpw6[11]);  // ../RTL/cortexm0ds_logic.v(4272)
  and u2643 (n433, F3phu6, Nx5iu6);  // ../RTL/cortexm0ds_logic.v(4273)
  not u2644 (Sw5iu6, n433);  // ../RTL/cortexm0ds_logic.v(4273)
  not u2645 (Nx5iu6, Odgpw6[10]);  // ../RTL/cortexm0ds_logic.v(4274)
  and u2646 (Tt5iu6, Ux5iu6, By5iu6);  // ../RTL/cortexm0ds_logic.v(4275)
  and u2647 (By5iu6, Iy5iu6, Py5iu6);  // ../RTL/cortexm0ds_logic.v(4276)
  and u2648 (n434, M3phu6, Wy5iu6);  // ../RTL/cortexm0ds_logic.v(4277)
  not u2649 (Py5iu6, n434);  // ../RTL/cortexm0ds_logic.v(4277)
  buf u265 (vis_r5_o[21], Ljppw6);  // ../RTL/cortexm0ds_logic.v(1909)
  not u2650 (Wy5iu6, Odgpw6[7]);  // ../RTL/cortexm0ds_logic.v(4278)
  and u2651 (n435, T3phu6, Dz5iu6);  // ../RTL/cortexm0ds_logic.v(4279)
  not u2652 (Iy5iu6, n435);  // ../RTL/cortexm0ds_logic.v(4279)
  not u2653 (Dz5iu6, Odgpw6[6]);  // ../RTL/cortexm0ds_logic.v(4280)
  and u2654 (Ux5iu6, Kz5iu6, Rz5iu6);  // ../RTL/cortexm0ds_logic.v(4281)
  and u2655 (n436, A4phu6, Yz5iu6);  // ../RTL/cortexm0ds_logic.v(4282)
  not u2656 (Rz5iu6, n436);  // ../RTL/cortexm0ds_logic.v(4282)
  not u2657 (Yz5iu6, Odgpw6[5]);  // ../RTL/cortexm0ds_logic.v(4283)
  and u2658 (n437, H4phu6, F06iu6);  // ../RTL/cortexm0ds_logic.v(4284)
  not u2659 (Kz5iu6, n437);  // ../RTL/cortexm0ds_logic.v(4284)
  buf u266 (vis_psp_o[0], Ftypw6);  // ../RTL/cortexm0ds_logic.v(2085)
  not u2660 (F06iu6, Odgpw6[4]);  // ../RTL/cortexm0ds_logic.v(4285)
  and u2661 (Ft5iu6, M06iu6, T06iu6);  // ../RTL/cortexm0ds_logic.v(4286)
  and u2662 (T06iu6, A16iu6, H16iu6);  // ../RTL/cortexm0ds_logic.v(4287)
  and u2663 (H16iu6, O16iu6, V16iu6);  // ../RTL/cortexm0ds_logic.v(4288)
  and u2664 (n438, C5phu6, C26iu6);  // ../RTL/cortexm0ds_logic.v(4289)
  not u2665 (V16iu6, n438);  // ../RTL/cortexm0ds_logic.v(4289)
  not u2666 (C26iu6, Odgpw6[1]);  // ../RTL/cortexm0ds_logic.v(4290)
  and u2667 (O16iu6, J26iu6, Q26iu6);  // ../RTL/cortexm0ds_logic.v(4291)
  and u2668 (n439, O4phu6, X26iu6);  // ../RTL/cortexm0ds_logic.v(4292)
  not u2669 (Q26iu6, n439);  // ../RTL/cortexm0ds_logic.v(4292)
  buf u267 (Vbgpw6[30], Rz0bx6);  // ../RTL/cortexm0ds_logic.v(3092)
  not u2670 (X26iu6, Odgpw6[3]);  // ../RTL/cortexm0ds_logic.v(4293)
  and u2671 (n440, V4phu6, E36iu6);  // ../RTL/cortexm0ds_logic.v(4294)
  not u2672 (J26iu6, n440);  // ../RTL/cortexm0ds_logic.v(4294)
  not u2673 (E36iu6, Odgpw6[2]);  // ../RTL/cortexm0ds_logic.v(4295)
  and u2674 (A16iu6, L36iu6, S36iu6);  // ../RTL/cortexm0ds_logic.v(4296)
  and u2675 (n441, J5phu6, Z36iu6);  // ../RTL/cortexm0ds_logic.v(4297)
  not u2676 (S36iu6, n441);  // ../RTL/cortexm0ds_logic.v(4297)
  not u2677 (Z36iu6, Odgpw6[0]);  // ../RTL/cortexm0ds_logic.v(4298)
  and u2678 (n442, Bxdpw6, G46iu6);  // ../RTL/cortexm0ds_logic.v(4299)
  not u2679 (L36iu6, n442);  // ../RTL/cortexm0ds_logic.v(4299)
  buf u268 (vis_r4_o[24], Wjuax6);  // ../RTL/cortexm0ds_logic.v(2626)
  not u2680 (G46iu6, Odgpw6[8]);  // ../RTL/cortexm0ds_logic.v(4300)
  and u2681 (Bxdpw6, N46iu6, U46iu6);  // ../RTL/cortexm0ds_logic.v(4301)
  and u2682 (n443, B56iu6, I56iu6);  // ../RTL/cortexm0ds_logic.v(4302)
  not u2683 (U46iu6, n443);  // ../RTL/cortexm0ds_logic.v(4302)
  and u2684 (n444, Sodpw6, IRQ[8]);  // ../RTL/cortexm0ds_logic.v(4303)
  not u2685 (I56iu6, n444);  // ../RTL/cortexm0ds_logic.v(4303)
  and u2686 (B56iu6, P56iu6, W56iu6);  // ../RTL/cortexm0ds_logic.v(4304)
  and u2687 (n445, Odgpw6[8], D66iu6);  // ../RTL/cortexm0ds_logic.v(4305)
  not u2688 (P56iu6, n445);  // ../RTL/cortexm0ds_logic.v(4305)
  and u2689 (n446, K66iu6, HWDATA[8]);  // ../RTL/cortexm0ds_logic.v(4306)
  buf u269 (vis_r14_o[24], Nfnax6);  // ../RTL/cortexm0ds_logic.v(2497)
  not u2690 (D66iu6, n446);  // ../RTL/cortexm0ds_logic.v(4306)
  and u2691 (M06iu6, R66iu6, Y66iu6);  // ../RTL/cortexm0ds_logic.v(4307)
  and u2692 (Y66iu6, F76iu6, M76iu6);  // ../RTL/cortexm0ds_logic.v(4308)
  and u2693 (n447, Uwdpw6, T76iu6);  // ../RTL/cortexm0ds_logic.v(4309)
  not u2694 (M76iu6, n447);  // ../RTL/cortexm0ds_logic.v(4309)
  not u2695 (T76iu6, Odgpw6[9]);  // ../RTL/cortexm0ds_logic.v(4310)
  and u2696 (Uwdpw6, A86iu6, H86iu6);  // ../RTL/cortexm0ds_logic.v(4311)
  and u2697 (n448, O86iu6, V86iu6);  // ../RTL/cortexm0ds_logic.v(4312)
  not u2698 (H86iu6, n448);  // ../RTL/cortexm0ds_logic.v(4312)
  and u2699 (n449, Cndpw6, IRQ[9]);  // ../RTL/cortexm0ds_logic.v(4313)
  buf u27 (vis_r0_o[0], N0lax6);  // ../RTL/cortexm0ds_logic.v(1875)
  buf u270 (A2nhu6, Dg2qw6);  // ../RTL/cortexm0ds_logic.v(2151)
  not u2700 (V86iu6, n449);  // ../RTL/cortexm0ds_logic.v(4313)
  and u2701 (O86iu6, C96iu6, J96iu6);  // ../RTL/cortexm0ds_logic.v(4314)
  and u2702 (n450, Odgpw6[9], Q96iu6);  // ../RTL/cortexm0ds_logic.v(4315)
  not u2703 (C96iu6, n450);  // ../RTL/cortexm0ds_logic.v(4315)
  and u2704 (n451, K66iu6, HWDATA[9]);  // ../RTL/cortexm0ds_logic.v(4316)
  not u2705 (Q96iu6, n451);  // ../RTL/cortexm0ds_logic.v(4316)
  and u2706 (n452, Nwdpw6, X96iu6);  // ../RTL/cortexm0ds_logic.v(4317)
  not u2707 (F76iu6, n452);  // ../RTL/cortexm0ds_logic.v(4317)
  not u2708 (X96iu6, Odgpw6[24]);  // ../RTL/cortexm0ds_logic.v(4318)
  and u2709 (Nwdpw6, Ea6iu6, La6iu6);  // ../RTL/cortexm0ds_logic.v(4319)
  buf u271 (R6hhu6, Uh2qw6);  // ../RTL/cortexm0ds_logic.v(2152)
  and u2710 (n453, Sa6iu6, Za6iu6);  // ../RTL/cortexm0ds_logic.v(4320)
  not u2711 (La6iu6, n453);  // ../RTL/cortexm0ds_logic.v(4320)
  and u2712 (n454, Wqdpw6, IRQ[24]);  // ../RTL/cortexm0ds_logic.v(4321)
  not u2713 (Za6iu6, n454);  // ../RTL/cortexm0ds_logic.v(4321)
  and u2714 (Sa6iu6, Gb6iu6, Nb6iu6);  // ../RTL/cortexm0ds_logic.v(4322)
  and u2715 (n455, Odgpw6[24], Ub6iu6);  // ../RTL/cortexm0ds_logic.v(4323)
  not u2716 (Gb6iu6, n455);  // ../RTL/cortexm0ds_logic.v(4323)
  and u2717 (n456, K66iu6, HWDATA[24]);  // ../RTL/cortexm0ds_logic.v(4324)
  not u2718 (Ub6iu6, n456);  // ../RTL/cortexm0ds_logic.v(4324)
  and u2719 (R66iu6, Bc6iu6, Ic6iu6);  // ../RTL/cortexm0ds_logic.v(4325)
  buf u272 (D8hhu6, Nj2qw6);  // ../RTL/cortexm0ds_logic.v(2153)
  and u2720 (n457, Gwdpw6, Pc6iu6);  // ../RTL/cortexm0ds_logic.v(4326)
  not u2721 (Ic6iu6, n457);  // ../RTL/cortexm0ds_logic.v(4326)
  not u2722 (Pc6iu6, Odgpw6[25]);  // ../RTL/cortexm0ds_logic.v(4327)
  and u2723 (Gwdpw6, Wc6iu6, Dd6iu6);  // ../RTL/cortexm0ds_logic.v(4328)
  and u2724 (n458, Kd6iu6, Rd6iu6);  // ../RTL/cortexm0ds_logic.v(4329)
  not u2725 (Dd6iu6, n458);  // ../RTL/cortexm0ds_logic.v(4329)
  and u2726 (n459, Krdpw6, IRQ[25]);  // ../RTL/cortexm0ds_logic.v(4330)
  not u2727 (Rd6iu6, n459);  // ../RTL/cortexm0ds_logic.v(4330)
  and u2728 (Kd6iu6, Yd6iu6, Fe6iu6);  // ../RTL/cortexm0ds_logic.v(4331)
  and u2729 (n460, Odgpw6[25], Me6iu6);  // ../RTL/cortexm0ds_logic.v(4332)
  buf u273 (Jfgpw6[2], W5ypw6);  // ../RTL/cortexm0ds_logic.v(2010)
  not u2730 (Yd6iu6, n460);  // ../RTL/cortexm0ds_logic.v(4332)
  and u2731 (n461, K66iu6, HWDATA[25]);  // ../RTL/cortexm0ds_logic.v(4333)
  not u2732 (Me6iu6, n461);  // ../RTL/cortexm0ds_logic.v(4333)
  and u2733 (n462, Npghu6, Te6iu6);  // ../RTL/cortexm0ds_logic.v(4334)
  not u2734 (Bc6iu6, n462);  // ../RTL/cortexm0ds_logic.v(4334)
  and u2735 (Npghu6, Af6iu6, Hf6iu6);  // ../RTL/cortexm0ds_logic.v(4335)
  and u2736 (n463, Of6iu6, Vf6iu6);  // ../RTL/cortexm0ds_logic.v(4336)
  not u2737 (Hf6iu6, n463);  // ../RTL/cortexm0ds_logic.v(4336)
  and u2738 (n464, Evdpw6, NMI);  // ../RTL/cortexm0ds_logic.v(4337)
  not u2739 (Vf6iu6, n464);  // ../RTL/cortexm0ds_logic.v(4337)
  buf u274 (vis_r5_o[26], X1upw6);  // ../RTL/cortexm0ds_logic.v(1909)
  and u2740 (Of6iu6, Cg6iu6, Jg6iu6);  // ../RTL/cortexm0ds_logic.v(4338)
  or u2741 (Cg6iu6, Te6iu6, Qg6iu6);  // ../RTL/cortexm0ds_logic.v(4339)
  AL_MUX u2742 (
    .i0(Xg6iu6),
    .i1(R0nhu6),
    .sel(Eh6iu6),
    .o(C4xhu6));  // ../RTL/cortexm0ds_logic.v(4340)
  and u2743 (n465, Lh6iu6, Sh6iu6);  // ../RTL/cortexm0ds_logic.v(4341)
  not u2744 (O3xhu6, n465);  // ../RTL/cortexm0ds_logic.v(4341)
  or u2745 (Sh6iu6, Zh6iu6, HREADY);  // ../RTL/cortexm0ds_logic.v(4342)
  and u2746 (Lh6iu6, Gi6iu6, Ni6iu6);  // ../RTL/cortexm0ds_logic.v(4343)
  and u2747 (n466, Ui6iu6, Nr4iu6);  // ../RTL/cortexm0ds_logic.v(4344)
  not u2748 (Gi6iu6, n466);  // ../RTL/cortexm0ds_logic.v(4344)
  xor u2749 (n467, Bj6iu6, Jshpw6[5]);  // ../RTL/cortexm0ds_logic.v(4345)
  buf u275 (vis_r8_o[4], Rgrax6);  // ../RTL/cortexm0ds_logic.v(2579)
  not u2750 (Ui6iu6, n467);  // ../RTL/cortexm0ds_logic.v(4345)
  and u2751 (n468, Ij6iu6, Pj6iu6);  // ../RTL/cortexm0ds_logic.v(4346)
  not u2752 (H3xhu6, n468);  // ../RTL/cortexm0ds_logic.v(4346)
  or u2753 (Pj6iu6, Wj6iu6, HREADY);  // ../RTL/cortexm0ds_logic.v(4347)
  and u2754 (Ij6iu6, Dk6iu6, Ni6iu6);  // ../RTL/cortexm0ds_logic.v(4348)
  and u2755 (n469, Kk6iu6, Nr4iu6);  // ../RTL/cortexm0ds_logic.v(4349)
  not u2756 (Dk6iu6, n469);  // ../RTL/cortexm0ds_logic.v(4349)
  xor u2757 (n470, Bj6iu6, Jshpw6[13]);  // ../RTL/cortexm0ds_logic.v(4350)
  not u2758 (Kk6iu6, n470);  // ../RTL/cortexm0ds_logic.v(4350)
  and u2759 (n471, Rk6iu6, Yk6iu6);  // ../RTL/cortexm0ds_logic.v(4351)
  buf u276 (Jehhu6, Gr2qw6);  // ../RTL/cortexm0ds_logic.v(2157)
  not u2760 (A3xhu6, n471);  // ../RTL/cortexm0ds_logic.v(4351)
  or u2761 (Yk6iu6, Fl6iu6, HREADY);  // ../RTL/cortexm0ds_logic.v(4352)
  and u2762 (Rk6iu6, Ml6iu6, Ni6iu6);  // ../RTL/cortexm0ds_logic.v(4353)
  and u2763 (n472, Tl6iu6, Nr4iu6);  // ../RTL/cortexm0ds_logic.v(4354)
  not u2764 (Ml6iu6, n472);  // ../RTL/cortexm0ds_logic.v(4354)
  xor u2765 (n473, Am6iu6, Jshpw6[4]);  // ../RTL/cortexm0ds_logic.v(4355)
  not u2766 (Tl6iu6, n473);  // ../RTL/cortexm0ds_logic.v(4355)
  and u2767 (n474, Hm6iu6, Om6iu6);  // ../RTL/cortexm0ds_logic.v(4356)
  not u2768 (T2xhu6, n474);  // ../RTL/cortexm0ds_logic.v(4356)
  or u2769 (Om6iu6, Vm6iu6, HREADY);  // ../RTL/cortexm0ds_logic.v(4357)
  buf u277 (P9hhu6, Bt2qw6);  // ../RTL/cortexm0ds_logic.v(2158)
  and u2770 (Hm6iu6, Cn6iu6, Ni6iu6);  // ../RTL/cortexm0ds_logic.v(4358)
  and u2771 (n475, Jn6iu6, Nr4iu6);  // ../RTL/cortexm0ds_logic.v(4359)
  not u2772 (Cn6iu6, n475);  // ../RTL/cortexm0ds_logic.v(4359)
  xor u2773 (n476, Am6iu6, Jshpw6[12]);  // ../RTL/cortexm0ds_logic.v(4360)
  not u2774 (Jn6iu6, n476);  // ../RTL/cortexm0ds_logic.v(4360)
  and u2775 (n477, Qn6iu6, Xn6iu6);  // ../RTL/cortexm0ds_logic.v(4361)
  not u2776 (M2xhu6, n477);  // ../RTL/cortexm0ds_logic.v(4361)
  or u2777 (Xn6iu6, Eo6iu6, HREADY);  // ../RTL/cortexm0ds_logic.v(4362)
  and u2778 (Qn6iu6, Lo6iu6, Ni6iu6);  // ../RTL/cortexm0ds_logic.v(4363)
  and u2779 (n478, Nr4iu6, So6iu6);  // ../RTL/cortexm0ds_logic.v(4364)
  buf u278 (vis_r4_o[20], Vxuax6);  // ../RTL/cortexm0ds_logic.v(2626)
  not u2780 (Lo6iu6, n478);  // ../RTL/cortexm0ds_logic.v(4364)
  xor u2781 (n479, Zo6iu6, Jshpw6[15]);  // ../RTL/cortexm0ds_logic.v(4365)
  not u2782 (So6iu6, n479);  // ../RTL/cortexm0ds_logic.v(4365)
  and u2783 (n480, Gp6iu6, Np6iu6);  // ../RTL/cortexm0ds_logic.v(4366)
  not u2784 (F2xhu6, n480);  // ../RTL/cortexm0ds_logic.v(4366)
  and u2785 (n481, X8hpw6[1], Eh6iu6);  // ../RTL/cortexm0ds_logic.v(4367)
  not u2786 (Np6iu6, n481);  // ../RTL/cortexm0ds_logic.v(4367)
  and u2787 (Gp6iu6, Up6iu6, Ni6iu6);  // ../RTL/cortexm0ds_logic.v(4368)
  or u2788 (Up6iu6, Bq6iu6, Iq6iu6);  // ../RTL/cortexm0ds_logic.v(4369)
  and u2789 (n482, Pq6iu6, Wq6iu6);  // ../RTL/cortexm0ds_logic.v(4370)
  buf u279 (vis_r14_o[17], Nxnax6);  // ../RTL/cortexm0ds_logic.v(2497)
  not u2790 (Y1xhu6, n482);  // ../RTL/cortexm0ds_logic.v(4370)
  or u2791 (Wq6iu6, Dr6iu6, HREADY);  // ../RTL/cortexm0ds_logic.v(4371)
  and u2792 (Pq6iu6, Kr6iu6, Ni6iu6);  // ../RTL/cortexm0ds_logic.v(4372)
  and u2793 (n483, Nr4iu6, Rr6iu6);  // ../RTL/cortexm0ds_logic.v(4373)
  not u2794 (Ni6iu6, n483);  // ../RTL/cortexm0ds_logic.v(4373)
  and u2795 (n484, Yr6iu6, Fs6iu6);  // ../RTL/cortexm0ds_logic.v(4374)
  not u2796 (Rr6iu6, n484);  // ../RTL/cortexm0ds_logic.v(4374)
  and u2797 (Yr6iu6, Ms6iu6, Ts6iu6);  // ../RTL/cortexm0ds_logic.v(4375)
  and u2798 (Ts6iu6, At6iu6, Ht6iu6);  // ../RTL/cortexm0ds_logic.v(4376)
  or u2799 (Ht6iu6, Wqzhu6, Aphpw6[2]);  // ../RTL/cortexm0ds_logic.v(4377)
  buf u28 (vis_r0_o[24], Ynspw6);  // ../RTL/cortexm0ds_logic.v(1875)
  buf u280 (Jdnhu6, Ry2qw6);  // ../RTL/cortexm0ds_logic.v(2161)
  and u2800 (Ms6iu6, Ot6iu6, Vt6iu6);  // ../RTL/cortexm0ds_logic.v(4378)
  or u2801 (Vt6iu6, Cu6iu6, Jshpw6[8]);  // ../RTL/cortexm0ds_logic.v(4379)
  not u2802 (Cu6iu6, Jshpw6[11]);  // ../RTL/cortexm0ds_logic.v(4380)
  AL_MUX u2803 (
    .i0(Ju6iu6),
    .i1(Qu6iu6),
    .sel(Jshpw6[10]),
    .o(Ot6iu6));  // ../RTL/cortexm0ds_logic.v(4381)
  and u2804 (Qu6iu6, Jshpw6[11], Xu6iu6);  // ../RTL/cortexm0ds_logic.v(4382)
  and u2805 (n485, Ev6iu6, Lv6iu6);  // ../RTL/cortexm0ds_logic.v(4383)
  not u2806 (Xu6iu6, n485);  // ../RTL/cortexm0ds_logic.v(4383)
  and u2807 (n486, Sv6iu6, Zv6iu6);  // ../RTL/cortexm0ds_logic.v(4384)
  not u2808 (Lv6iu6, n486);  // ../RTL/cortexm0ds_logic.v(4384)
  and u2809 (Zv6iu6, Gw6iu6, Nw6iu6);  // ../RTL/cortexm0ds_logic.v(4385)
  buf u281 (vis_r8_o[26], X3upw6);  // ../RTL/cortexm0ds_logic.v(2579)
  and u2810 (Gw6iu6, Uw6iu6, Bx6iu6);  // ../RTL/cortexm0ds_logic.v(4386)
  and u2811 (Sv6iu6, Ix6iu6, Px6iu6);  // ../RTL/cortexm0ds_logic.v(4387)
  AL_MUX u2812 (
    .i0(Wx6iu6),
    .i1(Dy6iu6),
    .sel(Jshpw6[6]),
    .o(Px6iu6));  // ../RTL/cortexm0ds_logic.v(4388)
  or u2813 (n487, Ky6iu6, Ry6iu6);  // ../RTL/cortexm0ds_logic.v(4389)
  not u2814 (Dy6iu6, n487);  // ../RTL/cortexm0ds_logic.v(4389)
  and u2815 (Wx6iu6, Yy6iu6, Bj6iu6);  // ../RTL/cortexm0ds_logic.v(4390)
  or u2816 (n488, Jshpw6[7], Jshpw6[9]);  // ../RTL/cortexm0ds_logic.v(4391)
  not u2817 (Yy6iu6, n488);  // ../RTL/cortexm0ds_logic.v(4391)
  and u2818 (Ix6iu6, Fz6iu6, Mz6iu6);  // ../RTL/cortexm0ds_logic.v(4392)
  xor u2819 (n489, Jshpw6[4], Jshpw6[5]);  // ../RTL/cortexm0ds_logic.v(4393)
  buf u282 (Mdhpw6[0], Krlpw6);  // ../RTL/cortexm0ds_logic.v(1838)
  not u2820 (Fz6iu6, n489);  // ../RTL/cortexm0ds_logic.v(4393)
  and u2821 (n490, Tz6iu6, A07iu6);  // ../RTL/cortexm0ds_logic.v(4394)
  not u2822 (Ev6iu6, n490);  // ../RTL/cortexm0ds_logic.v(4394)
  and u2823 (A07iu6, Jshpw6[6], H07iu6);  // ../RTL/cortexm0ds_logic.v(4395)
  and u2824 (n491, O07iu6, V07iu6);  // ../RTL/cortexm0ds_logic.v(4396)
  not u2825 (H07iu6, n491);  // ../RTL/cortexm0ds_logic.v(4396)
  and u2826 (n492, C17iu6, J17iu6);  // ../RTL/cortexm0ds_logic.v(4397)
  not u2827 (V07iu6, n492);  // ../RTL/cortexm0ds_logic.v(4397)
  or u2828 (V77iu6, Am6iu6, Bj6iu6);  // ../RTL/cortexm0ds_logic.v(4398)
  not u2829 (C17iu6, V77iu6);  // ../RTL/cortexm0ds_logic.v(4398)
  buf u283 (vis_r14_o[22], Tdfbx6);  // ../RTL/cortexm0ds_logic.v(2497)
  and u2830 (n493, Q17iu6, X17iu6);  // ../RTL/cortexm0ds_logic.v(4399)
  not u2831 (O07iu6, n493);  // ../RTL/cortexm0ds_logic.v(4399)
  and u2832 (n494, E27iu6, L27iu6);  // ../RTL/cortexm0ds_logic.v(4400)
  not u2833 (X17iu6, n494);  // ../RTL/cortexm0ds_logic.v(4400)
  and u2834 (n495, S27iu6, Z27iu6);  // ../RTL/cortexm0ds_logic.v(4401)
  not u2835 (E27iu6, n495);  // ../RTL/cortexm0ds_logic.v(4401)
  AL_MUX u2836 (
    .i0(G37iu6),
    .i1(Jshpw6[13]),
    .sel(Bx6iu6),
    .o(S27iu6));  // ../RTL/cortexm0ds_logic.v(4402)
  and u2837 (n496, N37iu6, U37iu6);  // ../RTL/cortexm0ds_logic.v(4403)
  not u2838 (Q17iu6, n496);  // ../RTL/cortexm0ds_logic.v(4403)
  and u2839 (n497, B47iu6, Jshpw6[4]);  // ../RTL/cortexm0ds_logic.v(4404)
  buf u284 (vis_r4_o[19], Vzuax6);  // ../RTL/cortexm0ds_logic.v(2626)
  not u2840 (N37iu6, n497);  // ../RTL/cortexm0ds_logic.v(4404)
  or u2841 (n498, I47iu6, P47iu6);  // ../RTL/cortexm0ds_logic.v(4405)
  not u2842 (B47iu6, n498);  // ../RTL/cortexm0ds_logic.v(4405)
  or u2843 (n499, Iq6iu6, Ky6iu6);  // ../RTL/cortexm0ds_logic.v(4406)
  not u2844 (Tz6iu6, n499);  // ../RTL/cortexm0ds_logic.v(4406)
  not u2845 (Iq6iu6, Jshpw6[9]);  // ../RTL/cortexm0ds_logic.v(4407)
  and u2846 (Ju6iu6, W47iu6, D57iu6);  // ../RTL/cortexm0ds_logic.v(4408)
  and u2847 (D57iu6, K57iu6, Ky6iu6);  // ../RTL/cortexm0ds_logic.v(4409)
  not u2848 (Ky6iu6, Jshpw6[7]);  // ../RTL/cortexm0ds_logic.v(4410)
  or u2849 (n500, Jshpw6[8], Jshpw6[9]);  // ../RTL/cortexm0ds_logic.v(4411)
  buf u285 (vis_r14_o[16], Nznax6);  // ../RTL/cortexm0ds_logic.v(2497)
  not u2850 (K57iu6, n500);  // ../RTL/cortexm0ds_logic.v(4411)
  and u2851 (W47iu6, R57iu6, Zo6iu6);  // ../RTL/cortexm0ds_logic.v(4412)
  not u2852 (Zo6iu6, Jshpw6[6]);  // ../RTL/cortexm0ds_logic.v(4413)
  and u2853 (n501, Y57iu6, F67iu6);  // ../RTL/cortexm0ds_logic.v(4414)
  not u2854 (R57iu6, n501);  // ../RTL/cortexm0ds_logic.v(4414)
  and u2855 (n502, M67iu6, T67iu6);  // ../RTL/cortexm0ds_logic.v(4415)
  not u2856 (F67iu6, n502);  // ../RTL/cortexm0ds_logic.v(4415)
  and u2857 (T67iu6, A77iu6, Mz6iu6);  // ../RTL/cortexm0ds_logic.v(4416)
  or u2858 (n503, Bx6iu6, Jshpw6[15]);  // ../RTL/cortexm0ds_logic.v(4417)
  not u2859 (A77iu6, n503);  // ../RTL/cortexm0ds_logic.v(4417)
  buf u286 (vis_r8_o[25], Osrax6);  // ../RTL/cortexm0ds_logic.v(2579)
  and u2860 (M67iu6, H77iu6, G37iu6);  // ../RTL/cortexm0ds_logic.v(4418)
  or u2861 (n504, Jshpw6[14], Jshpw6[13]);  // ../RTL/cortexm0ds_logic.v(4419)
  not u2862 (G37iu6, n504);  // ../RTL/cortexm0ds_logic.v(4419)
  AL_MUX u2863 (
    .i0(O77iu6),
    .i1(V77iu6),
    .sel(Jshpw6[5]),
    .o(H77iu6));  // ../RTL/cortexm0ds_logic.v(4420)
  buf u2864 (Kmehu6, Ozkbx6[26]);  // ../RTL/cortexm0ds_logic.v(3176)
  and u2865 (O77iu6, C87iu6, J87iu6);  // ../RTL/cortexm0ds_logic.v(4422)
  or u2866 (J87iu6, Bj6iu6, Jshpw6[4]);  // ../RTL/cortexm0ds_logic.v(4423)
  AL_MUX u2867 (
    .i0(Ry6iu6),
    .i1(P47iu6),
    .sel(I47iu6),
    .o(C87iu6));  // ../RTL/cortexm0ds_logic.v(4424)
  not u2868 (Ry6iu6, Jshpw6[4]);  // ../RTL/cortexm0ds_logic.v(4425)
  and u2869 (n505, U37iu6, Q87iu6);  // ../RTL/cortexm0ds_logic.v(4426)
  buf u287 (Cynhu6, Tb3qw6);  // ../RTL/cortexm0ds_logic.v(2168)
  not u2870 (Y57iu6, n505);  // ../RTL/cortexm0ds_logic.v(4426)
  or u2871 (Q87iu6, J17iu6, X87iu6);  // ../RTL/cortexm0ds_logic.v(4427)
  and u2872 (X87iu6, E97iu6, L97iu6);  // ../RTL/cortexm0ds_logic.v(4428)
  and u2873 (L97iu6, S97iu6, Jshpw6[13]);  // ../RTL/cortexm0ds_logic.v(4429)
  and u2874 (S97iu6, Z97iu6, Bx6iu6);  // ../RTL/cortexm0ds_logic.v(4430)
  and u2875 (n506, Jshpw6[14], Uw6iu6);  // ../RTL/cortexm0ds_logic.v(4431)
  not u2876 (Z97iu6, n506);  // ../RTL/cortexm0ds_logic.v(4431)
  or u2877 (Uw6iu6, Am6iu6, P47iu6);  // ../RTL/cortexm0ds_logic.v(4432)
  not u2878 (Am6iu6, I47iu6);  // ../RTL/cortexm0ds_logic.v(4433)
  or u2879 (n507, Ga7iu6, Na7iu6);  // ../RTL/cortexm0ds_logic.v(4434)
  buf u288 (Vbgpw6[16], Ih0bx6);  // ../RTL/cortexm0ds_logic.v(3092)
  not u2880 (E97iu6, n507);  // ../RTL/cortexm0ds_logic.v(4434)
  not u2881 (Na7iu6, Z27iu6);  // ../RTL/cortexm0ds_logic.v(4435)
  and u2882 (Z27iu6, Ua7iu6, Mz6iu6);  // ../RTL/cortexm0ds_logic.v(4436)
  xor u2883 (n508, Jshpw6[14], Jshpw6[15]);  // ../RTL/cortexm0ds_logic.v(4437)
  not u2884 (Ua7iu6, n508);  // ../RTL/cortexm0ds_logic.v(4437)
  AL_MUX u2885 (
    .i0(Bb7iu6),
    .i1(I47iu6),
    .sel(Jshpw6[4]),
    .o(Ga7iu6));  // ../RTL/cortexm0ds_logic.v(4438)
  or u2886 (n509, I47iu6, Bj6iu6);  // ../RTL/cortexm0ds_logic.v(4439)
  not u2887 (Bb7iu6, n509);  // ../RTL/cortexm0ds_logic.v(4439)
  not u2888 (Bj6iu6, P47iu6);  // ../RTL/cortexm0ds_logic.v(4440)
  or u2889 (n510, L27iu6, Jshpw6[4]);  // ../RTL/cortexm0ds_logic.v(4441)
  buf u289 (Vbgpw6[18], Kl0bx6);  // ../RTL/cortexm0ds_logic.v(3092)
  not u2890 (J17iu6, n510);  // ../RTL/cortexm0ds_logic.v(4441)
  and u2891 (n511, Ib7iu6, Pb7iu6);  // ../RTL/cortexm0ds_logic.v(4442)
  not u2892 (L27iu6, n511);  // ../RTL/cortexm0ds_logic.v(4442)
  and u2893 (Pb7iu6, Wb7iu6, Jshpw6[17]);  // ../RTL/cortexm0ds_logic.v(4443)
  and u2894 (Wb7iu6, Jshpw6[16], Jshpw6[12]);  // ../RTL/cortexm0ds_logic.v(4444)
  and u2895 (Ib7iu6, Dc7iu6, Nw6iu6);  // ../RTL/cortexm0ds_logic.v(4445)
  and u2896 (Nw6iu6, Kc7iu6, Jshpw6[15]);  // ../RTL/cortexm0ds_logic.v(4446)
  and u2897 (Dc7iu6, Jshpw6[19], Jshpw6[18]);  // ../RTL/cortexm0ds_logic.v(4447)
  not u2898 (U37iu6, Jshpw6[5]);  // ../RTL/cortexm0ds_logic.v(4448)
  not u2899 (Nr4iu6, Bq6iu6);  // ../RTL/cortexm0ds_logic.v(4449)
  buf u29 (vis_r0_o[26], Xttpw6);  // ../RTL/cortexm0ds_logic.v(1875)
  buf u290 (Vbgpw6[19], Ln0bx6);  // ../RTL/cortexm0ds_logic.v(3092)
  or u2900 (Kr6iu6, Bq6iu6, Bx6iu6);  // ../RTL/cortexm0ds_logic.v(4450)
  AL_MUX u2901 (
    .i0(D84iu6),
    .i1(E5hhu6),
    .sel(Rc7iu6),
    .o(R1xhu6));  // ../RTL/cortexm0ds_logic.v(4451)
  AL_MUX u2902 (
    .i0(T24iu6),
    .i1(H2hhu6),
    .sel(Rc7iu6),
    .o(K1xhu6));  // ../RTL/cortexm0ds_logic.v(4452)
  AL_MUX u2903 (
    .i0(J44iu6),
    .i1(S3hhu6),
    .sel(Rc7iu6),
    .o(D1xhu6));  // ../RTL/cortexm0ds_logic.v(4453)
  and u2904 (n512, Yc7iu6, A2nhu6);  // ../RTL/cortexm0ds_logic.v(4454)
  not u2905 (Rc7iu6, n512);  // ../RTL/cortexm0ds_logic.v(4454)
  AL_MUX u2906 (
    .i0(T24iu6),
    .i1(Jehhu6),
    .sel(Fd7iu6),
    .o(W0xhu6));  // ../RTL/cortexm0ds_logic.v(4455)
  AL_MUX u2907 (
    .i0(Ud4iu6),
    .i1(Hbhhu6),
    .sel(Fd7iu6),
    .o(P0xhu6));  // ../RTL/cortexm0ds_logic.v(4456)
  not u2908 (Fd7iu6, Tu4iu6);  // ../RTL/cortexm0ds_logic.v(4457)
  AL_MUX u2909 (
    .i0(P9hhu6),
    .i1(Df4iu6),
    .sel(Tu4iu6),
    .o(I0xhu6));  // ../RTL/cortexm0ds_logic.v(4458)
  buf u291 (vis_r14_o[21], Npnax6);  // ../RTL/cortexm0ds_logic.v(2497)
  AL_MUX u2910 (
    .i0(Ud4iu6),
    .i1(Togpw6[2]),
    .sel(Md7iu6),
    .o(B0xhu6));  // ../RTL/cortexm0ds_logic.v(4459)
  AL_MUX u2911 (
    .i0(Lm1iu6),
    .i1(Ligpw6[28]),
    .sel(Md7iu6),
    .o(Uzwhu6));  // ../RTL/cortexm0ds_logic.v(4460)
  AL_MUX u2912 (
    .i0(T94iu6),
    .i1(Ligpw6[27]),
    .sel(Md7iu6),
    .o(Nzwhu6));  // ../RTL/cortexm0ds_logic.v(4461)
  AL_MUX u2913 (
    .i0(F94iu6),
    .i1(Togpw6[28]),
    .sel(Md7iu6),
    .o(Gzwhu6));  // ../RTL/cortexm0ds_logic.v(4462)
  AL_MUX u2914 (
    .i0(Y84iu6),
    .i1(Togpw6[27]),
    .sel(Md7iu6),
    .o(Zywhu6));  // ../RTL/cortexm0ds_logic.v(4463)
  AL_MUX u2915 (
    .i0(R84iu6),
    .i1(Togpw6[26]),
    .sel(Md7iu6),
    .o(Sywhu6));  // ../RTL/cortexm0ds_logic.v(4464)
  AL_MUX u2916 (
    .i0(K84iu6),
    .i1(Togpw6[25]),
    .sel(Md7iu6),
    .o(Lywhu6));  // ../RTL/cortexm0ds_logic.v(4465)
  AL_MUX u2917 (
    .i0(D84iu6),
    .i1(Togpw6[24]),
    .sel(Md7iu6),
    .o(Eywhu6));  // ../RTL/cortexm0ds_logic.v(4466)
  AL_MUX u2918 (
    .i0(W74iu6),
    .i1(Togpw6[23]),
    .sel(Md7iu6),
    .o(Xxwhu6));  // ../RTL/cortexm0ds_logic.v(4467)
  AL_MUX u2919 (
    .i0(P74iu6),
    .i1(Togpw6[22]),
    .sel(Md7iu6),
    .o(Qxwhu6));  // ../RTL/cortexm0ds_logic.v(4468)
  buf u292 (Vbgpw6[23], Ot0bx6);  // ../RTL/cortexm0ds_logic.v(3092)
  AL_MUX u2920 (
    .i0(I74iu6),
    .i1(Togpw6[21]),
    .sel(Md7iu6),
    .o(Jxwhu6));  // ../RTL/cortexm0ds_logic.v(4469)
  AL_MUX u2921 (
    .i0(B74iu6),
    .i1(Togpw6[20]),
    .sel(Md7iu6),
    .o(Cxwhu6));  // ../RTL/cortexm0ds_logic.v(4470)
  AL_MUX u2922 (
    .i0(U64iu6),
    .i1(Togpw6[19]),
    .sel(Md7iu6),
    .o(Vwwhu6));  // ../RTL/cortexm0ds_logic.v(4471)
  AL_MUX u2923 (
    .i0(N64iu6),
    .i1(Togpw6[18]),
    .sel(Md7iu6),
    .o(Owwhu6));  // ../RTL/cortexm0ds_logic.v(4472)
  AL_MUX u2924 (
    .i0(G64iu6),
    .i1(Togpw6[17]),
    .sel(Md7iu6),
    .o(Hwwhu6));  // ../RTL/cortexm0ds_logic.v(4473)
  AL_MUX u2925 (
    .i0(Z54iu6),
    .i1(Togpw6[16]),
    .sel(Md7iu6),
    .o(Awwhu6));  // ../RTL/cortexm0ds_logic.v(4474)
  AL_MUX u2926 (
    .i0(S54iu6),
    .i1(Togpw6[15]),
    .sel(Md7iu6),
    .o(Tvwhu6));  // ../RTL/cortexm0ds_logic.v(4475)
  AL_MUX u2927 (
    .i0(L54iu6),
    .i1(Togpw6[14]),
    .sel(Md7iu6),
    .o(Mvwhu6));  // ../RTL/cortexm0ds_logic.v(4476)
  AL_MUX u2928 (
    .i0(E54iu6),
    .i1(Togpw6[13]),
    .sel(Md7iu6),
    .o(Fvwhu6));  // ../RTL/cortexm0ds_logic.v(4477)
  AL_MUX u2929 (
    .i0(X44iu6),
    .i1(Togpw6[12]),
    .sel(Md7iu6),
    .o(Yuwhu6));  // ../RTL/cortexm0ds_logic.v(4478)
  buf u293 (Vbgpw6[5], Czzax6);  // ../RTL/cortexm0ds_logic.v(3092)
  AL_MUX u2930 (
    .i0(Q44iu6),
    .i1(Togpw6[11]),
    .sel(Md7iu6),
    .o(Ruwhu6));  // ../RTL/cortexm0ds_logic.v(4479)
  AL_MUX u2931 (
    .i0(J44iu6),
    .i1(Togpw6[10]),
    .sel(Md7iu6),
    .o(Kuwhu6));  // ../RTL/cortexm0ds_logic.v(4480)
  AL_MUX u2932 (
    .i0(Ym4iu6),
    .i1(Togpw6[9]),
    .sel(Md7iu6),
    .o(Duwhu6));  // ../RTL/cortexm0ds_logic.v(4481)
  AL_MUX u2933 (
    .i0(Pl4iu6),
    .i1(Togpw6[8]),
    .sel(Md7iu6),
    .o(Wtwhu6));  // ../RTL/cortexm0ds_logic.v(4482)
  AL_MUX u2934 (
    .i0(Gk4iu6),
    .i1(Togpw6[7]),
    .sel(Md7iu6),
    .o(Ptwhu6));  // ../RTL/cortexm0ds_logic.v(4483)
  AL_MUX u2935 (
    .i0(Xi4iu6),
    .i1(Togpw6[6]),
    .sel(Md7iu6),
    .o(Itwhu6));  // ../RTL/cortexm0ds_logic.v(4484)
  AL_MUX u2936 (
    .i0(Oh4iu6),
    .i1(Togpw6[5]),
    .sel(Md7iu6),
    .o(Btwhu6));  // ../RTL/cortexm0ds_logic.v(4485)
  AL_MUX u2937 (
    .i0(H34iu6),
    .i1(Togpw6[4]),
    .sel(Md7iu6),
    .o(Uswhu6));  // ../RTL/cortexm0ds_logic.v(4486)
  AL_MUX u2938 (
    .i0(Df4iu6),
    .i1(Togpw6[3]),
    .sel(Md7iu6),
    .o(Nswhu6));  // ../RTL/cortexm0ds_logic.v(4487)
  AL_MUX u2939 (
    .i0(T24iu6),
    .i1(Qhhhu6),
    .sel(Md7iu6),
    .o(Gswhu6));  // ../RTL/cortexm0ds_logic.v(4488)
  buf u294 (Vbgpw6[4], Ikhbx6);  // ../RTL/cortexm0ds_logic.v(3092)
  and u2940 (n513, A2nhu6, Vr1iu6);  // ../RTL/cortexm0ds_logic.v(4489)
  not u2941 (Md7iu6, n513);  // ../RTL/cortexm0ds_logic.v(4489)
  AL_MUX u2942 (
    .i0(Ud4iu6),
    .i1(Gqgpw6[2]),
    .sel(Td7iu6),
    .o(Zrwhu6));  // ../RTL/cortexm0ds_logic.v(4490)
  AL_MUX u2943 (
    .i0(Lm1iu6),
    .i1(Akgpw6[28]),
    .sel(Td7iu6),
    .o(Srwhu6));  // ../RTL/cortexm0ds_logic.v(4491)
  AL_MUX u2944 (
    .i0(T94iu6),
    .i1(Akgpw6[27]),
    .sel(Td7iu6),
    .o(Lrwhu6));  // ../RTL/cortexm0ds_logic.v(4492)
  AL_MUX u2945 (
    .i0(F94iu6),
    .i1(Gqgpw6[28]),
    .sel(Td7iu6),
    .o(Erwhu6));  // ../RTL/cortexm0ds_logic.v(4493)
  AL_MUX u2946 (
    .i0(Y84iu6),
    .i1(Gqgpw6[27]),
    .sel(Td7iu6),
    .o(Xqwhu6));  // ../RTL/cortexm0ds_logic.v(4494)
  AL_MUX u2947 (
    .i0(R84iu6),
    .i1(Gqgpw6[26]),
    .sel(Td7iu6),
    .o(Qqwhu6));  // ../RTL/cortexm0ds_logic.v(4495)
  AL_MUX u2948 (
    .i0(K84iu6),
    .i1(Gqgpw6[25]),
    .sel(Td7iu6),
    .o(Jqwhu6));  // ../RTL/cortexm0ds_logic.v(4496)
  AL_MUX u2949 (
    .i0(D84iu6),
    .i1(Gqgpw6[24]),
    .sel(Td7iu6),
    .o(Cqwhu6));  // ../RTL/cortexm0ds_logic.v(4497)
  buf u295 (vis_r4_o[30], B6uax6);  // ../RTL/cortexm0ds_logic.v(2626)
  AL_MUX u2950 (
    .i0(W74iu6),
    .i1(Gqgpw6[23]),
    .sel(Td7iu6),
    .o(Vpwhu6));  // ../RTL/cortexm0ds_logic.v(4498)
  AL_MUX u2951 (
    .i0(P74iu6),
    .i1(Gqgpw6[22]),
    .sel(Td7iu6),
    .o(Opwhu6));  // ../RTL/cortexm0ds_logic.v(4499)
  AL_MUX u2952 (
    .i0(I74iu6),
    .i1(Gqgpw6[21]),
    .sel(Td7iu6),
    .o(Hpwhu6));  // ../RTL/cortexm0ds_logic.v(4500)
  AL_MUX u2953 (
    .i0(B74iu6),
    .i1(Gqgpw6[20]),
    .sel(Td7iu6),
    .o(Apwhu6));  // ../RTL/cortexm0ds_logic.v(4501)
  AL_MUX u2954 (
    .i0(U64iu6),
    .i1(Gqgpw6[19]),
    .sel(Td7iu6),
    .o(Towhu6));  // ../RTL/cortexm0ds_logic.v(4502)
  AL_MUX u2955 (
    .i0(N64iu6),
    .i1(Gqgpw6[18]),
    .sel(Td7iu6),
    .o(Mowhu6));  // ../RTL/cortexm0ds_logic.v(4503)
  AL_MUX u2956 (
    .i0(G64iu6),
    .i1(Gqgpw6[17]),
    .sel(Td7iu6),
    .o(Fowhu6));  // ../RTL/cortexm0ds_logic.v(4504)
  AL_MUX u2957 (
    .i0(Z54iu6),
    .i1(Gqgpw6[16]),
    .sel(Td7iu6),
    .o(Ynwhu6));  // ../RTL/cortexm0ds_logic.v(4505)
  AL_MUX u2958 (
    .i0(S54iu6),
    .i1(Gqgpw6[15]),
    .sel(Td7iu6),
    .o(Rnwhu6));  // ../RTL/cortexm0ds_logic.v(4506)
  AL_MUX u2959 (
    .i0(L54iu6),
    .i1(Gqgpw6[14]),
    .sel(Td7iu6),
    .o(Knwhu6));  // ../RTL/cortexm0ds_logic.v(4507)
  buf u296 (vis_r4_o[25], Vtuax6);  // ../RTL/cortexm0ds_logic.v(2626)
  AL_MUX u2960 (
    .i0(E54iu6),
    .i1(Gqgpw6[13]),
    .sel(Td7iu6),
    .o(Dnwhu6));  // ../RTL/cortexm0ds_logic.v(4508)
  AL_MUX u2961 (
    .i0(X44iu6),
    .i1(Gqgpw6[12]),
    .sel(Td7iu6),
    .o(Wmwhu6));  // ../RTL/cortexm0ds_logic.v(4509)
  AL_MUX u2962 (
    .i0(Q44iu6),
    .i1(Gqgpw6[11]),
    .sel(Td7iu6),
    .o(Pmwhu6));  // ../RTL/cortexm0ds_logic.v(4510)
  AL_MUX u2963 (
    .i0(J44iu6),
    .i1(Gqgpw6[10]),
    .sel(Td7iu6),
    .o(Imwhu6));  // ../RTL/cortexm0ds_logic.v(4511)
  AL_MUX u2964 (
    .i0(Ym4iu6),
    .i1(Gqgpw6[9]),
    .sel(Td7iu6),
    .o(Bmwhu6));  // ../RTL/cortexm0ds_logic.v(4512)
  AL_MUX u2965 (
    .i0(Pl4iu6),
    .i1(Gqgpw6[8]),
    .sel(Td7iu6),
    .o(Ulwhu6));  // ../RTL/cortexm0ds_logic.v(4513)
  AL_MUX u2966 (
    .i0(Gk4iu6),
    .i1(Gqgpw6[7]),
    .sel(Td7iu6),
    .o(Nlwhu6));  // ../RTL/cortexm0ds_logic.v(4514)
  AL_MUX u2967 (
    .i0(Xi4iu6),
    .i1(Gqgpw6[6]),
    .sel(Td7iu6),
    .o(Glwhu6));  // ../RTL/cortexm0ds_logic.v(4515)
  AL_MUX u2968 (
    .i0(Oh4iu6),
    .i1(Gqgpw6[5]),
    .sel(Td7iu6),
    .o(Zkwhu6));  // ../RTL/cortexm0ds_logic.v(4516)
  AL_MUX u2969 (
    .i0(H34iu6),
    .i1(Gqgpw6[4]),
    .sel(Td7iu6),
    .o(Skwhu6));  // ../RTL/cortexm0ds_logic.v(4517)
  buf u297 (R4gpw6[61], Yt4bx6);  // ../RTL/cortexm0ds_logic.v(2815)
  AL_MUX u2970 (
    .i0(Df4iu6),
    .i1(Gqgpw6[3]),
    .sel(Td7iu6),
    .o(Lkwhu6));  // ../RTL/cortexm0ds_logic.v(4518)
  AL_MUX u2971 (
    .i0(T24iu6),
    .i1(Ijhhu6),
    .sel(Td7iu6),
    .o(Ekwhu6));  // ../RTL/cortexm0ds_logic.v(4519)
  and u2972 (n514, A2nhu6, Xs1iu6);  // ../RTL/cortexm0ds_logic.v(4520)
  not u2973 (Td7iu6, n514);  // ../RTL/cortexm0ds_logic.v(4520)
  AL_MUX u2974 (
    .i0(Ud4iu6),
    .i1(Trgpw6[2]),
    .sel(Ae7iu6),
    .o(Xjwhu6));  // ../RTL/cortexm0ds_logic.v(4521)
  AL_MUX u2975 (
    .i0(Lm1iu6),
    .i1(Plgpw6[28]),
    .sel(Ae7iu6),
    .o(Qjwhu6));  // ../RTL/cortexm0ds_logic.v(4522)
  AL_MUX u2976 (
    .i0(T94iu6),
    .i1(Plgpw6[27]),
    .sel(Ae7iu6),
    .o(Jjwhu6));  // ../RTL/cortexm0ds_logic.v(4523)
  AL_MUX u2977 (
    .i0(F94iu6),
    .i1(Trgpw6[28]),
    .sel(Ae7iu6),
    .o(Cjwhu6));  // ../RTL/cortexm0ds_logic.v(4524)
  AL_MUX u2978 (
    .i0(Y84iu6),
    .i1(Trgpw6[27]),
    .sel(Ae7iu6),
    .o(Viwhu6));  // ../RTL/cortexm0ds_logic.v(4525)
  AL_MUX u2979 (
    .i0(R84iu6),
    .i1(Trgpw6[26]),
    .sel(Ae7iu6),
    .o(Oiwhu6));  // ../RTL/cortexm0ds_logic.v(4526)
  buf u298 (vis_r5_o[22], T5fbx6);  // ../RTL/cortexm0ds_logic.v(1909)
  AL_MUX u2980 (
    .i0(K84iu6),
    .i1(Trgpw6[25]),
    .sel(Ae7iu6),
    .o(Hiwhu6));  // ../RTL/cortexm0ds_logic.v(4527)
  AL_MUX u2981 (
    .i0(D84iu6),
    .i1(Trgpw6[24]),
    .sel(Ae7iu6),
    .o(Aiwhu6));  // ../RTL/cortexm0ds_logic.v(4528)
  AL_MUX u2982 (
    .i0(W74iu6),
    .i1(Trgpw6[23]),
    .sel(Ae7iu6),
    .o(Thwhu6));  // ../RTL/cortexm0ds_logic.v(4529)
  AL_MUX u2983 (
    .i0(P74iu6),
    .i1(Trgpw6[22]),
    .sel(Ae7iu6),
    .o(Mhwhu6));  // ../RTL/cortexm0ds_logic.v(4530)
  AL_MUX u2984 (
    .i0(I74iu6),
    .i1(Trgpw6[21]),
    .sel(Ae7iu6),
    .o(Fhwhu6));  // ../RTL/cortexm0ds_logic.v(4531)
  AL_MUX u2985 (
    .i0(B74iu6),
    .i1(Trgpw6[20]),
    .sel(Ae7iu6),
    .o(Ygwhu6));  // ../RTL/cortexm0ds_logic.v(4532)
  AL_MUX u2986 (
    .i0(U64iu6),
    .i1(Trgpw6[19]),
    .sel(Ae7iu6),
    .o(Rgwhu6));  // ../RTL/cortexm0ds_logic.v(4533)
  AL_MUX u2987 (
    .i0(N64iu6),
    .i1(Trgpw6[18]),
    .sel(Ae7iu6),
    .o(Kgwhu6));  // ../RTL/cortexm0ds_logic.v(4534)
  AL_MUX u2988 (
    .i0(G64iu6),
    .i1(Trgpw6[17]),
    .sel(Ae7iu6),
    .o(Dgwhu6));  // ../RTL/cortexm0ds_logic.v(4535)
  AL_MUX u2989 (
    .i0(Z54iu6),
    .i1(Trgpw6[16]),
    .sel(Ae7iu6),
    .o(Wfwhu6));  // ../RTL/cortexm0ds_logic.v(4536)
  buf u299 (Vbgpw6[31], S0kbx6);  // ../RTL/cortexm0ds_logic.v(3092)
  AL_MUX u2990 (
    .i0(S54iu6),
    .i1(Trgpw6[15]),
    .sel(Ae7iu6),
    .o(Pfwhu6));  // ../RTL/cortexm0ds_logic.v(4537)
  AL_MUX u2991 (
    .i0(L54iu6),
    .i1(Trgpw6[14]),
    .sel(Ae7iu6),
    .o(Ifwhu6));  // ../RTL/cortexm0ds_logic.v(4538)
  AL_MUX u2992 (
    .i0(E54iu6),
    .i1(Trgpw6[13]),
    .sel(Ae7iu6),
    .o(Bfwhu6));  // ../RTL/cortexm0ds_logic.v(4539)
  AL_MUX u2993 (
    .i0(X44iu6),
    .i1(Trgpw6[12]),
    .sel(Ae7iu6),
    .o(Uewhu6));  // ../RTL/cortexm0ds_logic.v(4540)
  AL_MUX u2994 (
    .i0(Q44iu6),
    .i1(Trgpw6[11]),
    .sel(Ae7iu6),
    .o(Newhu6));  // ../RTL/cortexm0ds_logic.v(4541)
  AL_MUX u2995 (
    .i0(J44iu6),
    .i1(Trgpw6[10]),
    .sel(Ae7iu6),
    .o(Gewhu6));  // ../RTL/cortexm0ds_logic.v(4542)
  AL_MUX u2996 (
    .i0(Ym4iu6),
    .i1(Trgpw6[9]),
    .sel(Ae7iu6),
    .o(Zdwhu6));  // ../RTL/cortexm0ds_logic.v(4543)
  AL_MUX u2997 (
    .i0(Pl4iu6),
    .i1(Trgpw6[8]),
    .sel(Ae7iu6),
    .o(Sdwhu6));  // ../RTL/cortexm0ds_logic.v(4544)
  AL_MUX u2998 (
    .i0(Gk4iu6),
    .i1(Trgpw6[7]),
    .sel(Ae7iu6),
    .o(Ldwhu6));  // ../RTL/cortexm0ds_logic.v(4545)
  AL_MUX u2999 (
    .i0(Xi4iu6),
    .i1(Trgpw6[6]),
    .sel(Ae7iu6),
    .o(Edwhu6));  // ../RTL/cortexm0ds_logic.v(4546)
  buf u3 (R4gpw6[35], L8zax6);  // ../RTL/cortexm0ds_logic.v(2815)
  buf u30 (Gtgpw6[9], F7jbx6);  // ../RTL/cortexm0ds_logic.v(2375)
  buf u300 (K7hpw6[28], Nfgax6);  // ../RTL/cortexm0ds_logic.v(2366)
  AL_MUX u3000 (
    .i0(Oh4iu6),
    .i1(Trgpw6[5]),
    .sel(Ae7iu6),
    .o(Xcwhu6));  // ../RTL/cortexm0ds_logic.v(4547)
  AL_MUX u3001 (
    .i0(H34iu6),
    .i1(Trgpw6[4]),
    .sel(Ae7iu6),
    .o(Qcwhu6));  // ../RTL/cortexm0ds_logic.v(4548)
  AL_MUX u3002 (
    .i0(Df4iu6),
    .i1(Trgpw6[3]),
    .sel(Ae7iu6),
    .o(Jcwhu6));  // ../RTL/cortexm0ds_logic.v(4549)
  AL_MUX u3003 (
    .i0(T24iu6),
    .i1(Alhhu6),
    .sel(Ae7iu6),
    .o(Ccwhu6));  // ../RTL/cortexm0ds_logic.v(4550)
  and u3004 (n515, A2nhu6, Dw1iu6);  // ../RTL/cortexm0ds_logic.v(4551)
  not u3005 (Ae7iu6, n515);  // ../RTL/cortexm0ds_logic.v(4551)
  AL_MUX u3006 (
    .i0(Ud4iu6),
    .i1(Gtgpw6[2]),
    .sel(He7iu6),
    .o(Vbwhu6));  // ../RTL/cortexm0ds_logic.v(4552)
  AL_MUX u3007 (
    .i0(Lm1iu6),
    .i1(Engpw6[28]),
    .sel(He7iu6),
    .o(Obwhu6));  // ../RTL/cortexm0ds_logic.v(4553)
  AL_MUX u3008 (
    .i0(T94iu6),
    .i1(Engpw6[27]),
    .sel(He7iu6),
    .o(Hbwhu6));  // ../RTL/cortexm0ds_logic.v(4554)
  AL_MUX u3009 (
    .i0(F94iu6),
    .i1(Gtgpw6[28]),
    .sel(He7iu6),
    .o(Abwhu6));  // ../RTL/cortexm0ds_logic.v(4555)
  buf u301 (Yyfhu6, Sz3qw6);  // ../RTL/cortexm0ds_logic.v(2182)
  AL_MUX u3010 (
    .i0(Y84iu6),
    .i1(Gtgpw6[27]),
    .sel(He7iu6),
    .o(Tawhu6));  // ../RTL/cortexm0ds_logic.v(4556)
  AL_MUX u3011 (
    .i0(R84iu6),
    .i1(Gtgpw6[26]),
    .sel(He7iu6),
    .o(Mawhu6));  // ../RTL/cortexm0ds_logic.v(4557)
  AL_MUX u3012 (
    .i0(K84iu6),
    .i1(Gtgpw6[25]),
    .sel(He7iu6),
    .o(Fawhu6));  // ../RTL/cortexm0ds_logic.v(4558)
  AL_MUX u3013 (
    .i0(D84iu6),
    .i1(Gtgpw6[24]),
    .sel(He7iu6),
    .o(Y9whu6));  // ../RTL/cortexm0ds_logic.v(4559)
  AL_MUX u3014 (
    .i0(W74iu6),
    .i1(Gtgpw6[23]),
    .sel(He7iu6),
    .o(R9whu6));  // ../RTL/cortexm0ds_logic.v(4560)
  AL_MUX u3015 (
    .i0(P74iu6),
    .i1(Gtgpw6[22]),
    .sel(He7iu6),
    .o(K9whu6));  // ../RTL/cortexm0ds_logic.v(4561)
  AL_MUX u3016 (
    .i0(I74iu6),
    .i1(Gtgpw6[21]),
    .sel(He7iu6),
    .o(D9whu6));  // ../RTL/cortexm0ds_logic.v(4562)
  AL_MUX u3017 (
    .i0(B74iu6),
    .i1(Gtgpw6[20]),
    .sel(He7iu6),
    .o(W8whu6));  // ../RTL/cortexm0ds_logic.v(4563)
  AL_MUX u3018 (
    .i0(U64iu6),
    .i1(Gtgpw6[19]),
    .sel(He7iu6),
    .o(P8whu6));  // ../RTL/cortexm0ds_logic.v(4564)
  AL_MUX u3019 (
    .i0(N64iu6),
    .i1(Gtgpw6[18]),
    .sel(He7iu6),
    .o(I8whu6));  // ../RTL/cortexm0ds_logic.v(4565)
  buf u302 (vis_r2_o[17], Uyqax6);  // ../RTL/cortexm0ds_logic.v(2551)
  AL_MUX u3020 (
    .i0(G64iu6),
    .i1(Gtgpw6[17]),
    .sel(He7iu6),
    .o(B8whu6));  // ../RTL/cortexm0ds_logic.v(4566)
  AL_MUX u3021 (
    .i0(Z54iu6),
    .i1(Gtgpw6[16]),
    .sel(He7iu6),
    .o(U7whu6));  // ../RTL/cortexm0ds_logic.v(4567)
  AL_MUX u3022 (
    .i0(S54iu6),
    .i1(Gtgpw6[15]),
    .sel(He7iu6),
    .o(N7whu6));  // ../RTL/cortexm0ds_logic.v(4568)
  AL_MUX u3023 (
    .i0(L54iu6),
    .i1(Gtgpw6[14]),
    .sel(He7iu6),
    .o(G7whu6));  // ../RTL/cortexm0ds_logic.v(4569)
  AL_MUX u3024 (
    .i0(E54iu6),
    .i1(Gtgpw6[13]),
    .sel(He7iu6),
    .o(Z6whu6));  // ../RTL/cortexm0ds_logic.v(4570)
  AL_MUX u3025 (
    .i0(X44iu6),
    .i1(Gtgpw6[12]),
    .sel(He7iu6),
    .o(S6whu6));  // ../RTL/cortexm0ds_logic.v(4571)
  AL_MUX u3026 (
    .i0(Q44iu6),
    .i1(Gtgpw6[11]),
    .sel(He7iu6),
    .o(L6whu6));  // ../RTL/cortexm0ds_logic.v(4572)
  AL_MUX u3027 (
    .i0(J44iu6),
    .i1(Gtgpw6[10]),
    .sel(He7iu6),
    .o(E6whu6));  // ../RTL/cortexm0ds_logic.v(4573)
  AL_MUX u3028 (
    .i0(Ym4iu6),
    .i1(Gtgpw6[9]),
    .sel(He7iu6),
    .o(X5whu6));  // ../RTL/cortexm0ds_logic.v(4574)
  AL_MUX u3029 (
    .i0(Pl4iu6),
    .i1(Gtgpw6[8]),
    .sel(He7iu6),
    .o(Q5whu6));  // ../RTL/cortexm0ds_logic.v(4575)
  buf u303 (vis_r0_o[31], Ehnpw6);  // ../RTL/cortexm0ds_logic.v(1875)
  AL_MUX u3030 (
    .i0(Gk4iu6),
    .i1(Gtgpw6[7]),
    .sel(He7iu6),
    .o(J5whu6));  // ../RTL/cortexm0ds_logic.v(4576)
  AL_MUX u3031 (
    .i0(Xi4iu6),
    .i1(Gtgpw6[6]),
    .sel(He7iu6),
    .o(C5whu6));  // ../RTL/cortexm0ds_logic.v(4577)
  AL_MUX u3032 (
    .i0(Oh4iu6),
    .i1(Gtgpw6[5]),
    .sel(He7iu6),
    .o(V4whu6));  // ../RTL/cortexm0ds_logic.v(4578)
  AL_MUX u3033 (
    .i0(H34iu6),
    .i1(Gtgpw6[4]),
    .sel(He7iu6),
    .o(O4whu6));  // ../RTL/cortexm0ds_logic.v(4579)
  AL_MUX u3034 (
    .i0(Df4iu6),
    .i1(Gtgpw6[3]),
    .sel(He7iu6),
    .o(H4whu6));  // ../RTL/cortexm0ds_logic.v(4580)
  AL_MUX u3035 (
    .i0(T24iu6),
    .i1(Smhhu6),
    .sel(He7iu6),
    .o(A4whu6));  // ../RTL/cortexm0ds_logic.v(4581)
  and u3036 (n516, A2nhu6, Cs1iu6);  // ../RTL/cortexm0ds_logic.v(4582)
  not u3037 (He7iu6, n516);  // ../RTL/cortexm0ds_logic.v(4582)
  AL_MUX u3038 (
    .i0(Kohhu6),
    .i1(T24iu6),
    .sel(Oe7iu6),
    .o(T3whu6));  // ../RTL/cortexm0ds_logic.v(4583)
  and u3039 (Oe7iu6, Ve7iu6, A2nhu6);  // ../RTL/cortexm0ds_logic.v(4584)
  buf u304 (Shhpw6[18], Gwwpw6);  // ../RTL/cortexm0ds_logic.v(1941)
  AL_MUX u3040 (
    .i0(T24iu6),
    .i1(Aygpw6[0]),
    .sel(Cf7iu6),
    .o(M3whu6));  // ../RTL/cortexm0ds_logic.v(4585)
  AL_MUX u3041 (
    .i0(H34iu6),
    .i1(Aygpw6[4]),
    .sel(Cf7iu6),
    .o(F3whu6));  // ../RTL/cortexm0ds_logic.v(4586)
  AL_MUX u3042 (
    .i0(Df4iu6),
    .i1(Aygpw6[3]),
    .sel(Cf7iu6),
    .o(Y2whu6));  // ../RTL/cortexm0ds_logic.v(4587)
  AL_MUX u3043 (
    .i0(Ud4iu6),
    .i1(Aygpw6[2]),
    .sel(Cf7iu6),
    .o(R2whu6));  // ../RTL/cortexm0ds_logic.v(4588)
  AL_MUX u3044 (
    .i0(O34iu6),
    .i1(Aygpw6[1]),
    .sel(Cf7iu6),
    .o(K2whu6));  // ../RTL/cortexm0ds_logic.v(4589)
  and u3045 (n517, Jf7iu6, A2nhu6);  // ../RTL/cortexm0ds_logic.v(4590)
  not u3046 (Cf7iu6, n517);  // ../RTL/cortexm0ds_logic.v(4590)
  AL_MUX u3047 (
    .i0(T24iu6),
    .i1(Pzgpw6[0]),
    .sel(Qf7iu6),
    .o(D2whu6));  // ../RTL/cortexm0ds_logic.v(4591)
  AL_MUX u3048 (
    .i0(Lm1iu6),
    .i1(E1hpw6[31]),
    .sel(Qf7iu6),
    .o(W1whu6));  // ../RTL/cortexm0ds_logic.v(4592)
  AL_MUX u3049 (
    .i0(T94iu6),
    .i1(E1hpw6[30]),
    .sel(Qf7iu6),
    .o(P1whu6));  // ../RTL/cortexm0ds_logic.v(4593)
  buf u305 (vis_r12_o[20], Egtax6);  // ../RTL/cortexm0ds_logic.v(2599)
  AL_MUX u3050 (
    .i0(M94iu6),
    .i1(E1hpw6[29]),
    .sel(Qf7iu6),
    .o(I1whu6));  // ../RTL/cortexm0ds_logic.v(4594)
  AL_MUX u3051 (
    .i0(F94iu6),
    .i1(E1hpw6[28]),
    .sel(Qf7iu6),
    .o(B1whu6));  // ../RTL/cortexm0ds_logic.v(4595)
  AL_MUX u3052 (
    .i0(Y84iu6),
    .i1(E1hpw6[27]),
    .sel(Qf7iu6),
    .o(U0whu6));  // ../RTL/cortexm0ds_logic.v(4596)
  AL_MUX u3053 (
    .i0(R84iu6),
    .i1(E1hpw6[26]),
    .sel(Qf7iu6),
    .o(N0whu6));  // ../RTL/cortexm0ds_logic.v(4597)
  AL_MUX u3054 (
    .i0(K84iu6),
    .i1(E1hpw6[25]),
    .sel(Qf7iu6),
    .o(G0whu6));  // ../RTL/cortexm0ds_logic.v(4598)
  AL_MUX u3055 (
    .i0(D84iu6),
    .i1(E1hpw6[24]),
    .sel(Qf7iu6),
    .o(Zzvhu6));  // ../RTL/cortexm0ds_logic.v(4599)
  AL_MUX u3056 (
    .i0(W74iu6),
    .i1(E1hpw6[23]),
    .sel(Qf7iu6),
    .o(Szvhu6));  // ../RTL/cortexm0ds_logic.v(4600)
  AL_MUX u3057 (
    .i0(P74iu6),
    .i1(E1hpw6[22]),
    .sel(Qf7iu6),
    .o(Lzvhu6));  // ../RTL/cortexm0ds_logic.v(4601)
  AL_MUX u3058 (
    .i0(I74iu6),
    .i1(E1hpw6[21]),
    .sel(Qf7iu6),
    .o(Ezvhu6));  // ../RTL/cortexm0ds_logic.v(4602)
  AL_MUX u3059 (
    .i0(B74iu6),
    .i1(E1hpw6[20]),
    .sel(Qf7iu6),
    .o(Xyvhu6));  // ../RTL/cortexm0ds_logic.v(4603)
  buf u306 (Aphpw6[1], Ksgax6);  // ../RTL/cortexm0ds_logic.v(2381)
  AL_MUX u3060 (
    .i0(U64iu6),
    .i1(E1hpw6[19]),
    .sel(Qf7iu6),
    .o(Qyvhu6));  // ../RTL/cortexm0ds_logic.v(4604)
  AL_MUX u3061 (
    .i0(N64iu6),
    .i1(E1hpw6[18]),
    .sel(Qf7iu6),
    .o(Jyvhu6));  // ../RTL/cortexm0ds_logic.v(4605)
  AL_MUX u3062 (
    .i0(G64iu6),
    .i1(E1hpw6[17]),
    .sel(Qf7iu6),
    .o(Cyvhu6));  // ../RTL/cortexm0ds_logic.v(4606)
  AL_MUX u3063 (
    .i0(Z54iu6),
    .i1(E1hpw6[16]),
    .sel(Qf7iu6),
    .o(Vxvhu6));  // ../RTL/cortexm0ds_logic.v(4607)
  AL_MUX u3064 (
    .i0(S54iu6),
    .i1(E1hpw6[15]),
    .sel(Qf7iu6),
    .o(Oxvhu6));  // ../RTL/cortexm0ds_logic.v(4608)
  AL_MUX u3065 (
    .i0(L54iu6),
    .i1(E1hpw6[14]),
    .sel(Qf7iu6),
    .o(Hxvhu6));  // ../RTL/cortexm0ds_logic.v(4609)
  AL_MUX u3066 (
    .i0(E54iu6),
    .i1(E1hpw6[13]),
    .sel(Qf7iu6),
    .o(Axvhu6));  // ../RTL/cortexm0ds_logic.v(4610)
  AL_MUX u3067 (
    .i0(X44iu6),
    .i1(E1hpw6[12]),
    .sel(Qf7iu6),
    .o(Twvhu6));  // ../RTL/cortexm0ds_logic.v(4611)
  AL_MUX u3068 (
    .i0(Q44iu6),
    .i1(E1hpw6[11]),
    .sel(Qf7iu6),
    .o(Mwvhu6));  // ../RTL/cortexm0ds_logic.v(4612)
  AL_MUX u3069 (
    .i0(J44iu6),
    .i1(E1hpw6[10]),
    .sel(Qf7iu6),
    .o(Fwvhu6));  // ../RTL/cortexm0ds_logic.v(4613)
  buf u307 (Zlghu6, F17ax6);  // ../RTL/cortexm0ds_logic.v(2192)
  AL_MUX u3070 (
    .i0(Ym4iu6),
    .i1(E1hpw6[9]),
    .sel(Qf7iu6),
    .o(Yvvhu6));  // ../RTL/cortexm0ds_logic.v(4614)
  AL_MUX u3071 (
    .i0(Pl4iu6),
    .i1(E1hpw6[8]),
    .sel(Qf7iu6),
    .o(Rvvhu6));  // ../RTL/cortexm0ds_logic.v(4615)
  AL_MUX u3072 (
    .i0(Gk4iu6),
    .i1(E1hpw6[7]),
    .sel(Qf7iu6),
    .o(Kvvhu6));  // ../RTL/cortexm0ds_logic.v(4616)
  AL_MUX u3073 (
    .i0(Xi4iu6),
    .i1(E1hpw6[6]),
    .sel(Qf7iu6),
    .o(Dvvhu6));  // ../RTL/cortexm0ds_logic.v(4617)
  AL_MUX u3074 (
    .i0(Oh4iu6),
    .i1(E1hpw6[5]),
    .sel(Qf7iu6),
    .o(Wuvhu6));  // ../RTL/cortexm0ds_logic.v(4618)
  AL_MUX u3075 (
    .i0(H34iu6),
    .i1(E1hpw6[4]),
    .sel(Qf7iu6),
    .o(Puvhu6));  // ../RTL/cortexm0ds_logic.v(4619)
  AL_MUX u3076 (
    .i0(Df4iu6),
    .i1(E1hpw6[3]),
    .sel(Qf7iu6),
    .o(Iuvhu6));  // ../RTL/cortexm0ds_logic.v(4620)
  AL_MUX u3077 (
    .i0(Ud4iu6),
    .i1(E1hpw6[2]),
    .sel(Qf7iu6),
    .o(Buvhu6));  // ../RTL/cortexm0ds_logic.v(4621)
  AL_MUX u3078 (
    .i0(O34iu6),
    .i1(Pzgpw6[1]),
    .sel(Qf7iu6),
    .o(Utvhu6));  // ../RTL/cortexm0ds_logic.v(4622)
  and u3079 (n518, A2nhu6, Zt1iu6);  // ../RTL/cortexm0ds_logic.v(4623)
  buf u308 (vis_r1_o[21], I1qpw6);  // ../RTL/cortexm0ds_logic.v(1876)
  not u3080 (Qf7iu6, n518);  // ../RTL/cortexm0ds_logic.v(4623)
  AL_MUX u3081 (
    .i0(T24iu6),
    .i1(R2hpw6[0]),
    .sel(Xf7iu6),
    .o(Ntvhu6));  // ../RTL/cortexm0ds_logic.v(4624)
  AL_MUX u3082 (
    .i0(Ud4iu6),
    .i1(R2hpw6[2]),
    .sel(Xf7iu6),
    .o(Gtvhu6));  // ../RTL/cortexm0ds_logic.v(4625)
  AL_MUX u3083 (
    .i0(O34iu6),
    .i1(R2hpw6[1]),
    .sel(Xf7iu6),
    .o(Zsvhu6));  // ../RTL/cortexm0ds_logic.v(4626)
  and u3084 (n519, Eg7iu6, A2nhu6);  // ../RTL/cortexm0ds_logic.v(4627)
  not u3085 (Xf7iu6, n519);  // ../RTL/cortexm0ds_logic.v(4627)
  AL_MUX u3086 (
    .i0(T24iu6),
    .i1(G4hpw6[0]),
    .sel(Lg7iu6),
    .o(Ssvhu6));  // ../RTL/cortexm0ds_logic.v(4628)
  AL_MUX u3087 (
    .i0(H34iu6),
    .i1(G4hpw6[4]),
    .sel(Lg7iu6),
    .o(Lsvhu6));  // ../RTL/cortexm0ds_logic.v(4629)
  AL_MUX u3088 (
    .i0(Df4iu6),
    .i1(G4hpw6[3]),
    .sel(Lg7iu6),
    .o(Esvhu6));  // ../RTL/cortexm0ds_logic.v(4630)
  AL_MUX u3089 (
    .i0(Ud4iu6),
    .i1(G4hpw6[2]),
    .sel(Lg7iu6),
    .o(Xrvhu6));  // ../RTL/cortexm0ds_logic.v(4631)
  buf u309 (vis_psp_o[2], Ezypw6);  // ../RTL/cortexm0ds_logic.v(2085)
  AL_MUX u3090 (
    .i0(O34iu6),
    .i1(G4hpw6[1]),
    .sel(Lg7iu6),
    .o(Qrvhu6));  // ../RTL/cortexm0ds_logic.v(4632)
  and u3091 (n520, Sg7iu6, A2nhu6);  // ../RTL/cortexm0ds_logic.v(4633)
  not u3092 (Lg7iu6, n520);  // ../RTL/cortexm0ds_logic.v(4633)
  AL_MUX u3093 (
    .i0(T24iu6),
    .i1(V5hpw6[0]),
    .sel(Zg7iu6),
    .o(Jrvhu6));  // ../RTL/cortexm0ds_logic.v(4634)
  AL_MUX u3094 (
    .i0(Lm1iu6),
    .i1(K7hpw6[31]),
    .sel(Zg7iu6),
    .o(Crvhu6));  // ../RTL/cortexm0ds_logic.v(4635)
  AL_MUX u3095 (
    .i0(T94iu6),
    .i1(K7hpw6[30]),
    .sel(Zg7iu6),
    .o(Vqvhu6));  // ../RTL/cortexm0ds_logic.v(4636)
  AL_MUX u3096 (
    .i0(M94iu6),
    .i1(K7hpw6[29]),
    .sel(Zg7iu6),
    .o(Oqvhu6));  // ../RTL/cortexm0ds_logic.v(4637)
  AL_MUX u3097 (
    .i0(F94iu6),
    .i1(K7hpw6[28]),
    .sel(Zg7iu6),
    .o(Hqvhu6));  // ../RTL/cortexm0ds_logic.v(4638)
  AL_MUX u3098 (
    .i0(Y84iu6),
    .i1(K7hpw6[27]),
    .sel(Zg7iu6),
    .o(Aqvhu6));  // ../RTL/cortexm0ds_logic.v(4639)
  AL_MUX u3099 (
    .i0(R84iu6),
    .i1(K7hpw6[26]),
    .sel(Zg7iu6),
    .o(Tpvhu6));  // ../RTL/cortexm0ds_logic.v(4640)
  buf u31 (Uthpw6[8], M81qw6);  // ../RTL/cortexm0ds_logic.v(1882)
  buf u310 (vis_r4_o[8], Uhvax6);  // ../RTL/cortexm0ds_logic.v(2626)
  AL_MUX u3100 (
    .i0(K84iu6),
    .i1(K7hpw6[25]),
    .sel(Zg7iu6),
    .o(Mpvhu6));  // ../RTL/cortexm0ds_logic.v(4641)
  AL_MUX u3101 (
    .i0(D84iu6),
    .i1(K7hpw6[24]),
    .sel(Zg7iu6),
    .o(Fpvhu6));  // ../RTL/cortexm0ds_logic.v(4642)
  AL_MUX u3102 (
    .i0(W74iu6),
    .i1(K7hpw6[23]),
    .sel(Zg7iu6),
    .o(Yovhu6));  // ../RTL/cortexm0ds_logic.v(4643)
  AL_MUX u3103 (
    .i0(P74iu6),
    .i1(K7hpw6[22]),
    .sel(Zg7iu6),
    .o(Rovhu6));  // ../RTL/cortexm0ds_logic.v(4644)
  AL_MUX u3104 (
    .i0(I74iu6),
    .i1(K7hpw6[21]),
    .sel(Zg7iu6),
    .o(Kovhu6));  // ../RTL/cortexm0ds_logic.v(4645)
  AL_MUX u3105 (
    .i0(B74iu6),
    .i1(K7hpw6[20]),
    .sel(Zg7iu6),
    .o(Dovhu6));  // ../RTL/cortexm0ds_logic.v(4646)
  AL_MUX u3106 (
    .i0(U64iu6),
    .i1(K7hpw6[19]),
    .sel(Zg7iu6),
    .o(Wnvhu6));  // ../RTL/cortexm0ds_logic.v(4647)
  AL_MUX u3107 (
    .i0(N64iu6),
    .i1(K7hpw6[18]),
    .sel(Zg7iu6),
    .o(Pnvhu6));  // ../RTL/cortexm0ds_logic.v(4648)
  AL_MUX u3108 (
    .i0(G64iu6),
    .i1(K7hpw6[17]),
    .sel(Zg7iu6),
    .o(Invhu6));  // ../RTL/cortexm0ds_logic.v(4649)
  AL_MUX u3109 (
    .i0(Z54iu6),
    .i1(K7hpw6[16]),
    .sel(Zg7iu6),
    .o(Bnvhu6));  // ../RTL/cortexm0ds_logic.v(4650)
  buf u311 (vis_r14_o[5], Q9nax6);  // ../RTL/cortexm0ds_logic.v(2497)
  AL_MUX u3110 (
    .i0(S54iu6),
    .i1(K7hpw6[15]),
    .sel(Zg7iu6),
    .o(Umvhu6));  // ../RTL/cortexm0ds_logic.v(4651)
  AL_MUX u3111 (
    .i0(L54iu6),
    .i1(K7hpw6[14]),
    .sel(Zg7iu6),
    .o(Nmvhu6));  // ../RTL/cortexm0ds_logic.v(4652)
  AL_MUX u3112 (
    .i0(E54iu6),
    .i1(K7hpw6[13]),
    .sel(Zg7iu6),
    .o(Gmvhu6));  // ../RTL/cortexm0ds_logic.v(4653)
  AL_MUX u3113 (
    .i0(X44iu6),
    .i1(K7hpw6[12]),
    .sel(Zg7iu6),
    .o(Zlvhu6));  // ../RTL/cortexm0ds_logic.v(4654)
  AL_MUX u3114 (
    .i0(Q44iu6),
    .i1(K7hpw6[11]),
    .sel(Zg7iu6),
    .o(Slvhu6));  // ../RTL/cortexm0ds_logic.v(4655)
  AL_MUX u3115 (
    .i0(J44iu6),
    .i1(K7hpw6[10]),
    .sel(Zg7iu6),
    .o(Llvhu6));  // ../RTL/cortexm0ds_logic.v(4656)
  AL_MUX u3116 (
    .i0(Ym4iu6),
    .i1(K7hpw6[9]),
    .sel(Zg7iu6),
    .o(Elvhu6));  // ../RTL/cortexm0ds_logic.v(4657)
  AL_MUX u3117 (
    .i0(Pl4iu6),
    .i1(K7hpw6[8]),
    .sel(Zg7iu6),
    .o(Xkvhu6));  // ../RTL/cortexm0ds_logic.v(4658)
  AL_MUX u3118 (
    .i0(Gk4iu6),
    .i1(K7hpw6[7]),
    .sel(Zg7iu6),
    .o(Qkvhu6));  // ../RTL/cortexm0ds_logic.v(4659)
  AL_MUX u3119 (
    .i0(Xi4iu6),
    .i1(K7hpw6[6]),
    .sel(Zg7iu6),
    .o(Jkvhu6));  // ../RTL/cortexm0ds_logic.v(4660)
  buf u312 (vis_r8_o[14], O6sax6);  // ../RTL/cortexm0ds_logic.v(2579)
  AL_MUX u3120 (
    .i0(Oh4iu6),
    .i1(K7hpw6[5]),
    .sel(Zg7iu6),
    .o(Ckvhu6));  // ../RTL/cortexm0ds_logic.v(4661)
  AL_MUX u3121 (
    .i0(H34iu6),
    .i1(K7hpw6[4]),
    .sel(Zg7iu6),
    .o(Vjvhu6));  // ../RTL/cortexm0ds_logic.v(4662)
  AL_MUX u3122 (
    .i0(Df4iu6),
    .i1(K7hpw6[3]),
    .sel(Zg7iu6),
    .o(Ojvhu6));  // ../RTL/cortexm0ds_logic.v(4663)
  AL_MUX u3123 (
    .i0(Ud4iu6),
    .i1(K7hpw6[2]),
    .sel(Zg7iu6),
    .o(Hjvhu6));  // ../RTL/cortexm0ds_logic.v(4664)
  AL_MUX u3124 (
    .i0(O34iu6),
    .i1(V5hpw6[1]),
    .sel(Zg7iu6),
    .o(Ajvhu6));  // ../RTL/cortexm0ds_logic.v(4665)
  and u3125 (n521, A2nhu6, Kw1iu6);  // ../RTL/cortexm0ds_logic.v(4666)
  not u3126 (Zg7iu6, n521);  // ../RTL/cortexm0ds_logic.v(4666)
  and u3127 (n522, Gh7iu6, Nh7iu6);  // ../RTL/cortexm0ds_logic.v(4667)
  not u3128 (Tivhu6, n522);  // ../RTL/cortexm0ds_logic.v(4667)
  or u3129 (Nh7iu6, Uh7iu6, HREADY);  // ../RTL/cortexm0ds_logic.v(4668)
  buf u313 (Vbgpw6[8], C30bx6);  // ../RTL/cortexm0ds_logic.v(3092)
  and u3130 (Gh7iu6, Bi7iu6, Ii7iu6);  // ../RTL/cortexm0ds_logic.v(4669)
  and u3131 (n523, Pi7iu6, Wi7iu6);  // ../RTL/cortexm0ds_logic.v(4670)
  not u3132 (Bi7iu6, n523);  // ../RTL/cortexm0ds_logic.v(4670)
  and u3133 (Mivhu6, Dj7iu6, Kj7iu6);  // ../RTL/cortexm0ds_logic.v(4671)
  and u3134 (Kj7iu6, Rj7iu6, Yj7iu6);  // ../RTL/cortexm0ds_logic.v(4672)
  and u3135 (n524, Xudpw6, Fk7iu6);  // ../RTL/cortexm0ds_logic.v(4673)
  not u3136 (Rj7iu6, n524);  // ../RTL/cortexm0ds_logic.v(4673)
  and u3137 (Dj7iu6, IRQ[0], Mk7iu6);  // ../RTL/cortexm0ds_logic.v(4674)
  and u3138 (n525, Tk7iu6, Al7iu6);  // ../RTL/cortexm0ds_logic.v(4675)
  not u3139 (Mk7iu6, n525);  // ../RTL/cortexm0ds_logic.v(4675)
  buf u314 (vis_r14_o[23], Szmax6);  // ../RTL/cortexm0ds_logic.v(2497)
  or u3140 (Al7iu6, Qg6iu6, Hl7iu6);  // ../RTL/cortexm0ds_logic.v(4676)
  or u3141 (Fivhu6, Ol7iu6, Vl7iu6);  // ../RTL/cortexm0ds_logic.v(4677)
  and u3142 (Vl7iu6, Ivfhu6, Cm7iu6);  // ../RTL/cortexm0ds_logic.v(4678)
  and u3143 (n526, Jm7iu6, Qm7iu6);  // ../RTL/cortexm0ds_logic.v(4679)
  not u3144 (Cm7iu6, n526);  // ../RTL/cortexm0ds_logic.v(4679)
  and u3145 (n527, Gc5iu6, Xm7iu6);  // ../RTL/cortexm0ds_logic.v(4680)
  not u3146 (Qm7iu6, n527);  // ../RTL/cortexm0ds_logic.v(4680)
  or u3147 (Xm7iu6, Sb5iu6, Eh6iu6);  // ../RTL/cortexm0ds_logic.v(4681)
  or u3148 (Yhvhu6, En7iu6, Ln7iu6);  // ../RTL/cortexm0ds_logic.v(4682)
  AL_MUX u3149 (
    .i0(Ppfpw6[15]),
    .i1(Sn7iu6),
    .sel(Zn7iu6),
    .o(En7iu6));  // ../RTL/cortexm0ds_logic.v(4683)
  buf u315 (vis_r4_o[21], Vvuax6);  // ../RTL/cortexm0ds_logic.v(2626)
  and u3150 (Sn7iu6, HRDATA[15], Go7iu6);  // ../RTL/cortexm0ds_logic.v(4684)
  and u3151 (n528, No7iu6, Uo7iu6);  // ../RTL/cortexm0ds_logic.v(4685)
  not u3152 (Rhvhu6, n528);  // ../RTL/cortexm0ds_logic.v(4685)
  and u3153 (Uo7iu6, Bp7iu6, Ip7iu6);  // ../RTL/cortexm0ds_logic.v(4686)
  and u3154 (n529, Pp7iu6, HRDATA[15]);  // ../RTL/cortexm0ds_logic.v(4687)
  not u3155 (Ip7iu6, n529);  // ../RTL/cortexm0ds_logic.v(4687)
  and u3156 (Bp7iu6, Wp7iu6, Dq7iu6);  // ../RTL/cortexm0ds_logic.v(4688)
  and u3157 (n530, Hrfpw6[15], Uy4iu6);  // ../RTL/cortexm0ds_logic.v(4689)
  not u3158 (Dq7iu6, n530);  // ../RTL/cortexm0ds_logic.v(4689)
  and u3159 (n531, Kq7iu6, HRDATA[31]);  // ../RTL/cortexm0ds_logic.v(4690)
  buf u316 (vis_r14_o[18], Nvnax6);  // ../RTL/cortexm0ds_logic.v(2497)
  not u3160 (Wp7iu6, n531);  // ../RTL/cortexm0ds_logic.v(4690)
  and u3161 (No7iu6, Rq7iu6, Yq7iu6);  // ../RTL/cortexm0ds_logic.v(4691)
  and u3162 (n532, Fr7iu6, Z54iu6);  // ../RTL/cortexm0ds_logic.v(4692)
  not u3163 (Yq7iu6, n532);  // ../RTL/cortexm0ds_logic.v(4692)
  and u3164 (Rq7iu6, Mr7iu6, Tr7iu6);  // ../RTL/cortexm0ds_logic.v(4693)
  and u3165 (n533, Ppfpw6[15], A25iu6);  // ../RTL/cortexm0ds_logic.v(4694)
  not u3166 (Tr7iu6, n533);  // ../RTL/cortexm0ds_logic.v(4694)
  and u3167 (n534, R05iu6, D7fpw6[15]);  // ../RTL/cortexm0ds_logic.v(4695)
  not u3168 (Mr7iu6, n534);  // ../RTL/cortexm0ds_logic.v(4695)
  not u3169 (Khvhu6, As7iu6);  // ../RTL/cortexm0ds_logic.v(4696)
  buf u317 (vis_r8_o[27], Mlmpw6);  // ../RTL/cortexm0ds_logic.v(2579)
  AL_MUX u3170 (
    .i0(Hs7iu6),
    .i1(Os7iu6),
    .sel(HREADY),
    .o(As7iu6));  // ../RTL/cortexm0ds_logic.v(4697)
  and u3171 (n535, Vs7iu6, Ct7iu6);  // ../RTL/cortexm0ds_logic.v(4698)
  not u3172 (Os7iu6, n535);  // ../RTL/cortexm0ds_logic.v(4698)
  and u3173 (n536, Jt7iu6, Qt7iu6);  // ../RTL/cortexm0ds_logic.v(4699)
  not u3174 (Ct7iu6, n536);  // ../RTL/cortexm0ds_logic.v(4699)
  and u3175 (Qt7iu6, Xt7iu6, Eu7iu6);  // ../RTL/cortexm0ds_logic.v(4700)
  and u3176 (n537, Lu7iu6, Rthhu6);  // ../RTL/cortexm0ds_logic.v(4701)
  not u3177 (Eu7iu6, n537);  // ../RTL/cortexm0ds_logic.v(4701)
  and u3178 (Lu7iu6, Smhhu6, Engpw6[28]);  // ../RTL/cortexm0ds_logic.v(4702)
  and u3179 (n538, Su7iu6, Kshhu6);  // ../RTL/cortexm0ds_logic.v(4703)
  buf u318 (Hbhhu6, Fm7ax6);  // ../RTL/cortexm0ds_logic.v(2203)
  not u3180 (Xt7iu6, n538);  // ../RTL/cortexm0ds_logic.v(4703)
  and u3181 (Su7iu6, Alhhu6, Plgpw6[28]);  // ../RTL/cortexm0ds_logic.v(4704)
  and u3182 (Jt7iu6, Zu7iu6, Gv7iu6);  // ../RTL/cortexm0ds_logic.v(4705)
  and u3183 (n539, Nv7iu6, Drhhu6);  // ../RTL/cortexm0ds_logic.v(4706)
  not u3184 (Gv7iu6, n539);  // ../RTL/cortexm0ds_logic.v(4706)
  and u3185 (Nv7iu6, Ijhhu6, Akgpw6[28]);  // ../RTL/cortexm0ds_logic.v(4707)
  and u3186 (n540, Uv7iu6, Wphhu6);  // ../RTL/cortexm0ds_logic.v(4708)
  not u3187 (Zu7iu6, n540);  // ../RTL/cortexm0ds_logic.v(4708)
  and u3188 (Uv7iu6, Qhhhu6, Ligpw6[28]);  // ../RTL/cortexm0ds_logic.v(4709)
  not u3189 (Dhvhu6, Bw7iu6);  // ../RTL/cortexm0ds_logic.v(4710)
  buf u319 (Vbgpw6[22], B3gbx6);  // ../RTL/cortexm0ds_logic.v(3092)
  AL_MUX u3190 (
    .i0(Svdpw6),
    .i1(Iw7iu6),
    .sel(HREADY),
    .o(Bw7iu6));  // ../RTL/cortexm0ds_logic.v(4711)
  and u3191 (n541, Vs7iu6, Pw7iu6);  // ../RTL/cortexm0ds_logic.v(4712)
  not u3192 (Iw7iu6, n541);  // ../RTL/cortexm0ds_logic.v(4712)
  and u3193 (n542, Ww7iu6, Dx7iu6);  // ../RTL/cortexm0ds_logic.v(4713)
  not u3194 (Pw7iu6, n542);  // ../RTL/cortexm0ds_logic.v(4713)
  and u3195 (Dx7iu6, Kx7iu6, Rx7iu6);  // ../RTL/cortexm0ds_logic.v(4714)
  and u3196 (n543, Yx7iu6, Rthhu6);  // ../RTL/cortexm0ds_logic.v(4715)
  not u3197 (Rx7iu6, n543);  // ../RTL/cortexm0ds_logic.v(4715)
  and u3198 (Yx7iu6, Smhhu6, Engpw6[27]);  // ../RTL/cortexm0ds_logic.v(4716)
  and u3199 (n544, Fy7iu6, Kshhu6);  // ../RTL/cortexm0ds_logic.v(4717)
  buf u32 (Ligpw6[28], Bcgax6);  // ../RTL/cortexm0ds_logic.v(2371)
  buf u320 (Ftghu6, Lp7ax6);  // ../RTL/cortexm0ds_logic.v(2205)
  not u3200 (Kx7iu6, n544);  // ../RTL/cortexm0ds_logic.v(4717)
  and u3201 (Fy7iu6, Alhhu6, Plgpw6[27]);  // ../RTL/cortexm0ds_logic.v(4718)
  and u3202 (Ww7iu6, My7iu6, Ty7iu6);  // ../RTL/cortexm0ds_logic.v(4719)
  and u3203 (n545, Az7iu6, Drhhu6);  // ../RTL/cortexm0ds_logic.v(4720)
  not u3204 (Ty7iu6, n545);  // ../RTL/cortexm0ds_logic.v(4720)
  and u3205 (Az7iu6, Ijhhu6, Akgpw6[27]);  // ../RTL/cortexm0ds_logic.v(4721)
  and u3206 (n546, Hz7iu6, Wphhu6);  // ../RTL/cortexm0ds_logic.v(4722)
  not u3207 (My7iu6, n546);  // ../RTL/cortexm0ds_logic.v(4722)
  and u3208 (Hz7iu6, Qhhhu6, Ligpw6[27]);  // ../RTL/cortexm0ds_logic.v(4723)
  and u3209 (Vs7iu6, Oz7iu6, Vz7iu6);  // ../RTL/cortexm0ds_logic.v(4724)
  buf u321 (Jshpw6[25], Q2ibx6);  // ../RTL/cortexm0ds_logic.v(2372)
  or u3210 (n547, C08iu6, Dx0iu6);  // ../RTL/cortexm0ds_logic.v(4725)
  not u3211 (Vz7iu6, n547);  // ../RTL/cortexm0ds_logic.v(4725)
  and u3212 (n548, Jehhu6, J08iu6);  // ../RTL/cortexm0ds_logic.v(4726)
  not u3213 (C08iu6, n548);  // ../RTL/cortexm0ds_logic.v(4726)
  and u3214 (n549, Q08iu6, X08iu6);  // ../RTL/cortexm0ds_logic.v(4727)
  not u3215 (J08iu6, n549);  // ../RTL/cortexm0ds_logic.v(4727)
  and u3216 (n550, E18iu6, L18iu6);  // ../RTL/cortexm0ds_logic.v(4728)
  not u3217 (X08iu6, n550);  // ../RTL/cortexm0ds_logic.v(4728)
  and u3218 (E18iu6, S18iu6, Z18iu6);  // ../RTL/cortexm0ds_logic.v(4729)
  or u3219 (n551, G28iu6, Ef1iu6);  // ../RTL/cortexm0ds_logic.v(4730)
  buf u322 (Pzgpw6[1], Xwaax6);  // ../RTL/cortexm0ds_logic.v(2266)
  not u3220 (Oz7iu6, n551);  // ../RTL/cortexm0ds_logic.v(4730)
  or u3221 (G28iu6, N28iu6, Rx0iu6);  // ../RTL/cortexm0ds_logic.v(4731)
  not u3222 (N28iu6, Kohhu6);  // ../RTL/cortexm0ds_logic.v(4732)
  and u3223 (n552, U28iu6, B38iu6);  // ../RTL/cortexm0ds_logic.v(4733)
  not u3224 (Wgvhu6, n552);  // ../RTL/cortexm0ds_logic.v(4733)
  and u3225 (B38iu6, I38iu6, P38iu6);  // ../RTL/cortexm0ds_logic.v(4734)
  and u3226 (n553, HRDATA[13], Pp7iu6);  // ../RTL/cortexm0ds_logic.v(4735)
  not u3227 (P38iu6, n553);  // ../RTL/cortexm0ds_logic.v(4735)
  and u3228 (I38iu6, W38iu6, D48iu6);  // ../RTL/cortexm0ds_logic.v(4736)
  and u3229 (n554, Hrfpw6[13], Uy4iu6);  // ../RTL/cortexm0ds_logic.v(4737)
  buf u323 (G4hpw6[4], Lbbax6);  // ../RTL/cortexm0ds_logic.v(2274)
  not u3230 (D48iu6, n554);  // ../RTL/cortexm0ds_logic.v(4737)
  and u3231 (n555, HRDATA[29], Kq7iu6);  // ../RTL/cortexm0ds_logic.v(4738)
  not u3232 (W38iu6, n555);  // ../RTL/cortexm0ds_logic.v(4738)
  and u3233 (U28iu6, K48iu6, R48iu6);  // ../RTL/cortexm0ds_logic.v(4739)
  and u3234 (n556, A25iu6, Ppfpw6[13]);  // ../RTL/cortexm0ds_logic.v(4740)
  not u3235 (R48iu6, n556);  // ../RTL/cortexm0ds_logic.v(4740)
  and u3236 (n557, R05iu6, D7fpw6[13]);  // ../RTL/cortexm0ds_logic.v(4741)
  not u3237 (K48iu6, n557);  // ../RTL/cortexm0ds_logic.v(4741)
  AL_MUX u3238 (
    .i0(Y48iu6),
    .i1(S8fpw6[0]),
    .sel(F58iu6),
    .o(Pgvhu6));  // ../RTL/cortexm0ds_logic.v(4742)
  and u3239 (n558, M58iu6, T58iu6);  // ../RTL/cortexm0ds_logic.v(4743)
  buf u324 (Shhpw6[27], Drcbx6);  // ../RTL/cortexm0ds_logic.v(1941)
  not u3240 (Y48iu6, n558);  // ../RTL/cortexm0ds_logic.v(4743)
  and u3241 (T58iu6, A68iu6, H68iu6);  // ../RTL/cortexm0ds_logic.v(4744)
  and u3242 (H68iu6, O68iu6, V68iu6);  // ../RTL/cortexm0ds_logic.v(4745)
  or u3243 (n559, C78iu6, Bi0iu6);  // ../RTL/cortexm0ds_logic.v(4746)
  not u3244 (O68iu6, n559);  // ../RTL/cortexm0ds_logic.v(4746)
  and u3245 (A68iu6, J78iu6, Q78iu6);  // ../RTL/cortexm0ds_logic.v(4747)
  and u3246 (n560, X78iu6, E88iu6);  // ../RTL/cortexm0ds_logic.v(4748)
  not u3247 (Q78iu6, n560);  // ../RTL/cortexm0ds_logic.v(4748)
  xor u3248 (X78iu6, L88iu6, S88iu6);  // ../RTL/cortexm0ds_logic.v(4749)
  and u3249 (J78iu6, Z88iu6, G98iu6);  // ../RTL/cortexm0ds_logic.v(4750)
  buf u325 (vis_r12_o[29], F8tax6);  // ../RTL/cortexm0ds_logic.v(2599)
  and u3250 (n561, N98iu6, U98iu6);  // ../RTL/cortexm0ds_logic.v(4751)
  not u3251 (G98iu6, n561);  // ../RTL/cortexm0ds_logic.v(4751)
  or u3252 (K8aju6, Tr0iu6, Cyfpw6[6]);  // ../RTL/cortexm0ds_logic.v(4752)
  not u3253 (N98iu6, K8aju6);  // ../RTL/cortexm0ds_logic.v(4752)
  and u3254 (n562, Ba8iu6, Ia8iu6);  // ../RTL/cortexm0ds_logic.v(4753)
  not u3255 (Z88iu6, n562);  // ../RTL/cortexm0ds_logic.v(4753)
  and u3256 (M58iu6, Pa8iu6, Wa8iu6);  // ../RTL/cortexm0ds_logic.v(4754)
  and u3257 (Wa8iu6, Db8iu6, Kb8iu6);  // ../RTL/cortexm0ds_logic.v(4755)
  or u3258 (Kb8iu6, Rb8iu6, Yb8iu6);  // ../RTL/cortexm0ds_logic.v(4756)
  and u3259 (Db8iu6, Fc8iu6, Mc8iu6);  // ../RTL/cortexm0ds_logic.v(4757)
  buf u326 (vis_psp_o[3], C3zpw6);  // ../RTL/cortexm0ds_logic.v(2085)
  and u3260 (n563, Tc8iu6, Ppfpw6[0]);  // ../RTL/cortexm0ds_logic.v(4758)
  not u3261 (Mc8iu6, n563);  // ../RTL/cortexm0ds_logic.v(4758)
  or u3262 (Fc8iu6, Ad8iu6, Hd8iu6);  // ../RTL/cortexm0ds_logic.v(4759)
  and u3263 (Pa8iu6, Od8iu6, Vd8iu6);  // ../RTL/cortexm0ds_logic.v(4760)
  and u3264 (n564, Ce8iu6, Je8iu6);  // ../RTL/cortexm0ds_logic.v(4761)
  not u3265 (Vd8iu6, n564);  // ../RTL/cortexm0ds_logic.v(4761)
  and u3266 (n565, Qe8iu6, Xe8iu6);  // ../RTL/cortexm0ds_logic.v(4762)
  not u3267 (Od8iu6, n565);  // ../RTL/cortexm0ds_logic.v(4762)
  AL_MUX u3268 (
    .i0(Ef8iu6),
    .i1(vis_r0_o[4]),
    .sel(Lf8iu6),
    .o(Igvhu6));  // ../RTL/cortexm0ds_logic.v(4763)
  AL_MUX u3269 (
    .i0(vis_apsr_o[1]),
    .i1(Sf8iu6),
    .sel(Zf8iu6),
    .o(Bgvhu6));  // ../RTL/cortexm0ds_logic.v(4764)
  buf u327 (vis_r4_o[9], Vfvax6);  // ../RTL/cortexm0ds_logic.v(2626)
  and u3270 (Zf8iu6, HREADY, Gg8iu6);  // ../RTL/cortexm0ds_logic.v(4765)
  and u3271 (n566, Ng8iu6, Ug8iu6);  // ../RTL/cortexm0ds_logic.v(4766)
  not u3272 (Gg8iu6, n566);  // ../RTL/cortexm0ds_logic.v(4766)
  and u3273 (n567, Bh8iu6, Ih8iu6);  // ../RTL/cortexm0ds_logic.v(4767)
  not u3274 (Sf8iu6, n567);  // ../RTL/cortexm0ds_logic.v(4767)
  and u3275 (n568, Ph8iu6, Wh8iu6);  // ../RTL/cortexm0ds_logic.v(4768)
  not u3276 (Ih8iu6, n568);  // ../RTL/cortexm0ds_logic.v(4768)
  and u3277 (Bh8iu6, Di8iu6, Ki8iu6);  // ../RTL/cortexm0ds_logic.v(4769)
  and u3278 (n569, Ug8iu6, Ri8iu6);  // ../RTL/cortexm0ds_logic.v(4770)
  not u3279 (Ki8iu6, n569);  // ../RTL/cortexm0ds_logic.v(4770)
  buf u328 (vis_r14_o[6], Pbnax6);  // ../RTL/cortexm0ds_logic.v(2497)
  and u3280 (n570, Yi8iu6, Fj8iu6);  // ../RTL/cortexm0ds_logic.v(4771)
  not u3281 (Di8iu6, n570);  // ../RTL/cortexm0ds_logic.v(4771)
  and u3282 (n571, Mj8iu6, Tj8iu6);  // ../RTL/cortexm0ds_logic.v(4772)
  not u3283 (Ufvhu6, n571);  // ../RTL/cortexm0ds_logic.v(4772)
  and u3284 (Tj8iu6, Ak8iu6, Hk8iu6);  // ../RTL/cortexm0ds_logic.v(4773)
  and u3285 (n572, Ok8iu6, vis_pc_o[28]);  // ../RTL/cortexm0ds_logic.v(4774)
  not u3286 (Hk8iu6, n572);  // ../RTL/cortexm0ds_logic.v(4774)
  and u3287 (Ak8iu6, Vk8iu6, Cl8iu6);  // ../RTL/cortexm0ds_logic.v(4775)
  and u3288 (n573, Jl8iu6, Dx0iu6);  // ../RTL/cortexm0ds_logic.v(4776)
  not u3289 (Cl8iu6, n573);  // ../RTL/cortexm0ds_logic.v(4776)
  buf u329 (vis_r14_o[7], Odnax6);  // ../RTL/cortexm0ds_logic.v(2497)
  and u3290 (n574, Ql8iu6, vis_apsr_o[1]);  // ../RTL/cortexm0ds_logic.v(4777)
  not u3291 (Vk8iu6, n574);  // ../RTL/cortexm0ds_logic.v(4777)
  and u3292 (Mj8iu6, Xl8iu6, Em8iu6);  // ../RTL/cortexm0ds_logic.v(4778)
  or u3293 (Em8iu6, Lm8iu6, Sm8iu6);  // ../RTL/cortexm0ds_logic.v(4779)
  and u3294 (n575, Zm8iu6, M94iu6);  // ../RTL/cortexm0ds_logic.v(4780)
  not u3295 (Xl8iu6, n575);  // ../RTL/cortexm0ds_logic.v(4780)
  AL_MUX u3296 (
    .i0(Gn8iu6),
    .i1(vis_tbit_o),
    .sel(Nn8iu6),
    .o(Nfvhu6));  // ../RTL/cortexm0ds_logic.v(4781)
  and u3297 (Nn8iu6, Un8iu6, Bo8iu6);  // ../RTL/cortexm0ds_logic.v(4782)
  and u3298 (n576, Io8iu6, Po8iu6);  // ../RTL/cortexm0ds_logic.v(4783)
  not u3299 (Bo8iu6, n576);  // ../RTL/cortexm0ds_logic.v(4783)
  buf u33 (vis_r12_o[23], Kmsax6);  // ../RTL/cortexm0ds_logic.v(2599)
  buf u330 (vis_r8_o[16], O4sax6);  // ../RTL/cortexm0ds_logic.v(2579)
  and u3300 (Po8iu6, Wo8iu6, Dp8iu6);  // ../RTL/cortexm0ds_logic.v(4784)
  and u3301 (n577, Kp8iu6, Rp8iu6);  // ../RTL/cortexm0ds_logic.v(4785)
  not u3302 (Wo8iu6, n577);  // ../RTL/cortexm0ds_logic.v(4785)
  or u3303 (n578, Yp8iu6, Fq8iu6);  // ../RTL/cortexm0ds_logic.v(4786)
  not u3304 (Rp8iu6, n578);  // ../RTL/cortexm0ds_logic.v(4786)
  and u3305 (Kp8iu6, Mq8iu6, Tq8iu6);  // ../RTL/cortexm0ds_logic.v(4787)
  buf u3306 (Ynehu6, Ozkbx6[25]);  // ../RTL/cortexm0ds_logic.v(3176)
  or u3307 (Mq8iu6, Cyfpw6[3], Y7ghu6);  // ../RTL/cortexm0ds_logic.v(4789)
  and u3308 (Io8iu6, Ar8iu6, Hr8iu6);  // ../RTL/cortexm0ds_logic.v(4790)
  and u3309 (n579, HREADY, Or8iu6);  // ../RTL/cortexm0ds_logic.v(4791)
  buf u331 (Vbgpw6[10], C50bx6);  // ../RTL/cortexm0ds_logic.v(3092)
  not u3310 (Un8iu6, n579);  // ../RTL/cortexm0ds_logic.v(4791)
  and u3311 (n580, Vr8iu6, Cs8iu6);  // ../RTL/cortexm0ds_logic.v(4792)
  not u3312 (Or8iu6, n580);  // ../RTL/cortexm0ds_logic.v(4792)
  AL_MUX u3313 (
    .i0(Fkfpw6[24]),
    .i1(Js8iu6),
    .sel(Vr8iu6),
    .o(Gn8iu6));  // ../RTL/cortexm0ds_logic.v(4793)
  and u3314 (n581, Qs8iu6, Xs8iu6);  // ../RTL/cortexm0ds_logic.v(4794)
  not u3315 (Js8iu6, n581);  // ../RTL/cortexm0ds_logic.v(4794)
  and u3316 (n582, Eafpw6[0], Et8iu6);  // ../RTL/cortexm0ds_logic.v(4795)
  not u3317 (Xs8iu6, n582);  // ../RTL/cortexm0ds_logic.v(4795)
  and u3318 (Qs8iu6, Lt8iu6, St8iu6);  // ../RTL/cortexm0ds_logic.v(4796)
  or u3319 (St8iu6, Zt8iu6, Gu8iu6);  // ../RTL/cortexm0ds_logic.v(4797)
  buf u332 (vis_r14_o[20], Nrnax6);  // ../RTL/cortexm0ds_logic.v(2497)
  and u3320 (n583, Yi8iu6, Nu8iu6);  // ../RTL/cortexm0ds_logic.v(4798)
  not u3321 (Lt8iu6, n583);  // ../RTL/cortexm0ds_logic.v(4798)
  and u3322 (n584, Uu8iu6, Bv8iu6);  // ../RTL/cortexm0ds_logic.v(4799)
  not u3323 (Gfvhu6, n584);  // ../RTL/cortexm0ds_logic.v(4799)
  and u3324 (Bv8iu6, Iv8iu6, Pv8iu6);  // ../RTL/cortexm0ds_logic.v(4800)
  and u3325 (n585, Hrfpw6[14], Uy4iu6);  // ../RTL/cortexm0ds_logic.v(4801)
  not u3326 (Pv8iu6, n585);  // ../RTL/cortexm0ds_logic.v(4801)
  and u3327 (Iv8iu6, Wv8iu6, Dw8iu6);  // ../RTL/cortexm0ds_logic.v(4802)
  and u3328 (n586, M15iu6, Kw8iu6);  // ../RTL/cortexm0ds_logic.v(4803)
  not u3329 (Dw8iu6, n586);  // ../RTL/cortexm0ds_logic.v(4803)
  buf u333 (vis_r4_o[11], Ci7bx6);  // ../RTL/cortexm0ds_logic.v(2626)
  and u3330 (n587, Pz4iu6, Rw8iu6);  // ../RTL/cortexm0ds_logic.v(4804)
  not u3331 (Wv8iu6, n587);  // ../RTL/cortexm0ds_logic.v(4804)
  and u3332 (Uu8iu6, Yw8iu6, Fx8iu6);  // ../RTL/cortexm0ds_logic.v(4805)
  and u3333 (n588, Ppfpw6[14], A25iu6);  // ../RTL/cortexm0ds_logic.v(4806)
  not u3334 (Fx8iu6, n588);  // ../RTL/cortexm0ds_logic.v(4806)
  and u3335 (n589, R05iu6, D7fpw6[14]);  // ../RTL/cortexm0ds_logic.v(4807)
  not u3336 (Yw8iu6, n589);  // ../RTL/cortexm0ds_logic.v(4807)
  AL_MUX u3337 (
    .i0(Ef8iu6),
    .i1(vis_r1_o[4]),
    .sel(Mx8iu6),
    .o(Zevhu6));  // ../RTL/cortexm0ds_logic.v(4808)
  AL_MUX u3338 (
    .i0(Tx8iu6),
    .i1(vis_r1_o[0]),
    .sel(Mx8iu6),
    .o(Sevhu6));  // ../RTL/cortexm0ds_logic.v(4809)
  AL_MUX u3339 (
    .i0(Iwfpw6[0]),
    .i1(Ay8iu6),
    .sel(Hy8iu6),
    .o(Levhu6));  // ../RTL/cortexm0ds_logic.v(4810)
  buf u334 (vis_r14_o[8], N9oax6);  // ../RTL/cortexm0ds_logic.v(2497)
  AL_MUX u3340 (
    .i0(Tx8iu6),
    .i1(vis_r0_o[0]),
    .sel(Lf8iu6),
    .o(Eevhu6));  // ../RTL/cortexm0ds_logic.v(4811)
  AL_MUX u3341 (
    .i0(Oy8iu6),
    .i1(vis_primask_o),
    .sel(n590),
    .o(Xdvhu6));  // ../RTL/cortexm0ds_logic.v(4812)
  or u3342 (n590, Eh6iu6, Cz8iu6);  // ../RTL/cortexm0ds_logic.v(4813)
  buf u3343 (Eafpw6[3], Nxkbx6[4]);  // ../RTL/cortexm0ds_logic.v(3167)
  and u3344 (n591, Jz8iu6, Qz8iu6);  // ../RTL/cortexm0ds_logic.v(4814)
  not u3345 (Qdvhu6, n591);  // ../RTL/cortexm0ds_logic.v(4814)
  and u3346 (Qz8iu6, Xz8iu6, E09iu6);  // ../RTL/cortexm0ds_logic.v(4815)
  and u3347 (n592, Ql8iu6, vis_ipsr_o[0]);  // ../RTL/cortexm0ds_logic.v(4816)
  not u3348 (E09iu6, n592);  // ../RTL/cortexm0ds_logic.v(4816)
  and u3349 (Xz8iu6, L09iu6, S09iu6);  // ../RTL/cortexm0ds_logic.v(4817)
  buf u335 (vis_r8_o[17], O2sax6);  // ../RTL/cortexm0ds_logic.v(2579)
  and u3350 (n593, Jl8iu6, Z09iu6);  // ../RTL/cortexm0ds_logic.v(4818)
  not u3351 (S09iu6, n593);  // ../RTL/cortexm0ds_logic.v(4818)
  or u3352 (Z09iu6, Ay8iu6, G19iu6);  // ../RTL/cortexm0ds_logic.v(4819)
  or u3353 (n594, N19iu6, U19iu6);  // ../RTL/cortexm0ds_logic.v(4820)
  not u3354 (G19iu6, n594);  // ../RTL/cortexm0ds_logic.v(4820)
  and u3355 (n595, B29iu6, vis_primask_o);  // ../RTL/cortexm0ds_logic.v(4821)
  not u3356 (L09iu6, n595);  // ../RTL/cortexm0ds_logic.v(4821)
  and u3357 (Jz8iu6, I29iu6, P29iu6);  // ../RTL/cortexm0ds_logic.v(4822)
  and u3358 (n596, W29iu6, Fkfpw6[0]);  // ../RTL/cortexm0ds_logic.v(4823)
  not u3359 (P29iu6, n596);  // ../RTL/cortexm0ds_logic.v(4823)
  buf u336 (Vbgpw6[11], D70bx6);  // ../RTL/cortexm0ds_logic.v(3092)
  and u3360 (n597, Zm8iu6, T24iu6);  // ../RTL/cortexm0ds_logic.v(4824)
  not u3361 (I29iu6, n597);  // ../RTL/cortexm0ds_logic.v(4824)
  AL_MUX u3362 (
    .i0(D39iu6),
    .i1(vis_r1_o[31]),
    .sel(Mx8iu6),
    .o(Jdvhu6));  // ../RTL/cortexm0ds_logic.v(4825)
  AL_MUX u3363 (
    .i0(D39iu6),
    .i1(vis_r0_o[31]),
    .sel(Lf8iu6),
    .o(Cdvhu6));  // ../RTL/cortexm0ds_logic.v(4826)
  AL_MUX u3364 (
    .i0(K39iu6),
    .i1(vis_r1_o[30]),
    .sel(Mx8iu6),
    .o(Vcvhu6));  // ../RTL/cortexm0ds_logic.v(4827)
  AL_MUX u3365 (
    .i0(K39iu6),
    .i1(vis_r0_o[30]),
    .sel(Lf8iu6),
    .o(Ocvhu6));  // ../RTL/cortexm0ds_logic.v(4828)
  and u3366 (n598, R39iu6, Y39iu6);  // ../RTL/cortexm0ds_logic.v(4829)
  not u3367 (Hcvhu6, n598);  // ../RTL/cortexm0ds_logic.v(4829)
  and u3368 (n599, Jfgpw6[1], Eh6iu6);  // ../RTL/cortexm0ds_logic.v(4830)
  not u3369 (Y39iu6, n599);  // ../RTL/cortexm0ds_logic.v(4830)
  buf u337 (vis_r14_o[25], Nnnax6);  // ../RTL/cortexm0ds_logic.v(2497)
  and u3370 (R39iu6, F49iu6, Ii7iu6);  // ../RTL/cortexm0ds_logic.v(4831)
  and u3371 (n600, M49iu6, Wi7iu6);  // ../RTL/cortexm0ds_logic.v(4832)
  not u3372 (F49iu6, n600);  // ../RTL/cortexm0ds_logic.v(4832)
  and u3373 (n601, T49iu6, A59iu6);  // ../RTL/cortexm0ds_logic.v(4833)
  not u3374 (Acvhu6, n601);  // ../RTL/cortexm0ds_logic.v(4833)
  and u3375 (n602, Vbgpw6[31], H59iu6);  // ../RTL/cortexm0ds_logic.v(4834)
  not u3376 (A59iu6, n602);  // ../RTL/cortexm0ds_logic.v(4834)
  and u3377 (n603, HWDATA[31], O59iu6);  // ../RTL/cortexm0ds_logic.v(4835)
  not u3378 (H59iu6, n603);  // ../RTL/cortexm0ds_logic.v(4835)
  and u3379 (n604, V59iu6, HWDATA[31]);  // ../RTL/cortexm0ds_logic.v(4836)
  buf u338 (vis_r7_o[4], Slvax6);  // ../RTL/cortexm0ds_logic.v(2654)
  not u3380 (T49iu6, n604);  // ../RTL/cortexm0ds_logic.v(4836)
  and u3381 (n605, C69iu6, J69iu6);  // ../RTL/cortexm0ds_logic.v(4837)
  not u3382 (Tbvhu6, n605);  // ../RTL/cortexm0ds_logic.v(4837)
  and u3383 (n606, Vbgpw6[0], Q69iu6);  // ../RTL/cortexm0ds_logic.v(4838)
  not u3384 (J69iu6, n606);  // ../RTL/cortexm0ds_logic.v(4838)
  and u3385 (n607, HWDATA[0], O59iu6);  // ../RTL/cortexm0ds_logic.v(4839)
  not u3386 (Q69iu6, n607);  // ../RTL/cortexm0ds_logic.v(4839)
  and u3387 (n608, V59iu6, HWDATA[0]);  // ../RTL/cortexm0ds_logic.v(4840)
  not u3388 (C69iu6, n608);  // ../RTL/cortexm0ds_logic.v(4840)
  and u3389 (n609, X69iu6, E79iu6);  // ../RTL/cortexm0ds_logic.v(4841)
  buf u339 (B3gpw6[0], Tl4bx6);  // ../RTL/cortexm0ds_logic.v(2808)
  not u3390 (Mbvhu6, n609);  // ../RTL/cortexm0ds_logic.v(4841)
  and u3391 (n610, Jfgpw6[3], Eh6iu6);  // ../RTL/cortexm0ds_logic.v(4842)
  not u3392 (E79iu6, n610);  // ../RTL/cortexm0ds_logic.v(4842)
  and u3393 (X69iu6, L79iu6, Ii7iu6);  // ../RTL/cortexm0ds_logic.v(4843)
  and u3394 (n611, S79iu6, Wi7iu6);  // ../RTL/cortexm0ds_logic.v(4844)
  not u3395 (L79iu6, n611);  // ../RTL/cortexm0ds_logic.v(4844)
  xor u3396 (n612, HADDR[3], Z79iu6);  // ../RTL/cortexm0ds_logic.v(4845)
  not u3397 (S79iu6, n612);  // ../RTL/cortexm0ds_logic.v(4845)
  and u3398 (n613, G89iu6, N89iu6);  // ../RTL/cortexm0ds_logic.v(4846)
  not u3399 (Fbvhu6, n613);  // ../RTL/cortexm0ds_logic.v(4846)
  not u34 (Tugpw6[13], n1272[12]);  // ../RTL/cortexm0ds_logic.v(16030)
  buf u340 (vis_r7_o[3], Qvvax6);  // ../RTL/cortexm0ds_logic.v(2654)
  or u3400 (N89iu6, U89iu6, HREADY);  // ../RTL/cortexm0ds_logic.v(4847)
  and u3401 (G89iu6, B99iu6, Ii7iu6);  // ../RTL/cortexm0ds_logic.v(4848)
  and u3402 (n614, I99iu6, Wi7iu6);  // ../RTL/cortexm0ds_logic.v(4849)
  not u3403 (B99iu6, n614);  // ../RTL/cortexm0ds_logic.v(4849)
  xor u3404 (n615, HADDR[2], P99iu6);  // ../RTL/cortexm0ds_logic.v(4850)
  not u3405 (I99iu6, n615);  // ../RTL/cortexm0ds_logic.v(4850)
  and u3406 (n616, W99iu6, Da9iu6);  // ../RTL/cortexm0ds_logic.v(4851)
  not u3407 (Yavhu6, n616);  // ../RTL/cortexm0ds_logic.v(4851)
  or u3408 (Da9iu6, Ka9iu6, HREADY);  // ../RTL/cortexm0ds_logic.v(4852)
  and u3409 (W99iu6, Ra9iu6, Ii7iu6);  // ../RTL/cortexm0ds_logic.v(4853)
  buf u341 (vis_r9_o[24], Yrspw6);  // ../RTL/cortexm0ds_logic.v(1898)
  and u3410 (n617, Wi7iu6, Ya9iu6);  // ../RTL/cortexm0ds_logic.v(4854)
  not u3411 (Ii7iu6, n617);  // ../RTL/cortexm0ds_logic.v(4854)
  and u3412 (n618, Fb9iu6, Mb9iu6);  // ../RTL/cortexm0ds_logic.v(4855)
  not u3413 (Ya9iu6, n618);  // ../RTL/cortexm0ds_logic.v(4855)
  and u3414 (Mb9iu6, HSIZE[1], Tb9iu6);  // ../RTL/cortexm0ds_logic.v(4856)
  and u3415 (n619, Ac9iu6, Hc9iu6);  // ../RTL/cortexm0ds_logic.v(4857)
  not u3416 (Tb9iu6, n619);  // ../RTL/cortexm0ds_logic.v(4857)
  and u3417 (n620, Oc9iu6, Vc9iu6);  // ../RTL/cortexm0ds_logic.v(4858)
  not u3418 (Hc9iu6, n620);  // ../RTL/cortexm0ds_logic.v(4858)
  or u3419 (n621, Cd9iu6, HADDR[9]);  // ../RTL/cortexm0ds_logic.v(4859)
  buf u342 (vis_r14_o[26], Nhnax6);  // ../RTL/cortexm0ds_logic.v(2497)
  not u3420 (Vc9iu6, n621);  // ../RTL/cortexm0ds_logic.v(4859)
  and u3421 (n622, Jd9iu6, Qd9iu6);  // ../RTL/cortexm0ds_logic.v(4860)
  not u3422 (Cd9iu6, n622);  // ../RTL/cortexm0ds_logic.v(4860)
  and u3423 (n623, HADDR[6], Xd9iu6);  // ../RTL/cortexm0ds_logic.v(4861)
  not u3424 (Qd9iu6, n623);  // ../RTL/cortexm0ds_logic.v(4861)
  and u3425 (n624, HADDR[7], Ee9iu6);  // ../RTL/cortexm0ds_logic.v(4862)
  not u3426 (Xd9iu6, n624);  // ../RTL/cortexm0ds_logic.v(4862)
  or u3427 (Ee9iu6, HADDR[3], HADDR[2]);  // ../RTL/cortexm0ds_logic.v(4863)
  and u3428 (n625, HADDR[7], Le9iu6);  // ../RTL/cortexm0ds_logic.v(4864)
  not u3429 (Jd9iu6, n625);  // ../RTL/cortexm0ds_logic.v(4864)
  buf u343 (vis_r14_o[31], S3nax6);  // ../RTL/cortexm0ds_logic.v(2497)
  and u3430 (n626, Se9iu6, HADDR[11]);  // ../RTL/cortexm0ds_logic.v(4865)
  not u3431 (Le9iu6, n626);  // ../RTL/cortexm0ds_logic.v(4865)
  or u3432 (n627, M49iu6, Ze9iu6);  // ../RTL/cortexm0ds_logic.v(4866)
  not u3433 (Se9iu6, n627);  // ../RTL/cortexm0ds_logic.v(4866)
  and u3434 (Oc9iu6, Gf9iu6, Nf9iu6);  // ../RTL/cortexm0ds_logic.v(4867)
  AL_MUX u3435 (
    .i0(Pi7iu6),
    .i1(Uf9iu6),
    .sel(HADDR[11]),
    .o(Nf9iu6));  // ../RTL/cortexm0ds_logic.v(4868)
  and u3436 (Uf9iu6, Bg9iu6, Ig9iu6);  // ../RTL/cortexm0ds_logic.v(4869)
  and u3437 (Ig9iu6, Pg9iu6, Wg9iu6);  // ../RTL/cortexm0ds_logic.v(4870)
  and u3438 (n628, HADDR[3], Dh9iu6);  // ../RTL/cortexm0ds_logic.v(4871)
  not u3439 (Wg9iu6, n628);  // ../RTL/cortexm0ds_logic.v(4871)
  buf u344 (vis_r9_o[1], Rhypw6);  // ../RTL/cortexm0ds_logic.v(1898)
  or u3440 (Dh9iu6, M49iu6, HADDR[2]);  // ../RTL/cortexm0ds_logic.v(4872)
  or u3441 (Pg9iu6, M49iu6, HADDR[6]);  // ../RTL/cortexm0ds_logic.v(4873)
  not u3442 (M49iu6, HADDR[4]);  // ../RTL/cortexm0ds_logic.v(4874)
  and u3443 (Bg9iu6, HADDR[5], Kh9iu6);  // ../RTL/cortexm0ds_logic.v(4875)
  or u3444 (Kh9iu6, Rh9iu6, Xg6iu6);  // ../RTL/cortexm0ds_logic.v(4876)
  not u3445 (Rh9iu6, HADDR[2]);  // ../RTL/cortexm0ds_logic.v(4877)
  and u3446 (Gf9iu6, HADDR[10], Yh9iu6);  // ../RTL/cortexm0ds_logic.v(4878)
  or u3447 (Yh9iu6, Z79iu6, HADDR[8]);  // ../RTL/cortexm0ds_logic.v(4879)
  AL_MUX u3448 (
    .i0(Fi9iu6),
    .i1(Mi9iu6),
    .sel(HADDR[11]),
    .o(Ac9iu6));  // ../RTL/cortexm0ds_logic.v(4880)
  and u3449 (n629, Ti9iu6, Aj9iu6);  // ../RTL/cortexm0ds_logic.v(4882)
  buf u345 (vis_r9_o[6], Z3spw6);  // ../RTL/cortexm0ds_logic.v(1898)
  not u3450 (Mi9iu6, n629);  // ../RTL/cortexm0ds_logic.v(4882)
  and u3451 (Aj9iu6, Hj9iu6, Oj9iu6);  // ../RTL/cortexm0ds_logic.v(4883)
  and u3452 (Oj9iu6, HADDR[10], Vj9iu6);  // ../RTL/cortexm0ds_logic.v(4884)
  or u3453 (Vj9iu6, Ck9iu6, HADDR[2]);  // ../RTL/cortexm0ds_logic.v(4885)
  or u3454 (n630, HADDR[6], Pi7iu6);  // ../RTL/cortexm0ds_logic.v(4886)
  not u3455 (Hj9iu6, n630);  // ../RTL/cortexm0ds_logic.v(4886)
  and u3456 (Ti9iu6, Jk9iu6, P99iu6);  // ../RTL/cortexm0ds_logic.v(4887)
  not u3457 (P99iu6, HADDR[7]);  // ../RTL/cortexm0ds_logic.v(4888)
  or u3458 (n631, HADDR[9], HADDR[5]);  // ../RTL/cortexm0ds_logic.v(4889)
  not u3459 (Jk9iu6, n631);  // ../RTL/cortexm0ds_logic.v(4889)
  buf u346 (vis_r9_o[7], Cqrpw6);  // ../RTL/cortexm0ds_logic.v(1898)
  and u3460 (n632, Qk9iu6, Z79iu6);  // ../RTL/cortexm0ds_logic.v(4890)
  not u3461 (Fi9iu6, n632);  // ../RTL/cortexm0ds_logic.v(4890)
  not u3462 (Z79iu6, HADDR[5]);  // ../RTL/cortexm0ds_logic.v(4891)
  and u3463 (Qk9iu6, Xk9iu6, El9iu6);  // ../RTL/cortexm0ds_logic.v(4893)
  not u3464 (El9iu6, HADDR[6]);  // ../RTL/cortexm0ds_logic.v(4894)
  AL_MUX u3465 (
    .i0(Sl9iu6),
    .i1(Ll9iu6),
    .sel(n633),
    .o(Xk9iu6));  // ../RTL/cortexm0ds_logic.v(4895)
  or u3466 (n633, HADDR[4], HADDR[3]);  // ../RTL/cortexm0ds_logic.v(4896)
  buf u3467 (Eafpw6[2], Nxkbx6[3]);  // ../RTL/cortexm0ds_logic.v(3167)
  and u3468 (Sl9iu6, Gm9iu6, Nm9iu6);  // ../RTL/cortexm0ds_logic.v(4898)
  xor u3469 (n634, HADDR[9], Pi7iu6);  // ../RTL/cortexm0ds_logic.v(4899)
  buf u347 (vis_r9_o[9], Ht1qw6);  // ../RTL/cortexm0ds_logic.v(1898)
  not u3470 (Nm9iu6, n634);  // ../RTL/cortexm0ds_logic.v(4899)
  or u3471 (n635, HADDR[2], HADDR[10]);  // ../RTL/cortexm0ds_logic.v(4900)
  not u3472 (Gm9iu6, n635);  // ../RTL/cortexm0ds_logic.v(4900)
  AL_MUX u3473 (
    .i0(Tnhpw6[2]),
    .i1(Vo4iu6),
    .sel(Wqzhu6),
    .o(P47iu6));  // ../RTL/cortexm0ds_logic.v(4902)
  and u3474 (Ll9iu6, Um9iu6, Pi7iu6);  // ../RTL/cortexm0ds_logic.v(4903)
  not u3475 (Pi7iu6, HADDR[8]);  // ../RTL/cortexm0ds_logic.v(4904)
  or u3476 (n636, HADDR[9], HADDR[7]);  // ../RTL/cortexm0ds_logic.v(4906)
  not u3477 (Um9iu6, n636);  // ../RTL/cortexm0ds_logic.v(4906)
  and u3478 (Fb9iu6, Bn9iu6, HADDR[15]);  // ../RTL/cortexm0ds_logic.v(4908)
  AL_MUX u3479 (
    .i0(In9iu6),
    .i1(Pn9iu6),
    .sel(Xg6iu6),
    .o(Bn9iu6));  // ../RTL/cortexm0ds_logic.v(4909)
  buf u348 (vis_r9_o[10], Hoxpw6);  // ../RTL/cortexm0ds_logic.v(1898)
  and u3480 (Pn9iu6, Wn9iu6, Fs6iu6);  // ../RTL/cortexm0ds_logic.v(4910)
  and u3481 (Fs6iu6, Do9iu6, Ko9iu6);  // ../RTL/cortexm0ds_logic.v(4911)
  and u3482 (Ko9iu6, Ro9iu6, Yo9iu6);  // ../RTL/cortexm0ds_logic.v(4912)
  not u3483 (Yo9iu6, Jshpw6[25]);  // ../RTL/cortexm0ds_logic.v(4913)
  or u3484 (n637, Jshpw6[26], Jshpw6[27]);  // ../RTL/cortexm0ds_logic.v(4914)
  not u3485 (Ro9iu6, n637);  // ../RTL/cortexm0ds_logic.v(4914)
  and u3486 (Do9iu6, Fp9iu6, Mp9iu6);  // ../RTL/cortexm0ds_logic.v(4915)
  not u3487 (Mp9iu6, Jshpw6[22]);  // ../RTL/cortexm0ds_logic.v(4916)
  or u3488 (n638, Jshpw6[23], Jshpw6[24]);  // ../RTL/cortexm0ds_logic.v(4917)
  not u3489 (Fp9iu6, n638);  // ../RTL/cortexm0ds_logic.v(4917)
  buf u349 (vis_r9_o[12], O3ppw6);  // ../RTL/cortexm0ds_logic.v(1898)
  and u3490 (Wn9iu6, Tp9iu6, Aq9iu6);  // ../RTL/cortexm0ds_logic.v(4918)
  and u3491 (Aq9iu6, At6iu6, Bx6iu6);  // ../RTL/cortexm0ds_logic.v(4919)
  not u3492 (Bx6iu6, Jshpw6[12]);  // ../RTL/cortexm0ds_logic.v(4920)
  or u3493 (n639, Jshpw6[20], Jshpw6[21]);  // ../RTL/cortexm0ds_logic.v(4921)
  not u3494 (At6iu6, n639);  // ../RTL/cortexm0ds_logic.v(4921)
  and u3495 (Tp9iu6, Kc7iu6, Mz6iu6);  // ../RTL/cortexm0ds_logic.v(4922)
  and u3496 (Mz6iu6, Hq9iu6, Oq9iu6);  // ../RTL/cortexm0ds_logic.v(4923)
  or u3497 (n640, Jshpw6[18], Jshpw6[19]);  // ../RTL/cortexm0ds_logic.v(4924)
  not u3498 (Oq9iu6, n640);  // ../RTL/cortexm0ds_logic.v(4924)
  or u3499 (n641, Jshpw6[16], Jshpw6[17]);  // ../RTL/cortexm0ds_logic.v(4925)
  buf u35 (Jshpw6[24], No3qw6);  // ../RTL/cortexm0ds_logic.v(2372)
  buf u350 (vis_r9_o[13], O1ppw6);  // ../RTL/cortexm0ds_logic.v(1898)
  not u3500 (Hq9iu6, n641);  // ../RTL/cortexm0ds_logic.v(4925)
  and u3501 (Kc7iu6, Jshpw6[14], Jshpw6[13]);  // ../RTL/cortexm0ds_logic.v(4926)
  and u3502 (In9iu6, Vq9iu6, Cr9iu6);  // ../RTL/cortexm0ds_logic.v(4927)
  and u3503 (Cr9iu6, Jr9iu6, Qr9iu6);  // ../RTL/cortexm0ds_logic.v(4928)
  and u3504 (Qr9iu6, Xr9iu6, Es9iu6);  // ../RTL/cortexm0ds_logic.v(4929)
  or u3505 (n642, Pxdpw6, Ixdpw6);  // ../RTL/cortexm0ds_logic.v(4930)
  not u3506 (Es9iu6, n642);  // ../RTL/cortexm0ds_logic.v(4930)
  or u3507 (n643, Dydpw6, Wxdpw6);  // ../RTL/cortexm0ds_logic.v(4931)
  not u3508 (Xr9iu6, n643);  // ../RTL/cortexm0ds_logic.v(4931)
  and u3509 (Jr9iu6, Ls9iu6, Ss9iu6);  // ../RTL/cortexm0ds_logic.v(4932)
  buf u351 (vis_r9_o[15], Z18bx6);  // ../RTL/cortexm0ds_logic.v(1898)
  or u3510 (n644, Rydpw6, Kydpw6);  // ../RTL/cortexm0ds_logic.v(4933)
  not u3511 (Ss9iu6, n644);  // ../RTL/cortexm0ds_logic.v(4933)
  or u3512 (n645, Fzdpw6, Yydpw6);  // ../RTL/cortexm0ds_logic.v(4934)
  not u3513 (Ls9iu6, n645);  // ../RTL/cortexm0ds_logic.v(4934)
  and u3514 (Vq9iu6, Zs9iu6, Gt9iu6);  // ../RTL/cortexm0ds_logic.v(4935)
  and u3515 (Gt9iu6, Nt9iu6, Ut9iu6);  // ../RTL/cortexm0ds_logic.v(4936)
  or u3516 (n646, Tzdpw6, Mzdpw6);  // ../RTL/cortexm0ds_logic.v(4937)
  not u3517 (Ut9iu6, n646);  // ../RTL/cortexm0ds_logic.v(4937)
  or u3518 (n647, H0epw6, A0epw6);  // ../RTL/cortexm0ds_logic.v(4938)
  not u3519 (Nt9iu6, n647);  // ../RTL/cortexm0ds_logic.v(4938)
  buf u352 (vis_r9_o[17], Ybupw6);  // ../RTL/cortexm0ds_logic.v(1898)
  and u3520 (Zs9iu6, Bu9iu6, Tugpw6[12]);  // ../RTL/cortexm0ds_logic.v(4939)
  or u3521 (n648, Iu9iu6, O0epw6);  // ../RTL/cortexm0ds_logic.v(4940)
  not u3522 (Bu9iu6, n648);  // ../RTL/cortexm0ds_logic.v(4940)
  and u3523 (n649, Pu9iu6, Wi7iu6);  // ../RTL/cortexm0ds_logic.v(4942)
  not u3524 (Ra9iu6, n649);  // ../RTL/cortexm0ds_logic.v(4942)
  xor u3525 (n650, HADDR[10], Ck9iu6);  // ../RTL/cortexm0ds_logic.v(4943)
  not u3526 (Pu9iu6, n650);  // ../RTL/cortexm0ds_logic.v(4943)
  not u3527 (Ck9iu6, HADDR[3]);  // ../RTL/cortexm0ds_logic.v(4944)
  AL_MUX u3528 (
    .i0(Tnhpw6[3]),
    .i1(Wu9iu6),
    .sel(Wqzhu6),
    .o(I47iu6));  // ../RTL/cortexm0ds_logic.v(4946)
  AL_MUX u3529 (
    .i0(HWDATA[31]),
    .i1(R4gpw6[7]),
    .sel(Dv9iu6),
    .o(Ravhu6));  // ../RTL/cortexm0ds_logic.v(4948)
  buf u353 (vis_r9_o[18], P6xpw6);  // ../RTL/cortexm0ds_logic.v(1898)
  and u3530 (n651, Kv9iu6, Rv9iu6);  // ../RTL/cortexm0ds_logic.v(4949)
  not u3531 (Kavhu6, n651);  // ../RTL/cortexm0ds_logic.v(4949)
  and u3532 (Rv9iu6, Yv9iu6, Fw9iu6);  // ../RTL/cortexm0ds_logic.v(4950)
  and u3533 (n652, Jl8iu6, Mzdpw6);  // ../RTL/cortexm0ds_logic.v(4951)
  not u3534 (Fw9iu6, n652);  // ../RTL/cortexm0ds_logic.v(4951)
  and u3535 (n653, vis_pc_o[22], Ok8iu6);  // ../RTL/cortexm0ds_logic.v(4952)
  not u3536 (Yv9iu6, n653);  // ../RTL/cortexm0ds_logic.v(4952)
  and u3537 (Kv9iu6, Mw9iu6, Tw9iu6);  // ../RTL/cortexm0ds_logic.v(4953)
  or u3538 (Tw9iu6, Lm8iu6, Ax9iu6);  // ../RTL/cortexm0ds_logic.v(4954)
  or u3539 (Mw9iu6, Hx9iu6, Ox9iu6);  // ../RTL/cortexm0ds_logic.v(4955)
  buf u354 (vis_r9_o[20], Ozopw6);  // ../RTL/cortexm0ds_logic.v(1898)
  AL_MUX u3540 (
    .i0(Vx9iu6),
    .i1(vis_r1_o[23]),
    .sel(Mx8iu6),
    .o(Davhu6));  // ../RTL/cortexm0ds_logic.v(4956)
  AL_MUX u3541 (
    .i0(Vx9iu6),
    .i1(vis_r0_o[23]),
    .sel(Lf8iu6),
    .o(W9vhu6));  // ../RTL/cortexm0ds_logic.v(4957)
  AL_MUX u3542 (
    .i0(Vrfhu6),
    .i1(Cy9iu6),
    .sel(Jy9iu6),
    .o(P9vhu6));  // ../RTL/cortexm0ds_logic.v(4958)
  and u3543 (Jy9iu6, HREADY, Qy9iu6);  // ../RTL/cortexm0ds_logic.v(4959)
  and u3544 (n654, Xy9iu6, Ez9iu6);  // ../RTL/cortexm0ds_logic.v(4960)
  not u3545 (Qy9iu6, n654);  // ../RTL/cortexm0ds_logic.v(4960)
  and u3546 (Ez9iu6, Lz9iu6, Sz9iu6);  // ../RTL/cortexm0ds_logic.v(4961)
  and u3547 (Sz9iu6, Zz9iu6, G0aiu6);  // ../RTL/cortexm0ds_logic.v(4962)
  and u3548 (n655, N0aiu6, U0aiu6);  // ../RTL/cortexm0ds_logic.v(4963)
  not u3549 (G0aiu6, n655);  // ../RTL/cortexm0ds_logic.v(4963)
  buf u355 (vis_r9_o[21], Oxopw6);  // ../RTL/cortexm0ds_logic.v(1898)
  or u3550 (n656, Cyfpw6[6], Y7ghu6);  // ../RTL/cortexm0ds_logic.v(4964)
  not u3551 (N0aiu6, n656);  // ../RTL/cortexm0ds_logic.v(4964)
  and u3552 (Zz9iu6, B1aiu6, I1aiu6);  // ../RTL/cortexm0ds_logic.v(4965)
  and u3553 (Lz9iu6, P1aiu6, W1aiu6);  // ../RTL/cortexm0ds_logic.v(4966)
  and u3554 (n657, D2aiu6, K2aiu6);  // ../RTL/cortexm0ds_logic.v(4967)
  not u3555 (W1aiu6, n657);  // ../RTL/cortexm0ds_logic.v(4967)
  or u3556 (n658, R2aiu6, Cyfpw6[4]);  // ../RTL/cortexm0ds_logic.v(4968)
  not u3557 (D2aiu6, n658);  // ../RTL/cortexm0ds_logic.v(4968)
  and u3558 (n659, Y2aiu6, F3aiu6);  // ../RTL/cortexm0ds_logic.v(4969)
  not u3559 (P1aiu6, n659);  // ../RTL/cortexm0ds_logic.v(4969)
  buf u356 (vis_r9_o[22], Txebx6);  // ../RTL/cortexm0ds_logic.v(1898)
  and u3560 (Xy9iu6, M3aiu6, T3aiu6);  // ../RTL/cortexm0ds_logic.v(4970)
  and u3561 (T3aiu6, A4aiu6, H4aiu6);  // ../RTL/cortexm0ds_logic.v(4971)
  or u3562 (H4aiu6, O4aiu6, V4aiu6);  // ../RTL/cortexm0ds_logic.v(4972)
  and u3563 (A4aiu6, C5aiu6, J5aiu6);  // ../RTL/cortexm0ds_logic.v(4973)
  or u3564 (C5aiu6, Q5aiu6, X5aiu6);  // ../RTL/cortexm0ds_logic.v(4974)
  and u3565 (M3aiu6, E6aiu6, L6aiu6);  // ../RTL/cortexm0ds_logic.v(4975)
  and u3566 (n660, S6aiu6, Z6aiu6);  // ../RTL/cortexm0ds_logic.v(4976)
  not u3567 (E6aiu6, n660);  // ../RTL/cortexm0ds_logic.v(4976)
  and u3568 (n661, G7aiu6, N7aiu6);  // ../RTL/cortexm0ds_logic.v(4977)
  not u3569 (Cy9iu6, n661);  // ../RTL/cortexm0ds_logic.v(4977)
  buf u357 (vis_r9_o[23], P34qw6);  // ../RTL/cortexm0ds_logic.v(1898)
  and u3570 (n662, U7aiu6, B8aiu6);  // ../RTL/cortexm0ds_logic.v(4978)
  not u3571 (N7aiu6, n662);  // ../RTL/cortexm0ds_logic.v(4978)
  or u3572 (B8aiu6, I8aiu6, P8aiu6);  // ../RTL/cortexm0ds_logic.v(4979)
  AL_MUX u3573 (
    .i0(W8aiu6),
    .i1(D9aiu6),
    .sel(Cyfpw6[3]),
    .o(P8aiu6));  // ../RTL/cortexm0ds_logic.v(4980)
  or u3574 (D9aiu6, K9aiu6, R9aiu6);  // ../RTL/cortexm0ds_logic.v(4981)
  and u3575 (n663, Y9aiu6, Faaiu6);  // ../RTL/cortexm0ds_logic.v(4982)
  not u3576 (I8aiu6, n663);  // ../RTL/cortexm0ds_logic.v(4982)
  AL_MUX u3577 (
    .i0(Cyfpw6[5]),
    .i1(D7fpw6[3]),
    .sel(Mr0iu6),
    .o(Y9aiu6));  // ../RTL/cortexm0ds_logic.v(4983)
  or u3578 (U7aiu6, vis_control_o, Maaiu6);  // ../RTL/cortexm0ds_logic.v(4984)
  or u3579 (n664, Taaiu6, Quzhu6);  // ../RTL/cortexm0ds_logic.v(4985)
  buf u358 (Aygpw6[0], Tikbx6);  // ../RTL/cortexm0ds_logic.v(2278)
  not u3580 (Maaiu6, n664);  // ../RTL/cortexm0ds_logic.v(4985)
  AL_MUX u3581 (
    .i0(Abaiu6),
    .i1(Hbaiu6),
    .sel(Cyfpw6[3]),
    .o(G7aiu6));  // ../RTL/cortexm0ds_logic.v(4986)
  and u3582 (n665, Obaiu6, Vbaiu6);  // ../RTL/cortexm0ds_logic.v(4987)
  not u3583 (Hbaiu6, n665);  // ../RTL/cortexm0ds_logic.v(4987)
  or u3584 (n666, R2aiu6, D7fpw6[0]);  // ../RTL/cortexm0ds_logic.v(4988)
  not u3585 (Vbaiu6, n666);  // ../RTL/cortexm0ds_logic.v(4988)
  or u3586 (n667, Ccaiu6, V4aiu6);  // ../RTL/cortexm0ds_logic.v(4989)
  not u3587 (Obaiu6, n667);  // ../RTL/cortexm0ds_logic.v(4989)
  or u3588 (Abaiu6, Rb8iu6, Jcaiu6);  // ../RTL/cortexm0ds_logic.v(4990)
  AL_MUX u3589 (
    .i0(Qcaiu6),
    .i1(vis_r1_o[2]),
    .sel(Mx8iu6),
    .o(I9vhu6));  // ../RTL/cortexm0ds_logic.v(4991)
  buf u359 (vis_r3_o[29], No5bx6);  // ../RTL/cortexm0ds_logic.v(2694)
  AL_MUX u3590 (
    .i0(Qcaiu6),
    .i1(vis_r0_o[2]),
    .sel(Lf8iu6),
    .o(B9vhu6));  // ../RTL/cortexm0ds_logic.v(4992)
  and u3591 (n668, Xcaiu6, Edaiu6);  // ../RTL/cortexm0ds_logic.v(4993)
  not u3592 (U8vhu6, n668);  // ../RTL/cortexm0ds_logic.v(4993)
  and u3593 (n669, Ldaiu6, Hy8iu6);  // ../RTL/cortexm0ds_logic.v(4994)
  not u3594 (Edaiu6, n669);  // ../RTL/cortexm0ds_logic.v(4994)
  or u3595 (n670, Z18iu6, Sdaiu6);  // ../RTL/cortexm0ds_logic.v(4995)
  not u3596 (Ldaiu6, n670);  // ../RTL/cortexm0ds_logic.v(4995)
  and u3597 (n671, Zdaiu6, Eh6iu6);  // ../RTL/cortexm0ds_logic.v(4996)
  not u3598 (Xcaiu6, n671);  // ../RTL/cortexm0ds_logic.v(4996)
  and u3599 (n672, Geaiu6, Neaiu6);  // ../RTL/cortexm0ds_logic.v(4997)
  buf u36 (vis_r12_o[31], Kqsax6);  // ../RTL/cortexm0ds_logic.v(2599)
  buf u360 (vis_r9_o[31], Qnopw6);  // ../RTL/cortexm0ds_logic.v(1898)
  not u3600 (Zdaiu6, n672);  // ../RTL/cortexm0ds_logic.v(4997)
  and u3601 (n673, V3xhu6, Ueaiu6);  // ../RTL/cortexm0ds_logic.v(4998)
  not u3602 (Neaiu6, n673);  // ../RTL/cortexm0ds_logic.v(4998)
  and u3603 (n674, Bfaiu6, Ifaiu6);  // ../RTL/cortexm0ds_logic.v(4999)
  not u3604 (Ueaiu6, n674);  // ../RTL/cortexm0ds_logic.v(4999)
  and u3605 (Ifaiu6, Pfaiu6, Wfaiu6);  // ../RTL/cortexm0ds_logic.v(5000)
  and u3606 (n675, K2aiu6, Dgaiu6);  // ../RTL/cortexm0ds_logic.v(5001)
  not u3607 (Wfaiu6, n675);  // ../RTL/cortexm0ds_logic.v(5001)
  and u3608 (n676, Kgaiu6, Rgaiu6);  // ../RTL/cortexm0ds_logic.v(5002)
  not u3609 (Dgaiu6, n676);  // ../RTL/cortexm0ds_logic.v(5002)
  buf u361 (vis_r3_o[5], S7yax6);  // ../RTL/cortexm0ds_logic.v(2694)
  and u3610 (n677, Ygaiu6, Fhaiu6);  // ../RTL/cortexm0ds_logic.v(5003)
  not u3611 (Rgaiu6, n677);  // ../RTL/cortexm0ds_logic.v(5003)
  or u3612 (n678, As0iu6, Y7ghu6);  // ../RTL/cortexm0ds_logic.v(5004)
  not u3613 (Ygaiu6, n678);  // ../RTL/cortexm0ds_logic.v(5004)
  and u3614 (Pfaiu6, Mhaiu6, Thaiu6);  // ../RTL/cortexm0ds_logic.v(5005)
  and u3615 (n679, Aiaiu6, Hiaiu6);  // ../RTL/cortexm0ds_logic.v(5006)
  not u3616 (Mhaiu6, n679);  // ../RTL/cortexm0ds_logic.v(5006)
  and u3617 (Aiaiu6, Oiaiu6, Viaiu6);  // ../RTL/cortexm0ds_logic.v(5007)
  and u3618 (n680, Cjaiu6, Jjaiu6);  // ../RTL/cortexm0ds_logic.v(5008)
  not u3619 (Viaiu6, n680);  // ../RTL/cortexm0ds_logic.v(5008)
  buf u362 (vis_r3_o[6], Pe5bx6);  // ../RTL/cortexm0ds_logic.v(2694)
  or u3620 (Jjaiu6, Qjaiu6, Cyfpw6[3]);  // ../RTL/cortexm0ds_logic.v(5009)
  and u3621 (Cjaiu6, Xjaiu6, Ekaiu6);  // ../RTL/cortexm0ds_logic.v(5010)
  or u3622 (Xjaiu6, As0iu6, Lkaiu6);  // ../RTL/cortexm0ds_logic.v(5011)
  and u3623 (Bfaiu6, Skaiu6, Zkaiu6);  // ../RTL/cortexm0ds_logic.v(5012)
  and u3624 (n681, Glaiu6, Nlaiu6);  // ../RTL/cortexm0ds_logic.v(5013)
  not u3625 (Zkaiu6, n681);  // ../RTL/cortexm0ds_logic.v(5013)
  and u3626 (Skaiu6, Ulaiu6, Bmaiu6);  // ../RTL/cortexm0ds_logic.v(5014)
  and u3627 (n682, Imaiu6, Pmaiu6);  // ../RTL/cortexm0ds_logic.v(5015)
  not u3628 (Bmaiu6, n682);  // ../RTL/cortexm0ds_logic.v(5015)
  and u3629 (n683, Wmaiu6, Dnaiu6);  // ../RTL/cortexm0ds_logic.v(5016)
  buf u363 (vis_r3_o[11], C87bx6);  // ../RTL/cortexm0ds_logic.v(2694)
  not u3630 (Pmaiu6, n683);  // ../RTL/cortexm0ds_logic.v(5016)
  or u3631 (Dnaiu6, Knaiu6, Cyfpw6[1]);  // ../RTL/cortexm0ds_logic.v(5017)
  and u3632 (n684, Cyfpw6[7], Rnaiu6);  // ../RTL/cortexm0ds_logic.v(5018)
  not u3633 (Ulaiu6, n684);  // ../RTL/cortexm0ds_logic.v(5018)
  and u3634 (n685, Ynaiu6, Foaiu6);  // ../RTL/cortexm0ds_logic.v(5019)
  not u3635 (Rnaiu6, n685);  // ../RTL/cortexm0ds_logic.v(5019)
  and u3636 (n686, Moaiu6, Ii0iu6);  // ../RTL/cortexm0ds_logic.v(5020)
  not u3637 (Foaiu6, n686);  // ../RTL/cortexm0ds_logic.v(5020)
  and u3638 (n687, Toaiu6, Apaiu6);  // ../RTL/cortexm0ds_logic.v(5021)
  not u3639 (Ynaiu6, n687);  // ../RTL/cortexm0ds_logic.v(5021)
  buf u364 (vis_r3_o[12], Dk6bx6);  // ../RTL/cortexm0ds_logic.v(2694)
  and u3640 (n688, Hpaiu6, Opaiu6);  // ../RTL/cortexm0ds_logic.v(5022)
  not u3641 (N8vhu6, n688);  // ../RTL/cortexm0ds_logic.v(5022)
  and u3642 (n689, Vpaiu6, Xbopw6);  // ../RTL/cortexm0ds_logic.v(5023)
  not u3643 (Opaiu6, n689);  // ../RTL/cortexm0ds_logic.v(5023)
  and u3644 (n690, Jqaiu6, Qqaiu6);  // ../RTL/cortexm0ds_logic.v(5024)
  not u3645 (Vpaiu6, n690);  // ../RTL/cortexm0ds_logic.v(5024)
  and u3646 (Qqaiu6, Xqaiu6, Eraiu6);  // ../RTL/cortexm0ds_logic.v(5025)
  and u3647 (n691, Lraiu6, Ja5iu6);  // ../RTL/cortexm0ds_logic.v(5026)
  not u3648 (Eraiu6, n691);  // ../RTL/cortexm0ds_logic.v(5026)
  and u3649 (Xqaiu6, Sraiu6, Zraiu6);  // ../RTL/cortexm0ds_logic.v(5027)
  buf u365 (vis_r3_o[14], Dg6bx6);  // ../RTL/cortexm0ds_logic.v(2694)
  and u3650 (n692, Gsaiu6, Nsaiu6);  // ../RTL/cortexm0ds_logic.v(5028)
  not u3651 (Sraiu6, n692);  // ../RTL/cortexm0ds_logic.v(5028)
  and u3652 (Jqaiu6, Usaiu6, HREADY);  // ../RTL/cortexm0ds_logic.v(5029)
  and u3653 (n693, SLEEPHOLDREQn, HREADY);  // ../RTL/cortexm0ds_logic.v(5030)
  not u3654 (Hpaiu6, n693);  // ../RTL/cortexm0ds_logic.v(5030)
  and u3655 (n694, Li5iu6, Btaiu6);  // ../RTL/cortexm0ds_logic.v(5031)
  not u3656 (G8vhu6, n694);  // ../RTL/cortexm0ds_logic.v(5031)
  and u3657 (n695, Itaiu6, Righu6);  // ../RTL/cortexm0ds_logic.v(5032)
  not u3658 (Btaiu6, n695);  // ../RTL/cortexm0ds_logic.v(5032)
  or u3659 (n696, Ptaiu6, Qg6iu6);  // ../RTL/cortexm0ds_logic.v(5033)
  buf u366 (vis_r3_o[15], Zx7bx6);  // ../RTL/cortexm0ds_logic.v(2694)
  not u3660 (Itaiu6, n696);  // ../RTL/cortexm0ds_logic.v(5033)
  and u3661 (Li5iu6, Wtaiu6, Duaiu6);  // ../RTL/cortexm0ds_logic.v(5034)
  and u3662 (n697, Kuaiu6, Ruaiu6);  // ../RTL/cortexm0ds_logic.v(5035)
  not u3663 (Duaiu6, n697);  // ../RTL/cortexm0ds_logic.v(5035)
  and u3664 (n698, Yuaiu6, Fvaiu6);  // ../RTL/cortexm0ds_logic.v(5036)
  not u3665 (Kuaiu6, n698);  // ../RTL/cortexm0ds_logic.v(5036)
  and u3666 (Fvaiu6, Mvaiu6, Tvaiu6);  // ../RTL/cortexm0ds_logic.v(5037)
  and u3667 (n699, Awaiu6, Hwaiu6);  // ../RTL/cortexm0ds_logic.v(5038)
  not u3668 (Tvaiu6, n699);  // ../RTL/cortexm0ds_logic.v(5038)
  or u3669 (n700, Owaiu6, Vwaiu6);  // ../RTL/cortexm0ds_logic.v(5039)
  buf u367 (vis_r3_o[17], Dc6bx6);  // ../RTL/cortexm0ds_logic.v(2694)
  not u3670 (Awaiu6, n700);  // ../RTL/cortexm0ds_logic.v(5039)
  and u3671 (n701, Cxaiu6, Jxaiu6);  // ../RTL/cortexm0ds_logic.v(5040)
  not u3672 (Mvaiu6, n701);  // ../RTL/cortexm0ds_logic.v(5040)
  or u3673 (n702, Qxaiu6, D7fpw6[14]);  // ../RTL/cortexm0ds_logic.v(5041)
  not u3674 (Cxaiu6, n702);  // ../RTL/cortexm0ds_logic.v(5041)
  and u3675 (Yuaiu6, Xxaiu6, Eyaiu6);  // ../RTL/cortexm0ds_logic.v(5042)
  and u3676 (n703, Lyaiu6, L3ehu6);  // ../RTL/cortexm0ds_logic.v(5043)
  not u3677 (Eyaiu6, n703);  // ../RTL/cortexm0ds_logic.v(5043)
  and u3678 (Wtaiu6, Syaiu6, Zyaiu6);  // ../RTL/cortexm0ds_logic.v(5044)
  and u3679 (n704, Lyaiu6, Gzaiu6);  // ../RTL/cortexm0ds_logic.v(5045)
  buf u368 (vis_r3_o[18], Da6bx6);  // ../RTL/cortexm0ds_logic.v(2694)
  not u3680 (Zyaiu6, n704);  // ../RTL/cortexm0ds_logic.v(5045)
  or u3681 (n705, Nzaiu6, L3ehu6);  // ../RTL/cortexm0ds_logic.v(5046)
  not u3682 (Gzaiu6, n705);  // ../RTL/cortexm0ds_logic.v(5046)
  and u3683 (Nzaiu6, Uzaiu6, B0biu6);  // ../RTL/cortexm0ds_logic.v(5047)
  or u3684 (n706, K9aiu6, Geaiu6);  // ../RTL/cortexm0ds_logic.v(5048)
  not u3685 (Lyaiu6, n706);  // ../RTL/cortexm0ds_logic.v(5048)
  or u3686 (Syaiu6, I0biu6, P0biu6);  // ../RTL/cortexm0ds_logic.v(5049)
  and u3687 (n707, W0biu6, D1biu6);  // ../RTL/cortexm0ds_logic.v(5050)
  not u3688 (Z7vhu6, n707);  // ../RTL/cortexm0ds_logic.v(5050)
  and u3689 (n708, K1biu6, R1biu6);  // ../RTL/cortexm0ds_logic.v(5051)
  buf u369 (vis_r3_o[20], D66bx6);  // ../RTL/cortexm0ds_logic.v(2694)
  not u3690 (D1biu6, n708);  // ../RTL/cortexm0ds_logic.v(5051)
  or u3691 (n709, Geaiu6, L3ehu6);  // ../RTL/cortexm0ds_logic.v(5052)
  not u3692 (R1biu6, n709);  // ../RTL/cortexm0ds_logic.v(5052)
  and u3693 (K1biu6, Y1biu6, F2biu6);  // ../RTL/cortexm0ds_logic.v(5053)
  AL_MUX u3694 (
    .i0(Quzhu6),
    .i1(M2biu6),
    .sel(Uzaiu6),
    .o(Y1biu6));  // ../RTL/cortexm0ds_logic.v(5054)
  and u3695 (n710, Qwdhu6, T2biu6);  // ../RTL/cortexm0ds_logic.v(5055)
  not u3696 (W0biu6, n710);  // ../RTL/cortexm0ds_logic.v(5055)
  and u3697 (n711, A3biu6, H3biu6);  // ../RTL/cortexm0ds_logic.v(5056)
  not u3698 (S7vhu6, n711);  // ../RTL/cortexm0ds_logic.v(5056)
  and u3699 (H3biu6, O3biu6, V3biu6);  // ../RTL/cortexm0ds_logic.v(5057)
  buf u37 (vis_r1_o[11], C47bx6);  // ../RTL/cortexm0ds_logic.v(1876)
  buf u370 (vis_r3_o[22], Ttebx6);  // ../RTL/cortexm0ds_logic.v(2694)
  and u3700 (n712, HRDATA[0], Pp7iu6);  // ../RTL/cortexm0ds_logic.v(5058)
  not u3701 (V3biu6, n712);  // ../RTL/cortexm0ds_logic.v(5058)
  and u3702 (O3biu6, C4biu6, J4biu6);  // ../RTL/cortexm0ds_logic.v(5059)
  and u3703 (n713, Hrfpw6[0], Uy4iu6);  // ../RTL/cortexm0ds_logic.v(5060)
  not u3704 (J4biu6, n713);  // ../RTL/cortexm0ds_logic.v(5060)
  and u3705 (n714, HRDATA[16], Kq7iu6);  // ../RTL/cortexm0ds_logic.v(5061)
  not u3706 (C4biu6, n714);  // ../RTL/cortexm0ds_logic.v(5061)
  and u3707 (A3biu6, Q4biu6, X4biu6);  // ../RTL/cortexm0ds_logic.v(5062)
  and u3708 (n715, Fr7iu6, T24iu6);  // ../RTL/cortexm0ds_logic.v(5063)
  not u3709 (X4biu6, n715);  // ../RTL/cortexm0ds_logic.v(5063)
  buf u371 (vis_r3_o[23], Vvxax6);  // ../RTL/cortexm0ds_logic.v(2694)
  and u3710 (Q4biu6, E5biu6, L5biu6);  // ../RTL/cortexm0ds_logic.v(5064)
  and u3711 (n716, Ppfpw6[0], A25iu6);  // ../RTL/cortexm0ds_logic.v(5065)
  not u3712 (L5biu6, n716);  // ../RTL/cortexm0ds_logic.v(5065)
  and u3713 (n717, R05iu6, D7fpw6[0]);  // ../RTL/cortexm0ds_logic.v(5066)
  not u3714 (E5biu6, n717);  // ../RTL/cortexm0ds_logic.v(5066)
  AL_MUX u3715 (
    .i0(S5biu6),
    .i1(S8fpw6[1]),
    .sel(F58iu6),
    .o(L7vhu6));  // ../RTL/cortexm0ds_logic.v(5067)
  and u3716 (n718, Z5biu6, G6biu6);  // ../RTL/cortexm0ds_logic.v(5068)
  not u3717 (S5biu6, n718);  // ../RTL/cortexm0ds_logic.v(5068)
  and u3718 (G6biu6, N6biu6, U6biu6);  // ../RTL/cortexm0ds_logic.v(5069)
  and u3719 (U6biu6, B7biu6, V68iu6);  // ../RTL/cortexm0ds_logic.v(5070)
  buf u372 (vis_r3_o[25], Jy5bx6);  // ../RTL/cortexm0ds_logic.v(2694)
  and u3720 (n719, I7biu6, E88iu6);  // ../RTL/cortexm0ds_logic.v(5071)
  not u3721 (B7biu6, n719);  // ../RTL/cortexm0ds_logic.v(5071)
  xor u3722 (I7biu6, P7biu6, W7biu6);  // ../RTL/cortexm0ds_logic.v(5072)
  and u3723 (N6biu6, D8biu6, K8biu6);  // ../RTL/cortexm0ds_logic.v(5073)
  and u3724 (n720, R8biu6, Ce8iu6);  // ../RTL/cortexm0ds_logic.v(5074)
  not u3725 (K8biu6, n720);  // ../RTL/cortexm0ds_logic.v(5074)
  xor u3726 (n721, Y8biu6, S8fpw6[0]);  // ../RTL/cortexm0ds_logic.v(5075)
  not u3727 (R8biu6, n721);  // ../RTL/cortexm0ds_logic.v(5075)
  and u3728 (n722, Tc8iu6, Ppfpw6[1]);  // ../RTL/cortexm0ds_logic.v(5076)
  not u3729 (D8biu6, n722);  // ../RTL/cortexm0ds_logic.v(5076)
  buf u373 (vis_r3_o[26], Nk5bx6);  // ../RTL/cortexm0ds_logic.v(2694)
  and u3730 (Z5biu6, F9biu6, M9biu6);  // ../RTL/cortexm0ds_logic.v(5077)
  and u3731 (M9biu6, T9biu6, Aabiu6);  // ../RTL/cortexm0ds_logic.v(5078)
  or u3732 (Aabiu6, O95iu6, Hd8iu6);  // ../RTL/cortexm0ds_logic.v(5079)
  and u3733 (n723, Habiu6, D7fpw6[0]);  // ../RTL/cortexm0ds_logic.v(5080)
  not u3734 (T9biu6, n723);  // ../RTL/cortexm0ds_logic.v(5080)
  and u3735 (F9biu6, Oabiu6, Vabiu6);  // ../RTL/cortexm0ds_logic.v(5081)
  or u3736 (Vabiu6, Ccaiu6, Yb8iu6);  // ../RTL/cortexm0ds_logic.v(5082)
  and u3737 (n724, Cbbiu6, D7fpw6[6]);  // ../RTL/cortexm0ds_logic.v(5083)
  not u3738 (Oabiu6, n724);  // ../RTL/cortexm0ds_logic.v(5083)
  and u3739 (n725, Jbbiu6, Qbbiu6);  // ../RTL/cortexm0ds_logic.v(5084)
  buf u374 (vis_r3_o[27], Nm5bx6);  // ../RTL/cortexm0ds_logic.v(2694)
  not u3740 (E7vhu6, n725);  // ../RTL/cortexm0ds_logic.v(5084)
  and u3741 (n726, D8hhu6, Xbbiu6);  // ../RTL/cortexm0ds_logic.v(5085)
  not u3742 (Qbbiu6, n726);  // ../RTL/cortexm0ds_logic.v(5085)
  and u3743 (n727, Qw4iu6, Ecbiu6);  // ../RTL/cortexm0ds_logic.v(5086)
  not u3744 (X6vhu6, n727);  // ../RTL/cortexm0ds_logic.v(5086)
  and u3745 (n728, Dhgpw6[1], Lcbiu6);  // ../RTL/cortexm0ds_logic.v(5087)
  not u3746 (Ecbiu6, n728);  // ../RTL/cortexm0ds_logic.v(5087)
  and u3747 (n729, Scbiu6, O34iu6);  // ../RTL/cortexm0ds_logic.v(5088)
  not u3748 (Lcbiu6, n729);  // ../RTL/cortexm0ds_logic.v(5088)
  and u3749 (n730, W8aiu6, Cyfpw6[0]);  // ../RTL/cortexm0ds_logic.v(5089)
  buf u375 (vis_r3_o[28], R9ibx6);  // ../RTL/cortexm0ds_logic.v(2694)
  not u3750 (Qw4iu6, n730);  // ../RTL/cortexm0ds_logic.v(5089)
  and u3751 (Q6vhu6, Zcbiu6, Gdbiu6);  // ../RTL/cortexm0ds_logic.v(5090)
  and u3752 (Gdbiu6, Ndbiu6, Udbiu6);  // ../RTL/cortexm0ds_logic.v(5091)
  and u3753 (n731, Npdpw6, Bebiu6);  // ../RTL/cortexm0ds_logic.v(5092)
  not u3754 (Ndbiu6, n731);  // ../RTL/cortexm0ds_logic.v(5092)
  and u3755 (Zcbiu6, IRQ[31], Iebiu6);  // ../RTL/cortexm0ds_logic.v(5093)
  and u3756 (n732, Tk7iu6, Pebiu6);  // ../RTL/cortexm0ds_logic.v(5094)
  not u3757 (Iebiu6, n732);  // ../RTL/cortexm0ds_logic.v(5094)
  or u3758 (Pebiu6, Webiu6, Qg6iu6);  // ../RTL/cortexm0ds_logic.v(5095)
  and u3759 (J6vhu6, Dfbiu6, Kfbiu6);  // ../RTL/cortexm0ds_logic.v(5096)
  buf u376 (K7hpw6[2], Lx9ax6);  // ../RTL/cortexm0ds_logic.v(2366)
  and u3760 (Kfbiu6, Rfbiu6, Yfbiu6);  // ../RTL/cortexm0ds_logic.v(5097)
  and u3761 (n733, Updpw6, Fgbiu6);  // ../RTL/cortexm0ds_logic.v(5098)
  not u3762 (Rfbiu6, n733);  // ../RTL/cortexm0ds_logic.v(5098)
  and u3763 (Dfbiu6, IRQ[29], Mgbiu6);  // ../RTL/cortexm0ds_logic.v(5099)
  and u3764 (n734, Tk7iu6, Tgbiu6);  // ../RTL/cortexm0ds_logic.v(5100)
  not u3765 (Mgbiu6, n734);  // ../RTL/cortexm0ds_logic.v(5100)
  or u3766 (Tgbiu6, Qg6iu6, Ahbiu6);  // ../RTL/cortexm0ds_logic.v(5101)
  and u3767 (n735, Hhbiu6, Ohbiu6);  // ../RTL/cortexm0ds_logic.v(5102)
  not u3768 (C6vhu6, n735);  // ../RTL/cortexm0ds_logic.v(5102)
  or u3769 (Ohbiu6, Vhbiu6, Cibiu6);  // ../RTL/cortexm0ds_logic.v(5103)
  buf u377 (vis_r9_o[30], Qlopw6);  // ../RTL/cortexm0ds_logic.v(1898)
  and u3770 (Hhbiu6, Jibiu6, Qibiu6);  // ../RTL/cortexm0ds_logic.v(5104)
  and u3771 (n736, Xibiu6, Ppfpw6[5]);  // ../RTL/cortexm0ds_logic.v(5105)
  not u3772 (Qibiu6, n736);  // ../RTL/cortexm0ds_logic.v(5105)
  or u3773 (Jibiu6, Ejbiu6, Ljbiu6);  // ../RTL/cortexm0ds_logic.v(5106)
  and u3774 (n737, Sjbiu6, Zjbiu6);  // ../RTL/cortexm0ds_logic.v(5107)
  not u3775 (V5vhu6, n737);  // ../RTL/cortexm0ds_logic.v(5107)
  and u3776 (Zjbiu6, Gkbiu6, Nkbiu6);  // ../RTL/cortexm0ds_logic.v(5108)
  and u3777 (n738, HRDATA[8], Pp7iu6);  // ../RTL/cortexm0ds_logic.v(5109)
  not u3778 (Nkbiu6, n738);  // ../RTL/cortexm0ds_logic.v(5109)
  and u3779 (Gkbiu6, Ukbiu6, Blbiu6);  // ../RTL/cortexm0ds_logic.v(5110)
  buf u378 (E1hpw6[2], Bvaax6);  // ../RTL/cortexm0ds_logic.v(2367)
  and u3780 (n739, Hrfpw6[8], Uy4iu6);  // ../RTL/cortexm0ds_logic.v(5111)
  not u3781 (Blbiu6, n739);  // ../RTL/cortexm0ds_logic.v(5111)
  and u3782 (n740, HRDATA[24], Kq7iu6);  // ../RTL/cortexm0ds_logic.v(5112)
  not u3783 (Ukbiu6, n740);  // ../RTL/cortexm0ds_logic.v(5112)
  and u3784 (Sjbiu6, Ilbiu6, Plbiu6);  // ../RTL/cortexm0ds_logic.v(5113)
  and u3785 (n741, A25iu6, Ppfpw6[8]);  // ../RTL/cortexm0ds_logic.v(5114)
  not u3786 (Plbiu6, n741);  // ../RTL/cortexm0ds_logic.v(5114)
  and u3787 (n742, D7fpw6[8], R05iu6);  // ../RTL/cortexm0ds_logic.v(5115)
  not u3788 (Ilbiu6, n742);  // ../RTL/cortexm0ds_logic.v(5115)
  and u3789 (n743, Wlbiu6, Dmbiu6);  // ../RTL/cortexm0ds_logic.v(5116)
  buf u379 (vis_r9_o[29], Ovopw6);  // ../RTL/cortexm0ds_logic.v(1898)
  not u3790 (O5vhu6, n743);  // ../RTL/cortexm0ds_logic.v(5116)
  or u3791 (Dmbiu6, Jm7iu6, Kmbiu6);  // ../RTL/cortexm0ds_logic.v(5117)
  and u3792 (Wlbiu6, Rmbiu6, Ymbiu6);  // ../RTL/cortexm0ds_logic.v(5118)
  and u3793 (n744, Ppfpw6[0], Fnbiu6);  // ../RTL/cortexm0ds_logic.v(5119)
  not u3794 (Ymbiu6, n744);  // ../RTL/cortexm0ds_logic.v(5119)
  and u3795 (n745, Mnbiu6, HRDATA[0]);  // ../RTL/cortexm0ds_logic.v(5120)
  not u3796 (Rmbiu6, n745);  // ../RTL/cortexm0ds_logic.v(5120)
  and u3797 (n746, Tnbiu6, Aobiu6);  // ../RTL/cortexm0ds_logic.v(5121)
  not u3798 (H5vhu6, n746);  // ../RTL/cortexm0ds_logic.v(5121)
  and u3799 (n747, Hobiu6, Kw8iu6);  // ../RTL/cortexm0ds_logic.v(5122)
  buf u38 (H6ghu6, Vgjpw6);  // ../RTL/cortexm0ds_logic.v(1799)
  buf u380 (Kohhu6, H4bax6);  // ../RTL/cortexm0ds_logic.v(2270)
  not u3800 (Aobiu6, n747);  // ../RTL/cortexm0ds_logic.v(5122)
  and u3801 (n748, Svdpw6, Oobiu6);  // ../RTL/cortexm0ds_logic.v(5123)
  not u3802 (Kw8iu6, n748);  // ../RTL/cortexm0ds_logic.v(5123)
  and u3803 (n749, HRDATA[14], Vobiu6);  // ../RTL/cortexm0ds_logic.v(5124)
  not u3804 (Oobiu6, n749);  // ../RTL/cortexm0ds_logic.v(5124)
  and u3805 (n750, Ppfpw6[14], Cpbiu6);  // ../RTL/cortexm0ds_logic.v(5125)
  not u3806 (Tnbiu6, n750);  // ../RTL/cortexm0ds_logic.v(5125)
  and u3807 (n751, Jpbiu6, Qpbiu6);  // ../RTL/cortexm0ds_logic.v(5126)
  not u3808 (A5vhu6, n751);  // ../RTL/cortexm0ds_logic.v(5126)
  and u3809 (Qpbiu6, Xpbiu6, Eqbiu6);  // ../RTL/cortexm0ds_logic.v(5127)
  buf u381 (vis_r9_o[27], Otopw6);  // ../RTL/cortexm0ds_logic.v(1898)
  and u3810 (n752, Xlfpw6[8], Lqbiu6);  // ../RTL/cortexm0ds_logic.v(5128)
  not u3811 (Eqbiu6, n752);  // ../RTL/cortexm0ds_logic.v(5128)
  and u3812 (n753, IRQLATENCY[7], Ol7iu6);  // ../RTL/cortexm0ds_logic.v(5129)
  not u3813 (Xpbiu6, n753);  // ../RTL/cortexm0ds_logic.v(5129)
  and u3814 (Jpbiu6, Sqbiu6, Zqbiu6);  // ../RTL/cortexm0ds_logic.v(5130)
  and u3815 (n754, Mnbiu6, HRDATA[13]);  // ../RTL/cortexm0ds_logic.v(5131)
  not u3816 (Zqbiu6, n754);  // ../RTL/cortexm0ds_logic.v(5131)
  and u3817 (n755, Cpbiu6, Ppfpw6[13]);  // ../RTL/cortexm0ds_logic.v(5132)
  not u3818 (Sqbiu6, n755);  // ../RTL/cortexm0ds_logic.v(5132)
  and u3819 (n756, Grbiu6, Nrbiu6);  // ../RTL/cortexm0ds_logic.v(5133)
  buf u382 (vis_r9_o[26], Xxtpw6);  // ../RTL/cortexm0ds_logic.v(1898)
  not u3820 (T4vhu6, n756);  // ../RTL/cortexm0ds_logic.v(5133)
  and u3821 (Nrbiu6, Urbiu6, Bsbiu6);  // ../RTL/cortexm0ds_logic.v(5134)
  and u3822 (n757, Xlfpw6[7], Lqbiu6);  // ../RTL/cortexm0ds_logic.v(5135)
  not u3823 (Bsbiu6, n757);  // ../RTL/cortexm0ds_logic.v(5135)
  and u3824 (n758, IRQLATENCY[6], Ol7iu6);  // ../RTL/cortexm0ds_logic.v(5136)
  not u3825 (Urbiu6, n758);  // ../RTL/cortexm0ds_logic.v(5136)
  and u3826 (Grbiu6, Isbiu6, Psbiu6);  // ../RTL/cortexm0ds_logic.v(5137)
  and u3827 (n759, Mnbiu6, HRDATA[12]);  // ../RTL/cortexm0ds_logic.v(5138)
  not u3828 (Psbiu6, n759);  // ../RTL/cortexm0ds_logic.v(5138)
  and u3829 (n760, Cpbiu6, Ppfpw6[12]);  // ../RTL/cortexm0ds_logic.v(5139)
  buf u383 (vis_r9_o[25], Z5tpw6);  // ../RTL/cortexm0ds_logic.v(1898)
  not u3830 (Isbiu6, n760);  // ../RTL/cortexm0ds_logic.v(5139)
  and u3831 (n761, Wsbiu6, Dtbiu6);  // ../RTL/cortexm0ds_logic.v(5140)
  not u3832 (M4vhu6, n761);  // ../RTL/cortexm0ds_logic.v(5140)
  and u3833 (Dtbiu6, Ktbiu6, Rtbiu6);  // ../RTL/cortexm0ds_logic.v(5141)
  and u3834 (n762, Xlfpw6[6], Lqbiu6);  // ../RTL/cortexm0ds_logic.v(5142)
  not u3835 (Rtbiu6, n762);  // ../RTL/cortexm0ds_logic.v(5142)
  and u3836 (n763, IRQLATENCY[5], Ol7iu6);  // ../RTL/cortexm0ds_logic.v(5143)
  not u3837 (Ktbiu6, n763);  // ../RTL/cortexm0ds_logic.v(5143)
  and u3838 (Wsbiu6, Ytbiu6, Fubiu6);  // ../RTL/cortexm0ds_logic.v(5144)
  and u3839 (n764, HRDATA[11], Mnbiu6);  // ../RTL/cortexm0ds_logic.v(5145)
  buf u384 (G4hpw6[0], Pkkbx6);  // ../RTL/cortexm0ds_logic.v(2274)
  not u3840 (Fubiu6, n764);  // ../RTL/cortexm0ds_logic.v(5145)
  and u3841 (n765, Cpbiu6, Ppfpw6[11]);  // ../RTL/cortexm0ds_logic.v(5146)
  not u3842 (Ytbiu6, n765);  // ../RTL/cortexm0ds_logic.v(5146)
  and u3843 (n766, Mubiu6, Tubiu6);  // ../RTL/cortexm0ds_logic.v(5147)
  not u3844 (F4vhu6, n766);  // ../RTL/cortexm0ds_logic.v(5147)
  and u3845 (Tubiu6, Avbiu6, Hvbiu6);  // ../RTL/cortexm0ds_logic.v(5148)
  and u3846 (n767, Xlfpw6[5], Lqbiu6);  // ../RTL/cortexm0ds_logic.v(5149)
  not u3847 (Hvbiu6, n767);  // ../RTL/cortexm0ds_logic.v(5149)
  and u3848 (n768, IRQLATENCY[4], Ol7iu6);  // ../RTL/cortexm0ds_logic.v(5150)
  not u3849 (Avbiu6, n768);  // ../RTL/cortexm0ds_logic.v(5150)
  buf u385 (vis_r7_o[1], Mbwax6);  // ../RTL/cortexm0ds_logic.v(2654)
  and u3850 (Mubiu6, Ovbiu6, Vvbiu6);  // ../RTL/cortexm0ds_logic.v(5151)
  and u3851 (n769, Mnbiu6, HRDATA[10]);  // ../RTL/cortexm0ds_logic.v(5152)
  not u3852 (Vvbiu6, n769);  // ../RTL/cortexm0ds_logic.v(5152)
  and u3853 (n770, Cpbiu6, Ppfpw6[10]);  // ../RTL/cortexm0ds_logic.v(5153)
  not u3854 (Ovbiu6, n770);  // ../RTL/cortexm0ds_logic.v(5153)
  and u3855 (n771, Cwbiu6, Jwbiu6);  // ../RTL/cortexm0ds_logic.v(5154)
  not u3856 (Y3vhu6, n771);  // ../RTL/cortexm0ds_logic.v(5154)
  and u3857 (Jwbiu6, Qwbiu6, Xwbiu6);  // ../RTL/cortexm0ds_logic.v(5155)
  and u3858 (n772, Xlfpw6[4], Lqbiu6);  // ../RTL/cortexm0ds_logic.v(5156)
  not u3859 (Xwbiu6, n772);  // ../RTL/cortexm0ds_logic.v(5156)
  buf u386 (vis_r3_o[31], Vzxax6);  // ../RTL/cortexm0ds_logic.v(2694)
  and u3860 (n773, IRQLATENCY[3], Ol7iu6);  // ../RTL/cortexm0ds_logic.v(5157)
  not u3861 (Qwbiu6, n773);  // ../RTL/cortexm0ds_logic.v(5157)
  and u3862 (Cwbiu6, Exbiu6, Lxbiu6);  // ../RTL/cortexm0ds_logic.v(5158)
  and u3863 (n774, HRDATA[9], Mnbiu6);  // ../RTL/cortexm0ds_logic.v(5159)
  not u3864 (Lxbiu6, n774);  // ../RTL/cortexm0ds_logic.v(5159)
  and u3865 (n775, Cpbiu6, Ppfpw6[9]);  // ../RTL/cortexm0ds_logic.v(5160)
  not u3866 (Exbiu6, n775);  // ../RTL/cortexm0ds_logic.v(5160)
  and u3867 (n776, Sxbiu6, Zxbiu6);  // ../RTL/cortexm0ds_logic.v(5161)
  not u3868 (R3vhu6, n776);  // ../RTL/cortexm0ds_logic.v(5161)
  and u3869 (Zxbiu6, Gybiu6, Nybiu6);  // ../RTL/cortexm0ds_logic.v(5162)
  buf u387 (vis_r3_o[30], Vxxax6);  // ../RTL/cortexm0ds_logic.v(2694)
  and u3870 (n777, Xlfpw6[3], Lqbiu6);  // ../RTL/cortexm0ds_logic.v(5163)
  not u3871 (Nybiu6, n777);  // ../RTL/cortexm0ds_logic.v(5163)
  and u3872 (n778, IRQLATENCY[2], Ol7iu6);  // ../RTL/cortexm0ds_logic.v(5164)
  not u3873 (Gybiu6, n778);  // ../RTL/cortexm0ds_logic.v(5164)
  and u3874 (Sxbiu6, Uybiu6, Bzbiu6);  // ../RTL/cortexm0ds_logic.v(5165)
  and u3875 (n779, Mnbiu6, HRDATA[8]);  // ../RTL/cortexm0ds_logic.v(5166)
  not u3876 (Bzbiu6, n779);  // ../RTL/cortexm0ds_logic.v(5166)
  and u3877 (n780, Cpbiu6, Ppfpw6[8]);  // ../RTL/cortexm0ds_logic.v(5167)
  not u3878 (Uybiu6, n780);  // ../RTL/cortexm0ds_logic.v(5167)
  and u3879 (n781, Izbiu6, Pzbiu6);  // ../RTL/cortexm0ds_logic.v(5168)
  buf u388 (V5hpw6[0], N39ax6);  // ../RTL/cortexm0ds_logic.v(2248)
  not u3880 (K3vhu6, n781);  // ../RTL/cortexm0ds_logic.v(5168)
  and u3881 (Pzbiu6, Wzbiu6, D0ciu6);  // ../RTL/cortexm0ds_logic.v(5169)
  and u3882 (n782, Xlfpw6[2], Lqbiu6);  // ../RTL/cortexm0ds_logic.v(5170)
  not u3883 (D0ciu6, n782);  // ../RTL/cortexm0ds_logic.v(5170)
  and u3884 (n783, IRQLATENCY[1], Ol7iu6);  // ../RTL/cortexm0ds_logic.v(5171)
  not u3885 (Wzbiu6, n783);  // ../RTL/cortexm0ds_logic.v(5171)
  and u3886 (Izbiu6, K0ciu6, R0ciu6);  // ../RTL/cortexm0ds_logic.v(5172)
  and u3887 (n784, Mnbiu6, HRDATA[7]);  // ../RTL/cortexm0ds_logic.v(5173)
  not u3888 (R0ciu6, n784);  // ../RTL/cortexm0ds_logic.v(5173)
  and u3889 (n785, Cpbiu6, Ppfpw6[7]);  // ../RTL/cortexm0ds_logic.v(5174)
  buf u389 (Gqgpw6[21], Acebx6);  // ../RTL/cortexm0ds_logic.v(2377)
  not u3890 (K0ciu6, n785);  // ../RTL/cortexm0ds_logic.v(5174)
  and u3891 (n786, Y0ciu6, F1ciu6);  // ../RTL/cortexm0ds_logic.v(5175)
  not u3892 (D3vhu6, n786);  // ../RTL/cortexm0ds_logic.v(5175)
  and u3893 (F1ciu6, M1ciu6, T1ciu6);  // ../RTL/cortexm0ds_logic.v(5176)
  and u3894 (n787, Xlfpw6[1], Lqbiu6);  // ../RTL/cortexm0ds_logic.v(5177)
  not u3895 (T1ciu6, n787);  // ../RTL/cortexm0ds_logic.v(5177)
  or u3896 (n788, Ol7iu6, A2ciu6);  // ../RTL/cortexm0ds_logic.v(5178)
  not u3897 (Lqbiu6, n788);  // ../RTL/cortexm0ds_logic.v(5178)
  and u3898 (n789, IRQLATENCY[0], Ol7iu6);  // ../RTL/cortexm0ds_logic.v(5179)
  not u3899 (M1ciu6, n789);  // ../RTL/cortexm0ds_logic.v(5179)
  buf u39 (vis_r1_o[12], I7qpw6);  // ../RTL/cortexm0ds_logic.v(1876)
  buf u390 (Pzgpw6[0], D1aax6);  // ../RTL/cortexm0ds_logic.v(2266)
  and u3900 (Ol7iu6, H2ciu6, O2ciu6);  // ../RTL/cortexm0ds_logic.v(5180)
  and u3901 (n790, V2ciu6, C3ciu6);  // ../RTL/cortexm0ds_logic.v(5181)
  not u3902 (O2ciu6, n790);  // ../RTL/cortexm0ds_logic.v(5181)
  and u3903 (C3ciu6, J3ciu6, Q3ciu6);  // ../RTL/cortexm0ds_logic.v(5182)
  and u3904 (Q3ciu6, Ivfhu6, X3ciu6);  // ../RTL/cortexm0ds_logic.v(5183)
  xor u3905 (n791, Ppfpw6[1], E4ciu6);  // ../RTL/cortexm0ds_logic.v(5184)
  not u3906 (X3ciu6, n791);  // ../RTL/cortexm0ds_logic.v(5184)
  and u3907 (J3ciu6, L4ciu6, S4ciu6);  // ../RTL/cortexm0ds_logic.v(5185)
  xor u3908 (S4ciu6, Z4ciu6, Ppfpw6[4]);  // ../RTL/cortexm0ds_logic.v(5186)
  xor u3909 (L4ciu6, Kmbiu6, Ppfpw6[0]);  // ../RTL/cortexm0ds_logic.v(5187)
  buf u391 (Gqgpw6[22], Hrfbx6);  // ../RTL/cortexm0ds_logic.v(2377)
  and u3910 (V2ciu6, G5ciu6, N5ciu6);  // ../RTL/cortexm0ds_logic.v(5188)
  xor u3911 (N5ciu6, U5ciu6, Ppfpw6[2]);  // ../RTL/cortexm0ds_logic.v(5189)
  and u3912 (G5ciu6, B6ciu6, I6ciu6);  // ../RTL/cortexm0ds_logic.v(5190)
  xor u3913 (I6ciu6, P6ciu6, Ppfpw6[3]);  // ../RTL/cortexm0ds_logic.v(5191)
  xor u3914 (B6ciu6, W6ciu6, Ppfpw6[5]);  // ../RTL/cortexm0ds_logic.v(5192)
  and u3915 (Y0ciu6, D7ciu6, K7ciu6);  // ../RTL/cortexm0ds_logic.v(5193)
  and u3916 (n792, Mnbiu6, HRDATA[6]);  // ../RTL/cortexm0ds_logic.v(5194)
  not u3917 (K7ciu6, n792);  // ../RTL/cortexm0ds_logic.v(5194)
  and u3918 (n793, Cpbiu6, Ppfpw6[6]);  // ../RTL/cortexm0ds_logic.v(5195)
  not u3919 (D7ciu6, n793);  // ../RTL/cortexm0ds_logic.v(5195)
  buf u392 (vis_msp_o[23], T40qw6);  // ../RTL/cortexm0ds_logic.v(2097)
  and u3920 (n794, R7ciu6, Y7ciu6);  // ../RTL/cortexm0ds_logic.v(5196)
  not u3921 (W2vhu6, n794);  // ../RTL/cortexm0ds_logic.v(5196)
  and u3922 (n795, vis_ipsr_o[0], F8ciu6);  // ../RTL/cortexm0ds_logic.v(5197)
  not u3923 (Y7ciu6, n795);  // ../RTL/cortexm0ds_logic.v(5197)
  and u3924 (R7ciu6, M8ciu6, T8ciu6);  // ../RTL/cortexm0ds_logic.v(5198)
  and u3925 (n796, Xibiu6, Ppfpw6[0]);  // ../RTL/cortexm0ds_logic.v(5199)
  not u3926 (T8ciu6, n796);  // ../RTL/cortexm0ds_logic.v(5199)
  or u3927 (M8ciu6, Ejbiu6, Zt8iu6);  // ../RTL/cortexm0ds_logic.v(5200)
  and u3928 (n797, A9ciu6, H9ciu6);  // ../RTL/cortexm0ds_logic.v(5201)
  not u3929 (P2vhu6, n797);  // ../RTL/cortexm0ds_logic.v(5201)
  buf u393 (Gqgpw6[16], Hsdax6);  // ../RTL/cortexm0ds_logic.v(2377)
  and u3930 (n798, O9ciu6, H2ciu6);  // ../RTL/cortexm0ds_logic.v(5202)
  not u3931 (H9ciu6, n798);  // ../RTL/cortexm0ds_logic.v(5202)
  and u3932 (O9ciu6, HREADY, V9ciu6);  // ../RTL/cortexm0ds_logic.v(5203)
  and u3933 (n799, Fvdhu6, Caciu6);  // ../RTL/cortexm0ds_logic.v(5204)
  not u3934 (A9ciu6, n799);  // ../RTL/cortexm0ds_logic.v(5204)
  and u3935 (n800, HREADY, Jaciu6);  // ../RTL/cortexm0ds_logic.v(5205)
  not u3936 (Caciu6, n800);  // ../RTL/cortexm0ds_logic.v(5205)
  and u3937 (n801, Gc5iu6, V9ciu6);  // ../RTL/cortexm0ds_logic.v(5206)
  not u3938 (Jaciu6, n801);  // ../RTL/cortexm0ds_logic.v(5206)
  or u3939 (V9ciu6, Uzaiu6, Qaciu6);  // ../RTL/cortexm0ds_logic.v(5207)
  buf u394 (vis_r7_o[31], Rrvax6);  // ../RTL/cortexm0ds_logic.v(2654)
  and u3940 (n802, Xaciu6, Ebciu6);  // ../RTL/cortexm0ds_logic.v(5208)
  not u3941 (I2vhu6, n802);  // ../RTL/cortexm0ds_logic.v(5208)
  or u3942 (Ebciu6, Jm7iu6, W6ciu6);  // ../RTL/cortexm0ds_logic.v(5209)
  and u3943 (Xaciu6, Lbciu6, Sbciu6);  // ../RTL/cortexm0ds_logic.v(5210)
  and u3944 (n803, Ppfpw6[5], Fnbiu6);  // ../RTL/cortexm0ds_logic.v(5211)
  not u3945 (Sbciu6, n803);  // ../RTL/cortexm0ds_logic.v(5211)
  and u3946 (n804, Mnbiu6, HRDATA[5]);  // ../RTL/cortexm0ds_logic.v(5212)
  not u3947 (Lbciu6, n804);  // ../RTL/cortexm0ds_logic.v(5212)
  and u3948 (n805, Zbciu6, Gcciu6);  // ../RTL/cortexm0ds_logic.v(5213)
  not u3949 (B2vhu6, n805);  // ../RTL/cortexm0ds_logic.v(5213)
  buf u395 (vis_msp_o[1], Xozpw6);  // ../RTL/cortexm0ds_logic.v(2097)
  or u3950 (Gcciu6, Jm7iu6, Z4ciu6);  // ../RTL/cortexm0ds_logic.v(5214)
  and u3951 (Zbciu6, Ncciu6, Ucciu6);  // ../RTL/cortexm0ds_logic.v(5215)
  and u3952 (n806, Ppfpw6[4], Fnbiu6);  // ../RTL/cortexm0ds_logic.v(5216)
  not u3953 (Ucciu6, n806);  // ../RTL/cortexm0ds_logic.v(5216)
  and u3954 (n807, Mnbiu6, HRDATA[4]);  // ../RTL/cortexm0ds_logic.v(5217)
  not u3955 (Ncciu6, n807);  // ../RTL/cortexm0ds_logic.v(5217)
  and u3956 (n808, Bdciu6, Idciu6);  // ../RTL/cortexm0ds_logic.v(5218)
  not u3957 (U1vhu6, n808);  // ../RTL/cortexm0ds_logic.v(5218)
  or u3958 (Idciu6, Jm7iu6, P6ciu6);  // ../RTL/cortexm0ds_logic.v(5219)
  and u3959 (Bdciu6, Pdciu6, Wdciu6);  // ../RTL/cortexm0ds_logic.v(5220)
  buf u396 (vis_msp_o[6], So0qw6);  // ../RTL/cortexm0ds_logic.v(2097)
  and u3960 (n809, Ppfpw6[3], Fnbiu6);  // ../RTL/cortexm0ds_logic.v(5221)
  not u3961 (Wdciu6, n809);  // ../RTL/cortexm0ds_logic.v(5221)
  and u3962 (n810, HRDATA[3], Mnbiu6);  // ../RTL/cortexm0ds_logic.v(5222)
  not u3963 (Pdciu6, n810);  // ../RTL/cortexm0ds_logic.v(5222)
  and u3964 (n811, Deciu6, Keciu6);  // ../RTL/cortexm0ds_logic.v(5223)
  not u3965 (N1vhu6, n811);  // ../RTL/cortexm0ds_logic.v(5223)
  or u3966 (Keciu6, Jm7iu6, U5ciu6);  // ../RTL/cortexm0ds_logic.v(5224)
  and u3967 (Deciu6, Reciu6, Yeciu6);  // ../RTL/cortexm0ds_logic.v(5225)
  and u3968 (n812, Ppfpw6[2], Fnbiu6);  // ../RTL/cortexm0ds_logic.v(5226)
  not u3969 (Yeciu6, n812);  // ../RTL/cortexm0ds_logic.v(5226)
  buf u397 (vis_msp_o[7], Pzibx6);  // ../RTL/cortexm0ds_logic.v(2097)
  and u3970 (n813, Mnbiu6, HRDATA[2]);  // ../RTL/cortexm0ds_logic.v(5227)
  not u3971 (Reciu6, n813);  // ../RTL/cortexm0ds_logic.v(5227)
  and u3972 (n814, Ffciu6, Mfciu6);  // ../RTL/cortexm0ds_logic.v(5228)
  not u3973 (G1vhu6, n814);  // ../RTL/cortexm0ds_logic.v(5228)
  or u3974 (Mfciu6, Tfciu6, Cibiu6);  // ../RTL/cortexm0ds_logic.v(5229)
  and u3975 (Ffciu6, Agciu6, Hgciu6);  // ../RTL/cortexm0ds_logic.v(5230)
  and u3976 (n815, Xibiu6, Ppfpw6[2]);  // ../RTL/cortexm0ds_logic.v(5231)
  not u3977 (Hgciu6, n815);  // ../RTL/cortexm0ds_logic.v(5231)
  or u3978 (Agciu6, Ejbiu6, Ogciu6);  // ../RTL/cortexm0ds_logic.v(5232)
  and u3979 (n816, Vgciu6, Chciu6);  // ../RTL/cortexm0ds_logic.v(5233)
  buf u398 (vis_msp_o[9], Zr8bx6);  // ../RTL/cortexm0ds_logic.v(2097)
  not u3980 (Z0vhu6, n816);  // ../RTL/cortexm0ds_logic.v(5233)
  and u3981 (n817, H2ciu6, E4ciu6);  // ../RTL/cortexm0ds_logic.v(5234)
  not u3982 (Chciu6, n817);  // ../RTL/cortexm0ds_logic.v(5234)
  and u3983 (Vgciu6, Jhciu6, Qhciu6);  // ../RTL/cortexm0ds_logic.v(5235)
  and u3984 (n818, Ppfpw6[1], Fnbiu6);  // ../RTL/cortexm0ds_logic.v(5236)
  not u3985 (Qhciu6, n818);  // ../RTL/cortexm0ds_logic.v(5236)
  and u3986 (n819, Zn7iu6, Xhciu6);  // ../RTL/cortexm0ds_logic.v(5237)
  not u3987 (Fnbiu6, n819);  // ../RTL/cortexm0ds_logic.v(5237)
  or u3988 (Xhciu6, A2ciu6, H2ciu6);  // ../RTL/cortexm0ds_logic.v(5238)
  and u3989 (n820, HRDATA[1], Mnbiu6);  // ../RTL/cortexm0ds_logic.v(5239)
  buf u399 (vis_msp_o[10], Tk0qw6);  // ../RTL/cortexm0ds_logic.v(2097)
  not u3990 (Jhciu6, n820);  // ../RTL/cortexm0ds_logic.v(5239)
  and u3991 (Mnbiu6, Hobiu6, Go7iu6);  // ../RTL/cortexm0ds_logic.v(5240)
  and u3992 (n821, Eiciu6, Liciu6);  // ../RTL/cortexm0ds_logic.v(5241)
  not u3993 (S0vhu6, n821);  // ../RTL/cortexm0ds_logic.v(5241)
  or u3994 (Liciu6, Siciu6, Cibiu6);  // ../RTL/cortexm0ds_logic.v(5242)
  and u3995 (Eiciu6, Ziciu6, Gjciu6);  // ../RTL/cortexm0ds_logic.v(5243)
  and u3996 (n822, Xibiu6, Ppfpw6[1]);  // ../RTL/cortexm0ds_logic.v(5244)
  not u3997 (Gjciu6, n822);  // ../RTL/cortexm0ds_logic.v(5244)
  or u3998 (Ziciu6, Ejbiu6, Njciu6);  // ../RTL/cortexm0ds_logic.v(5245)
  or u3999 (L0vhu6, Hobiu6, Ujciu6);  // ../RTL/cortexm0ds_logic.v(5246)
  buf u4 (HPROT[1], 1'b1);  // ../RTL/cortexm0ds_logic.v(1724)
  buf u40 (vis_r0_o[25], Z1tpw6);  // ../RTL/cortexm0ds_logic.v(1875)
  buf u400 (vis_msp_o[12], S78ax6);  // ../RTL/cortexm0ds_logic.v(2097)
  and u4000 (Ujciu6, Bkciu6, Ikciu6);  // ../RTL/cortexm0ds_logic.v(5247)
  and u4001 (Ikciu6, Ntfhu6, Pkciu6);  // ../RTL/cortexm0ds_logic.v(5248)
  and u4002 (Bkciu6, Cpbiu6, R05iu6);  // ../RTL/cortexm0ds_logic.v(5249)
  or u4003 (n823, Ln7iu6, Cpbiu6);  // ../RTL/cortexm0ds_logic.v(5250)
  not u4004 (Hobiu6, n823);  // ../RTL/cortexm0ds_logic.v(5250)
  and u4005 (n824, Wkciu6, Dlciu6);  // ../RTL/cortexm0ds_logic.v(5252)
  not u4006 (E0vhu6, n824);  // ../RTL/cortexm0ds_logic.v(5252)
  and u4007 (Dlciu6, Klciu6, Rlciu6);  // ../RTL/cortexm0ds_logic.v(5253)
  and u4008 (n825, HRDATA[12], Pp7iu6);  // ../RTL/cortexm0ds_logic.v(5254)
  not u4009 (Rlciu6, n825);  // ../RTL/cortexm0ds_logic.v(5254)
  buf u401 (vis_msp_o[13], Zj8bx6);  // ../RTL/cortexm0ds_logic.v(2097)
  and u4010 (Klciu6, Ylciu6, Fmciu6);  // ../RTL/cortexm0ds_logic.v(5255)
  and u4011 (n826, Hrfpw6[12], Uy4iu6);  // ../RTL/cortexm0ds_logic.v(5256)
  not u4012 (Fmciu6, n826);  // ../RTL/cortexm0ds_logic.v(5256)
  and u4013 (n827, HRDATA[28], Kq7iu6);  // ../RTL/cortexm0ds_logic.v(5257)
  not u4014 (Ylciu6, n827);  // ../RTL/cortexm0ds_logic.v(5257)
  and u4015 (Wkciu6, Mmciu6, Tmciu6);  // ../RTL/cortexm0ds_logic.v(5258)
  and u4016 (n828, A25iu6, Ppfpw6[12]);  // ../RTL/cortexm0ds_logic.v(5259)
  not u4017 (Tmciu6, n828);  // ../RTL/cortexm0ds_logic.v(5259)
  and u4018 (n829, R05iu6, D7fpw6[12]);  // ../RTL/cortexm0ds_logic.v(5260)
  not u4019 (Mmciu6, n829);  // ../RTL/cortexm0ds_logic.v(5260)
  buf u402 (vis_msp_o[15], Te0qw6);  // ../RTL/cortexm0ds_logic.v(2097)
  and u4020 (n830, Anciu6, Hnciu6);  // ../RTL/cortexm0ds_logic.v(5261)
  not u4021 (Xzuhu6, n830);  // ../RTL/cortexm0ds_logic.v(5261)
  and u4022 (Hnciu6, Onciu6, Vnciu6);  // ../RTL/cortexm0ds_logic.v(5262)
  and u4023 (n831, HRDATA[11], Pp7iu6);  // ../RTL/cortexm0ds_logic.v(5263)
  not u4024 (Vnciu6, n831);  // ../RTL/cortexm0ds_logic.v(5263)
  and u4025 (Onciu6, Cociu6, Jociu6);  // ../RTL/cortexm0ds_logic.v(5264)
  and u4026 (n832, Hrfpw6[11], Uy4iu6);  // ../RTL/cortexm0ds_logic.v(5265)
  not u4027 (Jociu6, n832);  // ../RTL/cortexm0ds_logic.v(5265)
  and u4028 (n833, HRDATA[27], Kq7iu6);  // ../RTL/cortexm0ds_logic.v(5266)
  not u4029 (Cociu6, n833);  // ../RTL/cortexm0ds_logic.v(5266)
  buf u403 (vis_msp_o[17], Ta0qw6);  // ../RTL/cortexm0ds_logic.v(2097)
  and u4030 (Anciu6, Qociu6, Xociu6);  // ../RTL/cortexm0ds_logic.v(5267)
  and u4031 (n834, A25iu6, Ppfpw6[11]);  // ../RTL/cortexm0ds_logic.v(5268)
  not u4032 (Xociu6, n834);  // ../RTL/cortexm0ds_logic.v(5268)
  and u4033 (n835, R05iu6, D7fpw6[11]);  // ../RTL/cortexm0ds_logic.v(5269)
  not u4034 (Qociu6, n835);  // ../RTL/cortexm0ds_logic.v(5269)
  and u4035 (n836, Epciu6, Lpciu6);  // ../RTL/cortexm0ds_logic.v(5270)
  not u4036 (Qzuhu6, n836);  // ../RTL/cortexm0ds_logic.v(5270)
  and u4037 (Lpciu6, Spciu6, Zpciu6);  // ../RTL/cortexm0ds_logic.v(5271)
  and u4038 (n837, HRDATA[10], Pp7iu6);  // ../RTL/cortexm0ds_logic.v(5272)
  not u4039 (Zpciu6, n837);  // ../RTL/cortexm0ds_logic.v(5272)
  buf u404 (vis_msp_o[18], T80qw6);  // ../RTL/cortexm0ds_logic.v(2097)
  and u4040 (Spciu6, Gqciu6, Nqciu6);  // ../RTL/cortexm0ds_logic.v(5273)
  and u4041 (n838, Hrfpw6[10], Uy4iu6);  // ../RTL/cortexm0ds_logic.v(5274)
  not u4042 (Nqciu6, n838);  // ../RTL/cortexm0ds_logic.v(5274)
  and u4043 (n839, HRDATA[26], Kq7iu6);  // ../RTL/cortexm0ds_logic.v(5275)
  not u4044 (Gqciu6, n839);  // ../RTL/cortexm0ds_logic.v(5275)
  and u4045 (Epciu6, Uqciu6, Brciu6);  // ../RTL/cortexm0ds_logic.v(5276)
  and u4046 (n840, A25iu6, Ppfpw6[10]);  // ../RTL/cortexm0ds_logic.v(5277)
  not u4047 (Brciu6, n840);  // ../RTL/cortexm0ds_logic.v(5277)
  and u4048 (n841, R05iu6, D7fpw6[10]);  // ../RTL/cortexm0ds_logic.v(5278)
  not u4049 (Uqciu6, n841);  // ../RTL/cortexm0ds_logic.v(5278)
  buf u405 (vis_msp_o[20], Tffbx6);  // ../RTL/cortexm0ds_logic.v(2097)
  and u4050 (n842, Irciu6, Prciu6);  // ../RTL/cortexm0ds_logic.v(5279)
  not u4051 (Jzuhu6, n842);  // ../RTL/cortexm0ds_logic.v(5279)
  and u4052 (Prciu6, Wrciu6, Dsciu6);  // ../RTL/cortexm0ds_logic.v(5280)
  and u4053 (n843, HRDATA[9], Pp7iu6);  // ../RTL/cortexm0ds_logic.v(5281)
  not u4054 (Dsciu6, n843);  // ../RTL/cortexm0ds_logic.v(5281)
  and u4055 (Wrciu6, Ksciu6, Rsciu6);  // ../RTL/cortexm0ds_logic.v(5282)
  and u4056 (n844, Hrfpw6[9], Uy4iu6);  // ../RTL/cortexm0ds_logic.v(5283)
  not u4057 (Rsciu6, n844);  // ../RTL/cortexm0ds_logic.v(5283)
  and u4058 (n845, HRDATA[25], Kq7iu6);  // ../RTL/cortexm0ds_logic.v(5284)
  not u4059 (Ksciu6, n845);  // ../RTL/cortexm0ds_logic.v(5284)
  buf u406 (vis_msp_o[21], Gp6ax6);  // ../RTL/cortexm0ds_logic.v(2097)
  and u4060 (Irciu6, Ysciu6, Ftciu6);  // ../RTL/cortexm0ds_logic.v(5285)
  and u4061 (n846, A25iu6, Ppfpw6[9]);  // ../RTL/cortexm0ds_logic.v(5286)
  not u4062 (Ftciu6, n846);  // ../RTL/cortexm0ds_logic.v(5286)
  and u4063 (n847, R05iu6, D7fpw6[9]);  // ../RTL/cortexm0ds_logic.v(5287)
  not u4064 (Ysciu6, n847);  // ../RTL/cortexm0ds_logic.v(5287)
  not u4065 (Czuhu6, Mtciu6);  // ../RTL/cortexm0ds_logic.v(5288)
  AL_MUX u4066 (
    .i0(Ttciu6),
    .i1(Auciu6),
    .sel(HREADY),
    .o(Mtciu6));  // ../RTL/cortexm0ds_logic.v(5289)
  and u4067 (n848, Huciu6, Ouciu6);  // ../RTL/cortexm0ds_logic.v(5290)
  not u4068 (Auciu6, n848);  // ../RTL/cortexm0ds_logic.v(5290)
  and u4069 (Ouciu6, Vuciu6, Cvciu6);  // ../RTL/cortexm0ds_logic.v(5291)
  buf u407 (vis_msp_o[22], Twzpw6);  // ../RTL/cortexm0ds_logic.v(2097)
  and u4070 (Huciu6, HALTED, A2nhu6);  // ../RTL/cortexm0ds_logic.v(5292)
  and u4071 (n849, Jvciu6, Qvciu6);  // ../RTL/cortexm0ds_logic.v(5293)
  not u4072 (Vyuhu6, n849);  // ../RTL/cortexm0ds_logic.v(5293)
  and u4073 (n850, Xvciu6, K7vpw6);  // ../RTL/cortexm0ds_logic.v(5294)
  not u4074 (Qvciu6, n850);  // ../RTL/cortexm0ds_logic.v(5294)
  and u4075 (n851, HALTED, HREADY);  // ../RTL/cortexm0ds_logic.v(5296)
  not u4076 (Xvciu6, n851);  // ../RTL/cortexm0ds_logic.v(5296)
  or u4077 (Jvciu6, Eh6iu6, DBGRESTART);  // ../RTL/cortexm0ds_logic.v(5297)
  and u4078 (n852, Jw4iu6, Ewciu6);  // ../RTL/cortexm0ds_logic.v(5298)
  not u4079 (Oyuhu6, n852);  // ../RTL/cortexm0ds_logic.v(5298)
  buf u408 (Smhhu6, Ljcax6);  // ../RTL/cortexm0ds_logic.v(2298)
  and u4080 (n853, Dhgpw6[4], Lwciu6);  // ../RTL/cortexm0ds_logic.v(5299)
  not u4081 (Ewciu6, n853);  // ../RTL/cortexm0ds_logic.v(5299)
  and u4082 (n854, Scbiu6, H34iu6);  // ../RTL/cortexm0ds_logic.v(5300)
  not u4083 (Lwciu6, n854);  // ../RTL/cortexm0ds_logic.v(5300)
  and u4084 (n855, Swciu6, EDBGRQ);  // ../RTL/cortexm0ds_logic.v(5301)
  not u4085 (Jw4iu6, n855);  // ../RTL/cortexm0ds_logic.v(5301)
  or u4086 (n856, Zwciu6, HALTED);  // ../RTL/cortexm0ds_logic.v(5302)
  not u4087 (Swciu6, n856);  // ../RTL/cortexm0ds_logic.v(5302)
  AL_MUX u4088 (
    .i0(Gxciu6),
    .i1(HWRITE),
    .sel(Wi7iu6),
    .o(Hyuhu6));  // ../RTL/cortexm0ds_logic.v(5303)
  and u4089 (n857, Bq6iu6, Nxciu6);  // ../RTL/cortexm0ds_logic.v(5304)
  buf u409 (Gqgpw6[15], Eudax6);  // ../RTL/cortexm0ds_logic.v(2377)
  not u4090 (Wi7iu6, n857);  // ../RTL/cortexm0ds_logic.v(5304)
  and u4091 (n858, Uxciu6, Byciu6);  // ../RTL/cortexm0ds_logic.v(5305)
  not u4092 (Nxciu6, n858);  // ../RTL/cortexm0ds_logic.v(5305)
  or u4093 (n859, Iyciu6, Pyciu6);  // ../RTL/cortexm0ds_logic.v(5306)
  not u4094 (Byciu6, n859);  // ../RTL/cortexm0ds_logic.v(5306)
  or u4095 (Iyciu6, Wyciu6, V0epw6);  // ../RTL/cortexm0ds_logic.v(5307)
  and u4096 (Uxciu6, S18iu6, Hy8iu6);  // ../RTL/cortexm0ds_logic.v(5309)
  or u4097 (Bq6iu6, Dzciu6, Kzciu6);  // ../RTL/cortexm0ds_logic.v(5310)
  and u4098 (n860, Xg6iu6, HREADY);  // ../RTL/cortexm0ds_logic.v(5311)
  not u4099 (Dzciu6, n860);  // ../RTL/cortexm0ds_logic.v(5311)
  buf u41 (Gtgpw6[8], Facax6);  // ../RTL/cortexm0ds_logic.v(2375)
  buf u410 (Gqgpw6[19], Nodax6);  // ../RTL/cortexm0ds_logic.v(2377)
  and u4100 (Gxciu6, Rzciu6, Yzciu6);  // ../RTL/cortexm0ds_logic.v(5312)
  and u4101 (n861, F0diu6, M0diu6);  // ../RTL/cortexm0ds_logic.v(5313)
  not u4102 (Ayuhu6, n861);  // ../RTL/cortexm0ds_logic.v(5313)
  and u4103 (n862, Vbgpw6[30], T0diu6);  // ../RTL/cortexm0ds_logic.v(5314)
  not u4104 (M0diu6, n862);  // ../RTL/cortexm0ds_logic.v(5314)
  and u4105 (n863, HWDATA[30], O59iu6);  // ../RTL/cortexm0ds_logic.v(5315)
  not u4106 (T0diu6, n863);  // ../RTL/cortexm0ds_logic.v(5315)
  and u4107 (n864, V59iu6, HWDATA[30]);  // ../RTL/cortexm0ds_logic.v(5316)
  not u4108 (F0diu6, n864);  // ../RTL/cortexm0ds_logic.v(5316)
  AL_MUX u4109 (
    .i0(HWDATA[30]),
    .i1(R4gpw6[6]),
    .sel(Dv9iu6),
    .o(Txuhu6));  // ../RTL/cortexm0ds_logic.v(5317)
  or u411 (Qbfpw6[26], U27ju6, M75ju6);  // ../RTL/cortexm0ds_logic.v(9482)
  and u4110 (n865, A1diu6, H1diu6);  // ../RTL/cortexm0ds_logic.v(5318)
  not u4111 (Mxuhu6, n865);  // ../RTL/cortexm0ds_logic.v(5318)
  and u4112 (n866, Vbgpw6[29], O1diu6);  // ../RTL/cortexm0ds_logic.v(5319)
  not u4113 (H1diu6, n866);  // ../RTL/cortexm0ds_logic.v(5319)
  and u4114 (n867, HWDATA[29], O59iu6);  // ../RTL/cortexm0ds_logic.v(5320)
  not u4115 (O1diu6, n867);  // ../RTL/cortexm0ds_logic.v(5320)
  and u4116 (n868, V59iu6, HWDATA[29]);  // ../RTL/cortexm0ds_logic.v(5321)
  not u4117 (A1diu6, n868);  // ../RTL/cortexm0ds_logic.v(5321)
  and u4118 (n869, V1diu6, C2diu6);  // ../RTL/cortexm0ds_logic.v(5322)
  not u4119 (Fxuhu6, n869);  // ../RTL/cortexm0ds_logic.v(5322)
  or u412 (Qbfpw6[27], V67ju6, M75ju6);  // ../RTL/cortexm0ds_logic.v(9482)
  and u4120 (n870, Vbgpw6[28], J2diu6);  // ../RTL/cortexm0ds_logic.v(5323)
  not u4121 (C2diu6, n870);  // ../RTL/cortexm0ds_logic.v(5323)
  and u4122 (n871, HWDATA[28], O59iu6);  // ../RTL/cortexm0ds_logic.v(5324)
  not u4123 (J2diu6, n871);  // ../RTL/cortexm0ds_logic.v(5324)
  and u4124 (n872, V59iu6, HWDATA[28]);  // ../RTL/cortexm0ds_logic.v(5325)
  not u4125 (V1diu6, n872);  // ../RTL/cortexm0ds_logic.v(5325)
  and u4126 (n873, Q2diu6, X2diu6);  // ../RTL/cortexm0ds_logic.v(5326)
  not u4127 (Ywuhu6, n873);  // ../RTL/cortexm0ds_logic.v(5326)
  and u4128 (n874, Vbgpw6[27], E3diu6);  // ../RTL/cortexm0ds_logic.v(5327)
  not u4129 (X2diu6, n874);  // ../RTL/cortexm0ds_logic.v(5327)
  buf u413 (X3fpw6[2], Htmpw6);  // ../RTL/cortexm0ds_logic.v(1784)
  and u4130 (n875, HWDATA[27], O59iu6);  // ../RTL/cortexm0ds_logic.v(5328)
  not u4131 (E3diu6, n875);  // ../RTL/cortexm0ds_logic.v(5328)
  and u4132 (n876, V59iu6, HWDATA[27]);  // ../RTL/cortexm0ds_logic.v(5329)
  not u4133 (Q2diu6, n876);  // ../RTL/cortexm0ds_logic.v(5329)
  and u4134 (n877, L3diu6, S3diu6);  // ../RTL/cortexm0ds_logic.v(5330)
  not u4135 (Rwuhu6, n877);  // ../RTL/cortexm0ds_logic.v(5330)
  and u4136 (n878, Vbgpw6[26], Z3diu6);  // ../RTL/cortexm0ds_logic.v(5331)
  not u4137 (S3diu6, n878);  // ../RTL/cortexm0ds_logic.v(5331)
  and u4138 (n879, HWDATA[26], O59iu6);  // ../RTL/cortexm0ds_logic.v(5332)
  not u4139 (Z3diu6, n879);  // ../RTL/cortexm0ds_logic.v(5332)
  buf u414 (X3fpw6[3], Vmipw6);  // ../RTL/cortexm0ds_logic.v(1784)
  and u4140 (n880, V59iu6, HWDATA[26]);  // ../RTL/cortexm0ds_logic.v(5333)
  not u4141 (L3diu6, n880);  // ../RTL/cortexm0ds_logic.v(5333)
  and u4142 (n881, G4diu6, N4diu6);  // ../RTL/cortexm0ds_logic.v(5334)
  not u4143 (Kwuhu6, n881);  // ../RTL/cortexm0ds_logic.v(5334)
  and u4144 (n882, Vbgpw6[25], U4diu6);  // ../RTL/cortexm0ds_logic.v(5335)
  not u4145 (N4diu6, n882);  // ../RTL/cortexm0ds_logic.v(5335)
  and u4146 (n883, HWDATA[25], O59iu6);  // ../RTL/cortexm0ds_logic.v(5336)
  not u4147 (U4diu6, n883);  // ../RTL/cortexm0ds_logic.v(5336)
  and u4148 (n884, V59iu6, HWDATA[25]);  // ../RTL/cortexm0ds_logic.v(5337)
  not u4149 (G4diu6, n884);  // ../RTL/cortexm0ds_logic.v(5337)
  buf u415 (Iwfpw6[1], Ms5bx6);  // ../RTL/cortexm0ds_logic.v(2830)
  and u4150 (n885, B5diu6, I5diu6);  // ../RTL/cortexm0ds_logic.v(5338)
  not u4151 (Dwuhu6, n885);  // ../RTL/cortexm0ds_logic.v(5338)
  and u4152 (n886, Vbgpw6[24], P5diu6);  // ../RTL/cortexm0ds_logic.v(5339)
  not u4153 (I5diu6, n886);  // ../RTL/cortexm0ds_logic.v(5339)
  and u4154 (n887, HWDATA[24], O59iu6);  // ../RTL/cortexm0ds_logic.v(5340)
  not u4155 (P5diu6, n887);  // ../RTL/cortexm0ds_logic.v(5340)
  and u4156 (n888, V59iu6, HWDATA[24]);  // ../RTL/cortexm0ds_logic.v(5341)
  not u4157 (B5diu6, n888);  // ../RTL/cortexm0ds_logic.v(5341)
  and u4158 (n889, W5diu6, D6diu6);  // ../RTL/cortexm0ds_logic.v(5342)
  not u4159 (Wvuhu6, n889);  // ../RTL/cortexm0ds_logic.v(5342)
  buf u416 (Sqhpw6[1], Uofax6);  // ../RTL/cortexm0ds_logic.v(2359)
  and u4160 (n890, Vbgpw6[23], K6diu6);  // ../RTL/cortexm0ds_logic.v(5343)
  not u4161 (D6diu6, n890);  // ../RTL/cortexm0ds_logic.v(5343)
  and u4162 (n891, HWDATA[23], O59iu6);  // ../RTL/cortexm0ds_logic.v(5344)
  not u4163 (K6diu6, n891);  // ../RTL/cortexm0ds_logic.v(5344)
  and u4164 (n892, V59iu6, HWDATA[23]);  // ../RTL/cortexm0ds_logic.v(5345)
  not u4165 (W5diu6, n892);  // ../RTL/cortexm0ds_logic.v(5345)
  and u4166 (Pvuhu6, R6diu6, Y6diu6);  // ../RTL/cortexm0ds_logic.v(5346)
  and u4167 (Y6diu6, F7diu6, M7diu6);  // ../RTL/cortexm0ds_logic.v(5347)
  and u4168 (n893, Drdpw6, T7diu6);  // ../RTL/cortexm0ds_logic.v(5348)
  not u4169 (F7diu6, n893);  // ../RTL/cortexm0ds_logic.v(5348)
  buf u417 (Gqgpw6[4], F7eax6);  // ../RTL/cortexm0ds_logic.v(2377)
  and u4170 (R6diu6, IRQ[23], A8diu6);  // ../RTL/cortexm0ds_logic.v(5349)
  and u4171 (n894, Tk7iu6, H8diu6);  // ../RTL/cortexm0ds_logic.v(5350)
  not u4172 (A8diu6, n894);  // ../RTL/cortexm0ds_logic.v(5350)
  or u4173 (H8diu6, O8diu6, Qg6iu6);  // ../RTL/cortexm0ds_logic.v(5351)
  AL_MUX u4174 (
    .i0(HWDATA[23]),
    .i1(R4gpw6[5]),
    .sel(Dv9iu6),
    .o(Ivuhu6));  // ../RTL/cortexm0ds_logic.v(5352)
  and u4175 (n895, V8diu6, C9diu6);  // ../RTL/cortexm0ds_logic.v(5353)
  not u4176 (Bvuhu6, n895);  // ../RTL/cortexm0ds_logic.v(5353)
  and u4177 (n896, Vbgpw6[22], J9diu6);  // ../RTL/cortexm0ds_logic.v(5354)
  not u4178 (C9diu6, n896);  // ../RTL/cortexm0ds_logic.v(5354)
  and u4179 (n897, HWDATA[22], O59iu6);  // ../RTL/cortexm0ds_logic.v(5355)
  buf u418 (Gqgpw6[5], J5eax6);  // ../RTL/cortexm0ds_logic.v(2377)
  not u4180 (J9diu6, n897);  // ../RTL/cortexm0ds_logic.v(5355)
  and u4181 (n898, V59iu6, HWDATA[22]);  // ../RTL/cortexm0ds_logic.v(5356)
  not u4182 (V8diu6, n898);  // ../RTL/cortexm0ds_logic.v(5356)
  and u4183 (Uuuhu6, Q9diu6, X9diu6);  // ../RTL/cortexm0ds_logic.v(5357)
  and u4184 (X9diu6, Eadiu6, Ladiu6);  // ../RTL/cortexm0ds_logic.v(5358)
  and u4185 (n899, Xndpw6, Sadiu6);  // ../RTL/cortexm0ds_logic.v(5359)
  not u4186 (Eadiu6, n899);  // ../RTL/cortexm0ds_logic.v(5359)
  and u4187 (Q9diu6, IRQ[22], Zadiu6);  // ../RTL/cortexm0ds_logic.v(5360)
  and u4188 (n900, Tk7iu6, Gbdiu6);  // ../RTL/cortexm0ds_logic.v(5361)
  not u4189 (Zadiu6, n900);  // ../RTL/cortexm0ds_logic.v(5361)
  buf u419 (Gqgpw6[7], N3eax6);  // ../RTL/cortexm0ds_logic.v(2377)
  or u4190 (Gbdiu6, Qg6iu6, Nbdiu6);  // ../RTL/cortexm0ds_logic.v(5362)
  AL_MUX u4191 (
    .i0(HWDATA[22]),
    .i1(R4gpw6[4]),
    .sel(Dv9iu6),
    .o(Nuuhu6));  // ../RTL/cortexm0ds_logic.v(5363)
  and u4192 (n901, Ubdiu6, Bcdiu6);  // ../RTL/cortexm0ds_logic.v(5364)
  not u4193 (Guuhu6, n901);  // ../RTL/cortexm0ds_logic.v(5364)
  and u4194 (n902, Vbgpw6[21], Icdiu6);  // ../RTL/cortexm0ds_logic.v(5365)
  not u4195 (Bcdiu6, n902);  // ../RTL/cortexm0ds_logic.v(5365)
  and u4196 (n903, HWDATA[21], O59iu6);  // ../RTL/cortexm0ds_logic.v(5366)
  not u4197 (Icdiu6, n903);  // ../RTL/cortexm0ds_logic.v(5366)
  and u4198 (n904, V59iu6, HWDATA[21]);  // ../RTL/cortexm0ds_logic.v(5367)
  not u4199 (Ubdiu6, n904);  // ../RTL/cortexm0ds_logic.v(5367)
  buf u42 (vis_r1_o[15], Zt7bx6);  // ../RTL/cortexm0ds_logic.v(1876)
  buf u420 (Gqgpw6[9], Xajbx6);  // ../RTL/cortexm0ds_logic.v(2377)
  and u4200 (Ztuhu6, Pcdiu6, Wcdiu6);  // ../RTL/cortexm0ds_logic.v(5368)
  and u4201 (Wcdiu6, Dddiu6, Kddiu6);  // ../RTL/cortexm0ds_logic.v(5369)
  and u4202 (n905, Rrdpw6, Rddiu6);  // ../RTL/cortexm0ds_logic.v(5370)
  not u4203 (Dddiu6, n905);  // ../RTL/cortexm0ds_logic.v(5370)
  and u4204 (Pcdiu6, IRQ[21], Yddiu6);  // ../RTL/cortexm0ds_logic.v(5371)
  and u4205 (n906, Tk7iu6, Fediu6);  // ../RTL/cortexm0ds_logic.v(5372)
  not u4206 (Yddiu6, n906);  // ../RTL/cortexm0ds_logic.v(5372)
  or u4207 (Fediu6, Mediu6, Qg6iu6);  // ../RTL/cortexm0ds_logic.v(5373)
  and u4208 (n907, Tediu6, Afdiu6);  // ../RTL/cortexm0ds_logic.v(5374)
  not u4209 (Stuhu6, n907);  // ../RTL/cortexm0ds_logic.v(5374)
  buf u421 (Gqgpw6[10], Vzdax6);  // ../RTL/cortexm0ds_logic.v(2377)
  and u4210 (n908, Vbgpw6[20], Hfdiu6);  // ../RTL/cortexm0ds_logic.v(5375)
  not u4211 (Afdiu6, n908);  // ../RTL/cortexm0ds_logic.v(5375)
  and u4212 (n909, HWDATA[20], O59iu6);  // ../RTL/cortexm0ds_logic.v(5376)
  not u4213 (Hfdiu6, n909);  // ../RTL/cortexm0ds_logic.v(5376)
  and u4214 (n910, V59iu6, HWDATA[20]);  // ../RTL/cortexm0ds_logic.v(5377)
  not u4215 (Tediu6, n910);  // ../RTL/cortexm0ds_logic.v(5377)
  and u4216 (Ltuhu6, Ofdiu6, Vfdiu6);  // ../RTL/cortexm0ds_logic.v(5378)
  and u4217 (Vfdiu6, Cgdiu6, Jgdiu6);  // ../RTL/cortexm0ds_logic.v(5379)
  and u4218 (n911, Yrdpw6, Qgdiu6);  // ../RTL/cortexm0ds_logic.v(5380)
  not u4219 (Cgdiu6, n911);  // ../RTL/cortexm0ds_logic.v(5380)
  buf u422 (Gqgpw6[12], Yxdax6);  // ../RTL/cortexm0ds_logic.v(2377)
  and u4220 (Ofdiu6, IRQ[20], Xgdiu6);  // ../RTL/cortexm0ds_logic.v(5381)
  and u4221 (n912, Tk7iu6, Ehdiu6);  // ../RTL/cortexm0ds_logic.v(5382)
  not u4222 (Xgdiu6, n912);  // ../RTL/cortexm0ds_logic.v(5382)
  or u4223 (Ehdiu6, Qg6iu6, Lhdiu6);  // ../RTL/cortexm0ds_logic.v(5383)
  and u4224 (n913, Shdiu6, Zhdiu6);  // ../RTL/cortexm0ds_logic.v(5384)
  not u4225 (Etuhu6, n913);  // ../RTL/cortexm0ds_logic.v(5384)
  and u4226 (n914, Vbgpw6[19], Gidiu6);  // ../RTL/cortexm0ds_logic.v(5385)
  not u4227 (Zhdiu6, n914);  // ../RTL/cortexm0ds_logic.v(5385)
  and u4228 (n915, HWDATA[19], O59iu6);  // ../RTL/cortexm0ds_logic.v(5386)
  not u4229 (Gidiu6, n915);  // ../RTL/cortexm0ds_logic.v(5386)
  buf u423 (Gqgpw6[13], Bwdax6);  // ../RTL/cortexm0ds_logic.v(2377)
  and u4230 (n916, V59iu6, HWDATA[19]);  // ../RTL/cortexm0ds_logic.v(5387)
  not u4231 (Shdiu6, n916);  // ../RTL/cortexm0ds_logic.v(5387)
  and u4232 (Xsuhu6, Nidiu6, Uidiu6);  // ../RTL/cortexm0ds_logic.v(5388)
  and u4233 (Uidiu6, Bjdiu6, Ijdiu6);  // ../RTL/cortexm0ds_logic.v(5389)
  and u4234 (n917, Msdpw6, Pjdiu6);  // ../RTL/cortexm0ds_logic.v(5390)
  not u4235 (Bjdiu6, n917);  // ../RTL/cortexm0ds_logic.v(5390)
  and u4236 (Nidiu6, IRQ[19], Wjdiu6);  // ../RTL/cortexm0ds_logic.v(5391)
  and u4237 (n918, Tk7iu6, Dkdiu6);  // ../RTL/cortexm0ds_logic.v(5392)
  not u4238 (Wjdiu6, n918);  // ../RTL/cortexm0ds_logic.v(5392)
  or u4239 (Dkdiu6, Qg6iu6, Kkdiu6);  // ../RTL/cortexm0ds_logic.v(5393)
  buf u424 (Gqgpw6[14], Esabx6);  // ../RTL/cortexm0ds_logic.v(2377)
  and u4240 (n919, Rkdiu6, Ykdiu6);  // ../RTL/cortexm0ds_logic.v(5394)
  not u4241 (Qsuhu6, n919);  // ../RTL/cortexm0ds_logic.v(5394)
  and u4242 (n920, Vbgpw6[18], Fldiu6);  // ../RTL/cortexm0ds_logic.v(5395)
  not u4243 (Ykdiu6, n920);  // ../RTL/cortexm0ds_logic.v(5395)
  and u4244 (n921, HWDATA[18], O59iu6);  // ../RTL/cortexm0ds_logic.v(5396)
  not u4245 (Fldiu6, n921);  // ../RTL/cortexm0ds_logic.v(5396)
  and u4246 (n922, V59iu6, HWDATA[18]);  // ../RTL/cortexm0ds_logic.v(5397)
  not u4247 (Rkdiu6, n922);  // ../RTL/cortexm0ds_logic.v(5397)
  and u4248 (Jsuhu6, Mldiu6, Tldiu6);  // ../RTL/cortexm0ds_logic.v(5398)
  and u4249 (Tldiu6, Amdiu6, Hmdiu6);  // ../RTL/cortexm0ds_logic.v(5399)
  buf u425 (Qhhhu6, Efdax6);  // ../RTL/cortexm0ds_logic.v(2315)
  and u4250 (n923, Tsdpw6, Omdiu6);  // ../RTL/cortexm0ds_logic.v(5400)
  not u4251 (Amdiu6, n923);  // ../RTL/cortexm0ds_logic.v(5400)
  and u4252 (Mldiu6, IRQ[18], Vmdiu6);  // ../RTL/cortexm0ds_logic.v(5401)
  and u4253 (n924, Tk7iu6, Cndiu6);  // ../RTL/cortexm0ds_logic.v(5402)
  not u4254 (Vmdiu6, n924);  // ../RTL/cortexm0ds_logic.v(5402)
  or u4255 (Cndiu6, Qg6iu6, Jndiu6);  // ../RTL/cortexm0ds_logic.v(5403)
  and u4256 (n925, Qndiu6, Xndiu6);  // ../RTL/cortexm0ds_logic.v(5404)
  not u4257 (Csuhu6, n925);  // ../RTL/cortexm0ds_logic.v(5404)
  and u4258 (n926, Vbgpw6[17], Eodiu6);  // ../RTL/cortexm0ds_logic.v(5405)
  not u4259 (Xndiu6, n926);  // ../RTL/cortexm0ds_logic.v(5405)
  buf u426 (Hrfpw6[15], Sejax6);  // ../RTL/cortexm0ds_logic.v(2428)
  and u4260 (n927, HWDATA[17], O59iu6);  // ../RTL/cortexm0ds_logic.v(5406)
  not u4261 (Eodiu6, n927);  // ../RTL/cortexm0ds_logic.v(5406)
  and u4262 (n928, V59iu6, HWDATA[17]);  // ../RTL/cortexm0ds_logic.v(5407)
  not u4263 (Qndiu6, n928);  // ../RTL/cortexm0ds_logic.v(5407)
  and u4264 (Vruhu6, Lodiu6, Sodiu6);  // ../RTL/cortexm0ds_logic.v(5408)
  and u4265 (Sodiu6, Zodiu6, Gpdiu6);  // ../RTL/cortexm0ds_logic.v(5409)
  and u4266 (n929, Htdpw6, Npdiu6);  // ../RTL/cortexm0ds_logic.v(5410)
  not u4267 (Zodiu6, n929);  // ../RTL/cortexm0ds_logic.v(5410)
  and u4268 (Lodiu6, IRQ[17], Updiu6);  // ../RTL/cortexm0ds_logic.v(5411)
  and u4269 (n930, Tk7iu6, Bqdiu6);  // ../RTL/cortexm0ds_logic.v(5412)
  buf u427 (Gqgpw6[18], Kqdax6);  // ../RTL/cortexm0ds_logic.v(2377)
  not u4270 (Updiu6, n930);  // ../RTL/cortexm0ds_logic.v(5412)
  or u4271 (Bqdiu6, Qg6iu6, Iqdiu6);  // ../RTL/cortexm0ds_logic.v(5413)
  and u4272 (n931, Pqdiu6, Wqdiu6);  // ../RTL/cortexm0ds_logic.v(5414)
  not u4273 (Oruhu6, n931);  // ../RTL/cortexm0ds_logic.v(5414)
  and u4274 (n932, Vbgpw6[16], Drdiu6);  // ../RTL/cortexm0ds_logic.v(5415)
  not u4275 (Wqdiu6, n932);  // ../RTL/cortexm0ds_logic.v(5415)
  and u4276 (n933, HWDATA[16], O59iu6);  // ../RTL/cortexm0ds_logic.v(5416)
  not u4277 (Drdiu6, n933);  // ../RTL/cortexm0ds_logic.v(5416)
  and u4278 (n934, V59iu6, HWDATA[16]);  // ../RTL/cortexm0ds_logic.v(5417)
  not u4279 (Pqdiu6, n934);  // ../RTL/cortexm0ds_logic.v(5417)
  buf u428 (vis_r11_o[23], P54qw6);  // ../RTL/cortexm0ds_logic.v(1874)
  and u4280 (n935, Krdiu6, Rrdiu6);  // ../RTL/cortexm0ds_logic.v(5418)
  not u4281 (Hruhu6, n935);  // ../RTL/cortexm0ds_logic.v(5418)
  and u4282 (n936, Vbgpw6[15], Yrdiu6);  // ../RTL/cortexm0ds_logic.v(5419)
  not u4283 (Rrdiu6, n936);  // ../RTL/cortexm0ds_logic.v(5419)
  and u4284 (n937, Fsdiu6, O59iu6);  // ../RTL/cortexm0ds_logic.v(5420)
  not u4285 (Yrdiu6, n937);  // ../RTL/cortexm0ds_logic.v(5420)
  and u4286 (n938, V59iu6, Fsdiu6);  // ../RTL/cortexm0ds_logic.v(5421)
  not u4287 (Krdiu6, n938);  // ../RTL/cortexm0ds_logic.v(5421)
  AL_MUX u4288 (
    .i0(Fsdiu6),
    .i1(R4gpw6[3]),
    .sel(Dv9iu6),
    .o(Aruhu6));  // ../RTL/cortexm0ds_logic.v(5422)
  and u4289 (n939, Msdiu6, Tsdiu6);  // ../RTL/cortexm0ds_logic.v(5423)
  buf u429 (vis_r11_o[24], Ytspw6);  // ../RTL/cortexm0ds_logic.v(1874)
  not u4290 (Tquhu6, n939);  // ../RTL/cortexm0ds_logic.v(5423)
  and u4291 (n940, Vbgpw6[14], Atdiu6);  // ../RTL/cortexm0ds_logic.v(5424)
  not u4292 (Tsdiu6, n940);  // ../RTL/cortexm0ds_logic.v(5424)
  and u4293 (n941, HWDATA[14], O59iu6);  // ../RTL/cortexm0ds_logic.v(5425)
  not u4294 (Atdiu6, n941);  // ../RTL/cortexm0ds_logic.v(5425)
  and u4295 (n942, V59iu6, HWDATA[14]);  // ../RTL/cortexm0ds_logic.v(5426)
  not u4296 (Msdiu6, n942);  // ../RTL/cortexm0ds_logic.v(5426)
  AL_MUX u4297 (
    .i0(HWDATA[14]),
    .i1(R4gpw6[2]),
    .sel(Dv9iu6),
    .o(Mquhu6));  // ../RTL/cortexm0ds_logic.v(5427)
  and u4298 (n943, Htdiu6, Otdiu6);  // ../RTL/cortexm0ds_logic.v(5428)
  not u4299 (Fquhu6, n943);  // ../RTL/cortexm0ds_logic.v(5428)
  buf u43 (Vchhu6, Isjpw6);  // ../RTL/cortexm0ds_logic.v(1805)
  buf u430 (vis_r11_o[29], Kkjpw6);  // ../RTL/cortexm0ds_logic.v(1874)
  and u4300 (n944, Vbgpw6[13], Vtdiu6);  // ../RTL/cortexm0ds_logic.v(5429)
  not u4301 (Otdiu6, n944);  // ../RTL/cortexm0ds_logic.v(5429)
  and u4302 (n945, HWDATA[13], O59iu6);  // ../RTL/cortexm0ds_logic.v(5430)
  not u4303 (Vtdiu6, n945);  // ../RTL/cortexm0ds_logic.v(5430)
  and u4304 (n946, V59iu6, HWDATA[13]);  // ../RTL/cortexm0ds_logic.v(5431)
  not u4305 (Htdiu6, n946);  // ../RTL/cortexm0ds_logic.v(5431)
  and u4306 (n947, Cudiu6, Judiu6);  // ../RTL/cortexm0ds_logic.v(5432)
  not u4307 (Ypuhu6, n947);  // ../RTL/cortexm0ds_logic.v(5432)
  and u4308 (n948, Vbgpw6[12], Qudiu6);  // ../RTL/cortexm0ds_logic.v(5433)
  not u4309 (Judiu6, n948);  // ../RTL/cortexm0ds_logic.v(5433)
  buf u431 (vis_r11_o[30], Uoipw6);  // ../RTL/cortexm0ds_logic.v(1874)
  and u4310 (n949, HWDATA[12], O59iu6);  // ../RTL/cortexm0ds_logic.v(5434)
  not u4311 (Qudiu6, n949);  // ../RTL/cortexm0ds_logic.v(5434)
  and u4312 (n950, V59iu6, HWDATA[12]);  // ../RTL/cortexm0ds_logic.v(5435)
  not u4313 (Cudiu6, n950);  // ../RTL/cortexm0ds_logic.v(5435)
  and u4314 (n951, Xudiu6, Evdiu6);  // ../RTL/cortexm0ds_logic.v(5436)
  not u4315 (Rpuhu6, n951);  // ../RTL/cortexm0ds_logic.v(5436)
  and u4316 (n952, Vbgpw6[11], Lvdiu6);  // ../RTL/cortexm0ds_logic.v(5437)
  not u4317 (Evdiu6, n952);  // ../RTL/cortexm0ds_logic.v(5437)
  and u4318 (n953, HWDATA[11], O59iu6);  // ../RTL/cortexm0ds_logic.v(5438)
  not u4319 (Lvdiu6, n953);  // ../RTL/cortexm0ds_logic.v(5438)
  buf u432 (Hrfpw6[1], Tujbx6);  // ../RTL/cortexm0ds_logic.v(2428)
  and u4320 (n954, V59iu6, HWDATA[11]);  // ../RTL/cortexm0ds_logic.v(5439)
  not u4321 (Xudiu6, n954);  // ../RTL/cortexm0ds_logic.v(5439)
  and u4322 (n955, Svdiu6, Zvdiu6);  // ../RTL/cortexm0ds_logic.v(5440)
  not u4323 (Kpuhu6, n955);  // ../RTL/cortexm0ds_logic.v(5440)
  and u4324 (n956, Vbgpw6[10], Gwdiu6);  // ../RTL/cortexm0ds_logic.v(5441)
  not u4325 (Zvdiu6, n956);  // ../RTL/cortexm0ds_logic.v(5441)
  and u4326 (n957, HWDATA[10], O59iu6);  // ../RTL/cortexm0ds_logic.v(5442)
  not u4327 (Gwdiu6, n957);  // ../RTL/cortexm0ds_logic.v(5442)
  and u4328 (n958, V59iu6, HWDATA[10]);  // ../RTL/cortexm0ds_logic.v(5443)
  not u4329 (Svdiu6, n958);  // ../RTL/cortexm0ds_logic.v(5443)
  buf u433 (Hrfpw6[2], Usjbx6);  // ../RTL/cortexm0ds_logic.v(2428)
  and u4330 (n959, Nwdiu6, Uwdiu6);  // ../RTL/cortexm0ds_logic.v(5444)
  not u4331 (Dpuhu6, n959);  // ../RTL/cortexm0ds_logic.v(5444)
  and u4332 (n960, Vbgpw6[9], Bxdiu6);  // ../RTL/cortexm0ds_logic.v(5445)
  not u4333 (Uwdiu6, n960);  // ../RTL/cortexm0ds_logic.v(5445)
  and u4334 (n961, HWDATA[9], O59iu6);  // ../RTL/cortexm0ds_logic.v(5446)
  not u4335 (Bxdiu6, n961);  // ../RTL/cortexm0ds_logic.v(5446)
  and u4336 (n962, V59iu6, HWDATA[9]);  // ../RTL/cortexm0ds_logic.v(5447)
  not u4337 (Nwdiu6, n962);  // ../RTL/cortexm0ds_logic.v(5447)
  and u4338 (n963, Ixdiu6, Pxdiu6);  // ../RTL/cortexm0ds_logic.v(5448)
  not u4339 (Wouhu6, n963);  // ../RTL/cortexm0ds_logic.v(5448)
  buf u434 (Hrfpw6[4], Tokax6);  // ../RTL/cortexm0ds_logic.v(2428)
  and u4340 (n964, Vbgpw6[8], Wxdiu6);  // ../RTL/cortexm0ds_logic.v(5449)
  not u4341 (Pxdiu6, n964);  // ../RTL/cortexm0ds_logic.v(5449)
  and u4342 (n965, HWDATA[8], O59iu6);  // ../RTL/cortexm0ds_logic.v(5450)
  not u4343 (Wxdiu6, n965);  // ../RTL/cortexm0ds_logic.v(5450)
  and u4344 (n966, V59iu6, HWDATA[8]);  // ../RTL/cortexm0ds_logic.v(5451)
  not u4345 (Ixdiu6, n966);  // ../RTL/cortexm0ds_logic.v(5451)
  and u4346 (n967, Dydiu6, Kydiu6);  // ../RTL/cortexm0ds_logic.v(5452)
  not u4347 (Pouhu6, n967);  // ../RTL/cortexm0ds_logic.v(5452)
  and u4348 (n968, Vbgpw6[7], Rydiu6);  // ../RTL/cortexm0ds_logic.v(5453)
  not u4349 (Kydiu6, n968);  // ../RTL/cortexm0ds_logic.v(5453)
  buf u435 (Hrfpw6[5], Kakax6);  // ../RTL/cortexm0ds_logic.v(2428)
  and u4350 (n969, HWDATA[7], O59iu6);  // ../RTL/cortexm0ds_logic.v(5454)
  not u4351 (Rydiu6, n969);  // ../RTL/cortexm0ds_logic.v(5454)
  and u4352 (n970, V59iu6, HWDATA[7]);  // ../RTL/cortexm0ds_logic.v(5455)
  not u4353 (Dydiu6, n970);  // ../RTL/cortexm0ds_logic.v(5455)
  AL_MUX u4354 (
    .i0(HWDATA[7]),
    .i1(R4gpw6[1]),
    .sel(Dv9iu6),
    .o(Iouhu6));  // ../RTL/cortexm0ds_logic.v(5456)
  and u4355 (n971, Yydiu6, Fzdiu6);  // ../RTL/cortexm0ds_logic.v(5457)
  not u4356 (Bouhu6, n971);  // ../RTL/cortexm0ds_logic.v(5457)
  and u4357 (n972, Vbgpw6[6], Mzdiu6);  // ../RTL/cortexm0ds_logic.v(5458)
  not u4358 (Fzdiu6, n972);  // ../RTL/cortexm0ds_logic.v(5458)
  and u4359 (n973, HWDATA[6], O59iu6);  // ../RTL/cortexm0ds_logic.v(5459)
  buf u436 (Hrfpw6[7], O2kax6);  // ../RTL/cortexm0ds_logic.v(2428)
  not u4360 (Mzdiu6, n973);  // ../RTL/cortexm0ds_logic.v(5459)
  and u4361 (n974, V59iu6, HWDATA[6]);  // ../RTL/cortexm0ds_logic.v(5460)
  not u4362 (Yydiu6, n974);  // ../RTL/cortexm0ds_logic.v(5460)
  AL_MUX u4363 (
    .i0(HWDATA[6]),
    .i1(R4gpw6[0]),
    .sel(Dv9iu6),
    .o(Unuhu6));  // ../RTL/cortexm0ds_logic.v(5461)
  and u4364 (n975, Tzdiu6, Npdhu6);  // ../RTL/cortexm0ds_logic.v(5462)
  not u4365 (Dv9iu6, n975);  // ../RTL/cortexm0ds_logic.v(5462)
  and u4366 (n976, A0eiu6, H0eiu6);  // ../RTL/cortexm0ds_logic.v(5463)
  not u4367 (Nnuhu6, n976);  // ../RTL/cortexm0ds_logic.v(5463)
  and u4368 (n977, Vbgpw6[5], O0eiu6);  // ../RTL/cortexm0ds_logic.v(5464)
  not u4369 (H0eiu6, n977);  // ../RTL/cortexm0ds_logic.v(5464)
  buf u437 (Hrfpw6[9], Sujax6);  // ../RTL/cortexm0ds_logic.v(2428)
  and u4370 (n978, HWDATA[5], O59iu6);  // ../RTL/cortexm0ds_logic.v(5465)
  not u4371 (O0eiu6, n978);  // ../RTL/cortexm0ds_logic.v(5465)
  and u4372 (n979, V59iu6, HWDATA[5]);  // ../RTL/cortexm0ds_logic.v(5466)
  not u4373 (A0eiu6, n979);  // ../RTL/cortexm0ds_logic.v(5466)
  and u4374 (n980, V0eiu6, C1eiu6);  // ../RTL/cortexm0ds_logic.v(5467)
  not u4375 (Gnuhu6, n980);  // ../RTL/cortexm0ds_logic.v(5467)
  and u4376 (n981, Vbgpw6[4], J1eiu6);  // ../RTL/cortexm0ds_logic.v(5468)
  not u4377 (C1eiu6, n981);  // ../RTL/cortexm0ds_logic.v(5468)
  and u4378 (n982, HWDATA[4], O59iu6);  // ../RTL/cortexm0ds_logic.v(5469)
  not u4379 (J1eiu6, n982);  // ../RTL/cortexm0ds_logic.v(5469)
  buf u438 (Hrfpw6[10], Sqjax6);  // ../RTL/cortexm0ds_logic.v(2428)
  and u4380 (n983, V59iu6, HWDATA[4]);  // ../RTL/cortexm0ds_logic.v(5470)
  not u4381 (V0eiu6, n983);  // ../RTL/cortexm0ds_logic.v(5470)
  and u4382 (n984, Q1eiu6, X1eiu6);  // ../RTL/cortexm0ds_logic.v(5471)
  not u4383 (Zmuhu6, n984);  // ../RTL/cortexm0ds_logic.v(5471)
  and u4384 (n985, Vbgpw6[3], E2eiu6);  // ../RTL/cortexm0ds_logic.v(5472)
  not u4385 (X1eiu6, n985);  // ../RTL/cortexm0ds_logic.v(5472)
  and u4386 (n986, HWDATA[3], O59iu6);  // ../RTL/cortexm0ds_logic.v(5473)
  not u4387 (E2eiu6, n986);  // ../RTL/cortexm0ds_logic.v(5473)
  and u4388 (n987, V59iu6, HWDATA[3]);  // ../RTL/cortexm0ds_logic.v(5474)
  not u4389 (Q1eiu6, n987);  // ../RTL/cortexm0ds_logic.v(5474)
  buf u439 (Hrfpw6[12], Sijax6);  // ../RTL/cortexm0ds_logic.v(2428)
  and u4390 (n988, L2eiu6, S2eiu6);  // ../RTL/cortexm0ds_logic.v(5475)
  not u4391 (Smuhu6, n988);  // ../RTL/cortexm0ds_logic.v(5475)
  and u4392 (n989, Vbgpw6[2], Z2eiu6);  // ../RTL/cortexm0ds_logic.v(5476)
  not u4393 (S2eiu6, n989);  // ../RTL/cortexm0ds_logic.v(5476)
  and u4394 (n990, G3eiu6, O59iu6);  // ../RTL/cortexm0ds_logic.v(5477)
  not u4395 (Z2eiu6, n990);  // ../RTL/cortexm0ds_logic.v(5477)
  and u4396 (n991, V59iu6, G3eiu6);  // ../RTL/cortexm0ds_logic.v(5478)
  not u4397 (L2eiu6, n991);  // ../RTL/cortexm0ds_logic.v(5478)
  and u4398 (n992, N3eiu6, U3eiu6);  // ../RTL/cortexm0ds_logic.v(5479)
  not u4399 (Lmuhu6, n992);  // ../RTL/cortexm0ds_logic.v(5479)
  buf u44 (E1hpw6[9], J5jbx6);  // ../RTL/cortexm0ds_logic.v(2367)
  buf u440 (Hrfpw6[13], Sgjax6);  // ../RTL/cortexm0ds_logic.v(2428)
  and u4400 (n993, Vbgpw6[1], B4eiu6);  // ../RTL/cortexm0ds_logic.v(5480)
  not u4401 (U3eiu6, n993);  // ../RTL/cortexm0ds_logic.v(5480)
  and u4402 (n994, I4eiu6, O59iu6);  // ../RTL/cortexm0ds_logic.v(5481)
  not u4403 (B4eiu6, n994);  // ../RTL/cortexm0ds_logic.v(5481)
  or u4404 (O59iu6, V59iu6, P4eiu6);  // ../RTL/cortexm0ds_logic.v(5482)
  and u4405 (P4eiu6, W4eiu6, D5eiu6);  // ../RTL/cortexm0ds_logic.v(5483)
  and u4406 (W4eiu6, Npdhu6, K5eiu6);  // ../RTL/cortexm0ds_logic.v(5484)
  and u4407 (n995, V59iu6, I4eiu6);  // ../RTL/cortexm0ds_logic.v(5485)
  not u4408 (N3eiu6, n995);  // ../RTL/cortexm0ds_logic.v(5485)
  and u4409 (V59iu6, Yzciu6, K5eiu6);  // ../RTL/cortexm0ds_logic.v(5486)
  buf u441 (Hrfpw6[14], Swjbx6);  // ../RTL/cortexm0ds_logic.v(2428)
  AL_MUX u4410 (
    .i0(HWDATA[0]),
    .i1(Bxghu6),
    .sel(R5eiu6),
    .o(Emuhu6));  // ../RTL/cortexm0ds_logic.v(5487)
  AL_MUX u4411 (
    .i0(G3eiu6),
    .i1(Ftghu6),
    .sel(R5eiu6),
    .o(Xluhu6));  // ../RTL/cortexm0ds_logic.v(5488)
  AL_MUX u4412 (
    .i0(I4eiu6),
    .i1(Dvghu6),
    .sel(R5eiu6),
    .o(Qluhu6));  // ../RTL/cortexm0ds_logic.v(5489)
  and u4413 (n996, Y5eiu6, Npdhu6);  // ../RTL/cortexm0ds_logic.v(5490)
  not u4414 (R5eiu6, n996);  // ../RTL/cortexm0ds_logic.v(5490)
  AL_MUX u4415 (
    .i0(HWDATA[0]),
    .i1(Bagpw6[0]),
    .sel(F6eiu6),
    .o(Jluhu6));  // ../RTL/cortexm0ds_logic.v(5491)
  AL_MUX u4416 (
    .i0(HWDATA[23]),
    .i1(Bagpw6[23]),
    .sel(F6eiu6),
    .o(Cluhu6));  // ../RTL/cortexm0ds_logic.v(5492)
  AL_MUX u4417 (
    .i0(HWDATA[22]),
    .i1(Bagpw6[22]),
    .sel(F6eiu6),
    .o(Vkuhu6));  // ../RTL/cortexm0ds_logic.v(5493)
  AL_MUX u4418 (
    .i0(HWDATA[21]),
    .i1(Bagpw6[21]),
    .sel(F6eiu6),
    .o(Okuhu6));  // ../RTL/cortexm0ds_logic.v(5494)
  AL_MUX u4419 (
    .i0(HWDATA[20]),
    .i1(Bagpw6[20]),
    .sel(F6eiu6),
    .o(Hkuhu6));  // ../RTL/cortexm0ds_logic.v(5495)
  buf u442 (Ijhhu6, Xaeax6);  // ../RTL/cortexm0ds_logic.v(2332)
  AL_MUX u4420 (
    .i0(HWDATA[19]),
    .i1(Bagpw6[19]),
    .sel(F6eiu6),
    .o(Akuhu6));  // ../RTL/cortexm0ds_logic.v(5496)
  AL_MUX u4421 (
    .i0(HWDATA[18]),
    .i1(Bagpw6[18]),
    .sel(F6eiu6),
    .o(Tjuhu6));  // ../RTL/cortexm0ds_logic.v(5497)
  AL_MUX u4422 (
    .i0(HWDATA[17]),
    .i1(Bagpw6[17]),
    .sel(F6eiu6),
    .o(Mjuhu6));  // ../RTL/cortexm0ds_logic.v(5498)
  AL_MUX u4423 (
    .i0(HWDATA[16]),
    .i1(Bagpw6[16]),
    .sel(F6eiu6),
    .o(Fjuhu6));  // ../RTL/cortexm0ds_logic.v(5499)
  AL_MUX u4424 (
    .i0(Fsdiu6),
    .i1(Bagpw6[15]),
    .sel(F6eiu6),
    .o(Yiuhu6));  // ../RTL/cortexm0ds_logic.v(5500)
  AL_MUX u4425 (
    .i0(HWDATA[14]),
    .i1(Bagpw6[14]),
    .sel(F6eiu6),
    .o(Riuhu6));  // ../RTL/cortexm0ds_logic.v(5501)
  AL_MUX u4426 (
    .i0(HWDATA[13]),
    .i1(Bagpw6[13]),
    .sel(F6eiu6),
    .o(Kiuhu6));  // ../RTL/cortexm0ds_logic.v(5502)
  AL_MUX u4427 (
    .i0(HWDATA[12]),
    .i1(Bagpw6[12]),
    .sel(F6eiu6),
    .o(Diuhu6));  // ../RTL/cortexm0ds_logic.v(5503)
  AL_MUX u4428 (
    .i0(HWDATA[11]),
    .i1(Bagpw6[11]),
    .sel(F6eiu6),
    .o(Whuhu6));  // ../RTL/cortexm0ds_logic.v(5504)
  AL_MUX u4429 (
    .i0(HWDATA[10]),
    .i1(Bagpw6[10]),
    .sel(F6eiu6),
    .o(Phuhu6));  // ../RTL/cortexm0ds_logic.v(5505)
  buf u443 (vis_r11_o[20], X2jpw6);  // ../RTL/cortexm0ds_logic.v(1874)
  AL_MUX u4430 (
    .i0(HWDATA[9]),
    .i1(Bagpw6[9]),
    .sel(F6eiu6),
    .o(Ihuhu6));  // ../RTL/cortexm0ds_logic.v(5506)
  AL_MUX u4431 (
    .i0(HWDATA[8]),
    .i1(Bagpw6[8]),
    .sel(F6eiu6),
    .o(Bhuhu6));  // ../RTL/cortexm0ds_logic.v(5507)
  AL_MUX u4432 (
    .i0(HWDATA[7]),
    .i1(Bagpw6[7]),
    .sel(F6eiu6),
    .o(Uguhu6));  // ../RTL/cortexm0ds_logic.v(5508)
  AL_MUX u4433 (
    .i0(HWDATA[6]),
    .i1(Bagpw6[6]),
    .sel(F6eiu6),
    .o(Nguhu6));  // ../RTL/cortexm0ds_logic.v(5509)
  AL_MUX u4434 (
    .i0(HWDATA[5]),
    .i1(Bagpw6[5]),
    .sel(F6eiu6),
    .o(Gguhu6));  // ../RTL/cortexm0ds_logic.v(5510)
  AL_MUX u4435 (
    .i0(HWDATA[4]),
    .i1(Bagpw6[4]),
    .sel(F6eiu6),
    .o(Zfuhu6));  // ../RTL/cortexm0ds_logic.v(5511)
  AL_MUX u4436 (
    .i0(HWDATA[3]),
    .i1(Bagpw6[3]),
    .sel(F6eiu6),
    .o(Sfuhu6));  // ../RTL/cortexm0ds_logic.v(5512)
  AL_MUX u4437 (
    .i0(G3eiu6),
    .i1(Bagpw6[2]),
    .sel(F6eiu6),
    .o(Lfuhu6));  // ../RTL/cortexm0ds_logic.v(5513)
  AL_MUX u4438 (
    .i0(I4eiu6),
    .i1(Bagpw6[1]),
    .sel(F6eiu6),
    .o(Efuhu6));  // ../RTL/cortexm0ds_logic.v(5514)
  and u4439 (n997, M6eiu6, Npdhu6);  // ../RTL/cortexm0ds_logic.v(5515)
  buf u444 (Gqgpw6[17], Erbbx6);  // ../RTL/cortexm0ds_logic.v(2377)
  not u4440 (F6eiu6, n997);  // ../RTL/cortexm0ds_logic.v(5515)
  and u4441 (n998, T6eiu6, A7eiu6);  // ../RTL/cortexm0ds_logic.v(5516)
  not u4442 (Xeuhu6, n998);  // ../RTL/cortexm0ds_logic.v(5516)
  or u4443 (A7eiu6, H7eiu6, O7eiu6);  // ../RTL/cortexm0ds_logic.v(5517)
  and u4444 (T6eiu6, V7eiu6, C8eiu6);  // ../RTL/cortexm0ds_logic.v(5518)
  and u4445 (n999, L6gpw6[0], J8eiu6);  // ../RTL/cortexm0ds_logic.v(5519)
  not u4446 (C8eiu6, n999);  // ../RTL/cortexm0ds_logic.v(5519)
  and u4447 (n1000, Q8eiu6, Bagpw6[0]);  // ../RTL/cortexm0ds_logic.v(5520)
  not u4448 (V7eiu6, n1000);  // ../RTL/cortexm0ds_logic.v(5520)
  and u4449 (n1001, X8eiu6, E9eiu6);  // ../RTL/cortexm0ds_logic.v(5521)
  buf u445 (vis_msp_o[26], Pejbx6);  // ../RTL/cortexm0ds_logic.v(2097)
  not u4450 (Qeuhu6, n1001);  // ../RTL/cortexm0ds_logic.v(5521)
  and u4451 (n1002, L9eiu6, Tzfpw6[1]);  // ../RTL/cortexm0ds_logic.v(5522)
  not u4452 (E9eiu6, n1002);  // ../RTL/cortexm0ds_logic.v(5522)
  and u4453 (X8eiu6, S9eiu6, Z9eiu6);  // ../RTL/cortexm0ds_logic.v(5523)
  and u4454 (n1003, L6gpw6[1], J8eiu6);  // ../RTL/cortexm0ds_logic.v(5524)
  not u4455 (Z9eiu6, n1003);  // ../RTL/cortexm0ds_logic.v(5524)
  and u4456 (n1004, Q8eiu6, Bagpw6[1]);  // ../RTL/cortexm0ds_logic.v(5525)
  not u4457 (S9eiu6, n1004);  // ../RTL/cortexm0ds_logic.v(5525)
  and u4458 (n1005, Gaeiu6, Naeiu6);  // ../RTL/cortexm0ds_logic.v(5526)
  not u4459 (Jeuhu6, n1005);  // ../RTL/cortexm0ds_logic.v(5526)
  buf u446 (vis_msp_o[27], T20qw6);  // ../RTL/cortexm0ds_logic.v(2097)
  and u4460 (n1006, L9eiu6, Tzfpw6[2]);  // ../RTL/cortexm0ds_logic.v(5527)
  not u4461 (Naeiu6, n1006);  // ../RTL/cortexm0ds_logic.v(5527)
  and u4462 (Gaeiu6, Uaeiu6, Bbeiu6);  // ../RTL/cortexm0ds_logic.v(5528)
  and u4463 (n1007, L6gpw6[2], J8eiu6);  // ../RTL/cortexm0ds_logic.v(5529)
  not u4464 (Bbeiu6, n1007);  // ../RTL/cortexm0ds_logic.v(5529)
  and u4465 (n1008, Q8eiu6, Bagpw6[2]);  // ../RTL/cortexm0ds_logic.v(5530)
  not u4466 (Uaeiu6, n1008);  // ../RTL/cortexm0ds_logic.v(5530)
  and u4467 (n1009, Ibeiu6, Pbeiu6);  // ../RTL/cortexm0ds_logic.v(5531)
  not u4468 (Ceuhu6, n1009);  // ../RTL/cortexm0ds_logic.v(5531)
  and u4469 (n1010, Tzfpw6[3], L9eiu6);  // ../RTL/cortexm0ds_logic.v(5532)
  buf u447 (vis_r11_o[3], Qbmpw6);  // ../RTL/cortexm0ds_logic.v(1874)
  not u4470 (Pbeiu6, n1010);  // ../RTL/cortexm0ds_logic.v(5532)
  and u4471 (Ibeiu6, Wbeiu6, Dceiu6);  // ../RTL/cortexm0ds_logic.v(5533)
  and u4472 (n1011, L6gpw6[3], J8eiu6);  // ../RTL/cortexm0ds_logic.v(5534)
  not u4473 (Dceiu6, n1011);  // ../RTL/cortexm0ds_logic.v(5534)
  and u4474 (n1012, Q8eiu6, Bagpw6[3]);  // ../RTL/cortexm0ds_logic.v(5535)
  not u4475 (Wbeiu6, n1012);  // ../RTL/cortexm0ds_logic.v(5535)
  and u4476 (n1013, Kceiu6, Rceiu6);  // ../RTL/cortexm0ds_logic.v(5536)
  not u4477 (Vduhu6, n1013);  // ../RTL/cortexm0ds_logic.v(5536)
  and u4478 (n1014, L9eiu6, Tzfpw6[4]);  // ../RTL/cortexm0ds_logic.v(5537)
  not u4479 (Rceiu6, n1014);  // ../RTL/cortexm0ds_logic.v(5537)
  buf u448 (vis_r11_o[4], Vuipw6);  // ../RTL/cortexm0ds_logic.v(1874)
  and u4480 (Kceiu6, Yceiu6, Fdeiu6);  // ../RTL/cortexm0ds_logic.v(5538)
  and u4481 (n1015, L6gpw6[4], J8eiu6);  // ../RTL/cortexm0ds_logic.v(5539)
  not u4482 (Fdeiu6, n1015);  // ../RTL/cortexm0ds_logic.v(5539)
  and u4483 (n1016, Q8eiu6, Bagpw6[4]);  // ../RTL/cortexm0ds_logic.v(5540)
  not u4484 (Yceiu6, n1016);  // ../RTL/cortexm0ds_logic.v(5540)
  and u4485 (n1017, Mdeiu6, Tdeiu6);  // ../RTL/cortexm0ds_logic.v(5541)
  not u4486 (Oduhu6, n1017);  // ../RTL/cortexm0ds_logic.v(5541)
  and u4487 (n1018, L9eiu6, Tzfpw6[5]);  // ../RTL/cortexm0ds_logic.v(5542)
  not u4488 (Tdeiu6, n1018);  // ../RTL/cortexm0ds_logic.v(5542)
  and u4489 (Mdeiu6, Aeeiu6, Heeiu6);  // ../RTL/cortexm0ds_logic.v(5543)
  buf u449 (vis_r11_o[6], Y5spw6);  // ../RTL/cortexm0ds_logic.v(1874)
  and u4490 (n1019, L6gpw6[5], J8eiu6);  // ../RTL/cortexm0ds_logic.v(5544)
  not u4491 (Heeiu6, n1019);  // ../RTL/cortexm0ds_logic.v(5544)
  and u4492 (n1020, Q8eiu6, Bagpw6[5]);  // ../RTL/cortexm0ds_logic.v(5545)
  not u4493 (Aeeiu6, n1020);  // ../RTL/cortexm0ds_logic.v(5545)
  and u4494 (n1021, Oeeiu6, Veeiu6);  // ../RTL/cortexm0ds_logic.v(5546)
  not u4495 (Hduhu6, n1021);  // ../RTL/cortexm0ds_logic.v(5546)
  and u4496 (n1022, L9eiu6, Tzfpw6[6]);  // ../RTL/cortexm0ds_logic.v(5547)
  not u4497 (Veeiu6, n1022);  // ../RTL/cortexm0ds_logic.v(5547)
  and u4498 (Oeeiu6, Cfeiu6, Jfeiu6);  // ../RTL/cortexm0ds_logic.v(5548)
  and u4499 (n1023, L6gpw6[6], J8eiu6);  // ../RTL/cortexm0ds_logic.v(5549)
  buf u45 (D7fpw6[0], Wfspw6);  // ../RTL/cortexm0ds_logic.v(2074)
  buf u450 (vis_r11_o[7], Bsrpw6);  // ../RTL/cortexm0ds_logic.v(1874)
  not u4500 (Jfeiu6, n1023);  // ../RTL/cortexm0ds_logic.v(5549)
  and u4501 (n1024, Q8eiu6, Bagpw6[6]);  // ../RTL/cortexm0ds_logic.v(5550)
  not u4502 (Cfeiu6, n1024);  // ../RTL/cortexm0ds_logic.v(5550)
  and u4503 (n1025, Qfeiu6, Xfeiu6);  // ../RTL/cortexm0ds_logic.v(5551)
  not u4504 (Aduhu6, n1025);  // ../RTL/cortexm0ds_logic.v(5551)
  and u4505 (n1026, L9eiu6, Tzfpw6[7]);  // ../RTL/cortexm0ds_logic.v(5552)
  not u4506 (Xfeiu6, n1026);  // ../RTL/cortexm0ds_logic.v(5552)
  and u4507 (Qfeiu6, Egeiu6, Lgeiu6);  // ../RTL/cortexm0ds_logic.v(5553)
  and u4508 (n1027, L6gpw6[7], J8eiu6);  // ../RTL/cortexm0ds_logic.v(5554)
  not u4509 (Lgeiu6, n1027);  // ../RTL/cortexm0ds_logic.v(5554)
  buf u451 (vis_r11_o[9], Gv1qw6);  // ../RTL/cortexm0ds_logic.v(1874)
  and u4510 (n1028, Q8eiu6, Bagpw6[7]);  // ../RTL/cortexm0ds_logic.v(5555)
  not u4511 (Egeiu6, n1028);  // ../RTL/cortexm0ds_logic.v(5555)
  and u4512 (n1029, Sgeiu6, Zgeiu6);  // ../RTL/cortexm0ds_logic.v(5556)
  not u4513 (Tcuhu6, n1029);  // ../RTL/cortexm0ds_logic.v(5556)
  and u4514 (n1030, L9eiu6, Tzfpw6[8]);  // ../RTL/cortexm0ds_logic.v(5557)
  not u4515 (Zgeiu6, n1030);  // ../RTL/cortexm0ds_logic.v(5557)
  and u4516 (Sgeiu6, Gheiu6, Nheiu6);  // ../RTL/cortexm0ds_logic.v(5558)
  and u4517 (n1031, L6gpw6[8], J8eiu6);  // ../RTL/cortexm0ds_logic.v(5559)
  not u4518 (Nheiu6, n1031);  // ../RTL/cortexm0ds_logic.v(5559)
  and u4519 (n1032, Q8eiu6, Bagpw6[8]);  // ../RTL/cortexm0ds_logic.v(5560)
  buf u452 (vis_r11_o[10], Hqxpw6);  // ../RTL/cortexm0ds_logic.v(1874)
  not u4520 (Gheiu6, n1032);  // ../RTL/cortexm0ds_logic.v(5560)
  and u4521 (n1033, Uheiu6, Bieiu6);  // ../RTL/cortexm0ds_logic.v(5561)
  not u4522 (Mcuhu6, n1033);  // ../RTL/cortexm0ds_logic.v(5561)
  and u4523 (n1034, L9eiu6, Tzfpw6[9]);  // ../RTL/cortexm0ds_logic.v(5562)
  not u4524 (Bieiu6, n1034);  // ../RTL/cortexm0ds_logic.v(5562)
  and u4525 (Uheiu6, Iieiu6, Pieiu6);  // ../RTL/cortexm0ds_logic.v(5563)
  and u4526 (n1035, L6gpw6[9], J8eiu6);  // ../RTL/cortexm0ds_logic.v(5564)
  not u4527 (Pieiu6, n1035);  // ../RTL/cortexm0ds_logic.v(5564)
  and u4528 (n1036, Q8eiu6, Bagpw6[9]);  // ../RTL/cortexm0ds_logic.v(5565)
  not u4529 (Iieiu6, n1036);  // ../RTL/cortexm0ds_logic.v(5565)
  buf u453 (vis_r11_o[12], Bbjpw6);  // ../RTL/cortexm0ds_logic.v(1874)
  and u4530 (n1037, Wieiu6, Djeiu6);  // ../RTL/cortexm0ds_logic.v(5566)
  not u4531 (Fcuhu6, n1037);  // ../RTL/cortexm0ds_logic.v(5566)
  and u4532 (n1038, L9eiu6, Tzfpw6[10]);  // ../RTL/cortexm0ds_logic.v(5567)
  not u4533 (Djeiu6, n1038);  // ../RTL/cortexm0ds_logic.v(5567)
  and u4534 (Wieiu6, Kjeiu6, Rjeiu6);  // ../RTL/cortexm0ds_logic.v(5568)
  and u4535 (n1039, L6gpw6[10], J8eiu6);  // ../RTL/cortexm0ds_logic.v(5569)
  not u4536 (Rjeiu6, n1039);  // ../RTL/cortexm0ds_logic.v(5569)
  and u4537 (n1040, Q8eiu6, Bagpw6[10]);  // ../RTL/cortexm0ds_logic.v(5570)
  not u4538 (Kjeiu6, n1040);  // ../RTL/cortexm0ds_logic.v(5570)
  and u4539 (n1041, Yjeiu6, Fkeiu6);  // ../RTL/cortexm0ds_logic.v(5571)
  buf u454 (vis_r11_o[14], S38ax6);  // ../RTL/cortexm0ds_logic.v(1874)
  not u4540 (Ybuhu6, n1041);  // ../RTL/cortexm0ds_logic.v(5571)
  and u4541 (n1042, Tzfpw6[11], L9eiu6);  // ../RTL/cortexm0ds_logic.v(5572)
  not u4542 (Fkeiu6, n1042);  // ../RTL/cortexm0ds_logic.v(5572)
  and u4543 (Yjeiu6, Mkeiu6, Tkeiu6);  // ../RTL/cortexm0ds_logic.v(5573)
  and u4544 (n1043, L6gpw6[11], J8eiu6);  // ../RTL/cortexm0ds_logic.v(5574)
  not u4545 (Tkeiu6, n1043);  // ../RTL/cortexm0ds_logic.v(5574)
  and u4546 (n1044, Q8eiu6, Bagpw6[11]);  // ../RTL/cortexm0ds_logic.v(5575)
  not u4547 (Mkeiu6, n1044);  // ../RTL/cortexm0ds_logic.v(5575)
  and u4548 (n1045, Aleiu6, Hleiu6);  // ../RTL/cortexm0ds_logic.v(5576)
  not u4549 (Rbuhu6, n1045);  // ../RTL/cortexm0ds_logic.v(5576)
  buf u455 (vis_r11_o[15], Z58bx6);  // ../RTL/cortexm0ds_logic.v(1874)
  and u4550 (n1046, L9eiu6, Tzfpw6[12]);  // ../RTL/cortexm0ds_logic.v(5577)
  not u4551 (Hleiu6, n1046);  // ../RTL/cortexm0ds_logic.v(5577)
  and u4552 (Aleiu6, Oleiu6, Vleiu6);  // ../RTL/cortexm0ds_logic.v(5578)
  and u4553 (n1047, L6gpw6[12], J8eiu6);  // ../RTL/cortexm0ds_logic.v(5579)
  not u4554 (Vleiu6, n1047);  // ../RTL/cortexm0ds_logic.v(5579)
  and u4555 (n1048, Q8eiu6, Bagpw6[12]);  // ../RTL/cortexm0ds_logic.v(5580)
  not u4556 (Oleiu6, n1048);  // ../RTL/cortexm0ds_logic.v(5580)
  and u4557 (n1049, Cmeiu6, Jmeiu6);  // ../RTL/cortexm0ds_logic.v(5581)
  not u4558 (Kbuhu6, n1049);  // ../RTL/cortexm0ds_logic.v(5581)
  and u4559 (n1050, L9eiu6, Tzfpw6[13]);  // ../RTL/cortexm0ds_logic.v(5582)
  buf u456 (vis_r11_o[17], Ydupw6);  // ../RTL/cortexm0ds_logic.v(1874)
  not u4560 (Jmeiu6, n1050);  // ../RTL/cortexm0ds_logic.v(5582)
  and u4561 (Cmeiu6, Qmeiu6, Xmeiu6);  // ../RTL/cortexm0ds_logic.v(5583)
  and u4562 (n1051, L6gpw6[13], J8eiu6);  // ../RTL/cortexm0ds_logic.v(5584)
  not u4563 (Xmeiu6, n1051);  // ../RTL/cortexm0ds_logic.v(5584)
  and u4564 (n1052, Q8eiu6, Bagpw6[13]);  // ../RTL/cortexm0ds_logic.v(5585)
  not u4565 (Qmeiu6, n1052);  // ../RTL/cortexm0ds_logic.v(5585)
  and u4566 (n1053, Eneiu6, Lneiu6);  // ../RTL/cortexm0ds_logic.v(5586)
  not u4567 (Dbuhu6, n1053);  // ../RTL/cortexm0ds_logic.v(5586)
  and u4568 (n1054, L9eiu6, Tzfpw6[14]);  // ../RTL/cortexm0ds_logic.v(5587)
  not u4569 (Lneiu6, n1054);  // ../RTL/cortexm0ds_logic.v(5587)
  buf u457 (vis_r11_o[18], P8xpw6);  // ../RTL/cortexm0ds_logic.v(1874)
  and u4570 (Eneiu6, Sneiu6, Zneiu6);  // ../RTL/cortexm0ds_logic.v(5588)
  and u4571 (n1055, L6gpw6[14], J8eiu6);  // ../RTL/cortexm0ds_logic.v(5589)
  not u4572 (Zneiu6, n1055);  // ../RTL/cortexm0ds_logic.v(5589)
  and u4573 (n1056, Q8eiu6, Bagpw6[14]);  // ../RTL/cortexm0ds_logic.v(5590)
  not u4574 (Sneiu6, n1056);  // ../RTL/cortexm0ds_logic.v(5590)
  and u4575 (n1057, Goeiu6, Noeiu6);  // ../RTL/cortexm0ds_logic.v(5591)
  not u4576 (Wauhu6, n1057);  // ../RTL/cortexm0ds_logic.v(5591)
  and u4577 (n1058, L9eiu6, Tzfpw6[15]);  // ../RTL/cortexm0ds_logic.v(5592)
  not u4578 (Noeiu6, n1058);  // ../RTL/cortexm0ds_logic.v(5592)
  and u4579 (Goeiu6, Uoeiu6, Bpeiu6);  // ../RTL/cortexm0ds_logic.v(5593)
  buf u458 (vis_r11_o[19], Jpvpw6);  // ../RTL/cortexm0ds_logic.v(1874)
  and u4580 (n1059, L6gpw6[15], J8eiu6);  // ../RTL/cortexm0ds_logic.v(5594)
  not u4581 (Bpeiu6, n1059);  // ../RTL/cortexm0ds_logic.v(5594)
  and u4582 (n1060, Q8eiu6, Bagpw6[15]);  // ../RTL/cortexm0ds_logic.v(5595)
  not u4583 (Uoeiu6, n1060);  // ../RTL/cortexm0ds_logic.v(5595)
  and u4584 (n1061, Ipeiu6, Ppeiu6);  // ../RTL/cortexm0ds_logic.v(5596)
  not u4585 (Pauhu6, n1061);  // ../RTL/cortexm0ds_logic.v(5596)
  and u4586 (n1062, L9eiu6, Tzfpw6[16]);  // ../RTL/cortexm0ds_logic.v(5597)
  not u4587 (Ppeiu6, n1062);  // ../RTL/cortexm0ds_logic.v(5597)
  and u4588 (Ipeiu6, Wpeiu6, Dqeiu6);  // ../RTL/cortexm0ds_logic.v(5598)
  and u4589 (n1063, L6gpw6[16], J8eiu6);  // ../RTL/cortexm0ds_logic.v(5599)
  buf u459 (Alhhu6, Q6fax6);  // ../RTL/cortexm0ds_logic.v(2349)
  not u4590 (Dqeiu6, n1063);  // ../RTL/cortexm0ds_logic.v(5599)
  and u4591 (n1064, Q8eiu6, Bagpw6[16]);  // ../RTL/cortexm0ds_logic.v(5600)
  not u4592 (Wpeiu6, n1064);  // ../RTL/cortexm0ds_logic.v(5600)
  and u4593 (n1065, Kqeiu6, Rqeiu6);  // ../RTL/cortexm0ds_logic.v(5601)
  not u4594 (Iauhu6, n1065);  // ../RTL/cortexm0ds_logic.v(5601)
  and u4595 (n1066, L9eiu6, Tzfpw6[17]);  // ../RTL/cortexm0ds_logic.v(5602)
  not u4596 (Rqeiu6, n1066);  // ../RTL/cortexm0ds_logic.v(5602)
  and u4597 (Kqeiu6, Yqeiu6, Freiu6);  // ../RTL/cortexm0ds_logic.v(5603)
  and u4598 (n1067, L6gpw6[17], J8eiu6);  // ../RTL/cortexm0ds_logic.v(5604)
  not u4599 (Freiu6, n1067);  // ../RTL/cortexm0ds_logic.v(5604)
  buf u46 (vis_r1_o[4], Lrppw6);  // ../RTL/cortexm0ds_logic.v(1876)
  buf u460 (T0hhu6, M8fax6);  // ../RTL/cortexm0ds_logic.v(2350)
  and u4600 (n1068, Q8eiu6, Bagpw6[17]);  // ../RTL/cortexm0ds_logic.v(5605)
  not u4601 (Yqeiu6, n1068);  // ../RTL/cortexm0ds_logic.v(5605)
  and u4602 (n1069, Mreiu6, Treiu6);  // ../RTL/cortexm0ds_logic.v(5606)
  not u4603 (Bauhu6, n1069);  // ../RTL/cortexm0ds_logic.v(5606)
  and u4604 (n1070, L9eiu6, Tzfpw6[18]);  // ../RTL/cortexm0ds_logic.v(5607)
  not u4605 (Treiu6, n1070);  // ../RTL/cortexm0ds_logic.v(5607)
  and u4606 (Mreiu6, Aseiu6, Hseiu6);  // ../RTL/cortexm0ds_logic.v(5608)
  and u4607 (n1071, L6gpw6[18], J8eiu6);  // ../RTL/cortexm0ds_logic.v(5609)
  not u4608 (Hseiu6, n1071);  // ../RTL/cortexm0ds_logic.v(5609)
  and u4609 (n1072, Q8eiu6, Bagpw6[18]);  // ../RTL/cortexm0ds_logic.v(5610)
  buf u461 (H2hhu6, Eafax6);  // ../RTL/cortexm0ds_logic.v(2351)
  not u4610 (Aseiu6, n1072);  // ../RTL/cortexm0ds_logic.v(5610)
  and u4611 (n1073, Oseiu6, Vseiu6);  // ../RTL/cortexm0ds_logic.v(5611)
  not u4612 (U9uhu6, n1073);  // ../RTL/cortexm0ds_logic.v(5611)
  and u4613 (n1074, Tzfpw6[19], L9eiu6);  // ../RTL/cortexm0ds_logic.v(5612)
  not u4614 (Vseiu6, n1074);  // ../RTL/cortexm0ds_logic.v(5612)
  and u4615 (Oseiu6, Cteiu6, Jteiu6);  // ../RTL/cortexm0ds_logic.v(5613)
  and u4616 (n1075, L6gpw6[19], J8eiu6);  // ../RTL/cortexm0ds_logic.v(5614)
  not u4617 (Jteiu6, n1075);  // ../RTL/cortexm0ds_logic.v(5614)
  and u4618 (n1076, Q8eiu6, Bagpw6[19]);  // ../RTL/cortexm0ds_logic.v(5615)
  not u4619 (Cteiu6, n1076);  // ../RTL/cortexm0ds_logic.v(5615)
  buf u462 (E5hhu6, Sbfax6);  // ../RTL/cortexm0ds_logic.v(2352)
  and u4620 (n1077, Qteiu6, Xteiu6);  // ../RTL/cortexm0ds_logic.v(5616)
  not u4621 (N9uhu6, n1077);  // ../RTL/cortexm0ds_logic.v(5616)
  and u4622 (n1078, L9eiu6, Tzfpw6[20]);  // ../RTL/cortexm0ds_logic.v(5617)
  not u4623 (Xteiu6, n1078);  // ../RTL/cortexm0ds_logic.v(5617)
  and u4624 (Qteiu6, Eueiu6, Lueiu6);  // ../RTL/cortexm0ds_logic.v(5618)
  and u4625 (n1079, L6gpw6[20], J8eiu6);  // ../RTL/cortexm0ds_logic.v(5619)
  not u4626 (Lueiu6, n1079);  // ../RTL/cortexm0ds_logic.v(5619)
  and u4627 (n1080, Q8eiu6, Bagpw6[20]);  // ../RTL/cortexm0ds_logic.v(5620)
  not u4628 (Eueiu6, n1080);  // ../RTL/cortexm0ds_logic.v(5620)
  and u4629 (n1081, Sueiu6, Zueiu6);  // ../RTL/cortexm0ds_logic.v(5621)
  buf u463 (S3hhu6, Hdfax6);  // ../RTL/cortexm0ds_logic.v(2353)
  not u4630 (G9uhu6, n1081);  // ../RTL/cortexm0ds_logic.v(5621)
  and u4631 (n1082, L9eiu6, Tzfpw6[21]);  // ../RTL/cortexm0ds_logic.v(5622)
  not u4632 (Zueiu6, n1082);  // ../RTL/cortexm0ds_logic.v(5622)
  and u4633 (Sueiu6, Gveiu6, Nveiu6);  // ../RTL/cortexm0ds_logic.v(5623)
  and u4634 (n1083, L6gpw6[21], J8eiu6);  // ../RTL/cortexm0ds_logic.v(5624)
  not u4635 (Nveiu6, n1083);  // ../RTL/cortexm0ds_logic.v(5624)
  and u4636 (n1084, Q8eiu6, Bagpw6[21]);  // ../RTL/cortexm0ds_logic.v(5625)
  not u4637 (Gveiu6, n1084);  // ../RTL/cortexm0ds_logic.v(5625)
  and u4638 (n1085, Uveiu6, Bweiu6);  // ../RTL/cortexm0ds_logic.v(5626)
  not u4639 (Z8uhu6, n1085);  // ../RTL/cortexm0ds_logic.v(5626)
  buf u464 (vis_r4_o[17], V3vax6);  // ../RTL/cortexm0ds_logic.v(2626)
  and u4640 (n1086, L9eiu6, Tzfpw6[22]);  // ../RTL/cortexm0ds_logic.v(5627)
  not u4641 (Bweiu6, n1086);  // ../RTL/cortexm0ds_logic.v(5627)
  and u4642 (Uveiu6, Iweiu6, Pweiu6);  // ../RTL/cortexm0ds_logic.v(5628)
  and u4643 (n1087, L6gpw6[22], J8eiu6);  // ../RTL/cortexm0ds_logic.v(5629)
  not u4644 (Pweiu6, n1087);  // ../RTL/cortexm0ds_logic.v(5629)
  and u4645 (n1088, Q8eiu6, Bagpw6[22]);  // ../RTL/cortexm0ds_logic.v(5630)
  not u4646 (Iweiu6, n1088);  // ../RTL/cortexm0ds_logic.v(5630)
  and u4647 (n1089, Wweiu6, Dxeiu6);  // ../RTL/cortexm0ds_logic.v(5631)
  not u4648 (S8uhu6, n1089);  // ../RTL/cortexm0ds_logic.v(5631)
  and u4649 (n1090, L9eiu6, Tzfpw6[23]);  // ../RTL/cortexm0ds_logic.v(5632)
  buf u465 (vis_r14_o[14], N1oax6);  // ../RTL/cortexm0ds_logic.v(2497)
  not u4650 (Dxeiu6, n1090);  // ../RTL/cortexm0ds_logic.v(5632)
  and u4651 (Wweiu6, Kxeiu6, Rxeiu6);  // ../RTL/cortexm0ds_logic.v(5633)
  and u4652 (n1091, L6gpw6[23], J8eiu6);  // ../RTL/cortexm0ds_logic.v(5634)
  not u4653 (Rxeiu6, n1091);  // ../RTL/cortexm0ds_logic.v(5634)
  and u4654 (J8eiu6, Yxeiu6, Fyeiu6);  // ../RTL/cortexm0ds_logic.v(5635)
  or u4655 (n1092, L9eiu6, Myeiu6);  // ../RTL/cortexm0ds_logic.v(5636)
  not u4656 (Yxeiu6, n1092);  // ../RTL/cortexm0ds_logic.v(5636)
  and u4657 (n1093, Q8eiu6, Bagpw6[23]);  // ../RTL/cortexm0ds_logic.v(5637)
  not u4658 (Kxeiu6, n1093);  // ../RTL/cortexm0ds_logic.v(5637)
  or u4659 (n1094, Tyeiu6, Fyeiu6);  // ../RTL/cortexm0ds_logic.v(5638)
  not u466 (Omdpw6, Pifax6);  // ../RTL/cortexm0ds_logic.v(2356)
  not u4660 (Q8eiu6, n1094);  // ../RTL/cortexm0ds_logic.v(5638)
  and u4661 (n1095, Azeiu6, O7eiu6);  // ../RTL/cortexm0ds_logic.v(5639)
  not u4662 (Fyeiu6, n1095);  // ../RTL/cortexm0ds_logic.v(5639)
  not u4663 (O7eiu6, Tzfpw6[0]);  // ../RTL/cortexm0ds_logic.v(5640)
  and u4664 (n1096, H7eiu6, Hzeiu6);  // ../RTL/cortexm0ds_logic.v(5641)
  not u4665 (Tyeiu6, n1096);  // ../RTL/cortexm0ds_logic.v(5641)
  or u4666 (H7eiu6, Ozeiu6, Myeiu6);  // ../RTL/cortexm0ds_logic.v(5643)
  not u4667 (L9eiu6, H7eiu6);  // ../RTL/cortexm0ds_logic.v(5643)
  AL_MUX u4668 (
    .i0(HWDATA[6]),
    .i1(R4gpw6[56]),
    .sel(Vzeiu6),
    .o(L8uhu6));  // ../RTL/cortexm0ds_logic.v(5645)
  AL_MUX u4669 (
    .i0(HWDATA[7]),
    .i1(R4gpw6[57]),
    .sel(Vzeiu6),
    .o(E8uhu6));  // ../RTL/cortexm0ds_logic.v(5646)
  buf u467 (N3nhu6, Okfax6);  // ../RTL/cortexm0ds_logic.v(2357)
  AL_MUX u4670 (
    .i0(HWDATA[14]),
    .i1(R4gpw6[58]),
    .sel(Vzeiu6),
    .o(X7uhu6));  // ../RTL/cortexm0ds_logic.v(5647)
  AL_MUX u4671 (
    .i0(Fsdiu6),
    .i1(R4gpw6[59]),
    .sel(Vzeiu6),
    .o(Q7uhu6));  // ../RTL/cortexm0ds_logic.v(5648)
  AL_MUX u4672 (
    .i0(HWDATA[22]),
    .i1(R4gpw6[60]),
    .sel(Vzeiu6),
    .o(J7uhu6));  // ../RTL/cortexm0ds_logic.v(5649)
  AL_MUX u4673 (
    .i0(HWDATA[23]),
    .i1(R4gpw6[61]),
    .sel(Vzeiu6),
    .o(C7uhu6));  // ../RTL/cortexm0ds_logic.v(5650)
  AL_MUX u4674 (
    .i0(HWDATA[30]),
    .i1(R4gpw6[62]),
    .sel(Vzeiu6),
    .o(V6uhu6));  // ../RTL/cortexm0ds_logic.v(5651)
  AL_MUX u4675 (
    .i0(HWDATA[31]),
    .i1(R4gpw6[63]),
    .sel(Vzeiu6),
    .o(O6uhu6));  // ../RTL/cortexm0ds_logic.v(5652)
  and u4676 (n1097, C0fiu6, Npdhu6);  // ../RTL/cortexm0ds_logic.v(5653)
  not u4677 (Vzeiu6, n1097);  // ../RTL/cortexm0ds_logic.v(5653)
  AL_MUX u4678 (
    .i0(HWDATA[6]),
    .i1(R4gpw6[48]),
    .sel(J0fiu6),
    .o(H6uhu6));  // ../RTL/cortexm0ds_logic.v(5654)
  AL_MUX u4679 (
    .i0(HWDATA[7]),
    .i1(R4gpw6[49]),
    .sel(J0fiu6),
    .o(A6uhu6));  // ../RTL/cortexm0ds_logic.v(5655)
  buf u468 (Vbgpw6[27], Qx0bx6);  // ../RTL/cortexm0ds_logic.v(3092)
  AL_MUX u4680 (
    .i0(HWDATA[14]),
    .i1(R4gpw6[50]),
    .sel(J0fiu6),
    .o(T5uhu6));  // ../RTL/cortexm0ds_logic.v(5656)
  AL_MUX u4681 (
    .i0(Fsdiu6),
    .i1(R4gpw6[51]),
    .sel(J0fiu6),
    .o(M5uhu6));  // ../RTL/cortexm0ds_logic.v(5657)
  AL_MUX u4682 (
    .i0(HWDATA[22]),
    .i1(R4gpw6[52]),
    .sel(J0fiu6),
    .o(F5uhu6));  // ../RTL/cortexm0ds_logic.v(5658)
  AL_MUX u4683 (
    .i0(HWDATA[23]),
    .i1(R4gpw6[53]),
    .sel(J0fiu6),
    .o(Y4uhu6));  // ../RTL/cortexm0ds_logic.v(5659)
  AL_MUX u4684 (
    .i0(HWDATA[30]),
    .i1(R4gpw6[54]),
    .sel(J0fiu6),
    .o(R4uhu6));  // ../RTL/cortexm0ds_logic.v(5660)
  AL_MUX u4685 (
    .i0(HWDATA[31]),
    .i1(R4gpw6[55]),
    .sel(J0fiu6),
    .o(K4uhu6));  // ../RTL/cortexm0ds_logic.v(5661)
  and u4686 (n1098, Q0fiu6, Npdhu6);  // ../RTL/cortexm0ds_logic.v(5662)
  not u4687 (J0fiu6, n1098);  // ../RTL/cortexm0ds_logic.v(5662)
  AL_MUX u4688 (
    .i0(HWDATA[6]),
    .i1(R4gpw6[40]),
    .sel(X0fiu6),
    .o(D4uhu6));  // ../RTL/cortexm0ds_logic.v(5663)
  AL_MUX u4689 (
    .i0(HWDATA[7]),
    .i1(R4gpw6[41]),
    .sel(X0fiu6),
    .o(W3uhu6));  // ../RTL/cortexm0ds_logic.v(5664)
  buf u469 (Ligpw6[27], Dncax6);  // ../RTL/cortexm0ds_logic.v(2371)
  AL_MUX u4690 (
    .i0(HWDATA[14]),
    .i1(R4gpw6[42]),
    .sel(X0fiu6),
    .o(P3uhu6));  // ../RTL/cortexm0ds_logic.v(5665)
  AL_MUX u4691 (
    .i0(Fsdiu6),
    .i1(R4gpw6[43]),
    .sel(X0fiu6),
    .o(I3uhu6));  // ../RTL/cortexm0ds_logic.v(5666)
  AL_MUX u4692 (
    .i0(HWDATA[22]),
    .i1(R4gpw6[44]),
    .sel(X0fiu6),
    .o(B3uhu6));  // ../RTL/cortexm0ds_logic.v(5667)
  AL_MUX u4693 (
    .i0(HWDATA[23]),
    .i1(R4gpw6[45]),
    .sel(X0fiu6),
    .o(U2uhu6));  // ../RTL/cortexm0ds_logic.v(5668)
  AL_MUX u4694 (
    .i0(HWDATA[30]),
    .i1(R4gpw6[46]),
    .sel(X0fiu6),
    .o(N2uhu6));  // ../RTL/cortexm0ds_logic.v(5669)
  AL_MUX u4695 (
    .i0(HWDATA[31]),
    .i1(R4gpw6[47]),
    .sel(X0fiu6),
    .o(G2uhu6));  // ../RTL/cortexm0ds_logic.v(5670)
  and u4696 (n1099, E1fiu6, Npdhu6);  // ../RTL/cortexm0ds_logic.v(5671)
  not u4697 (X0fiu6, n1099);  // ../RTL/cortexm0ds_logic.v(5671)
  AL_MUX u4698 (
    .i0(HWDATA[6]),
    .i1(R4gpw6[32]),
    .sel(L1fiu6),
    .o(Z1uhu6));  // ../RTL/cortexm0ds_logic.v(5672)
  AL_MUX u4699 (
    .i0(HWDATA[7]),
    .i1(R4gpw6[33]),
    .sel(L1fiu6),
    .o(S1uhu6));  // ../RTL/cortexm0ds_logic.v(5673)
  buf u47 (Ivfhu6, Vzjpw6);  // ../RTL/cortexm0ds_logic.v(1809)
  buf u470 (Vbgpw6[20], Mp0bx6);  // ../RTL/cortexm0ds_logic.v(3092)
  AL_MUX u4700 (
    .i0(HWDATA[14]),
    .i1(R4gpw6[34]),
    .sel(L1fiu6),
    .o(L1uhu6));  // ../RTL/cortexm0ds_logic.v(5674)
  AL_MUX u4701 (
    .i0(Fsdiu6),
    .i1(R4gpw6[35]),
    .sel(L1fiu6),
    .o(E1uhu6));  // ../RTL/cortexm0ds_logic.v(5675)
  AL_MUX u4702 (
    .i0(HWDATA[22]),
    .i1(R4gpw6[36]),
    .sel(L1fiu6),
    .o(X0uhu6));  // ../RTL/cortexm0ds_logic.v(5676)
  AL_MUX u4703 (
    .i0(HWDATA[23]),
    .i1(R4gpw6[37]),
    .sel(L1fiu6),
    .o(Q0uhu6));  // ../RTL/cortexm0ds_logic.v(5677)
  AL_MUX u4704 (
    .i0(HWDATA[30]),
    .i1(R4gpw6[38]),
    .sel(L1fiu6),
    .o(J0uhu6));  // ../RTL/cortexm0ds_logic.v(5678)
  AL_MUX u4705 (
    .i0(HWDATA[31]),
    .i1(R4gpw6[39]),
    .sel(L1fiu6),
    .o(C0uhu6));  // ../RTL/cortexm0ds_logic.v(5679)
  and u4706 (n1100, S1fiu6, Npdhu6);  // ../RTL/cortexm0ds_logic.v(5680)
  not u4707 (L1fiu6, n1100);  // ../RTL/cortexm0ds_logic.v(5680)
  AL_MUX u4708 (
    .i0(HWDATA[6]),
    .i1(R4gpw6[24]),
    .sel(Z1fiu6),
    .o(Vzthu6));  // ../RTL/cortexm0ds_logic.v(5681)
  AL_MUX u4709 (
    .i0(HWDATA[7]),
    .i1(R4gpw6[25]),
    .sel(Z1fiu6),
    .o(Ozthu6));  // ../RTL/cortexm0ds_logic.v(5682)
  buf u471 (Dtnhu6, Qsfax6);  // ../RTL/cortexm0ds_logic.v(2361)
  AL_MUX u4710 (
    .i0(HWDATA[14]),
    .i1(R4gpw6[26]),
    .sel(Z1fiu6),
    .o(Hzthu6));  // ../RTL/cortexm0ds_logic.v(5683)
  AL_MUX u4711 (
    .i0(Fsdiu6),
    .i1(R4gpw6[27]),
    .sel(Z1fiu6),
    .o(Azthu6));  // ../RTL/cortexm0ds_logic.v(5684)
  AL_MUX u4712 (
    .i0(HWDATA[22]),
    .i1(R4gpw6[28]),
    .sel(Z1fiu6),
    .o(Tythu6));  // ../RTL/cortexm0ds_logic.v(5685)
  AL_MUX u4713 (
    .i0(HWDATA[23]),
    .i1(R4gpw6[29]),
    .sel(Z1fiu6),
    .o(Mythu6));  // ../RTL/cortexm0ds_logic.v(5686)
  AL_MUX u4714 (
    .i0(HWDATA[30]),
    .i1(R4gpw6[30]),
    .sel(Z1fiu6),
    .o(Fythu6));  // ../RTL/cortexm0ds_logic.v(5687)
  AL_MUX u4715 (
    .i0(HWDATA[31]),
    .i1(R4gpw6[31]),
    .sel(Z1fiu6),
    .o(Yxthu6));  // ../RTL/cortexm0ds_logic.v(5688)
  and u4716 (n1101, G2fiu6, Npdhu6);  // ../RTL/cortexm0ds_logic.v(5689)
  not u4717 (Z1fiu6, n1101);  // ../RTL/cortexm0ds_logic.v(5689)
  AL_MUX u4718 (
    .i0(HWDATA[6]),
    .i1(R4gpw6[16]),
    .sel(N2fiu6),
    .o(Rxthu6));  // ../RTL/cortexm0ds_logic.v(5690)
  AL_MUX u4719 (
    .i0(HWDATA[7]),
    .i1(R4gpw6[17]),
    .sel(N2fiu6),
    .o(Kxthu6));  // ../RTL/cortexm0ds_logic.v(5691)
  buf u472 (S3ohu6, Qufax6);  // ../RTL/cortexm0ds_logic.v(2362)
  AL_MUX u4720 (
    .i0(HWDATA[14]),
    .i1(R4gpw6[18]),
    .sel(N2fiu6),
    .o(Dxthu6));  // ../RTL/cortexm0ds_logic.v(5692)
  AL_MUX u4721 (
    .i0(Fsdiu6),
    .i1(R4gpw6[19]),
    .sel(N2fiu6),
    .o(Wwthu6));  // ../RTL/cortexm0ds_logic.v(5693)
  AL_MUX u4722 (
    .i0(HWDATA[22]),
    .i1(R4gpw6[20]),
    .sel(N2fiu6),
    .o(Pwthu6));  // ../RTL/cortexm0ds_logic.v(5694)
  AL_MUX u4723 (
    .i0(HWDATA[23]),
    .i1(R4gpw6[21]),
    .sel(N2fiu6),
    .o(Iwthu6));  // ../RTL/cortexm0ds_logic.v(5695)
  AL_MUX u4724 (
    .i0(HWDATA[30]),
    .i1(R4gpw6[22]),
    .sel(N2fiu6),
    .o(Bwthu6));  // ../RTL/cortexm0ds_logic.v(5696)
  AL_MUX u4725 (
    .i0(HWDATA[31]),
    .i1(R4gpw6[23]),
    .sel(N2fiu6),
    .o(Uvthu6));  // ../RTL/cortexm0ds_logic.v(5697)
  and u4726 (n1102, U2fiu6, Npdhu6);  // ../RTL/cortexm0ds_logic.v(5698)
  not u4727 (N2fiu6, n1102);  // ../RTL/cortexm0ds_logic.v(5698)
  AL_MUX u4728 (
    .i0(HWDATA[6]),
    .i1(R4gpw6[8]),
    .sel(B3fiu6),
    .o(Nvthu6));  // ../RTL/cortexm0ds_logic.v(5699)
  AL_MUX u4729 (
    .i0(HWDATA[7]),
    .i1(R4gpw6[9]),
    .sel(B3fiu6),
    .o(Gvthu6));  // ../RTL/cortexm0ds_logic.v(5700)
  buf u473 (Rrnhu6, Qwfax6);  // ../RTL/cortexm0ds_logic.v(2363)
  AL_MUX u4730 (
    .i0(HWDATA[14]),
    .i1(R4gpw6[10]),
    .sel(B3fiu6),
    .o(Zuthu6));  // ../RTL/cortexm0ds_logic.v(5701)
  AL_MUX u4731 (
    .i0(Fsdiu6),
    .i1(R4gpw6[11]),
    .sel(B3fiu6),
    .o(Suthu6));  // ../RTL/cortexm0ds_logic.v(5702)
  AL_MUX u4732 (
    .i0(HWDATA[22]),
    .i1(R4gpw6[12]),
    .sel(B3fiu6),
    .o(Luthu6));  // ../RTL/cortexm0ds_logic.v(5703)
  AL_MUX u4733 (
    .i0(HWDATA[23]),
    .i1(R4gpw6[13]),
    .sel(B3fiu6),
    .o(Euthu6));  // ../RTL/cortexm0ds_logic.v(5704)
  AL_MUX u4734 (
    .i0(HWDATA[30]),
    .i1(R4gpw6[14]),
    .sel(B3fiu6),
    .o(Xtthu6));  // ../RTL/cortexm0ds_logic.v(5705)
  AL_MUX u4735 (
    .i0(HWDATA[31]),
    .i1(R4gpw6[15]),
    .sel(B3fiu6),
    .o(Qtthu6));  // ../RTL/cortexm0ds_logic.v(5706)
  and u4736 (n1103, I3fiu6, Npdhu6);  // ../RTL/cortexm0ds_logic.v(5707)
  not u4737 (B3fiu6, n1103);  // ../RTL/cortexm0ds_logic.v(5707)
  AL_MUX u4738 (
    .i0(HWDATA[4]),
    .i1(Gfghu6),
    .sel(P3fiu6),
    .o(Jtthu6));  // ../RTL/cortexm0ds_logic.v(5708)
  and u4739 (n1104, W3fiu6, D4fiu6);  // ../RTL/cortexm0ds_logic.v(5709)
  buf u474 (Rgnhu6, Ryfax6);  // ../RTL/cortexm0ds_logic.v(2364)
  not u4740 (Ctthu6, n1104);  // ../RTL/cortexm0ds_logic.v(5709)
  and u4741 (n1105, vis_ipsr_o[4], F8ciu6);  // ../RTL/cortexm0ds_logic.v(5710)
  not u4742 (D4fiu6, n1105);  // ../RTL/cortexm0ds_logic.v(5710)
  and u4743 (W3fiu6, K4fiu6, R4fiu6);  // ../RTL/cortexm0ds_logic.v(5711)
  and u4744 (n1106, Xibiu6, Ppfpw6[4]);  // ../RTL/cortexm0ds_logic.v(5712)
  not u4745 (R4fiu6, n1106);  // ../RTL/cortexm0ds_logic.v(5712)
  or u4746 (K4fiu6, Ejbiu6, Y4fiu6);  // ../RTL/cortexm0ds_logic.v(5713)
  and u4747 (Vsthu6, F5fiu6, M5fiu6);  // ../RTL/cortexm0ds_logic.v(5714)
  and u4748 (M5fiu6, T5fiu6, A6fiu6);  // ../RTL/cortexm0ds_logic.v(5715)
  and u4749 (n1107, Zodpw6, H6fiu6);  // ../RTL/cortexm0ds_logic.v(5716)
  buf u475 (Jshpw6[4], Pg3qw6);  // ../RTL/cortexm0ds_logic.v(2372)
  not u4750 (T5fiu6, n1107);  // ../RTL/cortexm0ds_logic.v(5716)
  and u4751 (F5fiu6, IRQ[7], O6fiu6);  // ../RTL/cortexm0ds_logic.v(5717)
  and u4752 (n1108, Tk7iu6, V6fiu6);  // ../RTL/cortexm0ds_logic.v(5718)
  not u4753 (O6fiu6, n1108);  // ../RTL/cortexm0ds_logic.v(5718)
  or u4754 (V6fiu6, Qg6iu6, C7fiu6);  // ../RTL/cortexm0ds_logic.v(5719)
  and u4755 (Osthu6, J7fiu6, Q7fiu6);  // ../RTL/cortexm0ds_logic.v(5720)
  and u4756 (Q7fiu6, X7fiu6, E8fiu6);  // ../RTL/cortexm0ds_logic.v(5721)
  and u4757 (n1109, Lodpw6, L8fiu6);  // ../RTL/cortexm0ds_logic.v(5722)
  not u4758 (X7fiu6, n1109);  // ../RTL/cortexm0ds_logic.v(5722)
  and u4759 (J7fiu6, IRQ[6], S8fiu6);  // ../RTL/cortexm0ds_logic.v(5723)
  not u476 (Pkhpw6[0], n101[0]);  // ../RTL/cortexm0ds_logic.v(3356)
  and u4760 (n1110, Tk7iu6, Z8fiu6);  // ../RTL/cortexm0ds_logic.v(5724)
  not u4761 (S8fiu6, n1110);  // ../RTL/cortexm0ds_logic.v(5724)
  or u4762 (Z8fiu6, G9fiu6, Qg6iu6);  // ../RTL/cortexm0ds_logic.v(5725)
  and u4763 (Hsthu6, N9fiu6, U9fiu6);  // ../RTL/cortexm0ds_logic.v(5726)
  and u4764 (U9fiu6, Bafiu6, Iafiu6);  // ../RTL/cortexm0ds_logic.v(5727)
  and u4765 (n1111, Gpdpw6, Pafiu6);  // ../RTL/cortexm0ds_logic.v(5728)
  not u4766 (Bafiu6, n1111);  // ../RTL/cortexm0ds_logic.v(5728)
  and u4767 (N9fiu6, IRQ[5], Wafiu6);  // ../RTL/cortexm0ds_logic.v(5729)
  and u4768 (n1112, Tk7iu6, Dbfiu6);  // ../RTL/cortexm0ds_logic.v(5730)
  not u4769 (Wafiu6, n1112);  // ../RTL/cortexm0ds_logic.v(5730)
  buf u477 (X8hpw6[0], Hw8ax6);  // ../RTL/cortexm0ds_logic.v(2046)
  or u4770 (Dbfiu6, Kbfiu6, Qg6iu6);  // ../RTL/cortexm0ds_logic.v(5731)
  and u4771 (Asthu6, Rbfiu6, Ybfiu6);  // ../RTL/cortexm0ds_logic.v(5732)
  and u4772 (Ybfiu6, Fcfiu6, Mcfiu6);  // ../RTL/cortexm0ds_logic.v(5733)
  and u4773 (n1113, Qndpw6, Tcfiu6);  // ../RTL/cortexm0ds_logic.v(5734)
  not u4774 (Fcfiu6, n1113);  // ../RTL/cortexm0ds_logic.v(5734)
  and u4775 (Rbfiu6, IRQ[4], Adfiu6);  // ../RTL/cortexm0ds_logic.v(5735)
  and u4776 (n1114, Tk7iu6, Hdfiu6);  // ../RTL/cortexm0ds_logic.v(5736)
  not u4777 (Adfiu6, n1114);  // ../RTL/cortexm0ds_logic.v(5736)
  or u4778 (Hdfiu6, Qg6iu6, Odfiu6);  // ../RTL/cortexm0ds_logic.v(5737)
  and u4779 (Trthu6, Vdfiu6, Cefiu6);  // ../RTL/cortexm0ds_logic.v(5738)
  buf u478 (R2hpw6[0], Tyaax6);  // ../RTL/cortexm0ds_logic.v(2268)
  and u4780 (Cefiu6, Jefiu6, Qefiu6);  // ../RTL/cortexm0ds_logic.v(5739)
  and u4781 (n1115, Jndpw6, Xefiu6);  // ../RTL/cortexm0ds_logic.v(5740)
  not u4782 (Jefiu6, n1115);  // ../RTL/cortexm0ds_logic.v(5740)
  and u4783 (Vdfiu6, IRQ[3], Effiu6);  // ../RTL/cortexm0ds_logic.v(5741)
  and u4784 (n1116, Tk7iu6, Lffiu6);  // ../RTL/cortexm0ds_logic.v(5742)
  not u4785 (Effiu6, n1116);  // ../RTL/cortexm0ds_logic.v(5742)
  or u4786 (Lffiu6, Sffiu6, Qg6iu6);  // ../RTL/cortexm0ds_logic.v(5743)
  and u4787 (n1117, Zffiu6, Ggfiu6);  // ../RTL/cortexm0ds_logic.v(5744)
  not u4788 (Mrthu6, n1117);  // ../RTL/cortexm0ds_logic.v(5744)
  or u4789 (Ggfiu6, Ngfiu6, Cibiu6);  // ../RTL/cortexm0ds_logic.v(5745)
  buf u479 (Togpw6[2], Hlcax6);  // ../RTL/cortexm0ds_logic.v(2378)
  and u4790 (Zffiu6, Ugfiu6, Bhfiu6);  // ../RTL/cortexm0ds_logic.v(5746)
  and u4791 (n1118, Xibiu6, Ppfpw6[3]);  // ../RTL/cortexm0ds_logic.v(5747)
  not u4792 (Bhfiu6, n1118);  // ../RTL/cortexm0ds_logic.v(5747)
  and u4793 (Xibiu6, Ihfiu6, Phfiu6);  // ../RTL/cortexm0ds_logic.v(5748)
  or u4794 (n1119, Qaciu6, Qg6iu6);  // ../RTL/cortexm0ds_logic.v(5749)
  not u4795 (Phfiu6, n1119);  // ../RTL/cortexm0ds_logic.v(5749)
  or u4796 (n1120, Whfiu6, Difiu6);  // ../RTL/cortexm0ds_logic.v(5750)
  not u4797 (Qaciu6, n1120);  // ../RTL/cortexm0ds_logic.v(5750)
  and u4798 (Ihfiu6, Cibiu6, Ivfhu6);  // ../RTL/cortexm0ds_logic.v(5751)
  or u4799 (Ugfiu6, Ejbiu6, Kifiu6);  // ../RTL/cortexm0ds_logic.v(5752)
  buf u48 (vis_r2_o[12], U6rax6);  // ../RTL/cortexm0ds_logic.v(2551)
  buf u480 (Engpw6[27], Krbax6);  // ../RTL/cortexm0ds_logic.v(2368)
  and u4800 (n1121, Rifiu6, Cibiu6);  // ../RTL/cortexm0ds_logic.v(5753)
  not u4801 (Ejbiu6, n1121);  // ../RTL/cortexm0ds_logic.v(5753)
  and u4802 (Cibiu6, HREADY, Yifiu6);  // ../RTL/cortexm0ds_logic.v(5755)
  not u4803 (F8ciu6, Cibiu6);  // ../RTL/cortexm0ds_logic.v(5755)
  and u4804 (n1122, Uzaiu6, Fjfiu6);  // ../RTL/cortexm0ds_logic.v(5756)
  not u4805 (Yifiu6, n1122);  // ../RTL/cortexm0ds_logic.v(5756)
  or u4806 (n1123, Mjfiu6, Qg6iu6);  // ../RTL/cortexm0ds_logic.v(5757)
  not u4807 (Rifiu6, n1123);  // ../RTL/cortexm0ds_logic.v(5757)
  and u4808 (n1124, Xw4iu6, Tjfiu6);  // ../RTL/cortexm0ds_logic.v(5758)
  not u4809 (Frthu6, n1124);  // ../RTL/cortexm0ds_logic.v(5758)
  buf u481 (Plgpw6[27], Peeax6);  // ../RTL/cortexm0ds_logic.v(2369)
  and u4810 (n1125, Dhgpw6[3], Akfiu6);  // ../RTL/cortexm0ds_logic.v(5759)
  not u4811 (Tjfiu6, n1125);  // ../RTL/cortexm0ds_logic.v(5759)
  and u4812 (n1126, Scbiu6, Df4iu6);  // ../RTL/cortexm0ds_logic.v(5760)
  not u4813 (Akfiu6, n1126);  // ../RTL/cortexm0ds_logic.v(5760)
  and u4814 (n1127, Jehhu6, Hkfiu6);  // ../RTL/cortexm0ds_logic.v(5761)
  not u4815 (Xw4iu6, n1127);  // ../RTL/cortexm0ds_logic.v(5761)
  and u4816 (n1128, Okfiu6, Vkfiu6);  // ../RTL/cortexm0ds_logic.v(5762)
  not u4817 (Hkfiu6, n1128);  // ../RTL/cortexm0ds_logic.v(5762)
  and u4818 (n1129, S3hhu6, Ptaiu6);  // ../RTL/cortexm0ds_logic.v(5763)
  not u4819 (Vkfiu6, n1129);  // ../RTL/cortexm0ds_logic.v(5763)
  buf u482 (Akgpw6[27], Widax6);  // ../RTL/cortexm0ds_logic.v(2370)
  and u4820 (Ptaiu6, M2biu6, Clfiu6);  // ../RTL/cortexm0ds_logic.v(5764)
  and u4821 (n1130, H2hhu6, Mu4iu6);  // ../RTL/cortexm0ds_logic.v(5765)
  not u4822 (Okfiu6, n1130);  // ../RTL/cortexm0ds_logic.v(5765)
  and u4823 (Yqthu6, Jlfiu6, Qlfiu6);  // ../RTL/cortexm0ds_logic.v(5766)
  and u4824 (Qlfiu6, Xlfiu6, Jg6iu6);  // ../RTL/cortexm0ds_logic.v(5767)
  and u4825 (n1131, Ch5iu6, HWDATA[31]);  // ../RTL/cortexm0ds_logic.v(5768)
  not u4826 (Jg6iu6, n1131);  // ../RTL/cortexm0ds_logic.v(5768)
  and u4827 (n1132, Evdpw6, Af6iu6);  // ../RTL/cortexm0ds_logic.v(5769)
  not u4828 (Xlfiu6, n1132);  // ../RTL/cortexm0ds_logic.v(5769)
  or u4829 (Af6iu6, Emfiu6, Sb5iu6);  // ../RTL/cortexm0ds_logic.v(5770)
  buf u483 (vis_r14_o[28], Rribx6);  // ../RTL/cortexm0ds_logic.v(2497)
  and u4830 (Jlfiu6, NMI, Lmfiu6);  // ../RTL/cortexm0ds_logic.v(5771)
  and u4831 (n1133, Tk7iu6, Smfiu6);  // ../RTL/cortexm0ds_logic.v(5772)
  not u4832 (Lmfiu6, n1133);  // ../RTL/cortexm0ds_logic.v(5772)
  or u4833 (Smfiu6, Qg6iu6, Zmfiu6);  // ../RTL/cortexm0ds_logic.v(5773)
  and u4834 (n1134, Gnfiu6, Nnfiu6);  // ../RTL/cortexm0ds_logic.v(5774)
  not u4835 (Rqthu6, n1134);  // ../RTL/cortexm0ds_logic.v(5774)
  or u4836 (Nnfiu6, Unfiu6, Bofiu6);  // ../RTL/cortexm0ds_logic.v(5775)
  AL_MUX u4837 (
    .i0(Iofiu6),
    .i1(Ruaiu6),
    .sel(L3ehu6),
    .o(Bofiu6));  // ../RTL/cortexm0ds_logic.v(5776)
  and u4838 (n1135, Uzaiu6, Zmfiu6);  // ../RTL/cortexm0ds_logic.v(5777)
  not u4839 (Iofiu6, n1135);  // ../RTL/cortexm0ds_logic.v(5777)
  buf u484 (vis_r3_o[2], K1xax6);  // ../RTL/cortexm0ds_logic.v(2694)
  and u4840 (n1136, F2biu6, Sbghu6);  // ../RTL/cortexm0ds_logic.v(5778)
  not u4841 (Unfiu6, n1136);  // ../RTL/cortexm0ds_logic.v(5778)
  and u4842 (n1137, Jydhu6, T2biu6);  // ../RTL/cortexm0ds_logic.v(5779)
  not u4843 (Gnfiu6, n1137);  // ../RTL/cortexm0ds_logic.v(5779)
  and u4844 (n1138, HREADY, Pofiu6);  // ../RTL/cortexm0ds_logic.v(5780)
  not u4845 (T2biu6, n1138);  // ../RTL/cortexm0ds_logic.v(5780)
  or u4846 (Pofiu6, Wofiu6, C0ehu6);  // ../RTL/cortexm0ds_logic.v(5781)
  and u4847 (Kqthu6, Dpfiu6, Kpfiu6);  // ../RTL/cortexm0ds_logic.v(5782)
  and u4848 (Kpfiu6, Rpfiu6, Ypfiu6);  // ../RTL/cortexm0ds_logic.v(5783)
  and u4849 (n1139, Bqdpw6, Fqfiu6);  // ../RTL/cortexm0ds_logic.v(5784)
  buf u485 (Uthpw6[0], H3lpw6);  // ../RTL/cortexm0ds_logic.v(1882)
  not u4850 (Rpfiu6, n1139);  // ../RTL/cortexm0ds_logic.v(5784)
  and u4851 (Dpfiu6, IRQ[28], Mqfiu6);  // ../RTL/cortexm0ds_logic.v(5785)
  and u4852 (n1140, Tk7iu6, Tqfiu6);  // ../RTL/cortexm0ds_logic.v(5786)
  not u4853 (Mqfiu6, n1140);  // ../RTL/cortexm0ds_logic.v(5786)
  or u4854 (Tqfiu6, Qg6iu6, Arfiu6);  // ../RTL/cortexm0ds_logic.v(5787)
  and u4855 (Dqthu6, Hrfiu6, Orfiu6);  // ../RTL/cortexm0ds_logic.v(5788)
  and u4856 (Orfiu6, Vrfiu6, Csfiu6);  // ../RTL/cortexm0ds_logic.v(5789)
  and u4857 (n1141, Iqdpw6, Jsfiu6);  // ../RTL/cortexm0ds_logic.v(5790)
  not u4858 (Vrfiu6, n1141);  // ../RTL/cortexm0ds_logic.v(5790)
  and u4859 (Hrfiu6, IRQ[27], Qsfiu6);  // ../RTL/cortexm0ds_logic.v(5791)
  not u486 (Tugpw6[0], n1272[0]);  // ../RTL/cortexm0ds_logic.v(16030)
  and u4860 (n1142, Tk7iu6, Xsfiu6);  // ../RTL/cortexm0ds_logic.v(5792)
  not u4861 (Qsfiu6, n1142);  // ../RTL/cortexm0ds_logic.v(5792)
  or u4862 (Xsfiu6, Etfiu6, Qg6iu6);  // ../RTL/cortexm0ds_logic.v(5793)
  and u4863 (Wpthu6, Ltfiu6, Stfiu6);  // ../RTL/cortexm0ds_logic.v(5794)
  and u4864 (Stfiu6, Ztfiu6, Gufiu6);  // ../RTL/cortexm0ds_logic.v(5795)
  and u4865 (n1143, Pqdpw6, Nufiu6);  // ../RTL/cortexm0ds_logic.v(5796)
  not u4866 (Ztfiu6, n1143);  // ../RTL/cortexm0ds_logic.v(5796)
  and u4867 (Ltfiu6, IRQ[26], Uufiu6);  // ../RTL/cortexm0ds_logic.v(5797)
  and u4868 (n1144, Tk7iu6, Bvfiu6);  // ../RTL/cortexm0ds_logic.v(5798)
  not u4869 (Uufiu6, n1144);  // ../RTL/cortexm0ds_logic.v(5798)
  buf u487 (Gtgpw6[2], Opbax6);  // ../RTL/cortexm0ds_logic.v(2375)
  or u4870 (Bvfiu6, Ivfiu6, Qg6iu6);  // ../RTL/cortexm0ds_logic.v(5799)
  and u4871 (Ppthu6, Pvfiu6, Wvfiu6);  // ../RTL/cortexm0ds_logic.v(5800)
  and u4872 (Wvfiu6, Dwfiu6, Fe6iu6);  // ../RTL/cortexm0ds_logic.v(5801)
  and u4873 (n1145, Kwfiu6, HWDATA[25]);  // ../RTL/cortexm0ds_logic.v(5802)
  not u4874 (Fe6iu6, n1145);  // ../RTL/cortexm0ds_logic.v(5802)
  and u4875 (n1146, Krdpw6, Wc6iu6);  // ../RTL/cortexm0ds_logic.v(5803)
  not u4876 (Dwfiu6, n1146);  // ../RTL/cortexm0ds_logic.v(5803)
  or u4877 (Wc6iu6, Sb5iu6, Rwfiu6);  // ../RTL/cortexm0ds_logic.v(5804)
  and u4878 (Pvfiu6, IRQ[25], Ywfiu6);  // ../RTL/cortexm0ds_logic.v(5805)
  and u4879 (n1147, Tk7iu6, Fxfiu6);  // ../RTL/cortexm0ds_logic.v(5806)
  buf u488 (Trgpw6[2], Tceax6);  // ../RTL/cortexm0ds_logic.v(2376)
  not u4880 (Ywfiu6, n1147);  // ../RTL/cortexm0ds_logic.v(5806)
  or u4881 (Fxfiu6, Mxfiu6, Qg6iu6);  // ../RTL/cortexm0ds_logic.v(5807)
  and u4882 (Ipthu6, Txfiu6, Ayfiu6);  // ../RTL/cortexm0ds_logic.v(5808)
  and u4883 (Ayfiu6, Hyfiu6, Nb6iu6);  // ../RTL/cortexm0ds_logic.v(5809)
  and u4884 (n1148, Kwfiu6, HWDATA[24]);  // ../RTL/cortexm0ds_logic.v(5810)
  not u4885 (Nb6iu6, n1148);  // ../RTL/cortexm0ds_logic.v(5810)
  and u4886 (n1149, Wqdpw6, Ea6iu6);  // ../RTL/cortexm0ds_logic.v(5811)
  not u4887 (Hyfiu6, n1149);  // ../RTL/cortexm0ds_logic.v(5811)
  or u4888 (Ea6iu6, Sb5iu6, Oyfiu6);  // ../RTL/cortexm0ds_logic.v(5812)
  and u4889 (Txfiu6, IRQ[24], Vyfiu6);  // ../RTL/cortexm0ds_logic.v(5813)
  buf u489 (vis_r4_o[26], Wluax6);  // ../RTL/cortexm0ds_logic.v(2626)
  and u4890 (n1150, Tk7iu6, Czfiu6);  // ../RTL/cortexm0ds_logic.v(5814)
  not u4891 (Vyfiu6, n1150);  // ../RTL/cortexm0ds_logic.v(5814)
  or u4892 (Czfiu6, Qg6iu6, Jzfiu6);  // ../RTL/cortexm0ds_logic.v(5815)
  and u4893 (Bpthu6, Qzfiu6, Xzfiu6);  // ../RTL/cortexm0ds_logic.v(5816)
  and u4894 (Xzfiu6, E0giu6, L0giu6);  // ../RTL/cortexm0ds_logic.v(5817)
  and u4895 (n1151, Lvdpw6, S0giu6);  // ../RTL/cortexm0ds_logic.v(5818)
  not u4896 (E0giu6, n1151);  // ../RTL/cortexm0ds_logic.v(5818)
  and u4897 (Qzfiu6, IRQ[15], Z0giu6);  // ../RTL/cortexm0ds_logic.v(5819)
  and u4898 (n1152, Tk7iu6, G1giu6);  // ../RTL/cortexm0ds_logic.v(5820)
  not u4899 (Z0giu6, n1152);  // ../RTL/cortexm0ds_logic.v(5820)
  buf u49 (Uthpw6[7], Nckbx6);  // ../RTL/cortexm0ds_logic.v(1882)
  buf u490 (Vbgpw6[21], Nr0bx6);  // ../RTL/cortexm0ds_logic.v(3092)
  or u4900 (G1giu6, N1giu6, Qg6iu6);  // ../RTL/cortexm0ds_logic.v(5821)
  and u4901 (Uothu6, U1giu6, B2giu6);  // ../RTL/cortexm0ds_logic.v(5822)
  and u4902 (B2giu6, I2giu6, P2giu6);  // ../RTL/cortexm0ds_logic.v(5823)
  and u4903 (n1153, Otdpw6, W2giu6);  // ../RTL/cortexm0ds_logic.v(5824)
  not u4904 (I2giu6, n1153);  // ../RTL/cortexm0ds_logic.v(5824)
  and u4905 (U1giu6, IRQ[14], D3giu6);  // ../RTL/cortexm0ds_logic.v(5825)
  and u4906 (n1154, Tk7iu6, K3giu6);  // ../RTL/cortexm0ds_logic.v(5826)
  not u4907 (D3giu6, n1154);  // ../RTL/cortexm0ds_logic.v(5826)
  or u4908 (K3giu6, R3giu6, Qg6iu6);  // ../RTL/cortexm0ds_logic.v(5827)
  and u4909 (Nothu6, Y3giu6, F4giu6);  // ../RTL/cortexm0ds_logic.v(5828)
  buf u491 (Gqgpw6[2], Ahdax6);  // ../RTL/cortexm0ds_logic.v(2377)
  and u4910 (F4giu6, M4giu6, T4giu6);  // ../RTL/cortexm0ds_logic.v(5829)
  and u4911 (n1155, Vtdpw6, A5giu6);  // ../RTL/cortexm0ds_logic.v(5830)
  not u4912 (M4giu6, n1155);  // ../RTL/cortexm0ds_logic.v(5830)
  and u4913 (Y3giu6, IRQ[13], H5giu6);  // ../RTL/cortexm0ds_logic.v(5831)
  and u4914 (n1156, Tk7iu6, O5giu6);  // ../RTL/cortexm0ds_logic.v(5832)
  not u4915 (H5giu6, n1156);  // ../RTL/cortexm0ds_logic.v(5832)
  or u4916 (O5giu6, Qg6iu6, V5giu6);  // ../RTL/cortexm0ds_logic.v(5833)
  and u4917 (Gothu6, C6giu6, J6giu6);  // ../RTL/cortexm0ds_logic.v(5834)
  and u4918 (J6giu6, Q6giu6, X6giu6);  // ../RTL/cortexm0ds_logic.v(5835)
  and u4919 (n1157, Qudpw6, E7giu6);  // ../RTL/cortexm0ds_logic.v(5836)
  buf u492 (R0nhu6, Wvgax6);  // ../RTL/cortexm0ds_logic.v(2382)
  not u4920 (Q6giu6, n1157);  // ../RTL/cortexm0ds_logic.v(5836)
  and u4921 (C6giu6, IRQ[12], L7giu6);  // ../RTL/cortexm0ds_logic.v(5837)
  and u4922 (n1158, Tk7iu6, S7giu6);  // ../RTL/cortexm0ds_logic.v(5838)
  not u4923 (L7giu6, n1158);  // ../RTL/cortexm0ds_logic.v(5838)
  or u4924 (S7giu6, Qg6iu6, Z7giu6);  // ../RTL/cortexm0ds_logic.v(5839)
  and u4925 (Znthu6, G8giu6, N8giu6);  // ../RTL/cortexm0ds_logic.v(5840)
  and u4926 (N8giu6, U8giu6, B9giu6);  // ../RTL/cortexm0ds_logic.v(5841)
  and u4927 (n1159, Cudpw6, I9giu6);  // ../RTL/cortexm0ds_logic.v(5842)
  not u4928 (U8giu6, n1159);  // ../RTL/cortexm0ds_logic.v(5842)
  and u4929 (G8giu6, IRQ[11], P9giu6);  // ../RTL/cortexm0ds_logic.v(5843)
  buf u493 (Jzmhu6, Jxgax6);  // ../RTL/cortexm0ds_logic.v(2383)
  and u4930 (n1160, Tk7iu6, W9giu6);  // ../RTL/cortexm0ds_logic.v(5844)
  not u4931 (P9giu6, n1160);  // ../RTL/cortexm0ds_logic.v(5844)
  or u4932 (W9giu6, Dagiu6, Qg6iu6);  // ../RTL/cortexm0ds_logic.v(5845)
  and u4933 (Snthu6, Kagiu6, Ragiu6);  // ../RTL/cortexm0ds_logic.v(5846)
  and u4934 (Ragiu6, Yagiu6, Fbgiu6);  // ../RTL/cortexm0ds_logic.v(5847)
  and u4935 (n1161, Judpw6, Mbgiu6);  // ../RTL/cortexm0ds_logic.v(5848)
  not u4936 (Yagiu6, n1161);  // ../RTL/cortexm0ds_logic.v(5848)
  and u4937 (Kagiu6, IRQ[10], Tbgiu6);  // ../RTL/cortexm0ds_logic.v(5849)
  and u4938 (n1162, Tk7iu6, Acgiu6);  // ../RTL/cortexm0ds_logic.v(5850)
  not u4939 (Tbgiu6, n1162);  // ../RTL/cortexm0ds_logic.v(5850)
  buf u494 (Sbghu6, Vygax6);  // ../RTL/cortexm0ds_logic.v(2384)
  or u4940 (Acgiu6, Hcgiu6, Qg6iu6);  // ../RTL/cortexm0ds_logic.v(5851)
  and u4941 (Lnthu6, Ocgiu6, Vcgiu6);  // ../RTL/cortexm0ds_logic.v(5852)
  and u4942 (Vcgiu6, Cdgiu6, J96iu6);  // ../RTL/cortexm0ds_logic.v(5853)
  and u4943 (n1163, Kwfiu6, HWDATA[9]);  // ../RTL/cortexm0ds_logic.v(5854)
  not u4944 (J96iu6, n1163);  // ../RTL/cortexm0ds_logic.v(5854)
  and u4945 (n1164, Cndpw6, A86iu6);  // ../RTL/cortexm0ds_logic.v(5855)
  not u4946 (Cdgiu6, n1164);  // ../RTL/cortexm0ds_logic.v(5855)
  or u4947 (A86iu6, Sb5iu6, Jdgiu6);  // ../RTL/cortexm0ds_logic.v(5856)
  and u4948 (Ocgiu6, IRQ[9], Qdgiu6);  // ../RTL/cortexm0ds_logic.v(5857)
  and u4949 (n1165, Tk7iu6, Xdgiu6);  // ../RTL/cortexm0ds_logic.v(5858)
  buf u495 (vis_r1_o[17], Y9upw6);  // ../RTL/cortexm0ds_logic.v(1876)
  not u4950 (Qdgiu6, n1165);  // ../RTL/cortexm0ds_logic.v(5858)
  or u4951 (Xdgiu6, Eegiu6, Qg6iu6);  // ../RTL/cortexm0ds_logic.v(5859)
  and u4952 (Enthu6, Legiu6, Segiu6);  // ../RTL/cortexm0ds_logic.v(5860)
  and u4953 (Segiu6, Zegiu6, W56iu6);  // ../RTL/cortexm0ds_logic.v(5861)
  and u4954 (n1166, Kwfiu6, HWDATA[8]);  // ../RTL/cortexm0ds_logic.v(5862)
  not u4955 (W56iu6, n1166);  // ../RTL/cortexm0ds_logic.v(5862)
  and u4956 (n1167, Sodpw6, N46iu6);  // ../RTL/cortexm0ds_logic.v(5863)
  not u4957 (Zegiu6, n1167);  // ../RTL/cortexm0ds_logic.v(5863)
  or u4958 (N46iu6, Sb5iu6, Gfgiu6);  // ../RTL/cortexm0ds_logic.v(5864)
  and u4959 (Legiu6, IRQ[8], Nfgiu6);  // ../RTL/cortexm0ds_logic.v(5865)
  buf u496 (vis_r1_o[18], P4xpw6);  // ../RTL/cortexm0ds_logic.v(1876)
  and u4960 (n1168, Tk7iu6, Ufgiu6);  // ../RTL/cortexm0ds_logic.v(5866)
  not u4961 (Nfgiu6, n1168);  // ../RTL/cortexm0ds_logic.v(5866)
  or u4962 (Ufgiu6, Qg6iu6, Bggiu6);  // ../RTL/cortexm0ds_logic.v(5867)
  and u4963 (n1169, Iggiu6, Pggiu6);  // ../RTL/cortexm0ds_logic.v(5868)
  not u4964 (Xmthu6, n1169);  // ../RTL/cortexm0ds_logic.v(5868)
  and u4965 (n1170, Ch5iu6, HWDATA[28]);  // ../RTL/cortexm0ds_logic.v(5869)
  not u4966 (Pggiu6, n1170);  // ../RTL/cortexm0ds_logic.v(5869)
  and u4967 (n1171, Wggiu6, Ikghu6);  // ../RTL/cortexm0ds_logic.v(5870)
  not u4968 (Iggiu6, n1171);  // ../RTL/cortexm0ds_logic.v(5870)
  and u4969 (Wggiu6, Dhgiu6, Khgiu6);  // ../RTL/cortexm0ds_logic.v(5871)
  buf u497 (vis_r1_o[19], Jlvpw6);  // ../RTL/cortexm0ds_logic.v(1876)
  and u4970 (n1172, Ch5iu6, HWDATA[27]);  // ../RTL/cortexm0ds_logic.v(5872)
  not u4971 (Khgiu6, n1172);  // ../RTL/cortexm0ds_logic.v(5872)
  and u4972 (n1173, Clfiu6, Rhgiu6);  // ../RTL/cortexm0ds_logic.v(5873)
  not u4973 (Dhgiu6, n1173);  // ../RTL/cortexm0ds_logic.v(5873)
  and u4974 (n1174, Ag5iu6, Yhgiu6);  // ../RTL/cortexm0ds_logic.v(5874)
  not u4975 (Qmthu6, n1174);  // ../RTL/cortexm0ds_logic.v(5874)
  and u4976 (n1175, Figiu6, Yyghu6);  // ../RTL/cortexm0ds_logic.v(5875)
  not u4977 (Yhgiu6, n1175);  // ../RTL/cortexm0ds_logic.v(5875)
  and u4978 (Figiu6, Migiu6, Tigiu6);  // ../RTL/cortexm0ds_logic.v(5876)
  and u4979 (n1176, Ch5iu6, HWDATA[25]);  // ../RTL/cortexm0ds_logic.v(5877)
  buf u498 (vis_r1_o[20], I3qpw6);  // ../RTL/cortexm0ds_logic.v(1876)
  not u4980 (Tigiu6, n1176);  // ../RTL/cortexm0ds_logic.v(5877)
  and u4981 (n1177, Clfiu6, Ajgiu6);  // ../RTL/cortexm0ds_logic.v(5878)
  not u4982 (Migiu6, n1177);  // ../RTL/cortexm0ds_logic.v(5878)
  and u4983 (Ag5iu6, Hjgiu6, Ojgiu6);  // ../RTL/cortexm0ds_logic.v(5879)
  and u4984 (n1178, Vjgiu6, Ckgiu6);  // ../RTL/cortexm0ds_logic.v(5880)
  not u4985 (Ojgiu6, n1178);  // ../RTL/cortexm0ds_logic.v(5880)
  and u4986 (Vjgiu6, Dvghu6, Tzfpw6[0]);  // ../RTL/cortexm0ds_logic.v(5881)
  and u4987 (n1179, Ch5iu6, HWDATA[26]);  // ../RTL/cortexm0ds_logic.v(5882)
  not u4988 (Hjgiu6, n1179);  // ../RTL/cortexm0ds_logic.v(5882)
  or u4989 (n1180, Jkgiu6, Qkgiu6);  // ../RTL/cortexm0ds_logic.v(5883)
  buf u499 (vis_r1_o[23], Gx6ax6);  // ../RTL/cortexm0ds_logic.v(1876)
  not u4990 (Ch5iu6, n1180);  // ../RTL/cortexm0ds_logic.v(5883)
  and u4991 (Jmthu6, Xkgiu6, Elgiu6);  // ../RTL/cortexm0ds_logic.v(5884)
  and u4992 (Elgiu6, Llgiu6, Slgiu6);  // ../RTL/cortexm0ds_logic.v(5885)
  and u4993 (n1181, Eodpw6, Zlgiu6);  // ../RTL/cortexm0ds_logic.v(5886)
  not u4994 (Llgiu6, n1181);  // ../RTL/cortexm0ds_logic.v(5886)
  and u4995 (Xkgiu6, IRQ[2], Gmgiu6);  // ../RTL/cortexm0ds_logic.v(5887)
  and u4996 (n1182, Tk7iu6, Nmgiu6);  // ../RTL/cortexm0ds_logic.v(5888)
  not u4997 (Gmgiu6, n1182);  // ../RTL/cortexm0ds_logic.v(5888)
  or u4998 (Nmgiu6, Qg6iu6, Umgiu6);  // ../RTL/cortexm0ds_logic.v(5889)
  and u4999 (Cmthu6, Bngiu6, Ingiu6);  // ../RTL/cortexm0ds_logic.v(5890)
  buf u5 (HMASTLOCK, 1'b0);  // ../RTL/cortexm0ds_logic.v(1728)
  buf u50 (Jshpw6[31], Ydgax6);  // ../RTL/cortexm0ds_logic.v(2372)
  buf u500 (vis_r1_o[24], Ypspw6);  // ../RTL/cortexm0ds_logic.v(1876)
  and u5000 (Ingiu6, Pngiu6, Wngiu6);  // ../RTL/cortexm0ds_logic.v(5891)
  and u5001 (n1183, Fsdpw6, Dogiu6);  // ../RTL/cortexm0ds_logic.v(5892)
  not u5002 (Pngiu6, n1183);  // ../RTL/cortexm0ds_logic.v(5892)
  and u5003 (Bngiu6, IRQ[1], Kogiu6);  // ../RTL/cortexm0ds_logic.v(5893)
  and u5004 (n1184, Tk7iu6, Rogiu6);  // ../RTL/cortexm0ds_logic.v(5894)
  not u5005 (Kogiu6, n1184);  // ../RTL/cortexm0ds_logic.v(5894)
  or u5006 (Rogiu6, Qg6iu6, Yogiu6);  // ../RTL/cortexm0ds_logic.v(5895)
  AL_MUX u5007 (
    .i0(I4eiu6),
    .i1(Qqdhu6),
    .sel(P3fiu6),
    .o(Vlthu6));  // ../RTL/cortexm0ds_logic.v(5896)
  AL_MUX u5008 (
    .i0(G3eiu6),
    .i1(Ndghu6),
    .sel(P3fiu6),
    .o(Olthu6));  // ../RTL/cortexm0ds_logic.v(5897)
  and u5009 (n1185, Fpgiu6, Npdhu6);  // ../RTL/cortexm0ds_logic.v(5898)
  buf u501 (vis_r1_o[25], Z3tpw6);  // ../RTL/cortexm0ds_logic.v(1876)
  not u5010 (P3fiu6, n1185);  // ../RTL/cortexm0ds_logic.v(5898)
  AL_MUX u5011 (
    .i0(HWDATA[30]),
    .i1(B3gpw6[0]),
    .sel(Mpgiu6),
    .o(Hlthu6));  // ../RTL/cortexm0ds_logic.v(5899)
  AL_MUX u5012 (
    .i0(HWDATA[31]),
    .i1(B3gpw6[1]),
    .sel(Mpgiu6),
    .o(Althu6));  // ../RTL/cortexm0ds_logic.v(5900)
  or u5013 (Mpgiu6, Tpgiu6, Jkgiu6);  // ../RTL/cortexm0ds_logic.v(5901)
  AL_MUX u5014 (
    .i0(HWDATA[22]),
    .i1(L1gpw6[0]),
    .sel(Aqgiu6),
    .o(Tkthu6));  // ../RTL/cortexm0ds_logic.v(5902)
  AL_MUX u5015 (
    .i0(HWDATA[23]),
    .i1(L1gpw6[1]),
    .sel(Aqgiu6),
    .o(Mkthu6));  // ../RTL/cortexm0ds_logic.v(5903)
  AL_MUX u5016 (
    .i0(HWDATA[30]),
    .i1(H8gpw6[0]),
    .sel(Aqgiu6),
    .o(Fkthu6));  // ../RTL/cortexm0ds_logic.v(5904)
  AL_MUX u5017 (
    .i0(HWDATA[31]),
    .i1(H8gpw6[1]),
    .sel(Aqgiu6),
    .o(Yjthu6));  // ../RTL/cortexm0ds_logic.v(5905)
  and u5018 (n1186, Hqgiu6, Npdhu6);  // ../RTL/cortexm0ds_logic.v(5906)
  not u5019 (Aqgiu6, n1186);  // ../RTL/cortexm0ds_logic.v(5906)
  buf u502 (vis_r1_o[26], Xvtpw6);  // ../RTL/cortexm0ds_logic.v(1876)
  and u5020 (n1187, Qh5iu6, Oqgiu6);  // ../RTL/cortexm0ds_logic.v(5907)
  not u5021 (Rjthu6, n1187);  // ../RTL/cortexm0ds_logic.v(5907)
  and u5022 (n1188, Vqgiu6, Zlghu6);  // ../RTL/cortexm0ds_logic.v(5908)
  not u5023 (Oqgiu6, n1188);  // ../RTL/cortexm0ds_logic.v(5908)
  and u5024 (Vqgiu6, Crgiu6, Jrgiu6);  // ../RTL/cortexm0ds_logic.v(5909)
  and u5025 (n1189, Clfiu6, Qrgiu6);  // ../RTL/cortexm0ds_logic.v(5910)
  not u5026 (Jrgiu6, n1189);  // ../RTL/cortexm0ds_logic.v(5910)
  and u5027 (n1190, Xrgiu6, Npdhu6);  // ../RTL/cortexm0ds_logic.v(5911)
  not u5028 (Crgiu6, n1190);  // ../RTL/cortexm0ds_logic.v(5911)
  and u5029 (Qh5iu6, Esgiu6, Lsgiu6);  // ../RTL/cortexm0ds_logic.v(5912)
  buf u503 (vis_r1_o[27], Ixppw6);  // ../RTL/cortexm0ds_logic.v(1876)
  and u5030 (n1191, P0biu6, Ssgiu6);  // ../RTL/cortexm0ds_logic.v(5913)
  not u5031 (Lsgiu6, n1191);  // ../RTL/cortexm0ds_logic.v(5913)
  and u5032 (n1192, I0biu6, Zsgiu6);  // ../RTL/cortexm0ds_logic.v(5914)
  not u5033 (Ssgiu6, n1192);  // ../RTL/cortexm0ds_logic.v(5914)
  or u5034 (Zsgiu6, Gtgiu6, Ntgiu6);  // ../RTL/cortexm0ds_logic.v(5915)
  and u5035 (n1193, Utgiu6, Bugiu6);  // ../RTL/cortexm0ds_logic.v(5916)
  not u5036 (I0biu6, n1193);  // ../RTL/cortexm0ds_logic.v(5916)
  or u5037 (n1194, Ae0iu6, Cyfpw6[4]);  // ../RTL/cortexm0ds_logic.v(5917)
  not u5038 (Bugiu6, n1194);  // ../RTL/cortexm0ds_logic.v(5917)
  and u5039 (Utgiu6, Iugiu6, Pugiu6);  // ../RTL/cortexm0ds_logic.v(5918)
  buf u504 (vis_r1_o[28], I9qpw6);  // ../RTL/cortexm0ds_logic.v(1876)
  and u5040 (n1195, Xrgiu6, Fsdiu6);  // ../RTL/cortexm0ds_logic.v(5919)
  not u5041 (Esgiu6, n1195);  // ../RTL/cortexm0ds_logic.v(5919)
  and u5042 (n1196, Wugiu6, Dvgiu6);  // ../RTL/cortexm0ds_logic.v(5920)
  not u5043 (Kjthu6, n1196);  // ../RTL/cortexm0ds_logic.v(5920)
  and u5044 (n1197, Kvgiu6, Krghu6);  // ../RTL/cortexm0ds_logic.v(5921)
  not u5045 (Dvgiu6, n1197);  // ../RTL/cortexm0ds_logic.v(5921)
  and u5046 (Kvgiu6, Rvgiu6, Hzeiu6);  // ../RTL/cortexm0ds_logic.v(5922)
  and u5047 (Myeiu6, Yvgiu6, Npdhu6);  // ../RTL/cortexm0ds_logic.v(5923)
  not u5048 (Hzeiu6, Myeiu6);  // ../RTL/cortexm0ds_logic.v(5923)
  and u5049 (n1198, Fwgiu6, Y5eiu6);  // ../RTL/cortexm0ds_logic.v(5924)
  buf u505 (vis_r1_o[30], Weipw6);  // ../RTL/cortexm0ds_logic.v(1876)
  not u5050 (Rvgiu6, n1198);  // ../RTL/cortexm0ds_logic.v(5924)
  and u5051 (Fwgiu6, Ur4iu6, Jkgiu6);  // ../RTL/cortexm0ds_logic.v(5925)
  and u5052 (n1199, Ckgiu6, Tzfpw6[0]);  // ../RTL/cortexm0ds_logic.v(5926)
  not u5053 (Wugiu6, n1199);  // ../RTL/cortexm0ds_logic.v(5926)
  and u5054 (Ckgiu6, Ozeiu6, Azeiu6);  // ../RTL/cortexm0ds_logic.v(5927)
  and u5055 (Azeiu6, Mwgiu6, Twgiu6);  // ../RTL/cortexm0ds_logic.v(5928)
  and u5056 (Twgiu6, Axgiu6, Hxgiu6);  // ../RTL/cortexm0ds_logic.v(5929)
  and u5057 (Hxgiu6, Oxgiu6, Vxgiu6);  // ../RTL/cortexm0ds_logic.v(5930)
  or u5058 (n1200, Cygiu6, Tzfpw6[7]);  // ../RTL/cortexm0ds_logic.v(5931)
  not u5059 (Vxgiu6, n1200);  // ../RTL/cortexm0ds_logic.v(5931)
  buf u506 (vis_r1_o[31], Ejnpw6);  // ../RTL/cortexm0ds_logic.v(1876)
  or u5060 (Cygiu6, Tzfpw6[8], Tzfpw6[9]);  // ../RTL/cortexm0ds_logic.v(5932)
  or u5061 (n1201, Jygiu6, Tzfpw6[4]);  // ../RTL/cortexm0ds_logic.v(5933)
  not u5062 (Oxgiu6, n1201);  // ../RTL/cortexm0ds_logic.v(5933)
  or u5063 (Jygiu6, Tzfpw6[5], Tzfpw6[6]);  // ../RTL/cortexm0ds_logic.v(5934)
  and u5064 (Axgiu6, Qygiu6, Xygiu6);  // ../RTL/cortexm0ds_logic.v(5935)
  or u5065 (n1202, Ezgiu6, Tzfpw6[23]);  // ../RTL/cortexm0ds_logic.v(5936)
  not u5066 (Xygiu6, n1202);  // ../RTL/cortexm0ds_logic.v(5936)
  or u5067 (Ezgiu6, Tzfpw6[2], Tzfpw6[3]);  // ../RTL/cortexm0ds_logic.v(5937)
  or u5068 (n1203, Lzgiu6, Tzfpw6[20]);  // ../RTL/cortexm0ds_logic.v(5938)
  not u5069 (Qygiu6, n1203);  // ../RTL/cortexm0ds_logic.v(5938)
  buf u507 (vis_r12_o[1], Fatax6);  // ../RTL/cortexm0ds_logic.v(2599)
  or u5070 (Lzgiu6, Tzfpw6[21], Tzfpw6[22]);  // ../RTL/cortexm0ds_logic.v(5939)
  and u5071 (Mwgiu6, Szgiu6, Zzgiu6);  // ../RTL/cortexm0ds_logic.v(5940)
  and u5072 (Zzgiu6, G0hiu6, N0hiu6);  // ../RTL/cortexm0ds_logic.v(5941)
  or u5073 (n1204, U0hiu6, Tzfpw6[18]);  // ../RTL/cortexm0ds_logic.v(5942)
  not u5074 (N0hiu6, n1204);  // ../RTL/cortexm0ds_logic.v(5942)
  or u5075 (U0hiu6, Tzfpw6[19], Tzfpw6[1]);  // ../RTL/cortexm0ds_logic.v(5943)
  or u5076 (n1205, B1hiu6, Tzfpw6[15]);  // ../RTL/cortexm0ds_logic.v(5944)
  not u5077 (G0hiu6, n1205);  // ../RTL/cortexm0ds_logic.v(5944)
  or u5078 (B1hiu6, Tzfpw6[16], Tzfpw6[17]);  // ../RTL/cortexm0ds_logic.v(5945)
  and u5079 (Szgiu6, I1hiu6, P1hiu6);  // ../RTL/cortexm0ds_logic.v(5946)
  buf u508 (vis_r12_o[5], Iwsax6);  // ../RTL/cortexm0ds_logic.v(2599)
  or u5080 (n1206, W1hiu6, Tzfpw6[12]);  // ../RTL/cortexm0ds_logic.v(5947)
  not u5081 (P1hiu6, n1206);  // ../RTL/cortexm0ds_logic.v(5947)
  or u5082 (W1hiu6, Tzfpw6[13], Tzfpw6[14]);  // ../RTL/cortexm0ds_logic.v(5948)
  or u5083 (n1207, Tzfpw6[10], Tzfpw6[11]);  // ../RTL/cortexm0ds_logic.v(5949)
  not u5084 (I1hiu6, n1207);  // ../RTL/cortexm0ds_logic.v(5949)
  and u5085 (Ozeiu6, D2hiu6, Bxghu6);  // ../RTL/cortexm0ds_logic.v(5950)
  and u5086 (D2hiu6, Gc5iu6, K2hiu6);  // ../RTL/cortexm0ds_logic.v(5951)
  or u5087 (K2hiu6, R2hiu6, STCALIB[25]);  // ../RTL/cortexm0ds_logic.v(5952)
  or u5088 (R2hiu6, Ftghu6, STCLKEN);  // ../RTL/cortexm0ds_logic.v(5953)
  and u5089 (n1208, Y2hiu6, F3hiu6);  // ../RTL/cortexm0ds_logic.v(5954)
  buf u509 (vis_r12_o[7], G0tax6);  // ../RTL/cortexm0ds_logic.v(2599)
  not u5090 (Djthu6, n1208);  // ../RTL/cortexm0ds_logic.v(5954)
  and u5091 (F3hiu6, M3hiu6, T3hiu6);  // ../RTL/cortexm0ds_logic.v(5955)
  and u5092 (n1209, HRDATA[7], Pp7iu6);  // ../RTL/cortexm0ds_logic.v(5956)
  not u5093 (T3hiu6, n1209);  // ../RTL/cortexm0ds_logic.v(5956)
  and u5094 (M3hiu6, A4hiu6, H4hiu6);  // ../RTL/cortexm0ds_logic.v(5957)
  and u5095 (n1210, Hrfpw6[7], Uy4iu6);  // ../RTL/cortexm0ds_logic.v(5958)
  not u5096 (H4hiu6, n1210);  // ../RTL/cortexm0ds_logic.v(5958)
  and u5097 (n1211, HRDATA[23], Kq7iu6);  // ../RTL/cortexm0ds_logic.v(5959)
  not u5098 (A4hiu6, n1211);  // ../RTL/cortexm0ds_logic.v(5959)
  and u5099 (Y2hiu6, O4hiu6, V4hiu6);  // ../RTL/cortexm0ds_logic.v(5960)
  buf u51 (Tzfpw6[0], N8rpw6);  // ../RTL/cortexm0ds_logic.v(2007)
  buf u510 (vis_r12_o[8], Eytax6);  // ../RTL/cortexm0ds_logic.v(2599)
  and u5100 (n1212, Fr7iu6, Df4iu6);  // ../RTL/cortexm0ds_logic.v(5961)
  not u5101 (V4hiu6, n1212);  // ../RTL/cortexm0ds_logic.v(5961)
  and u5102 (O4hiu6, C5hiu6, J5hiu6);  // ../RTL/cortexm0ds_logic.v(5962)
  and u5103 (n1213, A25iu6, Ppfpw6[7]);  // ../RTL/cortexm0ds_logic.v(5963)
  not u5104 (J5hiu6, n1213);  // ../RTL/cortexm0ds_logic.v(5963)
  and u5105 (n1214, R05iu6, D7fpw6[7]);  // ../RTL/cortexm0ds_logic.v(5964)
  not u5106 (C5hiu6, n1214);  // ../RTL/cortexm0ds_logic.v(5964)
  and u5107 (n1215, Q5hiu6, X5hiu6);  // ../RTL/cortexm0ds_logic.v(5965)
  not u5108 (Withu6, n1215);  // ../RTL/cortexm0ds_logic.v(5965)
  and u5109 (X5hiu6, E6hiu6, L6hiu6);  // ../RTL/cortexm0ds_logic.v(5966)
  buf u511 (vis_r12_o[9], Rvibx6);  // ../RTL/cortexm0ds_logic.v(2599)
  and u5110 (n1216, HRDATA[6], Pp7iu6);  // ../RTL/cortexm0ds_logic.v(5967)
  not u5111 (L6hiu6, n1216);  // ../RTL/cortexm0ds_logic.v(5967)
  and u5112 (E6hiu6, S6hiu6, Z6hiu6);  // ../RTL/cortexm0ds_logic.v(5968)
  and u5113 (n1217, Hrfpw6[6], Uy4iu6);  // ../RTL/cortexm0ds_logic.v(5969)
  not u5114 (Z6hiu6, n1217);  // ../RTL/cortexm0ds_logic.v(5969)
  and u5115 (n1218, HRDATA[22], Kq7iu6);  // ../RTL/cortexm0ds_logic.v(5970)
  not u5116 (S6hiu6, n1218);  // ../RTL/cortexm0ds_logic.v(5970)
  and u5117 (Q5hiu6, G7hiu6, N7hiu6);  // ../RTL/cortexm0ds_logic.v(5971)
  and u5118 (n1219, A25iu6, Ppfpw6[6]);  // ../RTL/cortexm0ds_logic.v(5972)
  not u5119 (N7hiu6, n1219);  // ../RTL/cortexm0ds_logic.v(5972)
  buf u512 (vis_r12_o[10], Ewtax6);  // ../RTL/cortexm0ds_logic.v(2599)
  and u5120 (n1220, R05iu6, D7fpw6[6]);  // ../RTL/cortexm0ds_logic.v(5973)
  not u5121 (G7hiu6, n1220);  // ../RTL/cortexm0ds_logic.v(5973)
  and u5122 (n1221, U7hiu6, B8hiu6);  // ../RTL/cortexm0ds_logic.v(5974)
  not u5123 (Pithu6, n1221);  // ../RTL/cortexm0ds_logic.v(5974)
  and u5124 (B8hiu6, I8hiu6, P8hiu6);  // ../RTL/cortexm0ds_logic.v(5975)
  and u5125 (n1222, HRDATA[5], Pp7iu6);  // ../RTL/cortexm0ds_logic.v(5976)
  not u5126 (P8hiu6, n1222);  // ../RTL/cortexm0ds_logic.v(5976)
  and u5127 (I8hiu6, W8hiu6, D9hiu6);  // ../RTL/cortexm0ds_logic.v(5977)
  and u5128 (n1223, Hrfpw6[5], Uy4iu6);  // ../RTL/cortexm0ds_logic.v(5978)
  not u5129 (D9hiu6, n1223);  // ../RTL/cortexm0ds_logic.v(5978)
  buf u513 (vis_r12_o[11], Zn8bx6);  // ../RTL/cortexm0ds_logic.v(2599)
  and u5130 (n1224, HRDATA[21], Kq7iu6);  // ../RTL/cortexm0ds_logic.v(5979)
  not u5131 (W8hiu6, n1224);  // ../RTL/cortexm0ds_logic.v(5979)
  and u5132 (U7hiu6, K9hiu6, R9hiu6);  // ../RTL/cortexm0ds_logic.v(5980)
  and u5133 (n1225, Ppfpw6[5], A25iu6);  // ../RTL/cortexm0ds_logic.v(5981)
  not u5134 (R9hiu6, n1225);  // ../RTL/cortexm0ds_logic.v(5981)
  and u5135 (n1226, R05iu6, D7fpw6[5]);  // ../RTL/cortexm0ds_logic.v(5982)
  not u5136 (K9hiu6, n1226);  // ../RTL/cortexm0ds_logic.v(5982)
  and u5137 (n1227, Y9hiu6, Fahiu6);  // ../RTL/cortexm0ds_logic.v(5983)
  not u5138 (Iithu6, n1227);  // ../RTL/cortexm0ds_logic.v(5983)
  and u5139 (Fahiu6, Mahiu6, Tahiu6);  // ../RTL/cortexm0ds_logic.v(5984)
  buf u514 (Sqhpw6[0], Sqfax6);  // ../RTL/cortexm0ds_logic.v(2359)
  and u5140 (n1228, HRDATA[4], Pp7iu6);  // ../RTL/cortexm0ds_logic.v(5985)
  not u5141 (Tahiu6, n1228);  // ../RTL/cortexm0ds_logic.v(5985)
  and u5142 (Mahiu6, Abhiu6, Hbhiu6);  // ../RTL/cortexm0ds_logic.v(5986)
  and u5143 (n1229, Hrfpw6[4], Uy4iu6);  // ../RTL/cortexm0ds_logic.v(5987)
  not u5144 (Hbhiu6, n1229);  // ../RTL/cortexm0ds_logic.v(5987)
  and u5145 (n1230, HRDATA[20], Kq7iu6);  // ../RTL/cortexm0ds_logic.v(5988)
  not u5146 (Abhiu6, n1230);  // ../RTL/cortexm0ds_logic.v(5988)
  and u5147 (Y9hiu6, Obhiu6, Vbhiu6);  // ../RTL/cortexm0ds_logic.v(5989)
  and u5148 (n1231, Ppfpw6[4], A25iu6);  // ../RTL/cortexm0ds_logic.v(5990)
  not u5149 (Vbhiu6, n1231);  // ../RTL/cortexm0ds_logic.v(5990)
  buf u515 (K7hpw6[15], Rg9ax6);  // ../RTL/cortexm0ds_logic.v(2366)
  and u5150 (n1232, R05iu6, D7fpw6[4]);  // ../RTL/cortexm0ds_logic.v(5991)
  not u5151 (Obhiu6, n1232);  // ../RTL/cortexm0ds_logic.v(5991)
  and u5152 (n1233, Cchiu6, Jchiu6);  // ../RTL/cortexm0ds_logic.v(5992)
  not u5153 (Bithu6, n1233);  // ../RTL/cortexm0ds_logic.v(5992)
  and u5154 (Jchiu6, Qchiu6, Xchiu6);  // ../RTL/cortexm0ds_logic.v(5993)
  and u5155 (n1234, HRDATA[3], Pp7iu6);  // ../RTL/cortexm0ds_logic.v(5994)
  not u5156 (Xchiu6, n1234);  // ../RTL/cortexm0ds_logic.v(5994)
  and u5157 (Qchiu6, Edhiu6, Ldhiu6);  // ../RTL/cortexm0ds_logic.v(5995)
  and u5158 (n1235, Hrfpw6[3], Uy4iu6);  // ../RTL/cortexm0ds_logic.v(5996)
  not u5159 (Ldhiu6, n1235);  // ../RTL/cortexm0ds_logic.v(5996)
  buf u516 (K7hpw6[14], Qkabx6);  // ../RTL/cortexm0ds_logic.v(2366)
  and u5160 (n1236, HRDATA[19], Kq7iu6);  // ../RTL/cortexm0ds_logic.v(5997)
  not u5161 (Edhiu6, n1236);  // ../RTL/cortexm0ds_logic.v(5997)
  and u5162 (Cchiu6, Sdhiu6, Zdhiu6);  // ../RTL/cortexm0ds_logic.v(5998)
  and u5163 (n1237, Fr7iu6, H34iu6);  // ../RTL/cortexm0ds_logic.v(5999)
  not u5164 (Zdhiu6, n1237);  // ../RTL/cortexm0ds_logic.v(5999)
  and u5165 (Sdhiu6, Gehiu6, Nehiu6);  // ../RTL/cortexm0ds_logic.v(6000)
  and u5166 (n1238, Ppfpw6[3], A25iu6);  // ../RTL/cortexm0ds_logic.v(6001)
  not u5167 (Nehiu6, n1238);  // ../RTL/cortexm0ds_logic.v(6001)
  and u5168 (n1239, R05iu6, D7fpw6[3]);  // ../RTL/cortexm0ds_logic.v(6002)
  not u5169 (Gehiu6, n1239);  // ../RTL/cortexm0ds_logic.v(6002)
  buf u517 (K7hpw6[5], Xr9ax6);  // ../RTL/cortexm0ds_logic.v(2366)
  and u5170 (n1240, Uehiu6, Bfhiu6);  // ../RTL/cortexm0ds_logic.v(6003)
  not u5171 (Uhthu6, n1240);  // ../RTL/cortexm0ds_logic.v(6003)
  and u5172 (Bfhiu6, Ifhiu6, Pfhiu6);  // ../RTL/cortexm0ds_logic.v(6004)
  and u5173 (n1241, HRDATA[2], Pp7iu6);  // ../RTL/cortexm0ds_logic.v(6005)
  not u5174 (Pfhiu6, n1241);  // ../RTL/cortexm0ds_logic.v(6005)
  and u5175 (Ifhiu6, Wfhiu6, Dghiu6);  // ../RTL/cortexm0ds_logic.v(6006)
  and u5176 (n1242, Hrfpw6[2], Uy4iu6);  // ../RTL/cortexm0ds_logic.v(6007)
  not u5177 (Dghiu6, n1242);  // ../RTL/cortexm0ds_logic.v(6007)
  and u5178 (n1243, HRDATA[18], Kq7iu6);  // ../RTL/cortexm0ds_logic.v(6008)
  not u5179 (Wfhiu6, n1243);  // ../RTL/cortexm0ds_logic.v(6008)
  buf u518 (K7hpw6[13], Oi9ax6);  // ../RTL/cortexm0ds_logic.v(2366)
  and u5180 (Uehiu6, Kghiu6, Rghiu6);  // ../RTL/cortexm0ds_logic.v(6009)
  and u5181 (n1244, Fr7iu6, Ud4iu6);  // ../RTL/cortexm0ds_logic.v(6010)
  not u5182 (Rghiu6, n1244);  // ../RTL/cortexm0ds_logic.v(6010)
  and u5183 (Kghiu6, Yghiu6, Fhhiu6);  // ../RTL/cortexm0ds_logic.v(6011)
  and u5184 (n1245, Ppfpw6[2], A25iu6);  // ../RTL/cortexm0ds_logic.v(6012)
  not u5185 (Fhhiu6, n1245);  // ../RTL/cortexm0ds_logic.v(6012)
  and u5186 (n1246, R05iu6, D7fpw6[2]);  // ../RTL/cortexm0ds_logic.v(6013)
  not u5187 (Yghiu6, n1246);  // ../RTL/cortexm0ds_logic.v(6013)
  and u5188 (n1247, Mhhiu6, Thhiu6);  // ../RTL/cortexm0ds_logic.v(6014)
  not u5189 (Nhthu6, n1247);  // ../RTL/cortexm0ds_logic.v(6014)
  buf u519 (N2ghu6, Daiax6);  // ../RTL/cortexm0ds_logic.v(2409)
  and u5190 (Thhiu6, Aihiu6, Hihiu6);  // ../RTL/cortexm0ds_logic.v(6015)
  and u5191 (n1248, HRDATA[1], Pp7iu6);  // ../RTL/cortexm0ds_logic.v(6016)
  not u5192 (Hihiu6, n1248);  // ../RTL/cortexm0ds_logic.v(6016)
  and u5193 (Pp7iu6, Go7iu6, M15iu6);  // ../RTL/cortexm0ds_logic.v(6017)
  and u5194 (M15iu6, Oihiu6, Vihiu6);  // ../RTL/cortexm0ds_logic.v(6018)
  and u5195 (Oihiu6, Dxfhu6, Cjhiu6);  // ../RTL/cortexm0ds_logic.v(6019)
  and u5196 (Nlhiu6, vis_pc_o[0], Jjhiu6);  // ../RTL/cortexm0ds_logic.v(6020)
  not u5197 (Cjhiu6, Nlhiu6);  // ../RTL/cortexm0ds_logic.v(6020)
  and u5198 (Aihiu6, Qjhiu6, Xjhiu6);  // ../RTL/cortexm0ds_logic.v(6022)
  and u5199 (n1249, Hrfpw6[1], Uy4iu6);  // ../RTL/cortexm0ds_logic.v(6023)
  buf u52 (vis_r12_o[22], Tbfbx6);  // ../RTL/cortexm0ds_logic.v(2599)
  buf u520 (Fvdhu6, Bciax6);  // ../RTL/cortexm0ds_logic.v(2410)
  not u5200 (Xjhiu6, n1249);  // ../RTL/cortexm0ds_logic.v(6023)
  and u5201 (Uy4iu6, Ekhiu6, Vihiu6);  // ../RTL/cortexm0ds_logic.v(6024)
  or u5202 (n1250, Lkhiu6, Dxfhu6);  // ../RTL/cortexm0ds_logic.v(6025)
  not u5203 (Ekhiu6, n1250);  // ../RTL/cortexm0ds_logic.v(6025)
  and u5204 (Lkhiu6, Pkciu6, Skhiu6);  // ../RTL/cortexm0ds_logic.v(6026)
  or u5205 (Skhiu6, Zkhiu6, Ntfhu6);  // ../RTL/cortexm0ds_logic.v(6027)
  and u5206 (n1251, HRDATA[17], Kq7iu6);  // ../RTL/cortexm0ds_logic.v(6028)
  not u5207 (Qjhiu6, n1251);  // ../RTL/cortexm0ds_logic.v(6028)
  and u5208 (Kq7iu6, Glhiu6, Pz4iu6);  // ../RTL/cortexm0ds_logic.v(6029)
  and u5209 (Pz4iu6, Nlhiu6, Vihiu6);  // ../RTL/cortexm0ds_logic.v(6030)
  buf u521 (T6ehu6, Zdiax6);  // ../RTL/cortexm0ds_logic.v(2411)
  buf u5210 (Mpehu6, Ozkbx6[24]);  // ../RTL/cortexm0ds_logic.v(3176)
  and u5211 (Mhhiu6, Ulhiu6, Bmhiu6);  // ../RTL/cortexm0ds_logic.v(6032)
  or u5212 (Bmhiu6, Iz4iu6, A34iu6);  // ../RTL/cortexm0ds_logic.v(6033)
  and u5213 (Ulhiu6, Imhiu6, Pmhiu6);  // ../RTL/cortexm0ds_logic.v(6034)
  and u5214 (n1252, Ppfpw6[1], A25iu6);  // ../RTL/cortexm0ds_logic.v(6035)
  not u5215 (Pmhiu6, n1252);  // ../RTL/cortexm0ds_logic.v(6035)
  and u5216 (A25iu6, Ntfhu6, Vihiu6);  // ../RTL/cortexm0ds_logic.v(6036)
  or u5217 (n1253, Wofiu6, R05iu6);  // ../RTL/cortexm0ds_logic.v(6037)
  not u5218 (Vihiu6, n1253);  // ../RTL/cortexm0ds_logic.v(6037)
  and u5219 (n1254, R05iu6, D7fpw6[1]);  // ../RTL/cortexm0ds_logic.v(6038)
  buf u522 (vis_primask_o, Xfiax6);  // ../RTL/cortexm0ds_logic.v(2412)
  not u5220 (Imhiu6, n1254);  // ../RTL/cortexm0ds_logic.v(6038)
  and u5221 (R05iu6, Wmhiu6, Iz4iu6);  // ../RTL/cortexm0ds_logic.v(6039)
  not u5222 (Iz4iu6, Fr7iu6);  // ../RTL/cortexm0ds_logic.v(6040)
  and u5223 (Fr7iu6, Dnhiu6, Knhiu6);  // ../RTL/cortexm0ds_logic.v(6041)
  and u5224 (Knhiu6, Rnhiu6, Ynhiu6);  // ../RTL/cortexm0ds_logic.v(6042)
  or u5225 (n1255, Jkgiu6, Jfgpw6[4]);  // ../RTL/cortexm0ds_logic.v(6043)
  not u5226 (Rnhiu6, n1255);  // ../RTL/cortexm0ds_logic.v(6043)
  not u5227 (Jkgiu6, Npdhu6);  // ../RTL/cortexm0ds_logic.v(6044)
  and u5228 (Dnhiu6, HALTED, Rzciu6);  // ../RTL/cortexm0ds_logic.v(6045)
  and u5229 (n1256, Fohiu6, Mohiu6);  // ../RTL/cortexm0ds_logic.v(6046)
  buf u523 (Gqgpw6[20], Tsdbx6);  // ../RTL/cortexm0ds_logic.v(2377)
  not u5230 (Wmhiu6, n1256);  // ../RTL/cortexm0ds_logic.v(6046)
  and u5231 (Mohiu6, Tohiu6, Aphiu6);  // ../RTL/cortexm0ds_logic.v(6047)
  and u5232 (Tohiu6, Hphiu6, Ophiu6);  // ../RTL/cortexm0ds_logic.v(6048)
  and u5233 (n1257, Vphiu6, Cqhiu6);  // ../RTL/cortexm0ds_logic.v(6049)
  not u5234 (Hphiu6, n1257);  // ../RTL/cortexm0ds_logic.v(6049)
  or u5235 (Cqhiu6, Jqhiu6, Qqhiu6);  // ../RTL/cortexm0ds_logic.v(6050)
  and u5236 (n1258, Pkciu6, Juzhu6);  // ../RTL/cortexm0ds_logic.v(6051)
  not u5237 (Jqhiu6, n1258);  // ../RTL/cortexm0ds_logic.v(6051)
  or u5238 (Vphiu6, Eh6iu6, Jjhiu6);  // ../RTL/cortexm0ds_logic.v(6052)
  and u5239 (Fohiu6, Xqhiu6, Erhiu6);  // ../RTL/cortexm0ds_logic.v(6053)
  buf u524 (vis_r1_o[6], A2spw6);  // ../RTL/cortexm0ds_logic.v(1876)
  and u5240 (Xqhiu6, Lrhiu6, Srhiu6);  // ../RTL/cortexm0ds_logic.v(6054)
  and u5241 (n1259, Zrhiu6, Gshiu6);  // ../RTL/cortexm0ds_logic.v(6055)
  not u5242 (Ghthu6, n1259);  // ../RTL/cortexm0ds_logic.v(6055)
  and u5243 (n1260, Nshiu6, R6hhu6);  // ../RTL/cortexm0ds_logic.v(6056)
  not u5244 (Gshiu6, n1260);  // ../RTL/cortexm0ds_logic.v(6056)
  and u5245 (Nshiu6, Xbbiu6, Jbbiu6);  // ../RTL/cortexm0ds_logic.v(6057)
  not u5246 (Jbbiu6, Mu4iu6);  // ../RTL/cortexm0ds_logic.v(6058)
  and u5247 (Mu4iu6, Ushiu6, Bthiu6);  // ../RTL/cortexm0ds_logic.v(6059)
  and u5248 (Bthiu6, Ithiu6, Pthiu6);  // ../RTL/cortexm0ds_logic.v(6060)
  or u5249 (n1261, Cyfpw6[7], H4ghu6);  // ../RTL/cortexm0ds_logic.v(6061)
  buf u525 (vis_r1_o[10], Hmxpw6);  // ../RTL/cortexm0ds_logic.v(1876)
  not u5250 (Ithiu6, n1261);  // ../RTL/cortexm0ds_logic.v(6061)
  or u5251 (n1262, Wthiu6, Qjaiu6);  // ../RTL/cortexm0ds_logic.v(6062)
  not u5252 (Ushiu6, n1262);  // ../RTL/cortexm0ds_logic.v(6062)
  or u5253 (Xbbiu6, Duhiu6, A2nhu6);  // ../RTL/cortexm0ds_logic.v(6063)
  and u5254 (Zgthu6, Kuhiu6, Ruhiu6);  // ../RTL/cortexm0ds_logic.v(6064)
  and u5255 (Ruhiu6, Yuhiu6, Fvhiu6);  // ../RTL/cortexm0ds_logic.v(6065)
  and u5256 (n1263, Atdpw6, Mvhiu6);  // ../RTL/cortexm0ds_logic.v(6066)
  not u5257 (Yuhiu6, n1263);  // ../RTL/cortexm0ds_logic.v(6066)
  and u5258 (Kuhiu6, IRQ[16], Tvhiu6);  // ../RTL/cortexm0ds_logic.v(6067)
  and u5259 (n1264, Tk7iu6, Awhiu6);  // ../RTL/cortexm0ds_logic.v(6068)
  buf u526 (vis_r1_o[8], Sw0qw6);  // ../RTL/cortexm0ds_logic.v(1876)
  not u5260 (Tvhiu6, n1264);  // ../RTL/cortexm0ds_logic.v(6068)
  or u5261 (Awhiu6, Hwhiu6, Qg6iu6);  // ../RTL/cortexm0ds_logic.v(6069)
  and u5262 (Sgthu6, Owhiu6, Vwhiu6);  // ../RTL/cortexm0ds_logic.v(6070)
  and u5263 (Vwhiu6, Cxhiu6, Jxhiu6);  // ../RTL/cortexm0ds_logic.v(6071)
  and u5264 (n1265, Zvdpw6, Qxhiu6);  // ../RTL/cortexm0ds_logic.v(6072)
  not u5265 (Cxhiu6, n1265);  // ../RTL/cortexm0ds_logic.v(6072)
  and u5266 (Owhiu6, IRQ[30], Xxhiu6);  // ../RTL/cortexm0ds_logic.v(6073)
  and u5267 (n1266, Tk7iu6, Eyhiu6);  // ../RTL/cortexm0ds_logic.v(6074)
  not u5268 (Xxhiu6, n1266);  // ../RTL/cortexm0ds_logic.v(6074)
  or u5269 (Eyhiu6, Lyhiu6, Qg6iu6);  // ../RTL/cortexm0ds_logic.v(6075)
  not u527 (Lvdpw6, Woiax6);  // ../RTL/cortexm0ds_logic.v(2417)
  and u5270 (n1267, Uc5iu6, Fjfiu6);  // ../RTL/cortexm0ds_logic.v(6077)
  not u5271 (Tk7iu6, n1267);  // ../RTL/cortexm0ds_logic.v(6077)
  and u5272 (Qg6iu6, Syhiu6, Zyhiu6);  // ../RTL/cortexm0ds_logic.v(6078)
  not u5273 (Fjfiu6, Qg6iu6);  // ../RTL/cortexm0ds_logic.v(6078)
  and u5274 (Zyhiu6, Gzhiu6, Nzhiu6);  // ../RTL/cortexm0ds_logic.v(6079)
  or u5275 (n1268, Ur4iu6, Gc5iu6);  // ../RTL/cortexm0ds_logic.v(6080)
  not u5276 (Gzhiu6, n1268);  // ../RTL/cortexm0ds_logic.v(6080)
  and u5277 (Syhiu6, I4eiu6, Uzhiu6);  // ../RTL/cortexm0ds_logic.v(6081)
  and u5278 (n1269, B0iiu6, I0iiu6);  // ../RTL/cortexm0ds_logic.v(6082)
  not u5279 (Lgthu6, n1269);  // ../RTL/cortexm0ds_logic.v(6082)
  buf u528 (K7hpw6[12], Lk9ax6);  // ../RTL/cortexm0ds_logic.v(2366)
  and u5280 (I0iiu6, P0iiu6, W0iiu6);  // ../RTL/cortexm0ds_logic.v(6083)
  and u5281 (n1270, vis_pc_o[3], Ok8iu6);  // ../RTL/cortexm0ds_logic.v(6084)
  not u5282 (W0iiu6, n1270);  // ../RTL/cortexm0ds_logic.v(6084)
  and u5283 (P0iiu6, D1iiu6, K1iiu6);  // ../RTL/cortexm0ds_logic.v(6085)
  and u5284 (n1271, Jl8iu6, Tugpw6[2]);  // ../RTL/cortexm0ds_logic.v(6086)
  not u5285 (K1iiu6, n1271);  // ../RTL/cortexm0ds_logic.v(6086)
  buf u5286 (vis_r7_o[14], Lrwax6);  // ../RTL/cortexm0ds_logic.v(2654)
  buf u5287 (vis_r7_o[26], M5wax6);  // ../RTL/cortexm0ds_logic.v(2654)
  and u5288 (n1273, N5fpw6[3], Sdaiu6);  // ../RTL/cortexm0ds_logic.v(6088)
  not u5289 (Y1iiu6, n1273);  // ../RTL/cortexm0ds_logic.v(6088)
  buf u529 (K7hpw6[11], Xv8bx6);  // ../RTL/cortexm0ds_logic.v(2366)
  and u5290 (R1iiu6, F2iiu6, M2iiu6);  // ../RTL/cortexm0ds_logic.v(6089)
  or u5291 (M2iiu6, T2iiu6, Eg0iu6);  // ../RTL/cortexm0ds_logic.v(6090)
  and u5292 (n1274, Eafpw6[4], A3iiu6);  // ../RTL/cortexm0ds_logic.v(6091)
  not u5293 (F2iiu6, n1274);  // ../RTL/cortexm0ds_logic.v(6091)
  and u5294 (n1275, Ql8iu6, vis_ipsr_o[4]);  // ../RTL/cortexm0ds_logic.v(6092)
  not u5295 (D1iiu6, n1275);  // ../RTL/cortexm0ds_logic.v(6092)
  and u5296 (B0iiu6, H3iiu6, O3iiu6);  // ../RTL/cortexm0ds_logic.v(6093)
  or u5297 (O3iiu6, Lm8iu6, V3iiu6);  // ../RTL/cortexm0ds_logic.v(6094)
  and u5298 (n1276, Zm8iu6, H34iu6);  // ../RTL/cortexm0ds_logic.v(6095)
  not u5299 (H3iiu6, n1276);  // ../RTL/cortexm0ds_logic.v(6095)
  not u53 (Tugpw6[12], n1272[11]);  // ../RTL/cortexm0ds_logic.v(16030)
  buf u530 (K7hpw6[10], Im9ax6);  // ../RTL/cortexm0ds_logic.v(2366)
  and u5300 (n1277, C4iiu6, J4iiu6);  // ../RTL/cortexm0ds_logic.v(6096)
  not u5301 (Egthu6, n1277);  // ../RTL/cortexm0ds_logic.v(6096)
  and u5302 (J4iiu6, Q4iiu6, X4iiu6);  // ../RTL/cortexm0ds_logic.v(6097)
  and u5303 (n1278, Ok8iu6, vis_pc_o[1]);  // ../RTL/cortexm0ds_logic.v(6098)
  not u5304 (X4iiu6, n1278);  // ../RTL/cortexm0ds_logic.v(6098)
  and u5305 (Q4iiu6, E5iiu6, L5iiu6);  // ../RTL/cortexm0ds_logic.v(6099)
  and u5306 (n1279, Jl8iu6, Tugpw6[0]);  // ../RTL/cortexm0ds_logic.v(6100)
  not u5307 (L5iiu6, n1279);  // ../RTL/cortexm0ds_logic.v(6100)
  buf u5308 (vis_r7_o[16], Lpwax6);  // ../RTL/cortexm0ds_logic.v(2654)
  buf u5309 (vis_r7_o[28], Rnibx6);  // ../RTL/cortexm0ds_logic.v(2654)
  buf u531 (K7hpw6[9], N3jbx6);  // ../RTL/cortexm0ds_logic.v(2366)
  and u5310 (n1280, Eafpw6[2], A3iiu6);  // ../RTL/cortexm0ds_logic.v(6102)
  not u5311 (Z5iiu6, n1280);  // ../RTL/cortexm0ds_logic.v(6102)
  and u5312 (S5iiu6, G6iiu6, N6iiu6);  // ../RTL/cortexm0ds_logic.v(6103)
  and u5313 (n1281, Sdaiu6, U6iiu6);  // ../RTL/cortexm0ds_logic.v(6104)
  not u5314 (N6iiu6, n1281);  // ../RTL/cortexm0ds_logic.v(6104)
  xor u5315 (U6iiu6, Vtzhu6, Cuzhu6);  // ../RTL/cortexm0ds_logic.v(6105)
  xor u5316 (Cuzhu6, Juzhu6, Quzhu6);  // ../RTL/cortexm0ds_logic.v(6106)
  and u5317 (n1282, B7iiu6, Gh0iu6);  // ../RTL/cortexm0ds_logic.v(6107)
  not u5318 (G6iiu6, n1282);  // ../RTL/cortexm0ds_logic.v(6107)
  and u5319 (n1283, Ql8iu6, vis_ipsr_o[2]);  // ../RTL/cortexm0ds_logic.v(6108)
  buf u532 (K7hpw6[8], Fo9ax6);  // ../RTL/cortexm0ds_logic.v(2366)
  not u5320 (E5iiu6, n1283);  // ../RTL/cortexm0ds_logic.v(6108)
  and u5321 (C4iiu6, I7iiu6, P7iiu6);  // ../RTL/cortexm0ds_logic.v(6109)
  and u5322 (n1284, W29iu6, Fkfpw6[2]);  // ../RTL/cortexm0ds_logic.v(6110)
  not u5323 (P7iiu6, n1284);  // ../RTL/cortexm0ds_logic.v(6110)
  and u5324 (n1285, Zm8iu6, Ud4iu6);  // ../RTL/cortexm0ds_logic.v(6111)
  not u5325 (I7iiu6, n1285);  // ../RTL/cortexm0ds_logic.v(6111)
  AL_MUX u5326 (
    .i0(S8fpw6[8]),
    .i1(W7iiu6),
    .sel(D8iiu6),
    .o(Xfthu6));  // ../RTL/cortexm0ds_logic.v(6112)
  and u5327 (n1286, K8iiu6, R8iiu6);  // ../RTL/cortexm0ds_logic.v(6113)
  not u5328 (W7iiu6, n1286);  // ../RTL/cortexm0ds_logic.v(6113)
  and u5329 (R8iiu6, Y8iiu6, F9iiu6);  // ../RTL/cortexm0ds_logic.v(6114)
  buf u533 (K7hpw6[7], Bq9ax6);  // ../RTL/cortexm0ds_logic.v(2366)
  and u5330 (n1287, D7fpw6[0], M9iiu6);  // ../RTL/cortexm0ds_logic.v(6115)
  not u5331 (F9iiu6, n1287);  // ../RTL/cortexm0ds_logic.v(6115)
  and u5332 (n1288, D7fpw6[8], T9iiu6);  // ../RTL/cortexm0ds_logic.v(6116)
  not u5333 (Y8iiu6, n1288);  // ../RTL/cortexm0ds_logic.v(6116)
  and u5334 (K8iiu6, Aaiiu6, Haiiu6);  // ../RTL/cortexm0ds_logic.v(6117)
  or u5335 (Haiiu6, Oaiiu6, O95iu6);  // ../RTL/cortexm0ds_logic.v(6118)
  and u5336 (n1289, Vaiiu6, Cbiiu6);  // ../RTL/cortexm0ds_logic.v(6119)
  not u5337 (Qfthu6, n1289);  // ../RTL/cortexm0ds_logic.v(6119)
  and u5338 (n1290, Jbiiu6, Qbiiu6);  // ../RTL/cortexm0ds_logic.v(6120)
  not u5339 (Cbiiu6, n1290);  // ../RTL/cortexm0ds_logic.v(6120)
  buf u534 (K7hpw6[6], Tc9bx6);  // ../RTL/cortexm0ds_logic.v(2366)
  AL_MUX u5340 (
    .i0(P65iu6),
    .i1(Xbiiu6),
    .sel(D8iiu6),
    .o(Vaiiu6));  // ../RTL/cortexm0ds_logic.v(6121)
  and u5341 (Xbiiu6, Eciiu6, Lciiu6);  // ../RTL/cortexm0ds_logic.v(6122)
  and u5342 (Lciiu6, Sciiu6, Zciiu6);  // ../RTL/cortexm0ds_logic.v(6123)
  and u5343 (n1291, D7fpw6[1], M9iiu6);  // ../RTL/cortexm0ds_logic.v(6124)
  not u5344 (Zciiu6, n1291);  // ../RTL/cortexm0ds_logic.v(6124)
  and u5345 (n1292, D7fpw6[9], T9iiu6);  // ../RTL/cortexm0ds_logic.v(6125)
  not u5346 (Sciiu6, n1292);  // ../RTL/cortexm0ds_logic.v(6125)
  and u5347 (Eciiu6, Aaiiu6, Gdiiu6);  // ../RTL/cortexm0ds_logic.v(6126)
  or u5348 (Gdiiu6, Oaiiu6, Ndiiu6);  // ../RTL/cortexm0ds_logic.v(6127)
  and u5349 (n1293, Udiiu6, Beiiu6);  // ../RTL/cortexm0ds_logic.v(6128)
  buf u535 (vis_r2_o[24], Veqax6);  // ../RTL/cortexm0ds_logic.v(2551)
  not u5350 (Jfthu6, n1293);  // ../RTL/cortexm0ds_logic.v(6128)
  and u5351 (n1294, S8fpw6[10], Ieiiu6);  // ../RTL/cortexm0ds_logic.v(6129)
  not u5352 (Beiiu6, n1294);  // ../RTL/cortexm0ds_logic.v(6129)
  and u5353 (n1295, D8iiu6, Peiiu6);  // ../RTL/cortexm0ds_logic.v(6130)
  not u5354 (Ieiiu6, n1295);  // ../RTL/cortexm0ds_logic.v(6130)
  and u5355 (n1296, Jbiiu6, Weiiu6);  // ../RTL/cortexm0ds_logic.v(6131)
  not u5356 (Peiiu6, n1296);  // ../RTL/cortexm0ds_logic.v(6131)
  or u5357 (Ooiiu6, Dfiiu6, Kfiiu6);  // ../RTL/cortexm0ds_logic.v(6132)
  not u5358 (Jbiiu6, Ooiiu6);  // ../RTL/cortexm0ds_logic.v(6132)
  and u5359 (n1297, D8iiu6, Rfiiu6);  // ../RTL/cortexm0ds_logic.v(6133)
  buf u536 (vis_r2_o[8], Tcrax6);  // ../RTL/cortexm0ds_logic.v(2551)
  not u5360 (Udiiu6, n1297);  // ../RTL/cortexm0ds_logic.v(6133)
  and u5361 (n1298, Yfiiu6, Fgiiu6);  // ../RTL/cortexm0ds_logic.v(6134)
  not u5362 (Rfiiu6, n1298);  // ../RTL/cortexm0ds_logic.v(6134)
  and u5363 (Fgiiu6, Mgiiu6, Tgiiu6);  // ../RTL/cortexm0ds_logic.v(6135)
  and u5364 (n1299, D7fpw6[2], M9iiu6);  // ../RTL/cortexm0ds_logic.v(6136)
  not u5365 (Tgiiu6, n1299);  // ../RTL/cortexm0ds_logic.v(6136)
  and u5366 (n1300, Ahiiu6, Hhiiu6);  // ../RTL/cortexm0ds_logic.v(6137)
  not u5367 (M9iiu6, n1300);  // ../RTL/cortexm0ds_logic.v(6137)
  and u5368 (Hhiiu6, Ohiiu6, Vhiiu6);  // ../RTL/cortexm0ds_logic.v(6138)
  and u5369 (n1301, Ciiiu6, Jiiiu6);  // ../RTL/cortexm0ds_logic.v(6139)
  buf u537 (Dxfhu6, U8jax6);  // ../RTL/cortexm0ds_logic.v(2427)
  not u5370 (Ohiiu6, n1301);  // ../RTL/cortexm0ds_logic.v(6139)
  and u5371 (Ciiiu6, Qiiiu6, Zraiu6);  // ../RTL/cortexm0ds_logic.v(6140)
  or u5372 (Qiiiu6, Xiiiu6, Ejiiu6);  // ../RTL/cortexm0ds_logic.v(6141)
  and u5373 (Ahiiu6, Ljiiu6, Sjiiu6);  // ../RTL/cortexm0ds_logic.v(6142)
  or u5374 (Sjiiu6, Zjiiu6, Gkiiu6);  // ../RTL/cortexm0ds_logic.v(6143)
  and u5375 (n1302, D7fpw6[10], T9iiu6);  // ../RTL/cortexm0ds_logic.v(6144)
  not u5376 (Mgiiu6, n1302);  // ../RTL/cortexm0ds_logic.v(6144)
  and u5377 (n1303, Nkiiu6, Ukiiu6);  // ../RTL/cortexm0ds_logic.v(6145)
  not u5378 (T9iiu6, n1303);  // ../RTL/cortexm0ds_logic.v(6145)
  and u5379 (Ukiiu6, Bliiu6, Iliiu6);  // ../RTL/cortexm0ds_logic.v(6146)
  buf u538 (Iwfpw6[0], S4kbx6);  // ../RTL/cortexm0ds_logic.v(2830)
  and u5380 (n1304, Pliiu6, Wliiu6);  // ../RTL/cortexm0ds_logic.v(6147)
  not u5381 (Iliiu6, n1304);  // ../RTL/cortexm0ds_logic.v(6147)
  and u5382 (Pliiu6, Dmiiu6, Zraiu6);  // ../RTL/cortexm0ds_logic.v(6148)
  or u5383 (n1305, Kmiiu6, Rmiiu6);  // ../RTL/cortexm0ds_logic.v(6149)
  not u5384 (Bliiu6, n1305);  // ../RTL/cortexm0ds_logic.v(6149)
  and u5385 (Nkiiu6, Ymiiu6, Fniiu6);  // ../RTL/cortexm0ds_logic.v(6150)
  and u5386 (Yfiiu6, Aaiiu6, Mniiu6);  // ../RTL/cortexm0ds_logic.v(6151)
  or u5387 (Mniiu6, Oaiiu6, Tniiu6);  // ../RTL/cortexm0ds_logic.v(6152)
  or u5388 (Cfthu6, Aoiiu6, Hoiiu6);  // ../RTL/cortexm0ds_logic.v(6153)
  or u5389 (n1306, Ooiiu6, Voiiu6);  // ../RTL/cortexm0ds_logic.v(6154)
  buf u539 (K7hpw6[3], Pv9ax6);  // ../RTL/cortexm0ds_logic.v(2366)
  not u5390 (Hoiiu6, n1306);  // ../RTL/cortexm0ds_logic.v(6154)
  buf u5391 (Arehu6, Ozkbx6[23]);  // ../RTL/cortexm0ds_logic.v(3176)
  or u5392 (n1307, Y7ghu6, U98iu6);  // ../RTL/cortexm0ds_logic.v(6156)
  not u5393 (Dfiiu6, n1307);  // ../RTL/cortexm0ds_logic.v(6156)
  AL_MUX u5394 (
    .i0(S8fpw6[11]),
    .i1(Cpiiu6),
    .sel(D8iiu6),
    .o(Aoiiu6));  // ../RTL/cortexm0ds_logic.v(6157)
  and u5395 (D8iiu6, HREADY, Jpiiu6);  // ../RTL/cortexm0ds_logic.v(6158)
  and u5396 (n1308, Qpiiu6, Xpiiu6);  // ../RTL/cortexm0ds_logic.v(6159)
  not u5397 (Jpiiu6, n1308);  // ../RTL/cortexm0ds_logic.v(6159)
  and u5398 (Xpiiu6, Eqiiu6, Lqiiu6);  // ../RTL/cortexm0ds_logic.v(6160)
  and u5399 (Lqiiu6, Sqiiu6, Zqiiu6);  // ../RTL/cortexm0ds_logic.v(6161)
  buf u54 (Jshpw6[23], H7hbx6);  // ../RTL/cortexm0ds_logic.v(2372)
  buf u540 (E1hpw6[17], Nlbbx6);  // ../RTL/cortexm0ds_logic.v(2367)
  and u5400 (n1309, Griiu6, Nriiu6);  // ../RTL/cortexm0ds_logic.v(6162)
  not u5401 (Zqiiu6, n1309);  // ../RTL/cortexm0ds_logic.v(6162)
  or u5402 (n1310, Uriiu6, Y7ghu6);  // ../RTL/cortexm0ds_logic.v(6163)
  not u5403 (Griiu6, n1310);  // ../RTL/cortexm0ds_logic.v(6163)
  and u5404 (Sqiiu6, Bsiiu6, Isiiu6);  // ../RTL/cortexm0ds_logic.v(6164)
  and u5405 (n1311, Psiiu6, Ae0iu6);  // ../RTL/cortexm0ds_logic.v(6165)
  not u5406 (Bsiiu6, n1311);  // ../RTL/cortexm0ds_logic.v(6165)
  or u5407 (n1312, Mjfiu6, H4ghu6);  // ../RTL/cortexm0ds_logic.v(6166)
  not u5408 (Psiiu6, n1312);  // ../RTL/cortexm0ds_logic.v(6166)
  and u5409 (Eqiiu6, Wsiiu6, Dtiiu6);  // ../RTL/cortexm0ds_logic.v(6167)
  buf u541 (E1hpw6[19], Q8aax6);  // ../RTL/cortexm0ds_logic.v(2367)
  and u5410 (n1313, Ktiiu6, Ndiiu6);  // ../RTL/cortexm0ds_logic.v(6168)
  not u5411 (Dtiiu6, n1313);  // ../RTL/cortexm0ds_logic.v(6168)
  and u5412 (n1314, Rtiiu6, Ytiiu6);  // ../RTL/cortexm0ds_logic.v(6169)
  not u5413 (Ktiiu6, n1314);  // ../RTL/cortexm0ds_logic.v(6169)
  and u5414 (n1315, D7fpw6[10], Fuiiu6);  // ../RTL/cortexm0ds_logic.v(6170)
  not u5415 (Ytiiu6, n1315);  // ../RTL/cortexm0ds_logic.v(6170)
  and u5416 (n1316, Muiiu6, Tuiiu6);  // ../RTL/cortexm0ds_logic.v(6171)
  not u5417 (Fuiiu6, n1316);  // ../RTL/cortexm0ds_logic.v(6171)
  and u5418 (n1317, Aviiu6, Hviiu6);  // ../RTL/cortexm0ds_logic.v(6172)
  not u5419 (Tuiiu6, n1317);  // ../RTL/cortexm0ds_logic.v(6172)
  buf u542 (E1hpw6[20], Cndbx6);  // ../RTL/cortexm0ds_logic.v(2367)
  or u5420 (n1318, Oviiu6, Zwciu6);  // ../RTL/cortexm0ds_logic.v(6173)
  not u5421 (Aviiu6, n1318);  // ../RTL/cortexm0ds_logic.v(6173)
  and u5422 (n1319, Vviiu6, Cwiiu6);  // ../RTL/cortexm0ds_logic.v(6174)
  not u5423 (Muiiu6, n1319);  // ../RTL/cortexm0ds_logic.v(6174)
  and u5424 (n1320, Vviiu6, Jwiiu6);  // ../RTL/cortexm0ds_logic.v(6175)
  not u5425 (Rtiiu6, n1320);  // ../RTL/cortexm0ds_logic.v(6175)
  and u5426 (Wsiiu6, Qwiiu6, Xwiiu6);  // ../RTL/cortexm0ds_logic.v(6176)
  and u5427 (n1321, D7fpw6[14], Exiiu6);  // ../RTL/cortexm0ds_logic.v(6177)
  not u5428 (Xwiiu6, n1321);  // ../RTL/cortexm0ds_logic.v(6177)
  and u5429 (n1322, Lxiiu6, Sxiiu6);  // ../RTL/cortexm0ds_logic.v(6178)
  buf u543 (vis_r2_o[18], Uwqax6);  // ../RTL/cortexm0ds_logic.v(2551)
  not u5430 (Exiiu6, n1322);  // ../RTL/cortexm0ds_logic.v(6178)
  and u5431 (n1323, Zxiiu6, C0ehu6);  // ../RTL/cortexm0ds_logic.v(6179)
  not u5432 (Sxiiu6, n1323);  // ../RTL/cortexm0ds_logic.v(6179)
  and u5433 (Zxiiu6, Gyiiu6, Q5aiu6);  // ../RTL/cortexm0ds_logic.v(6180)
  or u5434 (Gyiiu6, S1ehu6, Nyiiu6);  // ../RTL/cortexm0ds_logic.v(6181)
  and u5435 (n1324, Ejiiu6, Uyiiu6);  // ../RTL/cortexm0ds_logic.v(6182)
  not u5436 (Lxiiu6, n1324);  // ../RTL/cortexm0ds_logic.v(6182)
  and u5437 (n1325, Bziiu6, Uyiiu6);  // ../RTL/cortexm0ds_logic.v(6183)
  not u5438 (Qwiiu6, n1325);  // ../RTL/cortexm0ds_logic.v(6183)
  and u5439 (Qpiiu6, Iziiu6, Pziiu6);  // ../RTL/cortexm0ds_logic.v(6184)
  buf u544 (E1hpw6[21], J6ebx6);  // ../RTL/cortexm0ds_logic.v(2367)
  and u5440 (Pziiu6, Wziiu6, D0jiu6);  // ../RTL/cortexm0ds_logic.v(6185)
  and u5441 (Wziiu6, K0jiu6, R0jiu6);  // ../RTL/cortexm0ds_logic.v(6186)
  and u5442 (n1326, Y0jiu6, F1jiu6);  // ../RTL/cortexm0ds_logic.v(6187)
  not u5443 (R0jiu6, n1326);  // ../RTL/cortexm0ds_logic.v(6187)
  and u5444 (Iziiu6, M1jiu6, T1jiu6);  // ../RTL/cortexm0ds_logic.v(6188)
  and u5445 (n1327, A2jiu6, H2jiu6);  // ../RTL/cortexm0ds_logic.v(6189)
  not u5446 (Cpiiu6, n1327);  // ../RTL/cortexm0ds_logic.v(6189)
  and u5447 (H2jiu6, O2jiu6, V2jiu6);  // ../RTL/cortexm0ds_logic.v(6190)
  and u5448 (n1328, D7fpw6[11], C3jiu6);  // ../RTL/cortexm0ds_logic.v(6191)
  not u5449 (V2jiu6, n1328);  // ../RTL/cortexm0ds_logic.v(6191)
  buf u545 (vis_r2_o[19], Uuqax6);  // ../RTL/cortexm0ds_logic.v(2551)
  or u5450 (C3jiu6, Kmiiu6, J3jiu6);  // ../RTL/cortexm0ds_logic.v(6192)
  and u5451 (J3jiu6, Rmiiu6, D7fpw6[12]);  // ../RTL/cortexm0ds_logic.v(6193)
  and u5452 (Kmiiu6, Zraiu6, Q3jiu6);  // ../RTL/cortexm0ds_logic.v(6194)
  and u5453 (n1329, X3jiu6, E4jiu6);  // ../RTL/cortexm0ds_logic.v(6195)
  not u5454 (Q3jiu6, n1329);  // ../RTL/cortexm0ds_logic.v(6195)
  or u5455 (O2jiu6, V4aiu6, Ljiiu6);  // ../RTL/cortexm0ds_logic.v(6196)
  and u5456 (Ljiiu6, L4jiu6, S4jiu6);  // ../RTL/cortexm0ds_logic.v(6197)
  and u5457 (n1330, Z4jiu6, G5jiu6);  // ../RTL/cortexm0ds_logic.v(6198)
  not u5458 (L4jiu6, n1330);  // ../RTL/cortexm0ds_logic.v(6198)
  and u5459 (G5jiu6, N5jiu6, U5jiu6);  // ../RTL/cortexm0ds_logic.v(6199)
  buf u546 (E1hpw6[22], Qlfbx6);  // ../RTL/cortexm0ds_logic.v(2367)
  or u5460 (N5jiu6, Oviiu6, Tniiu6);  // ../RTL/cortexm0ds_logic.v(6200)
  and u5461 (A2jiu6, Aaiiu6, B6jiu6);  // ../RTL/cortexm0ds_logic.v(6201)
  or u5462 (B6jiu6, Oaiiu6, I6jiu6);  // ../RTL/cortexm0ds_logic.v(6202)
  and u5463 (Aaiiu6, P6jiu6, W6jiu6);  // ../RTL/cortexm0ds_logic.v(6203)
  and u5464 (P6jiu6, D7jiu6, Faaiu6);  // ../RTL/cortexm0ds_logic.v(6204)
  and u5465 (n1331, K7jiu6, R7jiu6);  // ../RTL/cortexm0ds_logic.v(6205)
  not u5466 (D7jiu6, n1331);  // ../RTL/cortexm0ds_logic.v(6205)
  and u5467 (K7jiu6, Ia8iu6, D7fpw6[7]);  // ../RTL/cortexm0ds_logic.v(6206)
  AL_MUX u5468 (
    .i0(Y7jiu6),
    .i1(S8fpw6[3]),
    .sel(F58iu6),
    .o(Vethu6));  // ../RTL/cortexm0ds_logic.v(6207)
  and u5469 (n1332, F8jiu6, M8jiu6);  // ../RTL/cortexm0ds_logic.v(6208)
  buf u547 (vis_r2_o[20], Usqax6);  // ../RTL/cortexm0ds_logic.v(2551)
  not u5470 (Y7jiu6, n1332);  // ../RTL/cortexm0ds_logic.v(6208)
  and u5471 (M8jiu6, T8jiu6, A9jiu6);  // ../RTL/cortexm0ds_logic.v(6209)
  and u5472 (A9jiu6, H9jiu6, O9jiu6);  // ../RTL/cortexm0ds_logic.v(6210)
  and u5473 (n1333, V9jiu6, Ce8iu6);  // ../RTL/cortexm0ds_logic.v(6211)
  not u5474 (O9jiu6, n1333);  // ../RTL/cortexm0ds_logic.v(6211)
  xor u5475 (n1334, Cajiu6, Jajiu6);  // ../RTL/cortexm0ds_logic.v(6212)
  not u5476 (V9jiu6, n1334);  // ../RTL/cortexm0ds_logic.v(6212)
  and u5477 (Jajiu6, Qajiu6, S8fpw6[2]);  // ../RTL/cortexm0ds_logic.v(6213)
  and u5478 (H9jiu6, Xajiu6, Faaiu6);  // ../RTL/cortexm0ds_logic.v(6214)
  and u5479 (n1335, Ebjiu6, E88iu6);  // ../RTL/cortexm0ds_logic.v(6215)
  buf u548 (E1hpw6[23], Wxgbx6);  // ../RTL/cortexm0ds_logic.v(2367)
  not u5480 (Xajiu6, n1335);  // ../RTL/cortexm0ds_logic.v(6215)
  and u5481 (n1336, Lbjiu6, Sbjiu6);  // ../RTL/cortexm0ds_logic.v(6216)
  not u5482 (Ebjiu6, n1336);  // ../RTL/cortexm0ds_logic.v(6216)
  and u5483 (n1337, Zbjiu6, Gcjiu6);  // ../RTL/cortexm0ds_logic.v(6217)
  not u5484 (Sbjiu6, n1337);  // ../RTL/cortexm0ds_logic.v(6217)
  and u5485 (n1338, Ncjiu6, Ucjiu6);  // ../RTL/cortexm0ds_logic.v(6218)
  not u5486 (Lbjiu6, n1338);  // ../RTL/cortexm0ds_logic.v(6218)
  and u5487 (T8jiu6, Bdjiu6, Idjiu6);  // ../RTL/cortexm0ds_logic.v(6219)
  and u5488 (n1339, Tc8iu6, Ppfpw6[3]);  // ../RTL/cortexm0ds_logic.v(6220)
  not u5489 (Idjiu6, n1339);  // ../RTL/cortexm0ds_logic.v(6220)
  buf u549 (vis_r2_o[21], Uqqax6);  // ../RTL/cortexm0ds_logic.v(2551)
  and u5490 (n1340, D7fpw6[9], Pdjiu6);  // ../RTL/cortexm0ds_logic.v(6221)
  not u5491 (Bdjiu6, n1340);  // ../RTL/cortexm0ds_logic.v(6221)
  and u5492 (F8jiu6, Wdjiu6, Dejiu6);  // ../RTL/cortexm0ds_logic.v(6222)
  and u5493 (Dejiu6, Kejiu6, Rejiu6);  // ../RTL/cortexm0ds_logic.v(6223)
  and u5494 (n1341, Habiu6, D7fpw6[2]);  // ../RTL/cortexm0ds_logic.v(6224)
  not u5495 (Rejiu6, n1341);  // ../RTL/cortexm0ds_logic.v(6224)
  or u5496 (Kejiu6, V4aiu6, Yb8iu6);  // ../RTL/cortexm0ds_logic.v(6225)
  and u5497 (Wdjiu6, Yejiu6, Ffjiu6);  // ../RTL/cortexm0ds_logic.v(6226)
  and u5498 (n1342, Cbbiu6, D7fpw6[8]);  // ../RTL/cortexm0ds_logic.v(6227)
  not u5499 (Ffjiu6, n1342);  // ../RTL/cortexm0ds_logic.v(6227)
  buf u55 (vis_r12_o[30], Kosax6);  // ../RTL/cortexm0ds_logic.v(2599)
  buf u550 (E1hpw6[24], T6aax6);  // ../RTL/cortexm0ds_logic.v(2367)
  and u5500 (n1343, Mfjiu6, Tfjiu6);  // ../RTL/cortexm0ds_logic.v(6228)
  not u5501 (Yejiu6, n1343);  // ../RTL/cortexm0ds_logic.v(6228)
  AL_MUX u5502 (
    .i0(Agjiu6),
    .i1(S8fpw6[2]),
    .sel(F58iu6),
    .o(Oethu6));  // ../RTL/cortexm0ds_logic.v(6229)
  and u5503 (n1344, HREADY, Hgjiu6);  // ../RTL/cortexm0ds_logic.v(6230)
  not u5504 (F58iu6, n1344);  // ../RTL/cortexm0ds_logic.v(6230)
  and u5505 (n1345, Ogjiu6, Vgjiu6);  // ../RTL/cortexm0ds_logic.v(6231)
  not u5506 (Hgjiu6, n1345);  // ../RTL/cortexm0ds_logic.v(6231)
  and u5507 (Vgjiu6, Chjiu6, Jhjiu6);  // ../RTL/cortexm0ds_logic.v(6232)
  and u5508 (Jhjiu6, Qhjiu6, Xhjiu6);  // ../RTL/cortexm0ds_logic.v(6233)
  and u5509 (n1346, Eijiu6, Lijiu6);  // ../RTL/cortexm0ds_logic.v(6234)
  buf u551 (vis_r2_o[22], Trebx6);  // ../RTL/cortexm0ds_logic.v(2551)
  not u5510 (Xhjiu6, n1346);  // ../RTL/cortexm0ds_logic.v(6234)
  or u5511 (n1347, Sijiu6, Cyfpw6[0]);  // ../RTL/cortexm0ds_logic.v(6235)
  not u5512 (Eijiu6, n1347);  // ../RTL/cortexm0ds_logic.v(6235)
  and u5513 (Qhjiu6, Zijiu6, Gjjiu6);  // ../RTL/cortexm0ds_logic.v(6236)
  and u5514 (n1348, Njjiu6, Ujjiu6);  // ../RTL/cortexm0ds_logic.v(6237)
  not u5515 (Zijiu6, n1348);  // ../RTL/cortexm0ds_logic.v(6237)
  or u5516 (n1349, Q5aiu6, Bkjiu6);  // ../RTL/cortexm0ds_logic.v(6238)
  not u5517 (Njjiu6, n1349);  // ../RTL/cortexm0ds_logic.v(6238)
  and u5518 (Chjiu6, Ikjiu6, Pkjiu6);  // ../RTL/cortexm0ds_logic.v(6239)
  and u5519 (n1350, Wkjiu6, D7fpw6[10]);  // ../RTL/cortexm0ds_logic.v(6240)
  buf u552 (E1hpw6[25], W4aax6);  // ../RTL/cortexm0ds_logic.v(2367)
  not u5520 (Pkjiu6, n1350);  // ../RTL/cortexm0ds_logic.v(6240)
  and u5521 (Ikjiu6, Dljiu6, Kljiu6);  // ../RTL/cortexm0ds_logic.v(6241)
  and u5522 (n1351, Rljiu6, Yljiu6);  // ../RTL/cortexm0ds_logic.v(6242)
  not u5523 (Kljiu6, n1351);  // ../RTL/cortexm0ds_logic.v(6242)
  or u5524 (Dljiu6, Fmjiu6, Mmjiu6);  // ../RTL/cortexm0ds_logic.v(6243)
  and u5525 (Ogjiu6, Tmjiu6, Anjiu6);  // ../RTL/cortexm0ds_logic.v(6244)
  and u5526 (Anjiu6, Hnjiu6, Onjiu6);  // ../RTL/cortexm0ds_logic.v(6245)
  and u5527 (Hnjiu6, Vnjiu6, Cojiu6);  // ../RTL/cortexm0ds_logic.v(6246)
  or u5528 (Cojiu6, Wmaiu6, Jojiu6);  // ../RTL/cortexm0ds_logic.v(6247)
  or u5529 (Vnjiu6, Qojiu6, Xojiu6);  // ../RTL/cortexm0ds_logic.v(6248)
  buf u553 (vis_r2_o[23], Azpax6);  // ../RTL/cortexm0ds_logic.v(2551)
  and u5530 (Tmjiu6, Epjiu6, Lpjiu6);  // ../RTL/cortexm0ds_logic.v(6249)
  and u5531 (n1352, Ae0iu6, Pthiu6);  // ../RTL/cortexm0ds_logic.v(6250)
  not u5532 (Lpjiu6, n1352);  // ../RTL/cortexm0ds_logic.v(6250)
  and u5533 (n1353, Spjiu6, Zpjiu6);  // ../RTL/cortexm0ds_logic.v(6251)
  not u5534 (Agjiu6, n1353);  // ../RTL/cortexm0ds_logic.v(6251)
  and u5535 (Zpjiu6, Gqjiu6, Nqjiu6);  // ../RTL/cortexm0ds_logic.v(6252)
  and u5536 (Nqjiu6, Uqjiu6, V68iu6);  // ../RTL/cortexm0ds_logic.v(6253)
  and u5537 (n1354, W8aiu6, Brjiu6);  // ../RTL/cortexm0ds_logic.v(6254)
  not u5538 (V68iu6, n1354);  // ../RTL/cortexm0ds_logic.v(6254)
  and u5539 (n1355, Irjiu6, Wthiu6);  // ../RTL/cortexm0ds_logic.v(6255)
  buf u554 (Sufpw6[0], L6lax6);  // ../RTL/cortexm0ds_logic.v(2404)
  not u5540 (Brjiu6, n1355);  // ../RTL/cortexm0ds_logic.v(6255)
  or u5541 (Irjiu6, Prjiu6, Cyfpw6[5]);  // ../RTL/cortexm0ds_logic.v(6256)
  and u5542 (n1356, Wrjiu6, E88iu6);  // ../RTL/cortexm0ds_logic.v(6257)
  not u5543 (Uqjiu6, n1356);  // ../RTL/cortexm0ds_logic.v(6257)
  and u5544 (n1357, Dsjiu6, Ksjiu6);  // ../RTL/cortexm0ds_logic.v(6258)
  not u5545 (E88iu6, n1357);  // ../RTL/cortexm0ds_logic.v(6258)
  and u5546 (n1358, Rsjiu6, Ysjiu6);  // ../RTL/cortexm0ds_logic.v(6259)
  not u5547 (Ksjiu6, n1358);  // ../RTL/cortexm0ds_logic.v(6259)
  or u5548 (n1359, Oviiu6, Ftjiu6);  // ../RTL/cortexm0ds_logic.v(6260)
  not u5549 (Ysjiu6, n1359);  // ../RTL/cortexm0ds_logic.v(6260)
  buf u555 (E1hpw6[26], Cccbx6);  // ../RTL/cortexm0ds_logic.v(2367)
  and u5550 (Rsjiu6, Ia8iu6, Mtjiu6);  // ../RTL/cortexm0ds_logic.v(6261)
  and u5551 (n1360, Ttjiu6, Aujiu6);  // ../RTL/cortexm0ds_logic.v(6262)
  not u5552 (Dsjiu6, n1360);  // ../RTL/cortexm0ds_logic.v(6262)
  or u5553 (Foiow6, Hujiu6, I6jiu6);  // ../RTL/cortexm0ds_logic.v(6263)
  not u5554 (Ttjiu6, Foiow6);  // ../RTL/cortexm0ds_logic.v(6263)
  xor u5555 (Wrjiu6, Gcjiu6, Zbjiu6);  // ../RTL/cortexm0ds_logic.v(6264)
  and u5556 (Zbjiu6, W7biu6, P7biu6);  // ../RTL/cortexm0ds_logic.v(6265)
  or u5557 (n1361, Oujiu6, Ncjiu6);  // ../RTL/cortexm0ds_logic.v(6266)
  not u5558 (P7biu6, n1361);  // ../RTL/cortexm0ds_logic.v(6266)
  and u5559 (Oujiu6, Vujiu6, Cvjiu6);  // ../RTL/cortexm0ds_logic.v(6267)
  buf u556 (E1hpw6[27], Fvcbx6);  // ../RTL/cortexm0ds_logic.v(2367)
  and u5560 (W7biu6, L88iu6, S88iu6);  // ../RTL/cortexm0ds_logic.v(6268)
  xor u5561 (S88iu6, Jvjiu6, O95iu6);  // ../RTL/cortexm0ds_logic.v(6269)
  xor u5562 (Gcjiu6, Ucjiu6, Ncjiu6);  // ../RTL/cortexm0ds_logic.v(6270)
  or u5563 (n1362, Cvjiu6, Vujiu6);  // ../RTL/cortexm0ds_logic.v(6271)
  not u5564 (Ncjiu6, n1362);  // ../RTL/cortexm0ds_logic.v(6271)
  and u5565 (n1363, Qvjiu6, Xvjiu6);  // ../RTL/cortexm0ds_logic.v(6272)
  not u5566 (Vujiu6, n1363);  // ../RTL/cortexm0ds_logic.v(6272)
  or u5567 (Xvjiu6, Ewjiu6, Lwjiu6);  // ../RTL/cortexm0ds_logic.v(6273)
  or u5568 (Cvjiu6, O95iu6, Jvjiu6);  // ../RTL/cortexm0ds_logic.v(6274)
  xor u5569 (Jvjiu6, Swjiu6, D7fpw6[6]);  // ../RTL/cortexm0ds_logic.v(6275)
  buf u557 (vis_r2_o[25], Uoqax6);  // ../RTL/cortexm0ds_logic.v(2551)
  and u5570 (n1364, Zwjiu6, Gxjiu6);  // ../RTL/cortexm0ds_logic.v(6276)
  not u5571 (Ucjiu6, n1364);  // ../RTL/cortexm0ds_logic.v(6276)
  and u5572 (Gxjiu6, Nxjiu6, Qvjiu6);  // ../RTL/cortexm0ds_logic.v(6277)
  and u5573 (n1365, Lwjiu6, Ewjiu6);  // ../RTL/cortexm0ds_logic.v(6278)
  not u5574 (Qvjiu6, n1365);  // ../RTL/cortexm0ds_logic.v(6278)
  xor u5575 (Ewjiu6, Uxjiu6, Byjiu6);  // ../RTL/cortexm0ds_logic.v(6279)
  or u5576 (n1366, Ad8iu6, Swjiu6);  // ../RTL/cortexm0ds_logic.v(6280)
  not u5577 (Lwjiu6, n1366);  // ../RTL/cortexm0ds_logic.v(6280)
  xor u5578 (Swjiu6, Iyjiu6, D7fpw6[5]);  // ../RTL/cortexm0ds_logic.v(6281)
  and u5579 (n1367, Byjiu6, Uxjiu6);  // ../RTL/cortexm0ds_logic.v(6282)
  buf u558 (vis_r2_o[7], Wcqax6);  // ../RTL/cortexm0ds_logic.v(2551)
  not u5580 (Nxjiu6, n1367);  // ../RTL/cortexm0ds_logic.v(6282)
  xor u5581 (Uxjiu6, Pyjiu6, Wyjiu6);  // ../RTL/cortexm0ds_logic.v(6283)
  or u5582 (n1368, Dzjiu6, Iyjiu6);  // ../RTL/cortexm0ds_logic.v(6284)
  not u5583 (Byjiu6, n1368);  // ../RTL/cortexm0ds_logic.v(6284)
  xor u5584 (Iyjiu6, Kzjiu6, D7fpw6[4]);  // ../RTL/cortexm0ds_logic.v(6285)
  and u5585 (Zwjiu6, Rzjiu6, Yzjiu6);  // ../RTL/cortexm0ds_logic.v(6286)
  and u5586 (n1369, Wyjiu6, Pyjiu6);  // ../RTL/cortexm0ds_logic.v(6287)
  not u5587 (Yzjiu6, n1369);  // ../RTL/cortexm0ds_logic.v(6287)
  xor u5588 (n1370, F0kiu6, M0kiu6);  // ../RTL/cortexm0ds_logic.v(6288)
  not u5589 (Pyjiu6, n1370);  // ../RTL/cortexm0ds_logic.v(6288)
  buf u559 (vis_r2_o[6], Xaqax6);  // ../RTL/cortexm0ds_logic.v(2551)
  or u5590 (F0kiu6, V4aiu6, T0kiu6);  // ../RTL/cortexm0ds_logic.v(6289)
  or u5591 (n1371, A1kiu6, Kzjiu6);  // ../RTL/cortexm0ds_logic.v(6290)
  not u5592 (Wyjiu6, n1371);  // ../RTL/cortexm0ds_logic.v(6290)
  xor u5593 (Kzjiu6, H1kiu6, V4aiu6);  // ../RTL/cortexm0ds_logic.v(6291)
  and u5594 (n1372, O1kiu6, D7fpw6[3]);  // ../RTL/cortexm0ds_logic.v(6292)
  not u5595 (Rzjiu6, n1372);  // ../RTL/cortexm0ds_logic.v(6292)
  and u5596 (O1kiu6, H1kiu6, M0kiu6);  // ../RTL/cortexm0ds_logic.v(6293)
  and u5597 (n1373, V1kiu6, C2kiu6);  // ../RTL/cortexm0ds_logic.v(6294)
  not u5598 (M0kiu6, n1373);  // ../RTL/cortexm0ds_logic.v(6294)
  or u5599 (C2kiu6, Prjiu6, J2kiu6);  // ../RTL/cortexm0ds_logic.v(6295)
  buf u56 (Hwmhu6, Vpkpw6);  // ../RTL/cortexm0ds_logic.v(1822)
  buf u560 (vis_r2_o[5], Y8qax6);  // ../RTL/cortexm0ds_logic.v(2551)
  or u5600 (V1kiu6, Rb8iu6, Ccaiu6);  // ../RTL/cortexm0ds_logic.v(6296)
  not u5601 (H1kiu6, T0kiu6);  // ../RTL/cortexm0ds_logic.v(6297)
  xor u5602 (T0kiu6, J2kiu6, D7fpw6[2]);  // ../RTL/cortexm0ds_logic.v(6298)
  xor u5603 (n1374, D7fpw6[0], D7fpw6[1]);  // ../RTL/cortexm0ds_logic.v(6299)
  not u5604 (J2kiu6, n1374);  // ../RTL/cortexm0ds_logic.v(6299)
  and u5605 (Gqjiu6, Q2kiu6, X2kiu6);  // ../RTL/cortexm0ds_logic.v(6300)
  and u5606 (n1375, E3kiu6, Ce8iu6);  // ../RTL/cortexm0ds_logic.v(6301)
  not u5607 (X2kiu6, n1375);  // ../RTL/cortexm0ds_logic.v(6301)
  and u5608 (n1376, L3kiu6, S3kiu6);  // ../RTL/cortexm0ds_logic.v(6302)
  not u5609 (Ce8iu6, n1376);  // ../RTL/cortexm0ds_logic.v(6302)
  buf u561 (X3fpw6[0], Vhspw6);  // ../RTL/cortexm0ds_logic.v(1784)
  and u5610 (L3kiu6, Z3kiu6, G4kiu6);  // ../RTL/cortexm0ds_logic.v(6303)
  and u5611 (n1377, N4kiu6, Cyfpw6[5]);  // ../RTL/cortexm0ds_logic.v(6304)
  not u5612 (G4kiu6, n1377);  // ../RTL/cortexm0ds_logic.v(6304)
  and u5613 (n1378, U98iu6, U4kiu6);  // ../RTL/cortexm0ds_logic.v(6305)
  not u5614 (Z3kiu6, n1378);  // ../RTL/cortexm0ds_logic.v(6305)
  xor u5615 (n1379, B5kiu6, Qajiu6);  // ../RTL/cortexm0ds_logic.v(6306)
  not u5616 (E3kiu6, n1379);  // ../RTL/cortexm0ds_logic.v(6306)
  or u5617 (n1380, Je8iu6, Y8biu6);  // ../RTL/cortexm0ds_logic.v(6307)
  not u5618 (Qajiu6, n1380);  // ../RTL/cortexm0ds_logic.v(6307)
  and u5619 (n1381, Tc8iu6, Ppfpw6[2]);  // ../RTL/cortexm0ds_logic.v(6308)
  buf u562 (vis_r2_o[9], Uarax6);  // ../RTL/cortexm0ds_logic.v(2551)
  not u5620 (Q2kiu6, n1381);  // ../RTL/cortexm0ds_logic.v(6308)
  and u5621 (Tc8iu6, Ivfhu6, I5kiu6);  // ../RTL/cortexm0ds_logic.v(6309)
  and u5622 (n1382, P5kiu6, W5kiu6);  // ../RTL/cortexm0ds_logic.v(6310)
  not u5623 (I5kiu6, n1382);  // ../RTL/cortexm0ds_logic.v(6310)
  and u5624 (n1383, D6kiu6, Qjaiu6);  // ../RTL/cortexm0ds_logic.v(6311)
  not u5625 (W5kiu6, n1383);  // ../RTL/cortexm0ds_logic.v(6311)
  and u5626 (Spjiu6, K6kiu6, R6kiu6);  // ../RTL/cortexm0ds_logic.v(6312)
  and u5627 (R6kiu6, Y6kiu6, F7kiu6);  // ../RTL/cortexm0ds_logic.v(6313)
  or u5628 (F7kiu6, Ndiiu6, Hd8iu6);  // ../RTL/cortexm0ds_logic.v(6314)
  or u5629 (n1384, Pdjiu6, M7kiu6);  // ../RTL/cortexm0ds_logic.v(6315)
  buf u563 (E1hpw6[28], Khgax6);  // ../RTL/cortexm0ds_logic.v(2367)
  not u5630 (Hd8iu6, n1384);  // ../RTL/cortexm0ds_logic.v(6315)
  and u5631 (n1385, T7kiu6, A8kiu6);  // ../RTL/cortexm0ds_logic.v(6316)
  not u5632 (Pdjiu6, n1385);  // ../RTL/cortexm0ds_logic.v(6316)
  and u5633 (n1386, H8kiu6, Ftjiu6);  // ../RTL/cortexm0ds_logic.v(6317)
  not u5634 (A8kiu6, n1386);  // ../RTL/cortexm0ds_logic.v(6317)
  and u5635 (n1387, O8kiu6, Vhiiu6);  // ../RTL/cortexm0ds_logic.v(6318)
  not u5636 (H8kiu6, n1387);  // ../RTL/cortexm0ds_logic.v(6318)
  and u5637 (n1388, M7kiu6, Oviiu6);  // ../RTL/cortexm0ds_logic.v(6319)
  not u5638 (T7kiu6, n1388);  // ../RTL/cortexm0ds_logic.v(6319)
  and u5639 (n1389, Habiu6, D7fpw6[1]);  // ../RTL/cortexm0ds_logic.v(6320)
  buf u564 (vis_r2_o[15], Zv7bx6);  // ../RTL/cortexm0ds_logic.v(2551)
  not u5640 (Y6kiu6, n1389);  // ../RTL/cortexm0ds_logic.v(6320)
  and u5641 (Habiu6, Ia8iu6, V8kiu6);  // ../RTL/cortexm0ds_logic.v(6321)
  and u5642 (n1390, H95iu6, C9kiu6);  // ../RTL/cortexm0ds_logic.v(6322)
  not u5643 (V8kiu6, n1390);  // ../RTL/cortexm0ds_logic.v(6322)
  and u5644 (n1391, J9kiu6, Oviiu6);  // ../RTL/cortexm0ds_logic.v(6323)
  not u5645 (C9kiu6, n1391);  // ../RTL/cortexm0ds_logic.v(6323)
  and u5646 (K6kiu6, Q9kiu6, X9kiu6);  // ../RTL/cortexm0ds_logic.v(6324)
  or u5647 (X9kiu6, Prjiu6, Yb8iu6);  // ../RTL/cortexm0ds_logic.v(6325)
  and u5648 (Yb8iu6, Eakiu6, Lakiu6);  // ../RTL/cortexm0ds_logic.v(6326)
  and u5649 (Lakiu6, Sakiu6, Zjiiu6);  // ../RTL/cortexm0ds_logic.v(6327)
  buf u565 (vis_r2_o[13], U4rax6);  // ../RTL/cortexm0ds_logic.v(2551)
  not u5650 (Zjiiu6, Zakiu6);  // ../RTL/cortexm0ds_logic.v(6328)
  and u5651 (n1392, Gbkiu6, Nyiiu6);  // ../RTL/cortexm0ds_logic.v(6329)
  not u5652 (Sakiu6, n1392);  // ../RTL/cortexm0ds_logic.v(6329)
  and u5653 (Gbkiu6, Ia8iu6, Nbkiu6);  // ../RTL/cortexm0ds_logic.v(6330)
  and u5654 (Eakiu6, Ubkiu6, Bckiu6);  // ../RTL/cortexm0ds_logic.v(6331)
  or u5655 (Bckiu6, E4jiu6, Jcaiu6);  // ../RTL/cortexm0ds_logic.v(6332)
  and u5656 (n1393, Cbbiu6, D7fpw6[7]);  // ../RTL/cortexm0ds_logic.v(6333)
  not u5657 (Q9kiu6, n1393);  // ../RTL/cortexm0ds_logic.v(6333)
  AL_MUX u5658 (
    .i0(Qcaiu6),
    .i1(vis_r2_o[2]),
    .sel(Ickiu6),
    .o(Hethu6));  // ../RTL/cortexm0ds_logic.v(6334)
  AL_MUX u5659 (
    .i0(Ef8iu6),
    .i1(vis_r2_o[4]),
    .sel(Ickiu6),
    .o(Aethu6));  // ../RTL/cortexm0ds_logic.v(6335)
  or u566 (Qbfpw6[24], Hz6ju6, M75ju6);  // ../RTL/cortexm0ds_logic.v(9482)
  AL_MUX u5660 (
    .i0(Vx9iu6),
    .i1(vis_r2_o[23]),
    .sel(Ickiu6),
    .o(Tdthu6));  // ../RTL/cortexm0ds_logic.v(6336)
  AL_MUX u5661 (
    .i0(K39iu6),
    .i1(vis_r2_o[30]),
    .sel(Ickiu6),
    .o(Mdthu6));  // ../RTL/cortexm0ds_logic.v(6337)
  AL_MUX u5662 (
    .i0(D39iu6),
    .i1(vis_r2_o[31]),
    .sel(Ickiu6),
    .o(Fdthu6));  // ../RTL/cortexm0ds_logic.v(6338)
  AL_MUX u5663 (
    .i0(Tx8iu6),
    .i1(vis_r2_o[0]),
    .sel(Ickiu6),
    .o(Ycthu6));  // ../RTL/cortexm0ds_logic.v(6339)
  AL_MUX u5664 (
    .i0(Qcaiu6),
    .i1(vis_r3_o[2]),
    .sel(Pckiu6),
    .o(Rcthu6));  // ../RTL/cortexm0ds_logic.v(6340)
  AL_MUX u5665 (
    .i0(Ef8iu6),
    .i1(vis_r3_o[4]),
    .sel(Pckiu6),
    .o(Kcthu6));  // ../RTL/cortexm0ds_logic.v(6341)
  AL_MUX u5666 (
    .i0(Vx9iu6),
    .i1(vis_r3_o[23]),
    .sel(Pckiu6),
    .o(Dcthu6));  // ../RTL/cortexm0ds_logic.v(6342)
  AL_MUX u5667 (
    .i0(K39iu6),
    .i1(vis_r3_o[30]),
    .sel(Pckiu6),
    .o(Wbthu6));  // ../RTL/cortexm0ds_logic.v(6343)
  AL_MUX u5668 (
    .i0(D39iu6),
    .i1(vis_r3_o[31]),
    .sel(Pckiu6),
    .o(Pbthu6));  // ../RTL/cortexm0ds_logic.v(6344)
  AL_MUX u5669 (
    .i0(Tx8iu6),
    .i1(vis_r3_o[0]),
    .sel(Pckiu6),
    .o(Ibthu6));  // ../RTL/cortexm0ds_logic.v(6345)
  buf u567 (E1hpw6[16], Kcaax6);  // ../RTL/cortexm0ds_logic.v(2367)
  AL_MUX u5670 (
    .i0(Qcaiu6),
    .i1(vis_r4_o[2]),
    .sel(Wckiu6),
    .o(Bbthu6));  // ../RTL/cortexm0ds_logic.v(6346)
  AL_MUX u5671 (
    .i0(Ef8iu6),
    .i1(vis_r4_o[4]),
    .sel(Wckiu6),
    .o(Uathu6));  // ../RTL/cortexm0ds_logic.v(6347)
  AL_MUX u5672 (
    .i0(Vx9iu6),
    .i1(vis_r4_o[23]),
    .sel(Wckiu6),
    .o(Nathu6));  // ../RTL/cortexm0ds_logic.v(6348)
  AL_MUX u5673 (
    .i0(K39iu6),
    .i1(vis_r4_o[30]),
    .sel(Wckiu6),
    .o(Gathu6));  // ../RTL/cortexm0ds_logic.v(6349)
  AL_MUX u5674 (
    .i0(D39iu6),
    .i1(vis_r4_o[31]),
    .sel(Wckiu6),
    .o(Z9thu6));  // ../RTL/cortexm0ds_logic.v(6350)
  AL_MUX u5675 (
    .i0(Tx8iu6),
    .i1(vis_r4_o[0]),
    .sel(Wckiu6),
    .o(S9thu6));  // ../RTL/cortexm0ds_logic.v(6351)
  AL_MUX u5676 (
    .i0(Qcaiu6),
    .i1(vis_r5_o[2]),
    .sel(Ddkiu6),
    .o(L9thu6));  // ../RTL/cortexm0ds_logic.v(6352)
  AL_MUX u5677 (
    .i0(Ef8iu6),
    .i1(vis_r5_o[4]),
    .sel(Ddkiu6),
    .o(E9thu6));  // ../RTL/cortexm0ds_logic.v(6353)
  AL_MUX u5678 (
    .i0(Vx9iu6),
    .i1(vis_r5_o[23]),
    .sel(Ddkiu6),
    .o(X8thu6));  // ../RTL/cortexm0ds_logic.v(6354)
  AL_MUX u5679 (
    .i0(K39iu6),
    .i1(vis_r5_o[30]),
    .sel(Ddkiu6),
    .o(Q8thu6));  // ../RTL/cortexm0ds_logic.v(6355)
  buf u568 (L3ehu6, I8lax6);  // ../RTL/cortexm0ds_logic.v(2463)
  AL_MUX u5680 (
    .i0(D39iu6),
    .i1(vis_r5_o[31]),
    .sel(Ddkiu6),
    .o(J8thu6));  // ../RTL/cortexm0ds_logic.v(6356)
  AL_MUX u5681 (
    .i0(Tx8iu6),
    .i1(vis_r5_o[0]),
    .sel(Ddkiu6),
    .o(C8thu6));  // ../RTL/cortexm0ds_logic.v(6357)
  AL_MUX u5682 (
    .i0(Qcaiu6),
    .i1(vis_r6_o[2]),
    .sel(Kdkiu6),
    .o(V7thu6));  // ../RTL/cortexm0ds_logic.v(6358)
  AL_MUX u5683 (
    .i0(Ef8iu6),
    .i1(vis_r6_o[4]),
    .sel(Kdkiu6),
    .o(O7thu6));  // ../RTL/cortexm0ds_logic.v(6359)
  AL_MUX u5684 (
    .i0(Vx9iu6),
    .i1(vis_r6_o[23]),
    .sel(Kdkiu6),
    .o(H7thu6));  // ../RTL/cortexm0ds_logic.v(6360)
  AL_MUX u5685 (
    .i0(K39iu6),
    .i1(vis_r6_o[30]),
    .sel(Kdkiu6),
    .o(A7thu6));  // ../RTL/cortexm0ds_logic.v(6361)
  AL_MUX u5686 (
    .i0(D39iu6),
    .i1(vis_r6_o[31]),
    .sel(Kdkiu6),
    .o(T6thu6));  // ../RTL/cortexm0ds_logic.v(6362)
  AL_MUX u5687 (
    .i0(Tx8iu6),
    .i1(vis_r6_o[0]),
    .sel(Kdkiu6),
    .o(M6thu6));  // ../RTL/cortexm0ds_logic.v(6363)
  AL_MUX u5688 (
    .i0(Qcaiu6),
    .i1(vis_r7_o[2]),
    .sel(Rdkiu6),
    .o(F6thu6));  // ../RTL/cortexm0ds_logic.v(6364)
  AL_MUX u5689 (
    .i0(Ef8iu6),
    .i1(vis_r7_o[4]),
    .sel(Rdkiu6),
    .o(Y5thu6));  // ../RTL/cortexm0ds_logic.v(6365)
  buf u569 (Qwdhu6, Halax6);  // ../RTL/cortexm0ds_logic.v(2464)
  AL_MUX u5690 (
    .i0(Vx9iu6),
    .i1(vis_r7_o[23]),
    .sel(Rdkiu6),
    .o(R5thu6));  // ../RTL/cortexm0ds_logic.v(6366)
  AL_MUX u5691 (
    .i0(K39iu6),
    .i1(vis_r7_o[30]),
    .sel(Rdkiu6),
    .o(K5thu6));  // ../RTL/cortexm0ds_logic.v(6367)
  AL_MUX u5692 (
    .i0(D39iu6),
    .i1(vis_r7_o[31]),
    .sel(Rdkiu6),
    .o(D5thu6));  // ../RTL/cortexm0ds_logic.v(6368)
  AL_MUX u5693 (
    .i0(Tx8iu6),
    .i1(vis_r7_o[0]),
    .sel(Rdkiu6),
    .o(W4thu6));  // ../RTL/cortexm0ds_logic.v(6369)
  AL_MUX u5694 (
    .i0(vis_psp_o[0]),
    .i1(Qcaiu6),
    .sel(Ydkiu6),
    .o(P4thu6));  // ../RTL/cortexm0ds_logic.v(6370)
  AL_MUX u5695 (
    .i0(vis_psp_o[29]),
    .i1(D39iu6),
    .sel(Ydkiu6),
    .o(I4thu6));  // ../RTL/cortexm0ds_logic.v(6371)
  AL_MUX u5696 (
    .i0(vis_psp_o[28]),
    .i1(K39iu6),
    .sel(Ydkiu6),
    .o(B4thu6));  // ../RTL/cortexm0ds_logic.v(6372)
  AL_MUX u5697 (
    .i0(vis_psp_o[21]),
    .i1(Vx9iu6),
    .sel(Ydkiu6),
    .o(U3thu6));  // ../RTL/cortexm0ds_logic.v(6373)
  AL_MUX u5698 (
    .i0(vis_psp_o[2]),
    .i1(Ef8iu6),
    .sel(Ydkiu6),
    .o(N3thu6));  // ../RTL/cortexm0ds_logic.v(6374)
  AL_MUX u5699 (
    .i0(vis_msp_o[0]),
    .i1(Qcaiu6),
    .sel(Fekiu6),
    .o(G3thu6));  // ../RTL/cortexm0ds_logic.v(6375)
  buf u57 (Jfgpw6[3], R9yax6);  // ../RTL/cortexm0ds_logic.v(2010)
  buf u570 (Hrfpw6[0], Tcjax6);  // ../RTL/cortexm0ds_logic.v(2428)
  AL_MUX u5700 (
    .i0(vis_msp_o[29]),
    .i1(D39iu6),
    .sel(Fekiu6),
    .o(Z2thu6));  // ../RTL/cortexm0ds_logic.v(6376)
  AL_MUX u5701 (
    .i0(vis_msp_o[28]),
    .i1(K39iu6),
    .sel(Fekiu6),
    .o(S2thu6));  // ../RTL/cortexm0ds_logic.v(6377)
  AL_MUX u5702 (
    .i0(vis_msp_o[21]),
    .i1(Vx9iu6),
    .sel(Fekiu6),
    .o(L2thu6));  // ../RTL/cortexm0ds_logic.v(6378)
  AL_MUX u5703 (
    .i0(vis_msp_o[2]),
    .i1(Ef8iu6),
    .sel(Fekiu6),
    .o(E2thu6));  // ../RTL/cortexm0ds_logic.v(6379)
  AL_MUX u5704 (
    .i0(Qcaiu6),
    .i1(vis_r14_o[2]),
    .sel(Mekiu6),
    .o(X1thu6));  // ../RTL/cortexm0ds_logic.v(6380)
  AL_MUX u5705 (
    .i0(Ef8iu6),
    .i1(vis_r14_o[4]),
    .sel(Mekiu6),
    .o(Q1thu6));  // ../RTL/cortexm0ds_logic.v(6381)
  AL_MUX u5706 (
    .i0(Vx9iu6),
    .i1(vis_r14_o[23]),
    .sel(Mekiu6),
    .o(J1thu6));  // ../RTL/cortexm0ds_logic.v(6382)
  AL_MUX u5707 (
    .i0(K39iu6),
    .i1(vis_r14_o[30]),
    .sel(Mekiu6),
    .o(C1thu6));  // ../RTL/cortexm0ds_logic.v(6383)
  AL_MUX u5708 (
    .i0(D39iu6),
    .i1(vis_r14_o[31]),
    .sel(Mekiu6),
    .o(V0thu6));  // ../RTL/cortexm0ds_logic.v(6384)
  AL_MUX u5709 (
    .i0(Tx8iu6),
    .i1(vis_r14_o[0]),
    .sel(Mekiu6),
    .o(O0thu6));  // ../RTL/cortexm0ds_logic.v(6385)
  buf u571 (D7fpw6[5], Jckax6);  // ../RTL/cortexm0ds_logic.v(2074)
  AL_MUX u5710 (
    .i0(Qcaiu6),
    .i1(vis_r12_o[2]),
    .sel(Tekiu6),
    .o(H0thu6));  // ../RTL/cortexm0ds_logic.v(6386)
  AL_MUX u5711 (
    .i0(Ef8iu6),
    .i1(vis_r12_o[4]),
    .sel(Tekiu6),
    .o(A0thu6));  // ../RTL/cortexm0ds_logic.v(6387)
  AL_MUX u5712 (
    .i0(Vx9iu6),
    .i1(vis_r12_o[23]),
    .sel(Tekiu6),
    .o(Tzshu6));  // ../RTL/cortexm0ds_logic.v(6388)
  AL_MUX u5713 (
    .i0(K39iu6),
    .i1(vis_r12_o[30]),
    .sel(Tekiu6),
    .o(Mzshu6));  // ../RTL/cortexm0ds_logic.v(6389)
  AL_MUX u5714 (
    .i0(D39iu6),
    .i1(vis_r12_o[31]),
    .sel(Tekiu6),
    .o(Fzshu6));  // ../RTL/cortexm0ds_logic.v(6390)
  AL_MUX u5715 (
    .i0(Tx8iu6),
    .i1(vis_r12_o[0]),
    .sel(Tekiu6),
    .o(Yyshu6));  // ../RTL/cortexm0ds_logic.v(6391)
  AL_MUX u5716 (
    .i0(Qcaiu6),
    .i1(vis_r11_o[2]),
    .sel(Afkiu6),
    .o(Ryshu6));  // ../RTL/cortexm0ds_logic.v(6392)
  AL_MUX u5717 (
    .i0(Ef8iu6),
    .i1(vis_r11_o[4]),
    .sel(Afkiu6),
    .o(Kyshu6));  // ../RTL/cortexm0ds_logic.v(6393)
  AL_MUX u5718 (
    .i0(Vx9iu6),
    .i1(vis_r11_o[23]),
    .sel(Afkiu6),
    .o(Dyshu6));  // ../RTL/cortexm0ds_logic.v(6394)
  AL_MUX u5719 (
    .i0(K39iu6),
    .i1(vis_r11_o[30]),
    .sel(Afkiu6),
    .o(Wxshu6));  // ../RTL/cortexm0ds_logic.v(6395)
  buf u572 (D7fpw6[3], Wkipw6);  // ../RTL/cortexm0ds_logic.v(2074)
  AL_MUX u5720 (
    .i0(D39iu6),
    .i1(vis_r11_o[31]),
    .sel(Afkiu6),
    .o(Pxshu6));  // ../RTL/cortexm0ds_logic.v(6396)
  AL_MUX u5721 (
    .i0(Tx8iu6),
    .i1(vis_r11_o[0]),
    .sel(Afkiu6),
    .o(Ixshu6));  // ../RTL/cortexm0ds_logic.v(6397)
  AL_MUX u5722 (
    .i0(Qcaiu6),
    .i1(vis_r10_o[2]),
    .sel(Hfkiu6),
    .o(Bxshu6));  // ../RTL/cortexm0ds_logic.v(6398)
  AL_MUX u5723 (
    .i0(Ef8iu6),
    .i1(vis_r10_o[4]),
    .sel(Hfkiu6),
    .o(Uwshu6));  // ../RTL/cortexm0ds_logic.v(6399)
  AL_MUX u5724 (
    .i0(Vx9iu6),
    .i1(vis_r10_o[23]),
    .sel(Hfkiu6),
    .o(Nwshu6));  // ../RTL/cortexm0ds_logic.v(6400)
  AL_MUX u5725 (
    .i0(K39iu6),
    .i1(vis_r10_o[30]),
    .sel(Hfkiu6),
    .o(Gwshu6));  // ../RTL/cortexm0ds_logic.v(6401)
  AL_MUX u5726 (
    .i0(D39iu6),
    .i1(vis_r10_o[31]),
    .sel(Hfkiu6),
    .o(Zvshu6));  // ../RTL/cortexm0ds_logic.v(6402)
  AL_MUX u5727 (
    .i0(Tx8iu6),
    .i1(vis_r10_o[0]),
    .sel(Hfkiu6),
    .o(Svshu6));  // ../RTL/cortexm0ds_logic.v(6403)
  AL_MUX u5728 (
    .i0(Qcaiu6),
    .i1(vis_r9_o[2]),
    .sel(Ofkiu6),
    .o(Lvshu6));  // ../RTL/cortexm0ds_logic.v(6404)
  AL_MUX u5729 (
    .i0(Ef8iu6),
    .i1(vis_r9_o[4]),
    .sel(Ofkiu6),
    .o(Evshu6));  // ../RTL/cortexm0ds_logic.v(6405)
  buf u573 (Tzfpw6[7], Ujxax6);  // ../RTL/cortexm0ds_logic.v(2007)
  AL_MUX u5730 (
    .i0(Vx9iu6),
    .i1(vis_r9_o[23]),
    .sel(Ofkiu6),
    .o(Xushu6));  // ../RTL/cortexm0ds_logic.v(6406)
  AL_MUX u5731 (
    .i0(K39iu6),
    .i1(vis_r9_o[30]),
    .sel(Ofkiu6),
    .o(Qushu6));  // ../RTL/cortexm0ds_logic.v(6407)
  AL_MUX u5732 (
    .i0(D39iu6),
    .i1(vis_r9_o[31]),
    .sel(Ofkiu6),
    .o(Jushu6));  // ../RTL/cortexm0ds_logic.v(6408)
  AL_MUX u5733 (
    .i0(Tx8iu6),
    .i1(vis_r9_o[0]),
    .sel(Ofkiu6),
    .o(Cushu6));  // ../RTL/cortexm0ds_logic.v(6409)
  AL_MUX u5734 (
    .i0(Qcaiu6),
    .i1(vis_r8_o[2]),
    .sel(Vfkiu6),
    .o(Vtshu6));  // ../RTL/cortexm0ds_logic.v(6410)
  and u5735 (n1394, Ogciu6, Cgkiu6);  // ../RTL/cortexm0ds_logic.v(6411)
  not u5736 (Qcaiu6, n1394);  // ../RTL/cortexm0ds_logic.v(6411)
  AL_MUX u5737 (
    .i0(Jgkiu6),
    .i1(vis_r8_o[3]),
    .sel(Vfkiu6),
    .o(Otshu6));  // ../RTL/cortexm0ds_logic.v(6412)
  and u5738 (n1395, Qgkiu6, Xgkiu6);  // ../RTL/cortexm0ds_logic.v(6413)
  not u5739 (Htshu6, n1395);  // ../RTL/cortexm0ds_logic.v(6413)
  buf u574 (H2fpw6[3], M6kax6);  // ../RTL/cortexm0ds_logic.v(2444)
  and u5740 (Xgkiu6, Ehkiu6, Lhkiu6);  // ../RTL/cortexm0ds_logic.v(6414)
  and u5741 (n1396, Ok8iu6, vis_pc_o[2]);  // ../RTL/cortexm0ds_logic.v(6415)
  not u5742 (Lhkiu6, n1396);  // ../RTL/cortexm0ds_logic.v(6415)
  and u5743 (Ehkiu6, Shkiu6, Zhkiu6);  // ../RTL/cortexm0ds_logic.v(6416)
  and u5744 (n1397, Jl8iu6, Tugpw6[1]);  // ../RTL/cortexm0ds_logic.v(6417)
  not u5745 (Zhkiu6, n1397);  // ../RTL/cortexm0ds_logic.v(6417)
  buf u5746 (vis_r7_o[15], Zd8bx6);  // ../RTL/cortexm0ds_logic.v(2654)
  buf u5747 (vis_r7_o[27], M7wax6);  // ../RTL/cortexm0ds_logic.v(2654)
  and u5748 (n1398, N5fpw6[2], Sdaiu6);  // ../RTL/cortexm0ds_logic.v(6419)
  not u5749 (Nikiu6, n1398);  // ../RTL/cortexm0ds_logic.v(6419)
  buf u575 (vis_r11_o[0], Pwkax6);  // ../RTL/cortexm0ds_logic.v(1874)
  and u5750 (Gikiu6, Uikiu6, Bjkiu6);  // ../RTL/cortexm0ds_logic.v(6420)
  or u5751 (Bjkiu6, T2iiu6, Lg0iu6);  // ../RTL/cortexm0ds_logic.v(6421)
  and u5752 (n1399, Eafpw6[3], A3iiu6);  // ../RTL/cortexm0ds_logic.v(6422)
  not u5753 (Uikiu6, n1399);  // ../RTL/cortexm0ds_logic.v(6422)
  and u5754 (n1400, Ql8iu6, vis_ipsr_o[3]);  // ../RTL/cortexm0ds_logic.v(6423)
  not u5755 (Shkiu6, n1400);  // ../RTL/cortexm0ds_logic.v(6423)
  and u5756 (Qgkiu6, Ijkiu6, Pjkiu6);  // ../RTL/cortexm0ds_logic.v(6424)
  or u5757 (Pjkiu6, Lm8iu6, Wjkiu6);  // ../RTL/cortexm0ds_logic.v(6425)
  and u5758 (n1401, Zm8iu6, Df4iu6);  // ../RTL/cortexm0ds_logic.v(6426)
  not u5759 (Ijkiu6, n1401);  // ../RTL/cortexm0ds_logic.v(6426)
  buf u576 (D7fpw6[7], N4kax6);  // ../RTL/cortexm0ds_logic.v(2074)
  AL_MUX u5760 (
    .i0(vis_psp_o[1]),
    .i1(Jgkiu6),
    .sel(Ydkiu6),
    .o(Atshu6));  // ../RTL/cortexm0ds_logic.v(6427)
  AL_MUX u5761 (
    .i0(vis_msp_o[1]),
    .i1(Jgkiu6),
    .sel(Fekiu6),
    .o(Tsshu6));  // ../RTL/cortexm0ds_logic.v(6428)
  AL_MUX u5762 (
    .i0(Jgkiu6),
    .i1(vis_r14_o[3]),
    .sel(Mekiu6),
    .o(Msshu6));  // ../RTL/cortexm0ds_logic.v(6429)
  AL_MUX u5763 (
    .i0(Jgkiu6),
    .i1(vis_r12_o[3]),
    .sel(Tekiu6),
    .o(Fsshu6));  // ../RTL/cortexm0ds_logic.v(6430)
  AL_MUX u5764 (
    .i0(Jgkiu6),
    .i1(vis_r7_o[3]),
    .sel(Rdkiu6),
    .o(Yrshu6));  // ../RTL/cortexm0ds_logic.v(6431)
  AL_MUX u5765 (
    .i0(Jgkiu6),
    .i1(vis_r6_o[3]),
    .sel(Kdkiu6),
    .o(Rrshu6));  // ../RTL/cortexm0ds_logic.v(6432)
  AL_MUX u5766 (
    .i0(Jgkiu6),
    .i1(vis_r5_o[3]),
    .sel(Ddkiu6),
    .o(Krshu6));  // ../RTL/cortexm0ds_logic.v(6433)
  AL_MUX u5767 (
    .i0(Jgkiu6),
    .i1(vis_r4_o[3]),
    .sel(Wckiu6),
    .o(Drshu6));  // ../RTL/cortexm0ds_logic.v(6434)
  AL_MUX u5768 (
    .i0(Jgkiu6),
    .i1(vis_r11_o[3]),
    .sel(Afkiu6),
    .o(Wqshu6));  // ../RTL/cortexm0ds_logic.v(6435)
  AL_MUX u5769 (
    .i0(Jgkiu6),
    .i1(vis_r10_o[3]),
    .sel(Hfkiu6),
    .o(Pqshu6));  // ../RTL/cortexm0ds_logic.v(6436)
  buf u577 (D7fpw6[4], Jgxpw6);  // ../RTL/cortexm0ds_logic.v(2074)
  AL_MUX u5770 (
    .i0(Jgkiu6),
    .i1(vis_r9_o[3]),
    .sel(Ofkiu6),
    .o(Iqshu6));  // ../RTL/cortexm0ds_logic.v(6437)
  AL_MUX u5771 (
    .i0(Jgkiu6),
    .i1(vis_r3_o[3]),
    .sel(Pckiu6),
    .o(Bqshu6));  // ../RTL/cortexm0ds_logic.v(6438)
  AL_MUX u5772 (
    .i0(Jgkiu6),
    .i1(vis_r2_o[3]),
    .sel(Ickiu6),
    .o(Upshu6));  // ../RTL/cortexm0ds_logic.v(6439)
  AL_MUX u5773 (
    .i0(Jgkiu6),
    .i1(vis_r1_o[3]),
    .sel(Mx8iu6),
    .o(Npshu6));  // ../RTL/cortexm0ds_logic.v(6440)
  AL_MUX u5774 (
    .i0(Jgkiu6),
    .i1(vis_r0_o[3]),
    .sel(Lf8iu6),
    .o(Gpshu6));  // ../RTL/cortexm0ds_logic.v(6441)
  and u5775 (n1402, Kifiu6, Dkkiu6);  // ../RTL/cortexm0ds_logic.v(6442)
  not u5776 (Jgkiu6, n1402);  // ../RTL/cortexm0ds_logic.v(6442)
  AL_MUX u5777 (
    .i0(Ef8iu6),
    .i1(vis_r8_o[4]),
    .sel(Vfkiu6),
    .o(Zoshu6));  // ../RTL/cortexm0ds_logic.v(6443)
  and u5778 (n1403, Y4fiu6, Kkkiu6);  // ../RTL/cortexm0ds_logic.v(6444)
  not u5779 (Ef8iu6, n1403);  // ../RTL/cortexm0ds_logic.v(6444)
  buf u578 (D7fpw6[2], Irmpw6);  // ../RTL/cortexm0ds_logic.v(2074)
  AL_MUX u5780 (
    .i0(Rkkiu6),
    .i1(vis_r8_o[5]),
    .sel(Vfkiu6),
    .o(Soshu6));  // ../RTL/cortexm0ds_logic.v(6445)
  and u5781 (n1404, Ykkiu6, Flkiu6);  // ../RTL/cortexm0ds_logic.v(6446)
  not u5782 (Loshu6, n1404);  // ../RTL/cortexm0ds_logic.v(6446)
  and u5783 (Flkiu6, Mlkiu6, Tlkiu6);  // ../RTL/cortexm0ds_logic.v(6447)
  and u5784 (n1405, vis_pc_o[4], Ok8iu6);  // ../RTL/cortexm0ds_logic.v(6448)
  not u5785 (Tlkiu6, n1405);  // ../RTL/cortexm0ds_logic.v(6448)
  and u5786 (Mlkiu6, Amkiu6, Hmkiu6);  // ../RTL/cortexm0ds_logic.v(6449)
  and u5787 (n1406, Jl8iu6, Tugpw6[3]);  // ../RTL/cortexm0ds_logic.v(6450)
  not u5788 (Hmkiu6, n1406);  // ../RTL/cortexm0ds_logic.v(6450)
  buf u5789 (vis_r7_o[13], Ltwax6);  // ../RTL/cortexm0ds_logic.v(2654)
  buf u579 (D7fpw6[1], S7mpw6);  // ../RTL/cortexm0ds_logic.v(2074)
  buf u5790 (vis_r7_o[25], Ldwax6);  // ../RTL/cortexm0ds_logic.v(2654)
  and u5791 (n1407, N5fpw6[4], Sdaiu6);  // ../RTL/cortexm0ds_logic.v(6452)
  not u5792 (Vmkiu6, n1407);  // ../RTL/cortexm0ds_logic.v(6452)
  and u5793 (Omkiu6, Cnkiu6, Jnkiu6);  // ../RTL/cortexm0ds_logic.v(6453)
  or u5794 (Jnkiu6, T2iiu6, Xf0iu6);  // ../RTL/cortexm0ds_logic.v(6454)
  and u5795 (n1408, Eafpw6[5], A3iiu6);  // ../RTL/cortexm0ds_logic.v(6455)
  not u5796 (Cnkiu6, n1408);  // ../RTL/cortexm0ds_logic.v(6455)
  and u5797 (n1409, Ql8iu6, vis_ipsr_o[5]);  // ../RTL/cortexm0ds_logic.v(6456)
  not u5798 (Amkiu6, n1409);  // ../RTL/cortexm0ds_logic.v(6456)
  and u5799 (Ykkiu6, Qnkiu6, Xnkiu6);  // ../RTL/cortexm0ds_logic.v(6457)
  buf u58 (vis_r5_o[27], Lfppw6);  // ../RTL/cortexm0ds_logic.v(1909)
  buf u580 (Tzfpw6[23], Coupw6);  // ../RTL/cortexm0ds_logic.v(2007)
  or u5800 (Xnkiu6, Lm8iu6, Eokiu6);  // ../RTL/cortexm0ds_logic.v(6458)
  and u5801 (n1410, Zm8iu6, Oh4iu6);  // ../RTL/cortexm0ds_logic.v(6459)
  not u5802 (Qnkiu6, n1410);  // ../RTL/cortexm0ds_logic.v(6459)
  AL_MUX u5803 (
    .i0(vis_psp_o[3]),
    .i1(Rkkiu6),
    .sel(Ydkiu6),
    .o(Eoshu6));  // ../RTL/cortexm0ds_logic.v(6460)
  AL_MUX u5804 (
    .i0(vis_msp_o[3]),
    .i1(Rkkiu6),
    .sel(Fekiu6),
    .o(Xnshu6));  // ../RTL/cortexm0ds_logic.v(6461)
  AL_MUX u5805 (
    .i0(Rkkiu6),
    .i1(vis_r14_o[5]),
    .sel(Mekiu6),
    .o(Qnshu6));  // ../RTL/cortexm0ds_logic.v(6462)
  AL_MUX u5806 (
    .i0(Rkkiu6),
    .i1(vis_r12_o[5]),
    .sel(Tekiu6),
    .o(Jnshu6));  // ../RTL/cortexm0ds_logic.v(6463)
  AL_MUX u5807 (
    .i0(Rkkiu6),
    .i1(vis_r7_o[5]),
    .sel(Rdkiu6),
    .o(Cnshu6));  // ../RTL/cortexm0ds_logic.v(6464)
  AL_MUX u5808 (
    .i0(Rkkiu6),
    .i1(vis_r6_o[5]),
    .sel(Kdkiu6),
    .o(Vmshu6));  // ../RTL/cortexm0ds_logic.v(6465)
  AL_MUX u5809 (
    .i0(Rkkiu6),
    .i1(vis_r5_o[5]),
    .sel(Ddkiu6),
    .o(Omshu6));  // ../RTL/cortexm0ds_logic.v(6466)
  buf u581 (Tzfpw6[6], Rv7ax6);  // ../RTL/cortexm0ds_logic.v(2007)
  AL_MUX u5810 (
    .i0(Rkkiu6),
    .i1(vis_r4_o[5]),
    .sel(Wckiu6),
    .o(Hmshu6));  // ../RTL/cortexm0ds_logic.v(6467)
  AL_MUX u5811 (
    .i0(Rkkiu6),
    .i1(vis_r11_o[5]),
    .sel(Afkiu6),
    .o(Amshu6));  // ../RTL/cortexm0ds_logic.v(6468)
  AL_MUX u5812 (
    .i0(Rkkiu6),
    .i1(vis_r10_o[5]),
    .sel(Hfkiu6),
    .o(Tlshu6));  // ../RTL/cortexm0ds_logic.v(6469)
  AL_MUX u5813 (
    .i0(Rkkiu6),
    .i1(vis_r9_o[5]),
    .sel(Ofkiu6),
    .o(Mlshu6));  // ../RTL/cortexm0ds_logic.v(6470)
  AL_MUX u5814 (
    .i0(Rkkiu6),
    .i1(vis_r3_o[5]),
    .sel(Pckiu6),
    .o(Flshu6));  // ../RTL/cortexm0ds_logic.v(6471)
  AL_MUX u5815 (
    .i0(Rkkiu6),
    .i1(vis_r2_o[5]),
    .sel(Ickiu6),
    .o(Ykshu6));  // ../RTL/cortexm0ds_logic.v(6472)
  AL_MUX u5816 (
    .i0(Rkkiu6),
    .i1(vis_r1_o[5]),
    .sel(Mx8iu6),
    .o(Rkshu6));  // ../RTL/cortexm0ds_logic.v(6473)
  AL_MUX u5817 (
    .i0(Rkkiu6),
    .i1(vis_r0_o[5]),
    .sel(Lf8iu6),
    .o(Kkshu6));  // ../RTL/cortexm0ds_logic.v(6474)
  and u5818 (n1411, Ljbiu6, Lokiu6);  // ../RTL/cortexm0ds_logic.v(6475)
  not u5819 (Rkkiu6, n1411);  // ../RTL/cortexm0ds_logic.v(6475)
  buf u582 (Tzfpw6[4], Johbx6);  // ../RTL/cortexm0ds_logic.v(2007)
  AL_MUX u5820 (
    .i0(Sokiu6),
    .i1(vis_r8_o[6]),
    .sel(Vfkiu6),
    .o(Dkshu6));  // ../RTL/cortexm0ds_logic.v(6476)
  and u5821 (n1412, Zokiu6, Gpkiu6);  // ../RTL/cortexm0ds_logic.v(6477)
  not u5822 (Wjshu6, n1412);  // ../RTL/cortexm0ds_logic.v(6477)
  and u5823 (Gpkiu6, Npkiu6, Upkiu6);  // ../RTL/cortexm0ds_logic.v(6478)
  and u5824 (n1413, Jl8iu6, Tugpw6[4]);  // ../RTL/cortexm0ds_logic.v(6479)
  not u5825 (Upkiu6, n1413);  // ../RTL/cortexm0ds_logic.v(6479)
  and u5826 (n1414, vis_pc_o[5], Ok8iu6);  // ../RTL/cortexm0ds_logic.v(6480)
  not u5827 (Npkiu6, n1414);  // ../RTL/cortexm0ds_logic.v(6480)
  and u5828 (Zokiu6, Bqkiu6, Iqkiu6);  // ../RTL/cortexm0ds_logic.v(6481)
  and u5829 (n1415, W29iu6, Fkfpw6[6]);  // ../RTL/cortexm0ds_logic.v(6482)
  buf u583 (Tzfpw6[3], P0ibx6);  // ../RTL/cortexm0ds_logic.v(2007)
  not u5830 (Iqkiu6, n1415);  // ../RTL/cortexm0ds_logic.v(6482)
  and u5831 (n1416, Zm8iu6, Xi4iu6);  // ../RTL/cortexm0ds_logic.v(6483)
  not u5832 (Bqkiu6, n1416);  // ../RTL/cortexm0ds_logic.v(6483)
  AL_MUX u5833 (
    .i0(vis_psp_o[4]),
    .i1(Sokiu6),
    .sel(Ydkiu6),
    .o(Pjshu6));  // ../RTL/cortexm0ds_logic.v(6484)
  AL_MUX u5834 (
    .i0(vis_msp_o[4]),
    .i1(Sokiu6),
    .sel(Fekiu6),
    .o(Ijshu6));  // ../RTL/cortexm0ds_logic.v(6485)
  AL_MUX u5835 (
    .i0(Sokiu6),
    .i1(vis_r14_o[6]),
    .sel(Mekiu6),
    .o(Bjshu6));  // ../RTL/cortexm0ds_logic.v(6486)
  AL_MUX u5836 (
    .i0(Sokiu6),
    .i1(vis_r12_o[6]),
    .sel(Tekiu6),
    .o(Uishu6));  // ../RTL/cortexm0ds_logic.v(6487)
  AL_MUX u5837 (
    .i0(Sokiu6),
    .i1(vis_r7_o[6]),
    .sel(Rdkiu6),
    .o(Nishu6));  // ../RTL/cortexm0ds_logic.v(6488)
  AL_MUX u5838 (
    .i0(Sokiu6),
    .i1(vis_r6_o[6]),
    .sel(Kdkiu6),
    .o(Gishu6));  // ../RTL/cortexm0ds_logic.v(6489)
  AL_MUX u5839 (
    .i0(Sokiu6),
    .i1(vis_r5_o[6]),
    .sel(Ddkiu6),
    .o(Zhshu6));  // ../RTL/cortexm0ds_logic.v(6490)
  buf u584 (Tzfpw6[1], Oarpw6);  // ../RTL/cortexm0ds_logic.v(2007)
  AL_MUX u5840 (
    .i0(Sokiu6),
    .i1(vis_r4_o[6]),
    .sel(Wckiu6),
    .o(Shshu6));  // ../RTL/cortexm0ds_logic.v(6491)
  AL_MUX u5841 (
    .i0(Sokiu6),
    .i1(vis_r11_o[6]),
    .sel(Afkiu6),
    .o(Lhshu6));  // ../RTL/cortexm0ds_logic.v(6492)
  AL_MUX u5842 (
    .i0(Sokiu6),
    .i1(vis_r10_o[6]),
    .sel(Hfkiu6),
    .o(Ehshu6));  // ../RTL/cortexm0ds_logic.v(6493)
  AL_MUX u5843 (
    .i0(Sokiu6),
    .i1(vis_r9_o[6]),
    .sel(Ofkiu6),
    .o(Xgshu6));  // ../RTL/cortexm0ds_logic.v(6494)
  AL_MUX u5844 (
    .i0(Sokiu6),
    .i1(vis_r3_o[6]),
    .sel(Pckiu6),
    .o(Qgshu6));  // ../RTL/cortexm0ds_logic.v(6495)
  AL_MUX u5845 (
    .i0(Sokiu6),
    .i1(vis_r2_o[6]),
    .sel(Ickiu6),
    .o(Jgshu6));  // ../RTL/cortexm0ds_logic.v(6496)
  AL_MUX u5846 (
    .i0(Sokiu6),
    .i1(vis_r1_o[6]),
    .sel(Mx8iu6),
    .o(Cgshu6));  // ../RTL/cortexm0ds_logic.v(6497)
  AL_MUX u5847 (
    .i0(Sokiu6),
    .i1(vis_r0_o[6]),
    .sel(Lf8iu6),
    .o(Vfshu6));  // ../RTL/cortexm0ds_logic.v(6498)
  or u5848 (Sokiu6, Pqkiu6, Wqkiu6);  // ../RTL/cortexm0ds_logic.v(6499)
  AL_MUX u5849 (
    .i0(Drkiu6),
    .i1(vis_r8_o[7]),
    .sel(Vfkiu6),
    .o(Ofshu6));  // ../RTL/cortexm0ds_logic.v(6500)
  buf u585 (Tzfpw6[5], Y7opw6);  // ../RTL/cortexm0ds_logic.v(2007)
  and u5850 (n1417, Krkiu6, Rrkiu6);  // ../RTL/cortexm0ds_logic.v(6501)
  not u5851 (Hfshu6, n1417);  // ../RTL/cortexm0ds_logic.v(6501)
  and u5852 (Rrkiu6, Yrkiu6, Fskiu6);  // ../RTL/cortexm0ds_logic.v(6502)
  and u5853 (n1418, Jl8iu6, Tugpw6[5]);  // ../RTL/cortexm0ds_logic.v(6503)
  not u5854 (Fskiu6, n1418);  // ../RTL/cortexm0ds_logic.v(6503)
  buf u5855 (vis_r7_o[11], Co7bx6);  // ../RTL/cortexm0ds_logic.v(2654)
  buf u5856 (vis_r7_o[23], Rnvax6);  // ../RTL/cortexm0ds_logic.v(2654)
  and u5857 (n1419, N5fpw6[6], Sdaiu6);  // ../RTL/cortexm0ds_logic.v(6505)
  not u5858 (Tskiu6, n1419);  // ../RTL/cortexm0ds_logic.v(6505)
  and u5859 (Mskiu6, Atkiu6, Htkiu6);  // ../RTL/cortexm0ds_logic.v(6506)
  buf u586 (Tzfpw6[9], Uojbx6);  // ../RTL/cortexm0ds_logic.v(2007)
  or u5860 (Htkiu6, T2iiu6, Jf0iu6);  // ../RTL/cortexm0ds_logic.v(6507)
  and u5861 (n1420, Eafpw6[7], A3iiu6);  // ../RTL/cortexm0ds_logic.v(6508)
  not u5862 (Atkiu6, n1420);  // ../RTL/cortexm0ds_logic.v(6508)
  and u5863 (n1421, vis_pc_o[6], Ok8iu6);  // ../RTL/cortexm0ds_logic.v(6509)
  not u5864 (Yrkiu6, n1421);  // ../RTL/cortexm0ds_logic.v(6509)
  and u5865 (Krkiu6, Otkiu6, Vtkiu6);  // ../RTL/cortexm0ds_logic.v(6510)
  or u5866 (Vtkiu6, Lm8iu6, Cukiu6);  // ../RTL/cortexm0ds_logic.v(6511)
  and u5867 (n1422, Zm8iu6, Gk4iu6);  // ../RTL/cortexm0ds_logic.v(6512)
  not u5868 (Otkiu6, n1422);  // ../RTL/cortexm0ds_logic.v(6512)
  AL_MUX u5869 (
    .i0(vis_psp_o[5]),
    .i1(Drkiu6),
    .sel(Ydkiu6),
    .o(Afshu6));  // ../RTL/cortexm0ds_logic.v(6513)
  buf u587 (Tzfpw6[10], Vrtpw6);  // ../RTL/cortexm0ds_logic.v(2007)
  AL_MUX u5870 (
    .i0(vis_msp_o[5]),
    .i1(Drkiu6),
    .sel(Fekiu6),
    .o(Teshu6));  // ../RTL/cortexm0ds_logic.v(6514)
  AL_MUX u5871 (
    .i0(Drkiu6),
    .i1(vis_r14_o[7]),
    .sel(Mekiu6),
    .o(Meshu6));  // ../RTL/cortexm0ds_logic.v(6515)
  AL_MUX u5872 (
    .i0(Drkiu6),
    .i1(vis_r12_o[7]),
    .sel(Tekiu6),
    .o(Feshu6));  // ../RTL/cortexm0ds_logic.v(6516)
  AL_MUX u5873 (
    .i0(Drkiu6),
    .i1(vis_r7_o[7]),
    .sel(Rdkiu6),
    .o(Ydshu6));  // ../RTL/cortexm0ds_logic.v(6517)
  AL_MUX u5874 (
    .i0(Drkiu6),
    .i1(vis_r6_o[7]),
    .sel(Kdkiu6),
    .o(Rdshu6));  // ../RTL/cortexm0ds_logic.v(6518)
  AL_MUX u5875 (
    .i0(Drkiu6),
    .i1(vis_r5_o[7]),
    .sel(Ddkiu6),
    .o(Kdshu6));  // ../RTL/cortexm0ds_logic.v(6519)
  AL_MUX u5876 (
    .i0(Drkiu6),
    .i1(vis_r4_o[7]),
    .sel(Wckiu6),
    .o(Ddshu6));  // ../RTL/cortexm0ds_logic.v(6520)
  AL_MUX u5877 (
    .i0(Drkiu6),
    .i1(vis_r11_o[7]),
    .sel(Afkiu6),
    .o(Wcshu6));  // ../RTL/cortexm0ds_logic.v(6521)
  AL_MUX u5878 (
    .i0(Drkiu6),
    .i1(vis_r10_o[7]),
    .sel(Hfkiu6),
    .o(Pcshu6));  // ../RTL/cortexm0ds_logic.v(6522)
  AL_MUX u5879 (
    .i0(Drkiu6),
    .i1(vis_r9_o[7]),
    .sel(Ofkiu6),
    .o(Icshu6));  // ../RTL/cortexm0ds_logic.v(6523)
  buf u588 (Tzfpw6[11], Pt7ax6);  // ../RTL/cortexm0ds_logic.v(2007)
  AL_MUX u5880 (
    .i0(Drkiu6),
    .i1(vis_r3_o[7]),
    .sel(Pckiu6),
    .o(Bcshu6));  // ../RTL/cortexm0ds_logic.v(6524)
  AL_MUX u5881 (
    .i0(Drkiu6),
    .i1(vis_r2_o[7]),
    .sel(Ickiu6),
    .o(Ubshu6));  // ../RTL/cortexm0ds_logic.v(6525)
  AL_MUX u5882 (
    .i0(Drkiu6),
    .i1(vis_r1_o[7]),
    .sel(Mx8iu6),
    .o(Nbshu6));  // ../RTL/cortexm0ds_logic.v(6526)
  AL_MUX u5883 (
    .i0(Drkiu6),
    .i1(vis_r0_o[7]),
    .sel(Lf8iu6),
    .o(Gbshu6));  // ../RTL/cortexm0ds_logic.v(6527)
  or u5884 (Drkiu6, Jukiu6, Qukiu6);  // ../RTL/cortexm0ds_logic.v(6528)
  AL_MUX u5885 (
    .i0(Vx9iu6),
    .i1(vis_r8_o[23]),
    .sel(Vfkiu6),
    .o(Zashu6));  // ../RTL/cortexm0ds_logic.v(6529)
  and u5886 (n1423, Xukiu6, Evkiu6);  // ../RTL/cortexm0ds_logic.v(6530)
  not u5887 (Vx9iu6, n1423);  // ../RTL/cortexm0ds_logic.v(6530)
  and u5888 (Xukiu6, Lvkiu6, Svkiu6);  // ../RTL/cortexm0ds_logic.v(6531)
  AL_MUX u5889 (
    .i0(Zvkiu6),
    .i1(vis_r8_o[24]),
    .sel(Vfkiu6),
    .o(Sashu6));  // ../RTL/cortexm0ds_logic.v(6532)
  buf u589 (Tzfpw6[12], V0jpw6);  // ../RTL/cortexm0ds_logic.v(2007)
  and u5890 (n1424, Gwkiu6, Nwkiu6);  // ../RTL/cortexm0ds_logic.v(6533)
  not u5891 (Lashu6, n1424);  // ../RTL/cortexm0ds_logic.v(6533)
  and u5892 (Nwkiu6, Uwkiu6, Bxkiu6);  // ../RTL/cortexm0ds_logic.v(6534)
  and u5893 (n1425, vis_pc_o[23], Ok8iu6);  // ../RTL/cortexm0ds_logic.v(6535)
  not u5894 (Bxkiu6, n1425);  // ../RTL/cortexm0ds_logic.v(6535)
  and u5895 (Uwkiu6, Ixkiu6, Pxkiu6);  // ../RTL/cortexm0ds_logic.v(6536)
  and u5896 (n1426, Jl8iu6, Tzdpw6);  // ../RTL/cortexm0ds_logic.v(6537)
  not u5897 (Pxkiu6, n1426);  // ../RTL/cortexm0ds_logic.v(6537)
  and u5898 (n1427, Ql8iu6, vis_tbit_o);  // ../RTL/cortexm0ds_logic.v(6538)
  not u5899 (Ixkiu6, n1427);  // ../RTL/cortexm0ds_logic.v(6538)
  buf u59 (vis_r8_o[5], S5kpw6);  // ../RTL/cortexm0ds_logic.v(2579)
  buf u590 (Tzfpw6[13], T9kpw6);  // ../RTL/cortexm0ds_logic.v(2007)
  and u5900 (Gwkiu6, Wxkiu6, Dykiu6);  // ../RTL/cortexm0ds_logic.v(6539)
  or u5901 (Dykiu6, Lm8iu6, Kykiu6);  // ../RTL/cortexm0ds_logic.v(6540)
  or u5902 (Wxkiu6, Hx9iu6, Rykiu6);  // ../RTL/cortexm0ds_logic.v(6541)
  AL_MUX u5903 (
    .i0(vis_psp_o[22]),
    .i1(Zvkiu6),
    .sel(Ydkiu6),
    .o(Eashu6));  // ../RTL/cortexm0ds_logic.v(6542)
  AL_MUX u5904 (
    .i0(vis_msp_o[22]),
    .i1(Zvkiu6),
    .sel(Fekiu6),
    .o(X9shu6));  // ../RTL/cortexm0ds_logic.v(6543)
  AL_MUX u5905 (
    .i0(Zvkiu6),
    .i1(vis_r14_o[24]),
    .sel(Mekiu6),
    .o(Q9shu6));  // ../RTL/cortexm0ds_logic.v(6544)
  AL_MUX u5906 (
    .i0(Zvkiu6),
    .i1(vis_r12_o[24]),
    .sel(Tekiu6),
    .o(J9shu6));  // ../RTL/cortexm0ds_logic.v(6545)
  AL_MUX u5907 (
    .i0(Zvkiu6),
    .i1(vis_r7_o[24]),
    .sel(Rdkiu6),
    .o(C9shu6));  // ../RTL/cortexm0ds_logic.v(6546)
  AL_MUX u5908 (
    .i0(Zvkiu6),
    .i1(vis_r6_o[24]),
    .sel(Kdkiu6),
    .o(V8shu6));  // ../RTL/cortexm0ds_logic.v(6547)
  AL_MUX u5909 (
    .i0(Zvkiu6),
    .i1(vis_r5_o[24]),
    .sel(Ddkiu6),
    .o(O8shu6));  // ../RTL/cortexm0ds_logic.v(6548)
  buf u591 (Tzfpw6[14], Rfxax6);  // ../RTL/cortexm0ds_logic.v(2007)
  AL_MUX u5910 (
    .i0(Zvkiu6),
    .i1(vis_r4_o[24]),
    .sel(Wckiu6),
    .o(H8shu6));  // ../RTL/cortexm0ds_logic.v(6549)
  AL_MUX u5911 (
    .i0(Zvkiu6),
    .i1(vis_r11_o[24]),
    .sel(Afkiu6),
    .o(A8shu6));  // ../RTL/cortexm0ds_logic.v(6550)
  AL_MUX u5912 (
    .i0(Zvkiu6),
    .i1(vis_r10_o[24]),
    .sel(Hfkiu6),
    .o(T7shu6));  // ../RTL/cortexm0ds_logic.v(6551)
  AL_MUX u5913 (
    .i0(Zvkiu6),
    .i1(vis_r9_o[24]),
    .sel(Ofkiu6),
    .o(M7shu6));  // ../RTL/cortexm0ds_logic.v(6552)
  AL_MUX u5914 (
    .i0(Zvkiu6),
    .i1(vis_r3_o[24]),
    .sel(Pckiu6),
    .o(F7shu6));  // ../RTL/cortexm0ds_logic.v(6553)
  AL_MUX u5915 (
    .i0(Zvkiu6),
    .i1(vis_r2_o[24]),
    .sel(Ickiu6),
    .o(Y6shu6));  // ../RTL/cortexm0ds_logic.v(6554)
  AL_MUX u5916 (
    .i0(Zvkiu6),
    .i1(vis_r1_o[24]),
    .sel(Mx8iu6),
    .o(R6shu6));  // ../RTL/cortexm0ds_logic.v(6555)
  AL_MUX u5917 (
    .i0(Zvkiu6),
    .i1(vis_r0_o[24]),
    .sel(Lf8iu6),
    .o(K6shu6));  // ../RTL/cortexm0ds_logic.v(6556)
  or u5918 (Zvkiu6, Nu8iu6, Yykiu6);  // ../RTL/cortexm0ds_logic.v(6557)
  AL_MUX u5919 (
    .i0(Fzkiu6),
    .i1(vis_r8_o[26]),
    .sel(Vfkiu6),
    .o(D6shu6));  // ../RTL/cortexm0ds_logic.v(6558)
  buf u592 (Tzfpw6[16], Wlspw6);  // ../RTL/cortexm0ds_logic.v(2007)
  and u5920 (n1428, Mzkiu6, Tzkiu6);  // ../RTL/cortexm0ds_logic.v(6559)
  not u5921 (W5shu6, n1428);  // ../RTL/cortexm0ds_logic.v(6559)
  and u5922 (Tzkiu6, A0liu6, H0liu6);  // ../RTL/cortexm0ds_logic.v(6560)
  and u5923 (n1429, Jl8iu6, H0epw6);  // ../RTL/cortexm0ds_logic.v(6561)
  not u5924 (H0liu6, n1429);  // ../RTL/cortexm0ds_logic.v(6561)
  and u5925 (n1430, vis_pc_o[25], Ok8iu6);  // ../RTL/cortexm0ds_logic.v(6562)
  not u5926 (A0liu6, n1430);  // ../RTL/cortexm0ds_logic.v(6562)
  and u5927 (Mzkiu6, O0liu6, V0liu6);  // ../RTL/cortexm0ds_logic.v(6563)
  and u5928 (n1431, W29iu6, Fkfpw6[26]);  // ../RTL/cortexm0ds_logic.v(6564)
  not u5929 (V0liu6, n1431);  // ../RTL/cortexm0ds_logic.v(6564)
  buf u593 (Tzfpw6[17], Amupw6);  // ../RTL/cortexm0ds_logic.v(2007)
  or u5930 (O0liu6, Hx9iu6, C1liu6);  // ../RTL/cortexm0ds_logic.v(6565)
  AL_MUX u5931 (
    .i0(vis_psp_o[24]),
    .i1(Fzkiu6),
    .sel(Ydkiu6),
    .o(P5shu6));  // ../RTL/cortexm0ds_logic.v(6566)
  AL_MUX u5932 (
    .i0(vis_msp_o[24]),
    .i1(Fzkiu6),
    .sel(Fekiu6),
    .o(I5shu6));  // ../RTL/cortexm0ds_logic.v(6567)
  AL_MUX u5933 (
    .i0(Fzkiu6),
    .i1(vis_r14_o[26]),
    .sel(Mekiu6),
    .o(B5shu6));  // ../RTL/cortexm0ds_logic.v(6568)
  AL_MUX u5934 (
    .i0(Fzkiu6),
    .i1(vis_r12_o[26]),
    .sel(Tekiu6),
    .o(U4shu6));  // ../RTL/cortexm0ds_logic.v(6569)
  AL_MUX u5935 (
    .i0(Fzkiu6),
    .i1(vis_r7_o[26]),
    .sel(Rdkiu6),
    .o(N4shu6));  // ../RTL/cortexm0ds_logic.v(6570)
  AL_MUX u5936 (
    .i0(Fzkiu6),
    .i1(vis_r6_o[26]),
    .sel(Kdkiu6),
    .o(G4shu6));  // ../RTL/cortexm0ds_logic.v(6571)
  AL_MUX u5937 (
    .i0(Fzkiu6),
    .i1(vis_r5_o[26]),
    .sel(Ddkiu6),
    .o(Z3shu6));  // ../RTL/cortexm0ds_logic.v(6572)
  AL_MUX u5938 (
    .i0(Fzkiu6),
    .i1(vis_r4_o[26]),
    .sel(Wckiu6),
    .o(S3shu6));  // ../RTL/cortexm0ds_logic.v(6573)
  AL_MUX u5939 (
    .i0(Fzkiu6),
    .i1(vis_r11_o[26]),
    .sel(Afkiu6),
    .o(L3shu6));  // ../RTL/cortexm0ds_logic.v(6574)
  buf u594 (Tzfpw6[18], N0xpw6);  // ../RTL/cortexm0ds_logic.v(2007)
  AL_MUX u5940 (
    .i0(Fzkiu6),
    .i1(vis_r10_o[26]),
    .sel(Hfkiu6),
    .o(E3shu6));  // ../RTL/cortexm0ds_logic.v(6575)
  AL_MUX u5941 (
    .i0(Fzkiu6),
    .i1(vis_r9_o[26]),
    .sel(Ofkiu6),
    .o(X2shu6));  // ../RTL/cortexm0ds_logic.v(6576)
  AL_MUX u5942 (
    .i0(Fzkiu6),
    .i1(vis_r3_o[26]),
    .sel(Pckiu6),
    .o(Q2shu6));  // ../RTL/cortexm0ds_logic.v(6577)
  AL_MUX u5943 (
    .i0(Fzkiu6),
    .i1(vis_r2_o[26]),
    .sel(Ickiu6),
    .o(J2shu6));  // ../RTL/cortexm0ds_logic.v(6578)
  AL_MUX u5944 (
    .i0(Fzkiu6),
    .i1(vis_r1_o[26]),
    .sel(Mx8iu6),
    .o(C2shu6));  // ../RTL/cortexm0ds_logic.v(6579)
  AL_MUX u5945 (
    .i0(Fzkiu6),
    .i1(vis_r0_o[26]),
    .sel(Lf8iu6),
    .o(V1shu6));  // ../RTL/cortexm0ds_logic.v(6580)
  or u5946 (Fzkiu6, J1liu6, Q1liu6);  // ../RTL/cortexm0ds_logic.v(6581)
  AL_MUX u5947 (
    .i0(X1liu6),
    .i1(vis_r8_o[27]),
    .sel(Vfkiu6),
    .o(O1shu6));  // ../RTL/cortexm0ds_logic.v(6582)
  and u5948 (n1432, E2liu6, L2liu6);  // ../RTL/cortexm0ds_logic.v(6583)
  not u5949 (H1shu6, n1432);  // ../RTL/cortexm0ds_logic.v(6583)
  buf u595 (Tzfpw6[20], Z8jpw6);  // ../RTL/cortexm0ds_logic.v(2007)
  and u5950 (L2liu6, S2liu6, Z2liu6);  // ../RTL/cortexm0ds_logic.v(6584)
  and u5951 (n1433, Jl8iu6, O0epw6);  // ../RTL/cortexm0ds_logic.v(6585)
  not u5952 (Z2liu6, n1433);  // ../RTL/cortexm0ds_logic.v(6585)
  and u5953 (n1434, vis_pc_o[26], Ok8iu6);  // ../RTL/cortexm0ds_logic.v(6586)
  not u5954 (S2liu6, n1434);  // ../RTL/cortexm0ds_logic.v(6586)
  and u5955 (E2liu6, G3liu6, N3liu6);  // ../RTL/cortexm0ds_logic.v(6587)
  and u5956 (n1435, W29iu6, Fkfpw6[27]);  // ../RTL/cortexm0ds_logic.v(6588)
  not u5957 (N3liu6, n1435);  // ../RTL/cortexm0ds_logic.v(6588)
  or u5958 (G3liu6, Hx9iu6, U3liu6);  // ../RTL/cortexm0ds_logic.v(6589)
  AL_MUX u5959 (
    .i0(vis_psp_o[25]),
    .i1(X1liu6),
    .sel(Ydkiu6),
    .o(A1shu6));  // ../RTL/cortexm0ds_logic.v(6590)
  buf u596 (Tzfpw6[22], F9gbx6);  // ../RTL/cortexm0ds_logic.v(2007)
  AL_MUX u5960 (
    .i0(vis_msp_o[25]),
    .i1(X1liu6),
    .sel(Fekiu6),
    .o(T0shu6));  // ../RTL/cortexm0ds_logic.v(6591)
  AL_MUX u5961 (
    .i0(X1liu6),
    .i1(vis_r14_o[27]),
    .sel(Mekiu6),
    .o(M0shu6));  // ../RTL/cortexm0ds_logic.v(6592)
  AL_MUX u5962 (
    .i0(X1liu6),
    .i1(vis_r12_o[27]),
    .sel(Tekiu6),
    .o(F0shu6));  // ../RTL/cortexm0ds_logic.v(6593)
  AL_MUX u5963 (
    .i0(X1liu6),
    .i1(vis_r7_o[27]),
    .sel(Rdkiu6),
    .o(Yzrhu6));  // ../RTL/cortexm0ds_logic.v(6594)
  AL_MUX u5964 (
    .i0(X1liu6),
    .i1(vis_r6_o[27]),
    .sel(Kdkiu6),
    .o(Rzrhu6));  // ../RTL/cortexm0ds_logic.v(6595)
  AL_MUX u5965 (
    .i0(X1liu6),
    .i1(vis_r5_o[27]),
    .sel(Ddkiu6),
    .o(Kzrhu6));  // ../RTL/cortexm0ds_logic.v(6596)
  AL_MUX u5966 (
    .i0(X1liu6),
    .i1(vis_r4_o[27]),
    .sel(Wckiu6),
    .o(Dzrhu6));  // ../RTL/cortexm0ds_logic.v(6597)
  AL_MUX u5967 (
    .i0(X1liu6),
    .i1(vis_r11_o[27]),
    .sel(Afkiu6),
    .o(Wyrhu6));  // ../RTL/cortexm0ds_logic.v(6598)
  AL_MUX u5968 (
    .i0(X1liu6),
    .i1(vis_r10_o[27]),
    .sel(Hfkiu6),
    .o(Pyrhu6));  // ../RTL/cortexm0ds_logic.v(6599)
  AL_MUX u5969 (
    .i0(X1liu6),
    .i1(vis_r9_o[27]),
    .sel(Ofkiu6),
    .o(Iyrhu6));  // ../RTL/cortexm0ds_logic.v(6600)
  buf u597 (vis_msp_o[0], Zgzpw6);  // ../RTL/cortexm0ds_logic.v(2097)
  AL_MUX u5970 (
    .i0(X1liu6),
    .i1(vis_r3_o[27]),
    .sel(Pckiu6),
    .o(Byrhu6));  // ../RTL/cortexm0ds_logic.v(6601)
  AL_MUX u5971 (
    .i0(X1liu6),
    .i1(vis_r2_o[27]),
    .sel(Ickiu6),
    .o(Uxrhu6));  // ../RTL/cortexm0ds_logic.v(6602)
  AL_MUX u5972 (
    .i0(X1liu6),
    .i1(vis_r1_o[27]),
    .sel(Mx8iu6),
    .o(Nxrhu6));  // ../RTL/cortexm0ds_logic.v(6603)
  AL_MUX u5973 (
    .i0(X1liu6),
    .i1(vis_r0_o[27]),
    .sel(Lf8iu6),
    .o(Gxrhu6));  // ../RTL/cortexm0ds_logic.v(6604)
  or u5974 (X1liu6, B4liu6, I4liu6);  // ../RTL/cortexm0ds_logic.v(6605)
  AL_MUX u5975 (
    .i0(P4liu6),
    .i1(vis_r8_o[29]),
    .sel(Vfkiu6),
    .o(Zwrhu6));  // ../RTL/cortexm0ds_logic.v(6606)
  AL_MUX u5976 (
    .i0(vis_psp_o[27]),
    .i1(P4liu6),
    .sel(Ydkiu6),
    .o(Swrhu6));  // ../RTL/cortexm0ds_logic.v(6607)
  AL_MUX u5977 (
    .i0(vis_msp_o[27]),
    .i1(P4liu6),
    .sel(Fekiu6),
    .o(Lwrhu6));  // ../RTL/cortexm0ds_logic.v(6608)
  AL_MUX u5978 (
    .i0(P4liu6),
    .i1(vis_r14_o[29]),
    .sel(Mekiu6),
    .o(Ewrhu6));  // ../RTL/cortexm0ds_logic.v(6609)
  AL_MUX u5979 (
    .i0(P4liu6),
    .i1(vis_r12_o[29]),
    .sel(Tekiu6),
    .o(Xvrhu6));  // ../RTL/cortexm0ds_logic.v(6610)
  buf u598 (vis_r7_o[0], Rtvax6);  // ../RTL/cortexm0ds_logic.v(2654)
  AL_MUX u5980 (
    .i0(P4liu6),
    .i1(vis_r7_o[29]),
    .sel(Rdkiu6),
    .o(Qvrhu6));  // ../RTL/cortexm0ds_logic.v(6611)
  AL_MUX u5981 (
    .i0(P4liu6),
    .i1(vis_r6_o[29]),
    .sel(Kdkiu6),
    .o(Jvrhu6));  // ../RTL/cortexm0ds_logic.v(6612)
  AL_MUX u5982 (
    .i0(P4liu6),
    .i1(vis_r5_o[29]),
    .sel(Ddkiu6),
    .o(Cvrhu6));  // ../RTL/cortexm0ds_logic.v(6613)
  AL_MUX u5983 (
    .i0(P4liu6),
    .i1(vis_r4_o[29]),
    .sel(Wckiu6),
    .o(Vurhu6));  // ../RTL/cortexm0ds_logic.v(6614)
  AL_MUX u5984 (
    .i0(P4liu6),
    .i1(vis_r11_o[29]),
    .sel(Afkiu6),
    .o(Ourhu6));  // ../RTL/cortexm0ds_logic.v(6615)
  AL_MUX u5985 (
    .i0(P4liu6),
    .i1(vis_r10_o[29]),
    .sel(Hfkiu6),
    .o(Hurhu6));  // ../RTL/cortexm0ds_logic.v(6616)
  AL_MUX u5986 (
    .i0(P4liu6),
    .i1(vis_r9_o[29]),
    .sel(Ofkiu6),
    .o(Aurhu6));  // ../RTL/cortexm0ds_logic.v(6617)
  AL_MUX u5987 (
    .i0(P4liu6),
    .i1(vis_r3_o[29]),
    .sel(Pckiu6),
    .o(Ttrhu6));  // ../RTL/cortexm0ds_logic.v(6618)
  AL_MUX u5988 (
    .i0(P4liu6),
    .i1(vis_r2_o[29]),
    .sel(Ickiu6),
    .o(Mtrhu6));  // ../RTL/cortexm0ds_logic.v(6619)
  AL_MUX u5989 (
    .i0(P4liu6),
    .i1(vis_r1_o[29]),
    .sel(Mx8iu6),
    .o(Ftrhu6));  // ../RTL/cortexm0ds_logic.v(6620)
  buf u599 (vis_r3_o[0], V1yax6);  // ../RTL/cortexm0ds_logic.v(2694)
  AL_MUX u5990 (
    .i0(P4liu6),
    .i1(vis_r0_o[29]),
    .sel(Lf8iu6),
    .o(Ysrhu6));  // ../RTL/cortexm0ds_logic.v(6621)
  or u5991 (P4liu6, Fj8iu6, W4liu6);  // ../RTL/cortexm0ds_logic.v(6622)
  AL_MUX u5992 (
    .i0(K39iu6),
    .i1(vis_r8_o[30]),
    .sel(Vfkiu6),
    .o(Rsrhu6));  // ../RTL/cortexm0ds_logic.v(6623)
  and u5993 (n1436, D5liu6, K5liu6);  // ../RTL/cortexm0ds_logic.v(6624)
  not u5994 (K39iu6, n1436);  // ../RTL/cortexm0ds_logic.v(6624)
  AL_MUX u5995 (
    .i0(vis_apsr_o[2]),
    .i1(R5liu6),
    .sel(Y5liu6),
    .o(Ksrhu6));  // ../RTL/cortexm0ds_logic.v(6625)
  and u5996 (n1437, F6liu6, M6liu6);  // ../RTL/cortexm0ds_logic.v(6626)
  not u5997 (R5liu6, n1437);  // ../RTL/cortexm0ds_logic.v(6626)
  and u5998 (n1438, Ph8iu6, T6liu6);  // ../RTL/cortexm0ds_logic.v(6627)
  not u5999 (M6liu6, n1438);  // ../RTL/cortexm0ds_logic.v(6627)
  buf u6 (HSIZE[2], 1'b0);  // ../RTL/cortexm0ds_logic.v(1729)
  buf u60 (Gtgpw6[13], P4cax6);  // ../RTL/cortexm0ds_logic.v(2375)
  buf u600 (vis_r0_o[21], E5npw6);  // ../RTL/cortexm0ds_logic.v(1875)
  and u6000 (F6liu6, A7liu6, H7liu6);  // ../RTL/cortexm0ds_logic.v(6628)
  or u6001 (H7liu6, O7liu6, V7liu6);  // ../RTL/cortexm0ds_logic.v(6629)
  or u6002 (A7liu6, Cs8iu6, D5liu6);  // ../RTL/cortexm0ds_logic.v(6630)
  and u6003 (n1439, C8liu6, J8liu6);  // ../RTL/cortexm0ds_logic.v(6631)
  not u6004 (Dsrhu6, n1439);  // ../RTL/cortexm0ds_logic.v(6631)
  and u6005 (J8liu6, Q8liu6, X8liu6);  // ../RTL/cortexm0ds_logic.v(6632)
  and u6006 (n1440, Ok8iu6, vis_pc_o[29]);  // ../RTL/cortexm0ds_logic.v(6633)
  not u6007 (X8liu6, n1440);  // ../RTL/cortexm0ds_logic.v(6633)
  and u6008 (Q8liu6, E9liu6, L9liu6);  // ../RTL/cortexm0ds_logic.v(6634)
  and u6009 (n1441, Jl8iu6, Rx0iu6);  // ../RTL/cortexm0ds_logic.v(6635)
  buf u601 (vis_r0_o[19], Jjvpw6);  // ../RTL/cortexm0ds_logic.v(1875)
  not u6010 (L9liu6, n1441);  // ../RTL/cortexm0ds_logic.v(6635)
  and u6011 (n1442, vis_apsr_o[2], Ql8iu6);  // ../RTL/cortexm0ds_logic.v(6636)
  not u6012 (E9liu6, n1442);  // ../RTL/cortexm0ds_logic.v(6636)
  and u6013 (C8liu6, S9liu6, Z9liu6);  // ../RTL/cortexm0ds_logic.v(6637)
  or u6014 (Z9liu6, Lm8iu6, Galiu6);  // ../RTL/cortexm0ds_logic.v(6638)
  or u6015 (S9liu6, Hx9iu6, Naliu6);  // ../RTL/cortexm0ds_logic.v(6639)
  AL_MUX u6016 (
    .i0(D39iu6),
    .i1(vis_r8_o[31]),
    .sel(Vfkiu6),
    .o(Wrrhu6));  // ../RTL/cortexm0ds_logic.v(6640)
  and u6017 (n1443, Ualiu6, Bbliu6);  // ../RTL/cortexm0ds_logic.v(6641)
  not u6018 (D39iu6, n1443);  // ../RTL/cortexm0ds_logic.v(6641)
  AL_MUX u6019 (
    .i0(Tx8iu6),
    .i1(vis_r8_o[0]),
    .sel(Vfkiu6),
    .o(Prrhu6));  // ../RTL/cortexm0ds_logic.v(6642)
  buf u602 (D7fpw6[15], U9ypw6);  // ../RTL/cortexm0ds_logic.v(2074)
  and u6020 (n1444, Zt8iu6, Ibliu6);  // ../RTL/cortexm0ds_logic.v(6643)
  not u6021 (Tx8iu6, n1444);  // ../RTL/cortexm0ds_logic.v(6643)
  and u6022 (Zt8iu6, Pbliu6, Wbliu6);  // ../RTL/cortexm0ds_logic.v(6644)
  and u6023 (Wbliu6, Dcliu6, Kcliu6);  // ../RTL/cortexm0ds_logic.v(6645)
  or u6024 (Kcliu6, Rcliu6, Ycliu6);  // ../RTL/cortexm0ds_logic.v(6646)
  and u6025 (Dcliu6, Fdliu6, Mdliu6);  // ../RTL/cortexm0ds_logic.v(6647)
  and u6026 (n1445, Tdliu6, Aeliu6);  // ../RTL/cortexm0ds_logic.v(6648)
  not u6027 (Fdliu6, n1445);  // ../RTL/cortexm0ds_logic.v(6648)
  and u6028 (Pbliu6, Heliu6, Oeliu6);  // ../RTL/cortexm0ds_logic.v(6649)
  or u6029 (Oeliu6, Veliu6, Cfliu6);  // ../RTL/cortexm0ds_logic.v(6650)
  buf u603 (D7fpw6[8], P0kax6);  // ../RTL/cortexm0ds_logic.v(2074)
  and u6030 (n1446, Jfliu6, Qfliu6);  // ../RTL/cortexm0ds_logic.v(6651)
  not u6031 (Heliu6, n1446);  // ../RTL/cortexm0ds_logic.v(6651)
  and u6032 (n1447, Xfliu6, Egliu6);  // ../RTL/cortexm0ds_logic.v(6652)
  not u6033 (Irrhu6, n1447);  // ../RTL/cortexm0ds_logic.v(6652)
  and u6034 (Egliu6, Lgliu6, Sgliu6);  // ../RTL/cortexm0ds_logic.v(6653)
  and u6035 (n1448, Ok8iu6, vis_pc_o[0]);  // ../RTL/cortexm0ds_logic.v(6654)
  not u6036 (Sgliu6, n1448);  // ../RTL/cortexm0ds_logic.v(6654)
  and u6037 (Lgliu6, Zgliu6, Ghliu6);  // ../RTL/cortexm0ds_logic.v(6655)
  and u6038 (n1449, Nhliu6, Uhliu6);  // ../RTL/cortexm0ds_logic.v(6656)
  not u6039 (Ghliu6, n1449);  // ../RTL/cortexm0ds_logic.v(6656)
  buf u604 (vis_r9_o[0], Qukax6);  // ../RTL/cortexm0ds_logic.v(1898)
  and u6040 (Uhliu6, Biliu6, Iiliu6);  // ../RTL/cortexm0ds_logic.v(6657)
  and u6041 (Nhliu6, Jl8iu6, Piliu6);  // ../RTL/cortexm0ds_logic.v(6658)
  or u6042 (Piliu6, Wiliu6, Oviiu6);  // ../RTL/cortexm0ds_logic.v(6659)
  and u6043 (n1450, Ql8iu6, vis_ipsr_o[1]);  // ../RTL/cortexm0ds_logic.v(6660)
  not u6044 (Zgliu6, n1450);  // ../RTL/cortexm0ds_logic.v(6660)
  and u6045 (Xfliu6, Djliu6, Kjliu6);  // ../RTL/cortexm0ds_logic.v(6661)
  or u6046 (Kjliu6, Lm8iu6, Rjliu6);  // ../RTL/cortexm0ds_logic.v(6662)
  or u6047 (Djliu6, Hx9iu6, A34iu6);  // ../RTL/cortexm0ds_logic.v(6663)
  AL_MUX u6048 (
    .i0(vis_control_o),
    .i1(Yjliu6),
    .sel(Fkliu6),
    .o(Brrhu6));  // ../RTL/cortexm0ds_logic.v(6664)
  and u6049 (Fkliu6, HREADY, Mkliu6);  // ../RTL/cortexm0ds_logic.v(6665)
  buf u605 (vis_r0_o[23], Gv6ax6);  // ../RTL/cortexm0ds_logic.v(1875)
  and u6050 (n1451, Tkliu6, Alliu6);  // ../RTL/cortexm0ds_logic.v(6666)
  not u6051 (Mkliu6, n1451);  // ../RTL/cortexm0ds_logic.v(6666)
  and u6052 (n1452, Hlliu6, Olliu6);  // ../RTL/cortexm0ds_logic.v(6667)
  not u6053 (Alliu6, n1452);  // ../RTL/cortexm0ds_logic.v(6667)
  and u6054 (n1453, Vlliu6, Cmliu6);  // ../RTL/cortexm0ds_logic.v(6668)
  not u6055 (Olliu6, n1453);  // ../RTL/cortexm0ds_logic.v(6668)
  and u6056 (n1454, Jmliu6, S8fpw6[2]);  // ../RTL/cortexm0ds_logic.v(6669)
  not u6057 (Cmliu6, n1454);  // ../RTL/cortexm0ds_logic.v(6669)
  and u6058 (Jmliu6, S8fpw6[4], Qmliu6);  // ../RTL/cortexm0ds_logic.v(6670)
  or u6059 (n1455, Clfiu6, Xmliu6);  // ../RTL/cortexm0ds_logic.v(6671)
  buf u606 (vis_r0_o[20], E7npw6);  // ../RTL/cortexm0ds_logic.v(1875)
  not u6060 (Tkliu6, n1455);  // ../RTL/cortexm0ds_logic.v(6671)
  and u6061 (n1456, Enliu6, Lnliu6);  // ../RTL/cortexm0ds_logic.v(6672)
  not u6062 (Yjliu6, n1456);  // ../RTL/cortexm0ds_logic.v(6672)
  and u6063 (n1457, Snliu6, Qmliu6);  // ../RTL/cortexm0ds_logic.v(6673)
  not u6064 (Lnliu6, n1457);  // ../RTL/cortexm0ds_logic.v(6673)
  AL_MUX u6065 (
    .i0(Znliu6),
    .i1(Goliu6),
    .sel(Wofiu6),
    .o(Snliu6));  // ../RTL/cortexm0ds_logic.v(6674)
  or u6066 (Enliu6, Quzhu6, Noliu6);  // ../RTL/cortexm0ds_logic.v(6675)
  AL_MUX u6067 (
    .i0(Uoliu6),
    .i1(vis_r14_o[1]),
    .sel(Mekiu6),
    .o(Uqrhu6));  // ../RTL/cortexm0ds_logic.v(6676)
  AL_MUX u6068 (
    .i0(Uoliu6),
    .i1(vis_r12_o[1]),
    .sel(Tekiu6),
    .o(Nqrhu6));  // ../RTL/cortexm0ds_logic.v(6677)
  AL_MUX u6069 (
    .i0(Uoliu6),
    .i1(vis_r7_o[1]),
    .sel(Rdkiu6),
    .o(Gqrhu6));  // ../RTL/cortexm0ds_logic.v(6678)
  buf u607 (vis_r0_o[18], P2xpw6);  // ../RTL/cortexm0ds_logic.v(1875)
  AL_MUX u6070 (
    .i0(Uoliu6),
    .i1(vis_r6_o[1]),
    .sel(Kdkiu6),
    .o(Zprhu6));  // ../RTL/cortexm0ds_logic.v(6679)
  AL_MUX u6071 (
    .i0(Uoliu6),
    .i1(vis_r5_o[1]),
    .sel(Ddkiu6),
    .o(Sprhu6));  // ../RTL/cortexm0ds_logic.v(6680)
  AL_MUX u6072 (
    .i0(Uoliu6),
    .i1(vis_r4_o[1]),
    .sel(Wckiu6),
    .o(Lprhu6));  // ../RTL/cortexm0ds_logic.v(6681)
  AL_MUX u6073 (
    .i0(Uoliu6),
    .i1(vis_r11_o[1]),
    .sel(Afkiu6),
    .o(Eprhu6));  // ../RTL/cortexm0ds_logic.v(6682)
  AL_MUX u6074 (
    .i0(Uoliu6),
    .i1(vis_r10_o[1]),
    .sel(Hfkiu6),
    .o(Xorhu6));  // ../RTL/cortexm0ds_logic.v(6683)
  AL_MUX u6075 (
    .i0(Uoliu6),
    .i1(vis_r9_o[1]),
    .sel(Ofkiu6),
    .o(Qorhu6));  // ../RTL/cortexm0ds_logic.v(6684)
  AL_MUX u6076 (
    .i0(Uoliu6),
    .i1(vis_r8_o[1]),
    .sel(Vfkiu6),
    .o(Jorhu6));  // ../RTL/cortexm0ds_logic.v(6685)
  AL_MUX u6077 (
    .i0(Uoliu6),
    .i1(vis_r3_o[1]),
    .sel(Pckiu6),
    .o(Corhu6));  // ../RTL/cortexm0ds_logic.v(6686)
  AL_MUX u6078 (
    .i0(Uoliu6),
    .i1(vis_r2_o[1]),
    .sel(Ickiu6),
    .o(Vnrhu6));  // ../RTL/cortexm0ds_logic.v(6687)
  AL_MUX u6079 (
    .i0(Uoliu6),
    .i1(vis_r1_o[1]),
    .sel(Mx8iu6),
    .o(Onrhu6));  // ../RTL/cortexm0ds_logic.v(6688)
  buf u608 (vis_r0_o[17], Y7upw6);  // ../RTL/cortexm0ds_logic.v(1875)
  AL_MUX u6080 (
    .i0(Uoliu6),
    .i1(vis_r0_o[1]),
    .sel(Lf8iu6),
    .o(Hnrhu6));  // ../RTL/cortexm0ds_logic.v(6689)
  and u6081 (n1458, Njciu6, Bpliu6);  // ../RTL/cortexm0ds_logic.v(6690)
  not u6082 (Uoliu6, n1458);  // ../RTL/cortexm0ds_logic.v(6690)
  and u6083 (n1459, Ipliu6, Ppliu6);  // ../RTL/cortexm0ds_logic.v(6691)
  not u6084 (Anrhu6, n1459);  // ../RTL/cortexm0ds_logic.v(6691)
  and u6085 (Ppliu6, Wpliu6, Dqliu6);  // ../RTL/cortexm0ds_logic.v(6692)
  and u6086 (n1460, vis_pc_o[24], Ok8iu6);  // ../RTL/cortexm0ds_logic.v(6693)
  not u6087 (Dqliu6, n1460);  // ../RTL/cortexm0ds_logic.v(6693)
  and u6088 (Wpliu6, Kqliu6, Rqliu6);  // ../RTL/cortexm0ds_logic.v(6694)
  and u6089 (n1461, vis_control_o, B29iu6);  // ../RTL/cortexm0ds_logic.v(6695)
  buf u609 (vis_r0_o[16], C5wpw6);  // ../RTL/cortexm0ds_logic.v(1875)
  not u6090 (Rqliu6, n1461);  // ../RTL/cortexm0ds_logic.v(6695)
  and u6091 (B29iu6, Yqliu6, Frliu6);  // ../RTL/cortexm0ds_logic.v(6696)
  or u6092 (n1462, U19iu6, W29iu6);  // ../RTL/cortexm0ds_logic.v(6697)
  not u6093 (Yqliu6, n1462);  // ../RTL/cortexm0ds_logic.v(6697)
  and u6094 (n1463, Jl8iu6, A0epw6);  // ../RTL/cortexm0ds_logic.v(6698)
  not u6095 (Kqliu6, n1463);  // ../RTL/cortexm0ds_logic.v(6698)
  and u6096 (Ipliu6, Mrliu6, Trliu6);  // ../RTL/cortexm0ds_logic.v(6699)
  and u6097 (n1464, W29iu6, Fkfpw6[25]);  // ../RTL/cortexm0ds_logic.v(6700)
  not u6098 (Trliu6, n1464);  // ../RTL/cortexm0ds_logic.v(6700)
  or u6099 (Mrliu6, Hx9iu6, Asliu6);  // ../RTL/cortexm0ds_logic.v(6701)
  buf u61 (vis_tbit_o, Pzkpw6);  // ../RTL/cortexm0ds_logic.v(1827)
  buf u610 (D7fpw6[14], Dxvpw6);  // ../RTL/cortexm0ds_logic.v(2074)
  AL_MUX u6100 (
    .i0(vis_psp_o[23]),
    .i1(Hsliu6),
    .sel(Ydkiu6),
    .o(Tmrhu6));  // ../RTL/cortexm0ds_logic.v(6702)
  AL_MUX u6101 (
    .i0(vis_msp_o[23]),
    .i1(Hsliu6),
    .sel(Fekiu6),
    .o(Mmrhu6));  // ../RTL/cortexm0ds_logic.v(6703)
  AL_MUX u6102 (
    .i0(Hsliu6),
    .i1(vis_r14_o[25]),
    .sel(Mekiu6),
    .o(Fmrhu6));  // ../RTL/cortexm0ds_logic.v(6704)
  AL_MUX u6103 (
    .i0(Hsliu6),
    .i1(vis_r12_o[25]),
    .sel(Tekiu6),
    .o(Ylrhu6));  // ../RTL/cortexm0ds_logic.v(6705)
  AL_MUX u6104 (
    .i0(Hsliu6),
    .i1(vis_r7_o[25]),
    .sel(Rdkiu6),
    .o(Rlrhu6));  // ../RTL/cortexm0ds_logic.v(6706)
  AL_MUX u6105 (
    .i0(Hsliu6),
    .i1(vis_r6_o[25]),
    .sel(Kdkiu6),
    .o(Klrhu6));  // ../RTL/cortexm0ds_logic.v(6707)
  AL_MUX u6106 (
    .i0(Hsliu6),
    .i1(vis_r5_o[25]),
    .sel(Ddkiu6),
    .o(Dlrhu6));  // ../RTL/cortexm0ds_logic.v(6708)
  AL_MUX u6107 (
    .i0(Hsliu6),
    .i1(vis_r4_o[25]),
    .sel(Wckiu6),
    .o(Wkrhu6));  // ../RTL/cortexm0ds_logic.v(6709)
  AL_MUX u6108 (
    .i0(Hsliu6),
    .i1(vis_r11_o[25]),
    .sel(Afkiu6),
    .o(Pkrhu6));  // ../RTL/cortexm0ds_logic.v(6710)
  AL_MUX u6109 (
    .i0(Hsliu6),
    .i1(vis_r10_o[25]),
    .sel(Hfkiu6),
    .o(Ikrhu6));  // ../RTL/cortexm0ds_logic.v(6711)
  buf u611 (D7fpw6[12], Skjax6);  // ../RTL/cortexm0ds_logic.v(2074)
  AL_MUX u6110 (
    .i0(Hsliu6),
    .i1(vis_r9_o[25]),
    .sel(Ofkiu6),
    .o(Bkrhu6));  // ../RTL/cortexm0ds_logic.v(6712)
  AL_MUX u6111 (
    .i0(Hsliu6),
    .i1(vis_r8_o[25]),
    .sel(Vfkiu6),
    .o(Ujrhu6));  // ../RTL/cortexm0ds_logic.v(6713)
  AL_MUX u6112 (
    .i0(Hsliu6),
    .i1(vis_r3_o[25]),
    .sel(Pckiu6),
    .o(Njrhu6));  // ../RTL/cortexm0ds_logic.v(6714)
  AL_MUX u6113 (
    .i0(Hsliu6),
    .i1(vis_r2_o[25]),
    .sel(Ickiu6),
    .o(Gjrhu6));  // ../RTL/cortexm0ds_logic.v(6715)
  AL_MUX u6114 (
    .i0(Hsliu6),
    .i1(vis_r1_o[25]),
    .sel(Mx8iu6),
    .o(Zirhu6));  // ../RTL/cortexm0ds_logic.v(6716)
  AL_MUX u6115 (
    .i0(Hsliu6),
    .i1(vis_r0_o[25]),
    .sel(Lf8iu6),
    .o(Sirhu6));  // ../RTL/cortexm0ds_logic.v(6717)
  or u6116 (Hsliu6, Osliu6, Vsliu6);  // ../RTL/cortexm0ds_logic.v(6718)
  AL_MUX u6117 (
    .i0(Iwfpw6[1]),
    .i1(Iiliu6),
    .sel(Hy8iu6),
    .o(Lirhu6));  // ../RTL/cortexm0ds_logic.v(6719)
  or u6118 (n1465, Eh6iu6, L18iu6);  // ../RTL/cortexm0ds_logic.v(6720)
  not u6119 (Hy8iu6, n1465);  // ../RTL/cortexm0ds_logic.v(6720)
  buf u612 (D7fpw6[11], Sojax6);  // ../RTL/cortexm0ds_logic.v(2074)
  and u6120 (n1466, Ctliu6, Jtliu6);  // ../RTL/cortexm0ds_logic.v(6721)
  not u6121 (Eirhu6, n1466);  // ../RTL/cortexm0ds_logic.v(6721)
  and u6122 (Jtliu6, Qtliu6, Xtliu6);  // ../RTL/cortexm0ds_logic.v(6722)
  and u6123 (n1467, Jl8iu6, Fzdpw6);  // ../RTL/cortexm0ds_logic.v(6723)
  not u6124 (Xtliu6, n1467);  // ../RTL/cortexm0ds_logic.v(6723)
  and u6125 (n1468, vis_pc_o[21], Ok8iu6);  // ../RTL/cortexm0ds_logic.v(6724)
  not u6126 (Qtliu6, n1468);  // ../RTL/cortexm0ds_logic.v(6724)
  and u6127 (Ctliu6, Euliu6, Luliu6);  // ../RTL/cortexm0ds_logic.v(6725)
  or u6128 (Luliu6, Lm8iu6, Suliu6);  // ../RTL/cortexm0ds_logic.v(6726)
  and u6129 (n1469, Zm8iu6, P74iu6);  // ../RTL/cortexm0ds_logic.v(6727)
  buf u613 (D7fpw6[9], Rwjax6);  // ../RTL/cortexm0ds_logic.v(2074)
  not u6130 (Euliu6, n1469);  // ../RTL/cortexm0ds_logic.v(6727)
  AL_MUX u6131 (
    .i0(vis_psp_o[20]),
    .i1(Zuliu6),
    .sel(Ydkiu6),
    .o(Xhrhu6));  // ../RTL/cortexm0ds_logic.v(6728)
  AL_MUX u6132 (
    .i0(vis_msp_o[20]),
    .i1(Zuliu6),
    .sel(Fekiu6),
    .o(Qhrhu6));  // ../RTL/cortexm0ds_logic.v(6729)
  AL_MUX u6133 (
    .i0(Zuliu6),
    .i1(vis_r14_o[22]),
    .sel(Mekiu6),
    .o(Jhrhu6));  // ../RTL/cortexm0ds_logic.v(6730)
  AL_MUX u6134 (
    .i0(Zuliu6),
    .i1(vis_r12_o[22]),
    .sel(Tekiu6),
    .o(Chrhu6));  // ../RTL/cortexm0ds_logic.v(6731)
  AL_MUX u6135 (
    .i0(Zuliu6),
    .i1(vis_r7_o[22]),
    .sel(Rdkiu6),
    .o(Vgrhu6));  // ../RTL/cortexm0ds_logic.v(6732)
  AL_MUX u6136 (
    .i0(Zuliu6),
    .i1(vis_r6_o[22]),
    .sel(Kdkiu6),
    .o(Ogrhu6));  // ../RTL/cortexm0ds_logic.v(6733)
  AL_MUX u6137 (
    .i0(Zuliu6),
    .i1(vis_r5_o[22]),
    .sel(Ddkiu6),
    .o(Hgrhu6));  // ../RTL/cortexm0ds_logic.v(6734)
  AL_MUX u6138 (
    .i0(Zuliu6),
    .i1(vis_r4_o[22]),
    .sel(Wckiu6),
    .o(Agrhu6));  // ../RTL/cortexm0ds_logic.v(6735)
  AL_MUX u6139 (
    .i0(Zuliu6),
    .i1(vis_r11_o[22]),
    .sel(Afkiu6),
    .o(Tfrhu6));  // ../RTL/cortexm0ds_logic.v(6736)
  buf u614 (vis_r0_o[22], Tnebx6);  // ../RTL/cortexm0ds_logic.v(1875)
  AL_MUX u6140 (
    .i0(Zuliu6),
    .i1(vis_r10_o[22]),
    .sel(Hfkiu6),
    .o(Mfrhu6));  // ../RTL/cortexm0ds_logic.v(6737)
  AL_MUX u6141 (
    .i0(Zuliu6),
    .i1(vis_r9_o[22]),
    .sel(Ofkiu6),
    .o(Ffrhu6));  // ../RTL/cortexm0ds_logic.v(6738)
  AL_MUX u6142 (
    .i0(Zuliu6),
    .i1(vis_r8_o[22]),
    .sel(Vfkiu6),
    .o(Yerhu6));  // ../RTL/cortexm0ds_logic.v(6739)
  AL_MUX u6143 (
    .i0(Zuliu6),
    .i1(vis_r3_o[22]),
    .sel(Pckiu6),
    .o(Rerhu6));  // ../RTL/cortexm0ds_logic.v(6740)
  AL_MUX u6144 (
    .i0(Zuliu6),
    .i1(vis_r2_o[22]),
    .sel(Ickiu6),
    .o(Kerhu6));  // ../RTL/cortexm0ds_logic.v(6741)
  AL_MUX u6145 (
    .i0(Zuliu6),
    .i1(vis_r1_o[22]),
    .sel(Mx8iu6),
    .o(Derhu6));  // ../RTL/cortexm0ds_logic.v(6742)
  AL_MUX u6146 (
    .i0(Zuliu6),
    .i1(vis_r0_o[22]),
    .sel(Lf8iu6),
    .o(Wdrhu6));  // ../RTL/cortexm0ds_logic.v(6743)
  and u6147 (n1470, Gvliu6, Nvliu6);  // ../RTL/cortexm0ds_logic.v(6744)
  not u6148 (Zuliu6, n1470);  // ../RTL/cortexm0ds_logic.v(6744)
  and u6149 (Gvliu6, Uvliu6, Svkiu6);  // ../RTL/cortexm0ds_logic.v(6745)
  buf u615 (D7fpw6[13], P14qw6);  // ../RTL/cortexm0ds_logic.v(2074)
  and u6150 (n1471, Bwliu6, Iwliu6);  // ../RTL/cortexm0ds_logic.v(6746)
  not u6151 (Pdrhu6, n1471);  // ../RTL/cortexm0ds_logic.v(6746)
  and u6152 (Iwliu6, Pwliu6, Wwliu6);  // ../RTL/cortexm0ds_logic.v(6747)
  and u6153 (n1472, Jl8iu6, Yydpw6);  // ../RTL/cortexm0ds_logic.v(6748)
  not u6154 (Wwliu6, n1472);  // ../RTL/cortexm0ds_logic.v(6748)
  and u6155 (n1473, vis_pc_o[20], Ok8iu6);  // ../RTL/cortexm0ds_logic.v(6749)
  not u6156 (Pwliu6, n1473);  // ../RTL/cortexm0ds_logic.v(6749)
  and u6157 (Bwliu6, Dxliu6, Kxliu6);  // ../RTL/cortexm0ds_logic.v(6750)
  or u6158 (Kxliu6, Lm8iu6, Rxliu6);  // ../RTL/cortexm0ds_logic.v(6751)
  or u6159 (Dxliu6, Hx9iu6, Yxliu6);  // ../RTL/cortexm0ds_logic.v(6752)
  buf u616 (vis_r0_o[2], Vltpw6);  // ../RTL/cortexm0ds_logic.v(1875)
  AL_MUX u6160 (
    .i0(vis_psp_o[19]),
    .i1(Fyliu6),
    .sel(Ydkiu6),
    .o(Idrhu6));  // ../RTL/cortexm0ds_logic.v(6753)
  AL_MUX u6161 (
    .i0(vis_msp_o[19]),
    .i1(Fyliu6),
    .sel(Fekiu6),
    .o(Bdrhu6));  // ../RTL/cortexm0ds_logic.v(6754)
  AL_MUX u6162 (
    .i0(Fyliu6),
    .i1(vis_r14_o[21]),
    .sel(Mekiu6),
    .o(Ucrhu6));  // ../RTL/cortexm0ds_logic.v(6755)
  AL_MUX u6163 (
    .i0(Fyliu6),
    .i1(vis_r12_o[21]),
    .sel(Tekiu6),
    .o(Ncrhu6));  // ../RTL/cortexm0ds_logic.v(6756)
  AL_MUX u6164 (
    .i0(Fyliu6),
    .i1(vis_r7_o[21]),
    .sel(Rdkiu6),
    .o(Gcrhu6));  // ../RTL/cortexm0ds_logic.v(6757)
  AL_MUX u6165 (
    .i0(Fyliu6),
    .i1(vis_r6_o[21]),
    .sel(Kdkiu6),
    .o(Zbrhu6));  // ../RTL/cortexm0ds_logic.v(6758)
  AL_MUX u6166 (
    .i0(Fyliu6),
    .i1(vis_r5_o[21]),
    .sel(Ddkiu6),
    .o(Sbrhu6));  // ../RTL/cortexm0ds_logic.v(6759)
  AL_MUX u6167 (
    .i0(Fyliu6),
    .i1(vis_r4_o[21]),
    .sel(Wckiu6),
    .o(Lbrhu6));  // ../RTL/cortexm0ds_logic.v(6760)
  AL_MUX u6168 (
    .i0(Fyliu6),
    .i1(vis_r11_o[21]),
    .sel(Afkiu6),
    .o(Ebrhu6));  // ../RTL/cortexm0ds_logic.v(6761)
  AL_MUX u6169 (
    .i0(Fyliu6),
    .i1(vis_r10_o[21]),
    .sel(Hfkiu6),
    .o(Xarhu6));  // ../RTL/cortexm0ds_logic.v(6762)
  buf u617 (vis_r0_o[3], Gxmpw6);  // ../RTL/cortexm0ds_logic.v(1875)
  AL_MUX u6170 (
    .i0(Fyliu6),
    .i1(vis_r9_o[21]),
    .sel(Ofkiu6),
    .o(Qarhu6));  // ../RTL/cortexm0ds_logic.v(6763)
  AL_MUX u6171 (
    .i0(Fyliu6),
    .i1(vis_r8_o[21]),
    .sel(Vfkiu6),
    .o(Jarhu6));  // ../RTL/cortexm0ds_logic.v(6764)
  AL_MUX u6172 (
    .i0(Fyliu6),
    .i1(vis_r3_o[21]),
    .sel(Pckiu6),
    .o(Carhu6));  // ../RTL/cortexm0ds_logic.v(6765)
  AL_MUX u6173 (
    .i0(Fyliu6),
    .i1(vis_r2_o[21]),
    .sel(Ickiu6),
    .o(V9rhu6));  // ../RTL/cortexm0ds_logic.v(6766)
  AL_MUX u6174 (
    .i0(Fyliu6),
    .i1(vis_r1_o[21]),
    .sel(Mx8iu6),
    .o(O9rhu6));  // ../RTL/cortexm0ds_logic.v(6767)
  AL_MUX u6175 (
    .i0(Fyliu6),
    .i1(vis_r0_o[21]),
    .sel(Lf8iu6),
    .o(H9rhu6));  // ../RTL/cortexm0ds_logic.v(6768)
  and u6176 (n1474, Myliu6, Tyliu6);  // ../RTL/cortexm0ds_logic.v(6769)
  not u6177 (Fyliu6, n1474);  // ../RTL/cortexm0ds_logic.v(6769)
  and u6178 (Myliu6, Azliu6, Svkiu6);  // ../RTL/cortexm0ds_logic.v(6770)
  and u6179 (n1475, Hzliu6, Ozliu6);  // ../RTL/cortexm0ds_logic.v(6771)
  buf u618 (vis_r0_o[4], Uwipw6);  // ../RTL/cortexm0ds_logic.v(1875)
  not u6180 (A9rhu6, n1475);  // ../RTL/cortexm0ds_logic.v(6771)
  and u6181 (Ozliu6, Vzliu6, C0miu6);  // ../RTL/cortexm0ds_logic.v(6772)
  and u6182 (n1476, Jl8iu6, Rydpw6);  // ../RTL/cortexm0ds_logic.v(6773)
  not u6183 (C0miu6, n1476);  // ../RTL/cortexm0ds_logic.v(6773)
  and u6184 (n1477, vis_pc_o[19], Ok8iu6);  // ../RTL/cortexm0ds_logic.v(6774)
  not u6185 (Vzliu6, n1477);  // ../RTL/cortexm0ds_logic.v(6774)
  and u6186 (Hzliu6, J0miu6, Q0miu6);  // ../RTL/cortexm0ds_logic.v(6775)
  or u6187 (Q0miu6, Lm8iu6, X0miu6);  // ../RTL/cortexm0ds_logic.v(6776)
  and u6188 (n1478, Zm8iu6, B74iu6);  // ../RTL/cortexm0ds_logic.v(6777)
  not u6189 (J0miu6, n1478);  // ../RTL/cortexm0ds_logic.v(6777)
  buf u619 (vis_r0_o[5], Fzmpw6);  // ../RTL/cortexm0ds_logic.v(1875)
  AL_MUX u6190 (
    .i0(vis_psp_o[18]),
    .i1(E1miu6),
    .sel(Ydkiu6),
    .o(T8rhu6));  // ../RTL/cortexm0ds_logic.v(6778)
  AL_MUX u6191 (
    .i0(vis_msp_o[18]),
    .i1(E1miu6),
    .sel(Fekiu6),
    .o(M8rhu6));  // ../RTL/cortexm0ds_logic.v(6779)
  AL_MUX u6192 (
    .i0(E1miu6),
    .i1(vis_r14_o[20]),
    .sel(Mekiu6),
    .o(F8rhu6));  // ../RTL/cortexm0ds_logic.v(6780)
  AL_MUX u6193 (
    .i0(E1miu6),
    .i1(vis_r12_o[20]),
    .sel(Tekiu6),
    .o(Y7rhu6));  // ../RTL/cortexm0ds_logic.v(6781)
  AL_MUX u6194 (
    .i0(E1miu6),
    .i1(vis_r7_o[20]),
    .sel(Rdkiu6),
    .o(R7rhu6));  // ../RTL/cortexm0ds_logic.v(6782)
  AL_MUX u6195 (
    .i0(E1miu6),
    .i1(vis_r6_o[20]),
    .sel(Kdkiu6),
    .o(K7rhu6));  // ../RTL/cortexm0ds_logic.v(6783)
  AL_MUX u6196 (
    .i0(E1miu6),
    .i1(vis_r5_o[20]),
    .sel(Ddkiu6),
    .o(D7rhu6));  // ../RTL/cortexm0ds_logic.v(6784)
  AL_MUX u6197 (
    .i0(E1miu6),
    .i1(vis_r4_o[20]),
    .sel(Wckiu6),
    .o(W6rhu6));  // ../RTL/cortexm0ds_logic.v(6785)
  AL_MUX u6198 (
    .i0(E1miu6),
    .i1(vis_r11_o[20]),
    .sel(Afkiu6),
    .o(P6rhu6));  // ../RTL/cortexm0ds_logic.v(6786)
  AL_MUX u6199 (
    .i0(E1miu6),
    .i1(vis_r10_o[20]),
    .sel(Hfkiu6),
    .o(I6rhu6));  // ../RTL/cortexm0ds_logic.v(6787)
  buf u62 (vis_psp_o[17], Jtvpw6);  // ../RTL/cortexm0ds_logic.v(2085)
  buf u620 (vis_r0_o[6], B0spw6);  // ../RTL/cortexm0ds_logic.v(1875)
  AL_MUX u6200 (
    .i0(E1miu6),
    .i1(vis_r9_o[20]),
    .sel(Ofkiu6),
    .o(B6rhu6));  // ../RTL/cortexm0ds_logic.v(6788)
  AL_MUX u6201 (
    .i0(E1miu6),
    .i1(vis_r8_o[20]),
    .sel(Vfkiu6),
    .o(U5rhu6));  // ../RTL/cortexm0ds_logic.v(6789)
  AL_MUX u6202 (
    .i0(E1miu6),
    .i1(vis_r3_o[20]),
    .sel(Pckiu6),
    .o(N5rhu6));  // ../RTL/cortexm0ds_logic.v(6790)
  AL_MUX u6203 (
    .i0(E1miu6),
    .i1(vis_r2_o[20]),
    .sel(Ickiu6),
    .o(G5rhu6));  // ../RTL/cortexm0ds_logic.v(6791)
  AL_MUX u6204 (
    .i0(E1miu6),
    .i1(vis_r1_o[20]),
    .sel(Mx8iu6),
    .o(Z4rhu6));  // ../RTL/cortexm0ds_logic.v(6792)
  AL_MUX u6205 (
    .i0(E1miu6),
    .i1(vis_r0_o[20]),
    .sel(Lf8iu6),
    .o(S4rhu6));  // ../RTL/cortexm0ds_logic.v(6793)
  and u6206 (n1479, L1miu6, S1miu6);  // ../RTL/cortexm0ds_logic.v(6794)
  not u6207 (E1miu6, n1479);  // ../RTL/cortexm0ds_logic.v(6794)
  and u6208 (L1miu6, Z1miu6, Svkiu6);  // ../RTL/cortexm0ds_logic.v(6795)
  and u6209 (n1480, G2miu6, N2miu6);  // ../RTL/cortexm0ds_logic.v(6796)
  buf u621 (vis_r0_o[7], Emrpw6);  // ../RTL/cortexm0ds_logic.v(1875)
  not u6210 (L4rhu6, n1480);  // ../RTL/cortexm0ds_logic.v(6796)
  and u6211 (N2miu6, U2miu6, B3miu6);  // ../RTL/cortexm0ds_logic.v(6797)
  and u6212 (n1481, Jl8iu6, Kydpw6);  // ../RTL/cortexm0ds_logic.v(6798)
  not u6213 (B3miu6, n1481);  // ../RTL/cortexm0ds_logic.v(6798)
  and u6214 (n1482, vis_pc_o[18], Ok8iu6);  // ../RTL/cortexm0ds_logic.v(6799)
  not u6215 (U2miu6, n1482);  // ../RTL/cortexm0ds_logic.v(6799)
  and u6216 (G2miu6, I3miu6, P3miu6);  // ../RTL/cortexm0ds_logic.v(6800)
  or u6217 (P3miu6, Lm8iu6, W3miu6);  // ../RTL/cortexm0ds_logic.v(6801)
  and u6218 (n1483, Zm8iu6, U64iu6);  // ../RTL/cortexm0ds_logic.v(6802)
  not u6219 (I3miu6, n1483);  // ../RTL/cortexm0ds_logic.v(6802)
  buf u622 (vis_r0_o[9], Jp1qw6);  // ../RTL/cortexm0ds_logic.v(1875)
  AL_MUX u6220 (
    .i0(vis_psp_o[17]),
    .i1(D4miu6),
    .sel(Ydkiu6),
    .o(E4rhu6));  // ../RTL/cortexm0ds_logic.v(6803)
  AL_MUX u6221 (
    .i0(vis_msp_o[17]),
    .i1(D4miu6),
    .sel(Fekiu6),
    .o(X3rhu6));  // ../RTL/cortexm0ds_logic.v(6804)
  AL_MUX u6222 (
    .i0(D4miu6),
    .i1(vis_r14_o[19]),
    .sel(Mekiu6),
    .o(Q3rhu6));  // ../RTL/cortexm0ds_logic.v(6805)
  AL_MUX u6223 (
    .i0(D4miu6),
    .i1(vis_r12_o[19]),
    .sel(Tekiu6),
    .o(J3rhu6));  // ../RTL/cortexm0ds_logic.v(6806)
  AL_MUX u6224 (
    .i0(D4miu6),
    .i1(vis_r7_o[19]),
    .sel(Rdkiu6),
    .o(C3rhu6));  // ../RTL/cortexm0ds_logic.v(6807)
  AL_MUX u6225 (
    .i0(D4miu6),
    .i1(vis_r6_o[19]),
    .sel(Kdkiu6),
    .o(V2rhu6));  // ../RTL/cortexm0ds_logic.v(6808)
  AL_MUX u6226 (
    .i0(D4miu6),
    .i1(vis_r5_o[19]),
    .sel(Ddkiu6),
    .o(O2rhu6));  // ../RTL/cortexm0ds_logic.v(6809)
  AL_MUX u6227 (
    .i0(D4miu6),
    .i1(vis_r4_o[19]),
    .sel(Wckiu6),
    .o(H2rhu6));  // ../RTL/cortexm0ds_logic.v(6810)
  AL_MUX u6228 (
    .i0(D4miu6),
    .i1(vis_r11_o[19]),
    .sel(Afkiu6),
    .o(A2rhu6));  // ../RTL/cortexm0ds_logic.v(6811)
  AL_MUX u6229 (
    .i0(D4miu6),
    .i1(vis_r10_o[19]),
    .sel(Hfkiu6),
    .o(T1rhu6));  // ../RTL/cortexm0ds_logic.v(6812)
  buf u623 (vis_r0_o[10], Hkxpw6);  // ../RTL/cortexm0ds_logic.v(1875)
  AL_MUX u6230 (
    .i0(D4miu6),
    .i1(vis_r9_o[19]),
    .sel(Ofkiu6),
    .o(M1rhu6));  // ../RTL/cortexm0ds_logic.v(6813)
  AL_MUX u6231 (
    .i0(D4miu6),
    .i1(vis_r8_o[19]),
    .sel(Vfkiu6),
    .o(F1rhu6));  // ../RTL/cortexm0ds_logic.v(6814)
  AL_MUX u6232 (
    .i0(D4miu6),
    .i1(vis_r3_o[19]),
    .sel(Pckiu6),
    .o(Y0rhu6));  // ../RTL/cortexm0ds_logic.v(6815)
  AL_MUX u6233 (
    .i0(D4miu6),
    .i1(vis_r2_o[19]),
    .sel(Ickiu6),
    .o(R0rhu6));  // ../RTL/cortexm0ds_logic.v(6816)
  AL_MUX u6234 (
    .i0(D4miu6),
    .i1(vis_r1_o[19]),
    .sel(Mx8iu6),
    .o(K0rhu6));  // ../RTL/cortexm0ds_logic.v(6817)
  AL_MUX u6235 (
    .i0(D4miu6),
    .i1(vis_r0_o[19]),
    .sel(Lf8iu6),
    .o(D0rhu6));  // ../RTL/cortexm0ds_logic.v(6818)
  and u6236 (n1484, K4miu6, R4miu6);  // ../RTL/cortexm0ds_logic.v(6819)
  not u6237 (D4miu6, n1484);  // ../RTL/cortexm0ds_logic.v(6819)
  and u6238 (K4miu6, Y4miu6, Svkiu6);  // ../RTL/cortexm0ds_logic.v(6820)
  and u6239 (n1485, F5miu6, M5miu6);  // ../RTL/cortexm0ds_logic.v(6821)
  buf u624 (vis_r0_o[11], C27bx6);  // ../RTL/cortexm0ds_logic.v(1875)
  not u6240 (Wzqhu6, n1485);  // ../RTL/cortexm0ds_logic.v(6821)
  and u6241 (M5miu6, T5miu6, A6miu6);  // ../RTL/cortexm0ds_logic.v(6822)
  and u6242 (n1486, Jl8iu6, Dydpw6);  // ../RTL/cortexm0ds_logic.v(6823)
  not u6243 (A6miu6, n1486);  // ../RTL/cortexm0ds_logic.v(6823)
  and u6244 (n1487, vis_pc_o[17], Ok8iu6);  // ../RTL/cortexm0ds_logic.v(6824)
  not u6245 (T5miu6, n1487);  // ../RTL/cortexm0ds_logic.v(6824)
  and u6246 (F5miu6, H6miu6, O6miu6);  // ../RTL/cortexm0ds_logic.v(6825)
  or u6247 (O6miu6, Lm8iu6, V6miu6);  // ../RTL/cortexm0ds_logic.v(6826)
  and u6248 (n1488, Zm8iu6, N64iu6);  // ../RTL/cortexm0ds_logic.v(6827)
  not u6249 (H6miu6, n1488);  // ../RTL/cortexm0ds_logic.v(6827)
  buf u625 (vis_r0_o[13], E9npw6);  // ../RTL/cortexm0ds_logic.v(1875)
  AL_MUX u6250 (
    .i0(vis_psp_o[16]),
    .i1(C7miu6),
    .sel(Ydkiu6),
    .o(Pzqhu6));  // ../RTL/cortexm0ds_logic.v(6828)
  AL_MUX u6251 (
    .i0(vis_msp_o[16]),
    .i1(C7miu6),
    .sel(Fekiu6),
    .o(Izqhu6));  // ../RTL/cortexm0ds_logic.v(6829)
  AL_MUX u6252 (
    .i0(C7miu6),
    .i1(vis_r14_o[18]),
    .sel(Mekiu6),
    .o(Bzqhu6));  // ../RTL/cortexm0ds_logic.v(6830)
  AL_MUX u6253 (
    .i0(C7miu6),
    .i1(vis_r12_o[18]),
    .sel(Tekiu6),
    .o(Uyqhu6));  // ../RTL/cortexm0ds_logic.v(6831)
  AL_MUX u6254 (
    .i0(C7miu6),
    .i1(vis_r7_o[18]),
    .sel(Rdkiu6),
    .o(Nyqhu6));  // ../RTL/cortexm0ds_logic.v(6832)
  AL_MUX u6255 (
    .i0(C7miu6),
    .i1(vis_r6_o[18]),
    .sel(Kdkiu6),
    .o(Gyqhu6));  // ../RTL/cortexm0ds_logic.v(6833)
  AL_MUX u6256 (
    .i0(C7miu6),
    .i1(vis_r5_o[18]),
    .sel(Ddkiu6),
    .o(Zxqhu6));  // ../RTL/cortexm0ds_logic.v(6834)
  AL_MUX u6257 (
    .i0(C7miu6),
    .i1(vis_r4_o[18]),
    .sel(Wckiu6),
    .o(Sxqhu6));  // ../RTL/cortexm0ds_logic.v(6835)
  AL_MUX u6258 (
    .i0(C7miu6),
    .i1(vis_r11_o[18]),
    .sel(Afkiu6),
    .o(Lxqhu6));  // ../RTL/cortexm0ds_logic.v(6836)
  AL_MUX u6259 (
    .i0(C7miu6),
    .i1(vis_r10_o[18]),
    .sel(Hfkiu6),
    .o(Exqhu6));  // ../RTL/cortexm0ds_logic.v(6837)
  buf u626 (vis_r0_o[15], Zr7bx6);  // ../RTL/cortexm0ds_logic.v(1875)
  AL_MUX u6260 (
    .i0(C7miu6),
    .i1(vis_r9_o[18]),
    .sel(Ofkiu6),
    .o(Xwqhu6));  // ../RTL/cortexm0ds_logic.v(6838)
  AL_MUX u6261 (
    .i0(C7miu6),
    .i1(vis_r8_o[18]),
    .sel(Vfkiu6),
    .o(Qwqhu6));  // ../RTL/cortexm0ds_logic.v(6839)
  AL_MUX u6262 (
    .i0(C7miu6),
    .i1(vis_r3_o[18]),
    .sel(Pckiu6),
    .o(Jwqhu6));  // ../RTL/cortexm0ds_logic.v(6840)
  AL_MUX u6263 (
    .i0(C7miu6),
    .i1(vis_r2_o[18]),
    .sel(Ickiu6),
    .o(Cwqhu6));  // ../RTL/cortexm0ds_logic.v(6841)
  AL_MUX u6264 (
    .i0(C7miu6),
    .i1(vis_r1_o[18]),
    .sel(Mx8iu6),
    .o(Vvqhu6));  // ../RTL/cortexm0ds_logic.v(6842)
  AL_MUX u6265 (
    .i0(C7miu6),
    .i1(vis_r0_o[18]),
    .sel(Lf8iu6),
    .o(Ovqhu6));  // ../RTL/cortexm0ds_logic.v(6843)
  and u6266 (n1489, J7miu6, Q7miu6);  // ../RTL/cortexm0ds_logic.v(6844)
  not u6267 (C7miu6, n1489);  // ../RTL/cortexm0ds_logic.v(6844)
  and u6268 (J7miu6, X7miu6, Svkiu6);  // ../RTL/cortexm0ds_logic.v(6845)
  and u6269 (n1490, E8miu6, L8miu6);  // ../RTL/cortexm0ds_logic.v(6846)
  buf u627 (vis_r14_o[0], S5nax6);  // ../RTL/cortexm0ds_logic.v(2497)
  not u6270 (Hvqhu6, n1490);  // ../RTL/cortexm0ds_logic.v(6846)
  and u6271 (L8miu6, S8miu6, Z8miu6);  // ../RTL/cortexm0ds_logic.v(6847)
  and u6272 (n1491, Jl8iu6, Wxdpw6);  // ../RTL/cortexm0ds_logic.v(6848)
  not u6273 (Z8miu6, n1491);  // ../RTL/cortexm0ds_logic.v(6848)
  and u6274 (n1492, vis_pc_o[16], Ok8iu6);  // ../RTL/cortexm0ds_logic.v(6849)
  not u6275 (S8miu6, n1492);  // ../RTL/cortexm0ds_logic.v(6849)
  and u6276 (E8miu6, G9miu6, N9miu6);  // ../RTL/cortexm0ds_logic.v(6850)
  or u6277 (N9miu6, Lm8iu6, U9miu6);  // ../RTL/cortexm0ds_logic.v(6851)
  and u6278 (n1493, Zm8iu6, G64iu6);  // ../RTL/cortexm0ds_logic.v(6852)
  not u6279 (G9miu6, n1493);  // ../RTL/cortexm0ds_logic.v(6852)
  buf u628 (vis_r5_o[0], Oykax6);  // ../RTL/cortexm0ds_logic.v(1909)
  AL_MUX u6280 (
    .i0(vis_psp_o[15]),
    .i1(Bamiu6),
    .sel(Ydkiu6),
    .o(Avqhu6));  // ../RTL/cortexm0ds_logic.v(6853)
  AL_MUX u6281 (
    .i0(vis_msp_o[15]),
    .i1(Bamiu6),
    .sel(Fekiu6),
    .o(Tuqhu6));  // ../RTL/cortexm0ds_logic.v(6854)
  AL_MUX u6282 (
    .i0(Bamiu6),
    .i1(vis_r14_o[17]),
    .sel(Mekiu6),
    .o(Muqhu6));  // ../RTL/cortexm0ds_logic.v(6855)
  AL_MUX u6283 (
    .i0(Bamiu6),
    .i1(vis_r12_o[17]),
    .sel(Tekiu6),
    .o(Fuqhu6));  // ../RTL/cortexm0ds_logic.v(6856)
  AL_MUX u6284 (
    .i0(Bamiu6),
    .i1(vis_r7_o[17]),
    .sel(Rdkiu6),
    .o(Ytqhu6));  // ../RTL/cortexm0ds_logic.v(6857)
  AL_MUX u6285 (
    .i0(Bamiu6),
    .i1(vis_r6_o[17]),
    .sel(Kdkiu6),
    .o(Rtqhu6));  // ../RTL/cortexm0ds_logic.v(6858)
  AL_MUX u6286 (
    .i0(Bamiu6),
    .i1(vis_r5_o[17]),
    .sel(Ddkiu6),
    .o(Ktqhu6));  // ../RTL/cortexm0ds_logic.v(6859)
  AL_MUX u6287 (
    .i0(Bamiu6),
    .i1(vis_r4_o[17]),
    .sel(Wckiu6),
    .o(Dtqhu6));  // ../RTL/cortexm0ds_logic.v(6860)
  AL_MUX u6288 (
    .i0(Bamiu6),
    .i1(vis_r11_o[17]),
    .sel(Afkiu6),
    .o(Wsqhu6));  // ../RTL/cortexm0ds_logic.v(6861)
  AL_MUX u6289 (
    .i0(Bamiu6),
    .i1(vis_r10_o[17]),
    .sel(Hfkiu6),
    .o(Psqhu6));  // ../RTL/cortexm0ds_logic.v(6862)
  buf u629 (Gqgpw6[26], Thcbx6);  // ../RTL/cortexm0ds_logic.v(2377)
  AL_MUX u6290 (
    .i0(Bamiu6),
    .i1(vis_r9_o[17]),
    .sel(Ofkiu6),
    .o(Isqhu6));  // ../RTL/cortexm0ds_logic.v(6863)
  AL_MUX u6291 (
    .i0(Bamiu6),
    .i1(vis_r8_o[17]),
    .sel(Vfkiu6),
    .o(Bsqhu6));  // ../RTL/cortexm0ds_logic.v(6864)
  AL_MUX u6292 (
    .i0(Bamiu6),
    .i1(vis_r3_o[17]),
    .sel(Pckiu6),
    .o(Urqhu6));  // ../RTL/cortexm0ds_logic.v(6865)
  AL_MUX u6293 (
    .i0(Bamiu6),
    .i1(vis_r2_o[17]),
    .sel(Ickiu6),
    .o(Nrqhu6));  // ../RTL/cortexm0ds_logic.v(6866)
  AL_MUX u6294 (
    .i0(Bamiu6),
    .i1(vis_r1_o[17]),
    .sel(Mx8iu6),
    .o(Grqhu6));  // ../RTL/cortexm0ds_logic.v(6867)
  AL_MUX u6295 (
    .i0(Bamiu6),
    .i1(vis_r0_o[17]),
    .sel(Lf8iu6),
    .o(Zqqhu6));  // ../RTL/cortexm0ds_logic.v(6868)
  and u6296 (n1494, Iamiu6, Pamiu6);  // ../RTL/cortexm0ds_logic.v(6869)
  not u6297 (Bamiu6, n1494);  // ../RTL/cortexm0ds_logic.v(6869)
  and u6298 (Iamiu6, Wamiu6, Svkiu6);  // ../RTL/cortexm0ds_logic.v(6870)
  and u6299 (n1495, Dbmiu6, Kbmiu6);  // ../RTL/cortexm0ds_logic.v(6871)
  buf u63 (vis_r4_o[23], B4uax6);  // ../RTL/cortexm0ds_logic.v(2626)
  buf u630 (vis_r8_o[0], Qorax6);  // ../RTL/cortexm0ds_logic.v(2579)
  not u6300 (Sqqhu6, n1495);  // ../RTL/cortexm0ds_logic.v(6871)
  and u6301 (Kbmiu6, Rbmiu6, Ybmiu6);  // ../RTL/cortexm0ds_logic.v(6872)
  and u6302 (n1496, Jl8iu6, Pxdpw6);  // ../RTL/cortexm0ds_logic.v(6873)
  not u6303 (Ybmiu6, n1496);  // ../RTL/cortexm0ds_logic.v(6873)
  and u6304 (n1497, vis_pc_o[15], Ok8iu6);  // ../RTL/cortexm0ds_logic.v(6874)
  not u6305 (Rbmiu6, n1497);  // ../RTL/cortexm0ds_logic.v(6874)
  and u6306 (Dbmiu6, Fcmiu6, Mcmiu6);  // ../RTL/cortexm0ds_logic.v(6875)
  or u6307 (Mcmiu6, Lm8iu6, Tcmiu6);  // ../RTL/cortexm0ds_logic.v(6876)
  and u6308 (n1498, Zm8iu6, Z54iu6);  // ../RTL/cortexm0ds_logic.v(6877)
  not u6309 (Fcmiu6, n1498);  // ../RTL/cortexm0ds_logic.v(6877)
  buf u631 (Uthpw6[5], Ceabx6);  // ../RTL/cortexm0ds_logic.v(1882)
  AL_MUX u6310 (
    .i0(vis_psp_o[14]),
    .i1(Admiu6),
    .sel(Ydkiu6),
    .o(Lqqhu6));  // ../RTL/cortexm0ds_logic.v(6878)
  AL_MUX u6311 (
    .i0(vis_msp_o[14]),
    .i1(Admiu6),
    .sel(Fekiu6),
    .o(Eqqhu6));  // ../RTL/cortexm0ds_logic.v(6879)
  AL_MUX u6312 (
    .i0(Admiu6),
    .i1(vis_r14_o[16]),
    .sel(Mekiu6),
    .o(Xpqhu6));  // ../RTL/cortexm0ds_logic.v(6880)
  AL_MUX u6313 (
    .i0(Admiu6),
    .i1(vis_r12_o[16]),
    .sel(Tekiu6),
    .o(Qpqhu6));  // ../RTL/cortexm0ds_logic.v(6881)
  AL_MUX u6314 (
    .i0(Admiu6),
    .i1(vis_r7_o[16]),
    .sel(Rdkiu6),
    .o(Jpqhu6));  // ../RTL/cortexm0ds_logic.v(6882)
  AL_MUX u6315 (
    .i0(Admiu6),
    .i1(vis_r6_o[16]),
    .sel(Kdkiu6),
    .o(Cpqhu6));  // ../RTL/cortexm0ds_logic.v(6883)
  AL_MUX u6316 (
    .i0(Admiu6),
    .i1(vis_r5_o[16]),
    .sel(Ddkiu6),
    .o(Voqhu6));  // ../RTL/cortexm0ds_logic.v(6884)
  AL_MUX u6317 (
    .i0(Admiu6),
    .i1(vis_r4_o[16]),
    .sel(Wckiu6),
    .o(Ooqhu6));  // ../RTL/cortexm0ds_logic.v(6885)
  AL_MUX u6318 (
    .i0(Admiu6),
    .i1(vis_r11_o[16]),
    .sel(Afkiu6),
    .o(Hoqhu6));  // ../RTL/cortexm0ds_logic.v(6886)
  AL_MUX u6319 (
    .i0(Admiu6),
    .i1(vis_r10_o[16]),
    .sel(Hfkiu6),
    .o(Aoqhu6));  // ../RTL/cortexm0ds_logic.v(6887)
  buf u632 (Jshpw6[29], Cq3qw6);  // ../RTL/cortexm0ds_logic.v(2372)
  AL_MUX u6320 (
    .i0(Admiu6),
    .i1(vis_r9_o[16]),
    .sel(Ofkiu6),
    .o(Tnqhu6));  // ../RTL/cortexm0ds_logic.v(6888)
  AL_MUX u6321 (
    .i0(Admiu6),
    .i1(vis_r8_o[16]),
    .sel(Vfkiu6),
    .o(Mnqhu6));  // ../RTL/cortexm0ds_logic.v(6889)
  AL_MUX u6322 (
    .i0(Admiu6),
    .i1(vis_r3_o[16]),
    .sel(Pckiu6),
    .o(Fnqhu6));  // ../RTL/cortexm0ds_logic.v(6890)
  AL_MUX u6323 (
    .i0(Admiu6),
    .i1(vis_r2_o[16]),
    .sel(Ickiu6),
    .o(Ymqhu6));  // ../RTL/cortexm0ds_logic.v(6891)
  AL_MUX u6324 (
    .i0(Admiu6),
    .i1(vis_r1_o[16]),
    .sel(Mx8iu6),
    .o(Rmqhu6));  // ../RTL/cortexm0ds_logic.v(6892)
  AL_MUX u6325 (
    .i0(Admiu6),
    .i1(vis_r0_o[16]),
    .sel(Lf8iu6),
    .o(Kmqhu6));  // ../RTL/cortexm0ds_logic.v(6893)
  and u6326 (n1499, Hdmiu6, Odmiu6);  // ../RTL/cortexm0ds_logic.v(6894)
  not u6327 (Admiu6, n1499);  // ../RTL/cortexm0ds_logic.v(6894)
  and u6328 (Hdmiu6, Vdmiu6, Svkiu6);  // ../RTL/cortexm0ds_logic.v(6895)
  and u6329 (n1500, Cemiu6, Jemiu6);  // ../RTL/cortexm0ds_logic.v(6896)
  buf u633 (Uthpw6[6], Vefax6);  // ../RTL/cortexm0ds_logic.v(1882)
  not u6330 (Dmqhu6, n1500);  // ../RTL/cortexm0ds_logic.v(6896)
  and u6331 (Jemiu6, Qemiu6, Xemiu6);  // ../RTL/cortexm0ds_logic.v(6897)
  and u6332 (n1501, Jl8iu6, Tugpw6[13]);  // ../RTL/cortexm0ds_logic.v(6898)
  not u6333 (Xemiu6, n1501);  // ../RTL/cortexm0ds_logic.v(6898)
  and u6334 (n1502, vis_pc_o[14], Ok8iu6);  // ../RTL/cortexm0ds_logic.v(6899)
  not u6335 (Qemiu6, n1502);  // ../RTL/cortexm0ds_logic.v(6899)
  and u6336 (Cemiu6, Efmiu6, Lfmiu6);  // ../RTL/cortexm0ds_logic.v(6900)
  or u6337 (Lfmiu6, Lm8iu6, Sfmiu6);  // ../RTL/cortexm0ds_logic.v(6901)
  and u6338 (n1503, Zm8iu6, S54iu6);  // ../RTL/cortexm0ds_logic.v(6902)
  not u6339 (Efmiu6, n1503);  // ../RTL/cortexm0ds_logic.v(6902)
  buf u634 (Jshpw6[30], Wc2qw6);  // ../RTL/cortexm0ds_logic.v(2372)
  AL_MUX u6340 (
    .i0(vis_psp_o[13]),
    .i1(Zfmiu6),
    .sel(Ydkiu6),
    .o(Wlqhu6));  // ../RTL/cortexm0ds_logic.v(6903)
  AL_MUX u6341 (
    .i0(vis_msp_o[13]),
    .i1(Zfmiu6),
    .sel(Fekiu6),
    .o(Plqhu6));  // ../RTL/cortexm0ds_logic.v(6904)
  AL_MUX u6342 (
    .i0(Zfmiu6),
    .i1(vis_r14_o[15]),
    .sel(Mekiu6),
    .o(Ilqhu6));  // ../RTL/cortexm0ds_logic.v(6905)
  AL_MUX u6343 (
    .i0(Zfmiu6),
    .i1(vis_r12_o[15]),
    .sel(Tekiu6),
    .o(Blqhu6));  // ../RTL/cortexm0ds_logic.v(6906)
  AL_MUX u6344 (
    .i0(Zfmiu6),
    .i1(vis_r7_o[15]),
    .sel(Rdkiu6),
    .o(Ukqhu6));  // ../RTL/cortexm0ds_logic.v(6907)
  AL_MUX u6345 (
    .i0(Zfmiu6),
    .i1(vis_r6_o[15]),
    .sel(Kdkiu6),
    .o(Nkqhu6));  // ../RTL/cortexm0ds_logic.v(6908)
  AL_MUX u6346 (
    .i0(Zfmiu6),
    .i1(vis_r5_o[15]),
    .sel(Ddkiu6),
    .o(Gkqhu6));  // ../RTL/cortexm0ds_logic.v(6909)
  AL_MUX u6347 (
    .i0(Zfmiu6),
    .i1(vis_r4_o[15]),
    .sel(Wckiu6),
    .o(Zjqhu6));  // ../RTL/cortexm0ds_logic.v(6910)
  AL_MUX u6348 (
    .i0(Zfmiu6),
    .i1(vis_r11_o[15]),
    .sel(Afkiu6),
    .o(Sjqhu6));  // ../RTL/cortexm0ds_logic.v(6911)
  AL_MUX u6349 (
    .i0(Zfmiu6),
    .i1(vis_r10_o[15]),
    .sel(Hfkiu6),
    .o(Ljqhu6));  // ../RTL/cortexm0ds_logic.v(6912)
  buf u635 (Uthpw6[13], Ggabx6);  // ../RTL/cortexm0ds_logic.v(1882)
  AL_MUX u6350 (
    .i0(Zfmiu6),
    .i1(vis_r9_o[15]),
    .sel(Ofkiu6),
    .o(Ejqhu6));  // ../RTL/cortexm0ds_logic.v(6913)
  AL_MUX u6351 (
    .i0(Zfmiu6),
    .i1(vis_r8_o[15]),
    .sel(Vfkiu6),
    .o(Xiqhu6));  // ../RTL/cortexm0ds_logic.v(6914)
  AL_MUX u6352 (
    .i0(Zfmiu6),
    .i1(vis_r3_o[15]),
    .sel(Pckiu6),
    .o(Qiqhu6));  // ../RTL/cortexm0ds_logic.v(6915)
  AL_MUX u6353 (
    .i0(Zfmiu6),
    .i1(vis_r2_o[15]),
    .sel(Ickiu6),
    .o(Jiqhu6));  // ../RTL/cortexm0ds_logic.v(6916)
  AL_MUX u6354 (
    .i0(Zfmiu6),
    .i1(vis_r1_o[15]),
    .sel(Mx8iu6),
    .o(Ciqhu6));  // ../RTL/cortexm0ds_logic.v(6917)
  AL_MUX u6355 (
    .i0(Zfmiu6),
    .i1(vis_r0_o[15]),
    .sel(Lf8iu6),
    .o(Vhqhu6));  // ../RTL/cortexm0ds_logic.v(6918)
  and u6356 (n1504, Ggmiu6, Ngmiu6);  // ../RTL/cortexm0ds_logic.v(6919)
  not u6357 (Zfmiu6, n1504);  // ../RTL/cortexm0ds_logic.v(6919)
  and u6358 (n1505, Ugmiu6, Bhmiu6);  // ../RTL/cortexm0ds_logic.v(6920)
  not u6359 (Ohqhu6, n1505);  // ../RTL/cortexm0ds_logic.v(6920)
  buf u636 (G4hpw6[3], P9bax6);  // ../RTL/cortexm0ds_logic.v(2274)
  and u6360 (Bhmiu6, Ihmiu6, Phmiu6);  // ../RTL/cortexm0ds_logic.v(6921)
  and u6361 (n1506, Jl8iu6, Tugpw6[12]);  // ../RTL/cortexm0ds_logic.v(6922)
  not u6362 (Phmiu6, n1506);  // ../RTL/cortexm0ds_logic.v(6922)
  and u6363 (n1507, vis_pc_o[13], Ok8iu6);  // ../RTL/cortexm0ds_logic.v(6923)
  not u6364 (Ihmiu6, n1507);  // ../RTL/cortexm0ds_logic.v(6923)
  and u6365 (Ugmiu6, Whmiu6, Dimiu6);  // ../RTL/cortexm0ds_logic.v(6924)
  or u6366 (Dimiu6, Lm8iu6, Kimiu6);  // ../RTL/cortexm0ds_logic.v(6925)
  and u6367 (n1508, Zm8iu6, L54iu6);  // ../RTL/cortexm0ds_logic.v(6926)
  not u6368 (Whmiu6, n1508);  // ../RTL/cortexm0ds_logic.v(6926)
  AL_MUX u6369 (
    .i0(vis_psp_o[12]),
    .i1(Rimiu6),
    .sel(Ydkiu6),
    .o(Hhqhu6));  // ../RTL/cortexm0ds_logic.v(6927)
  buf u637 (Uthpw6[18], Kswpw6);  // ../RTL/cortexm0ds_logic.v(1882)
  AL_MUX u6370 (
    .i0(vis_msp_o[12]),
    .i1(Rimiu6),
    .sel(Fekiu6),
    .o(Ahqhu6));  // ../RTL/cortexm0ds_logic.v(6928)
  AL_MUX u6371 (
    .i0(Rimiu6),
    .i1(vis_r14_o[14]),
    .sel(Mekiu6),
    .o(Tgqhu6));  // ../RTL/cortexm0ds_logic.v(6929)
  AL_MUX u6372 (
    .i0(Rimiu6),
    .i1(vis_r12_o[14]),
    .sel(Tekiu6),
    .o(Mgqhu6));  // ../RTL/cortexm0ds_logic.v(6930)
  AL_MUX u6373 (
    .i0(Rimiu6),
    .i1(vis_r7_o[14]),
    .sel(Rdkiu6),
    .o(Fgqhu6));  // ../RTL/cortexm0ds_logic.v(6931)
  AL_MUX u6374 (
    .i0(Rimiu6),
    .i1(vis_r6_o[14]),
    .sel(Kdkiu6),
    .o(Yfqhu6));  // ../RTL/cortexm0ds_logic.v(6932)
  AL_MUX u6375 (
    .i0(Rimiu6),
    .i1(vis_r5_o[14]),
    .sel(Ddkiu6),
    .o(Rfqhu6));  // ../RTL/cortexm0ds_logic.v(6933)
  AL_MUX u6376 (
    .i0(Rimiu6),
    .i1(vis_r4_o[14]),
    .sel(Wckiu6),
    .o(Kfqhu6));  // ../RTL/cortexm0ds_logic.v(6934)
  AL_MUX u6377 (
    .i0(Rimiu6),
    .i1(vis_r11_o[14]),
    .sel(Afkiu6),
    .o(Dfqhu6));  // ../RTL/cortexm0ds_logic.v(6935)
  AL_MUX u6378 (
    .i0(Rimiu6),
    .i1(vis_r10_o[14]),
    .sel(Hfkiu6),
    .o(Weqhu6));  // ../RTL/cortexm0ds_logic.v(6936)
  AL_MUX u6379 (
    .i0(Rimiu6),
    .i1(vis_r9_o[14]),
    .sel(Ofkiu6),
    .o(Peqhu6));  // ../RTL/cortexm0ds_logic.v(6937)
  buf u638 (Uthpw6[19], Gbvpw6);  // ../RTL/cortexm0ds_logic.v(1882)
  AL_MUX u6380 (
    .i0(Rimiu6),
    .i1(vis_r8_o[14]),
    .sel(Vfkiu6),
    .o(Ieqhu6));  // ../RTL/cortexm0ds_logic.v(6938)
  AL_MUX u6381 (
    .i0(Rimiu6),
    .i1(vis_r3_o[14]),
    .sel(Pckiu6),
    .o(Beqhu6));  // ../RTL/cortexm0ds_logic.v(6939)
  AL_MUX u6382 (
    .i0(Rimiu6),
    .i1(vis_r2_o[14]),
    .sel(Ickiu6),
    .o(Udqhu6));  // ../RTL/cortexm0ds_logic.v(6940)
  AL_MUX u6383 (
    .i0(Rimiu6),
    .i1(vis_r1_o[14]),
    .sel(Mx8iu6),
    .o(Ndqhu6));  // ../RTL/cortexm0ds_logic.v(6941)
  AL_MUX u6384 (
    .i0(Rimiu6),
    .i1(vis_r0_o[14]),
    .sel(Lf8iu6),
    .o(Gdqhu6));  // ../RTL/cortexm0ds_logic.v(6942)
  or u6385 (Rimiu6, Yimiu6, Fjmiu6);  // ../RTL/cortexm0ds_logic.v(6943)
  and u6386 (n1509, Mjmiu6, Tjmiu6);  // ../RTL/cortexm0ds_logic.v(6944)
  not u6387 (Zcqhu6, n1509);  // ../RTL/cortexm0ds_logic.v(6944)
  and u6388 (Tjmiu6, Akmiu6, Hkmiu6);  // ../RTL/cortexm0ds_logic.v(6945)
  and u6389 (n1510, Jl8iu6, Tugpw6[11]);  // ../RTL/cortexm0ds_logic.v(6946)
  buf u639 (vis_psp_o[4], B5zpw6);  // ../RTL/cortexm0ds_logic.v(2085)
  not u6390 (Hkmiu6, n1510);  // ../RTL/cortexm0ds_logic.v(6946)
  and u6391 (n1511, vis_pc_o[12], Ok8iu6);  // ../RTL/cortexm0ds_logic.v(6947)
  not u6392 (Akmiu6, n1511);  // ../RTL/cortexm0ds_logic.v(6947)
  and u6393 (Mjmiu6, Okmiu6, Vkmiu6);  // ../RTL/cortexm0ds_logic.v(6948)
  or u6394 (Vkmiu6, Lm8iu6, Clmiu6);  // ../RTL/cortexm0ds_logic.v(6949)
  and u6395 (n1512, Zm8iu6, E54iu6);  // ../RTL/cortexm0ds_logic.v(6950)
  not u6396 (Okmiu6, n1512);  // ../RTL/cortexm0ds_logic.v(6950)
  AL_MUX u6397 (
    .i0(vis_psp_o[11]),
    .i1(Jlmiu6),
    .sel(Ydkiu6),
    .o(Scqhu6));  // ../RTL/cortexm0ds_logic.v(6951)
  AL_MUX u6398 (
    .i0(vis_msp_o[11]),
    .i1(Jlmiu6),
    .sel(Fekiu6),
    .o(Lcqhu6));  // ../RTL/cortexm0ds_logic.v(6952)
  AL_MUX u6399 (
    .i0(Jlmiu6),
    .i1(vis_r14_o[13]),
    .sel(Mekiu6),
    .o(Ecqhu6));  // ../RTL/cortexm0ds_logic.v(6953)
  buf u64 (Tonhu6, L5lpw6);  // ../RTL/cortexm0ds_logic.v(1830)
  buf u640 (vis_psp_o[15], Yhupw6);  // ../RTL/cortexm0ds_logic.v(2085)
  AL_MUX u6400 (
    .i0(Jlmiu6),
    .i1(vis_r12_o[13]),
    .sel(Tekiu6),
    .o(Xbqhu6));  // ../RTL/cortexm0ds_logic.v(6954)
  AL_MUX u6401 (
    .i0(Jlmiu6),
    .i1(vis_r7_o[13]),
    .sel(Rdkiu6),
    .o(Qbqhu6));  // ../RTL/cortexm0ds_logic.v(6955)
  AL_MUX u6402 (
    .i0(Jlmiu6),
    .i1(vis_r6_o[13]),
    .sel(Kdkiu6),
    .o(Jbqhu6));  // ../RTL/cortexm0ds_logic.v(6956)
  AL_MUX u6403 (
    .i0(Jlmiu6),
    .i1(vis_r5_o[13]),
    .sel(Ddkiu6),
    .o(Cbqhu6));  // ../RTL/cortexm0ds_logic.v(6957)
  AL_MUX u6404 (
    .i0(Jlmiu6),
    .i1(vis_r4_o[13]),
    .sel(Wckiu6),
    .o(Vaqhu6));  // ../RTL/cortexm0ds_logic.v(6958)
  AL_MUX u6405 (
    .i0(Jlmiu6),
    .i1(vis_r11_o[13]),
    .sel(Afkiu6),
    .o(Oaqhu6));  // ../RTL/cortexm0ds_logic.v(6959)
  AL_MUX u6406 (
    .i0(Jlmiu6),
    .i1(vis_r10_o[13]),
    .sel(Hfkiu6),
    .o(Haqhu6));  // ../RTL/cortexm0ds_logic.v(6960)
  AL_MUX u6407 (
    .i0(Jlmiu6),
    .i1(vis_r9_o[13]),
    .sel(Ofkiu6),
    .o(Aaqhu6));  // ../RTL/cortexm0ds_logic.v(6961)
  AL_MUX u6408 (
    .i0(Jlmiu6),
    .i1(vis_r8_o[13]),
    .sel(Vfkiu6),
    .o(T9qhu6));  // ../RTL/cortexm0ds_logic.v(6962)
  AL_MUX u6409 (
    .i0(Jlmiu6),
    .i1(vis_r3_o[13]),
    .sel(Pckiu6),
    .o(M9qhu6));  // ../RTL/cortexm0ds_logic.v(6963)
  buf u641 (vis_psp_o[13], Zl8bx6);  // ../RTL/cortexm0ds_logic.v(2085)
  AL_MUX u6410 (
    .i0(Jlmiu6),
    .i1(vis_r2_o[13]),
    .sel(Ickiu6),
    .o(F9qhu6));  // ../RTL/cortexm0ds_logic.v(6964)
  AL_MUX u6411 (
    .i0(Jlmiu6),
    .i1(vis_r1_o[13]),
    .sel(Mx8iu6),
    .o(Y8qhu6));  // ../RTL/cortexm0ds_logic.v(6965)
  AL_MUX u6412 (
    .i0(Jlmiu6),
    .i1(vis_r0_o[13]),
    .sel(Lf8iu6),
    .o(R8qhu6));  // ../RTL/cortexm0ds_logic.v(6966)
  or u6413 (Jlmiu6, Qlmiu6, Xlmiu6);  // ../RTL/cortexm0ds_logic.v(6967)
  and u6414 (n1513, Emmiu6, Lmmiu6);  // ../RTL/cortexm0ds_logic.v(6968)
  not u6415 (K8qhu6, n1513);  // ../RTL/cortexm0ds_logic.v(6968)
  and u6416 (Lmmiu6, Smmiu6, Zmmiu6);  // ../RTL/cortexm0ds_logic.v(6969)
  and u6417 (n1514, Jl8iu6, Ixdpw6);  // ../RTL/cortexm0ds_logic.v(6970)
  not u6418 (Zmmiu6, n1514);  // ../RTL/cortexm0ds_logic.v(6970)
  and u6419 (n1515, vis_pc_o[11], Ok8iu6);  // ../RTL/cortexm0ds_logic.v(6971)
  buf u642 (Vbgpw6[0], C3wpw6);  // ../RTL/cortexm0ds_logic.v(3092)
  not u6420 (Smmiu6, n1515);  // ../RTL/cortexm0ds_logic.v(6971)
  and u6421 (Emmiu6, Gnmiu6, Nnmiu6);  // ../RTL/cortexm0ds_logic.v(6972)
  or u6422 (Nnmiu6, Lm8iu6, Unmiu6);  // ../RTL/cortexm0ds_logic.v(6973)
  and u6423 (n1516, Zm8iu6, X44iu6);  // ../RTL/cortexm0ds_logic.v(6974)
  not u6424 (Gnmiu6, n1516);  // ../RTL/cortexm0ds_logic.v(6974)
  AL_MUX u6425 (
    .i0(vis_psp_o[10]),
    .i1(Bomiu6),
    .sel(Ydkiu6),
    .o(D8qhu6));  // ../RTL/cortexm0ds_logic.v(6975)
  AL_MUX u6426 (
    .i0(vis_msp_o[10]),
    .i1(Bomiu6),
    .sel(Fekiu6),
    .o(W7qhu6));  // ../RTL/cortexm0ds_logic.v(6976)
  AL_MUX u6427 (
    .i0(Bomiu6),
    .i1(vis_r14_o[12]),
    .sel(Mekiu6),
    .o(P7qhu6));  // ../RTL/cortexm0ds_logic.v(6977)
  AL_MUX u6428 (
    .i0(Bomiu6),
    .i1(vis_r12_o[12]),
    .sel(Tekiu6),
    .o(I7qhu6));  // ../RTL/cortexm0ds_logic.v(6978)
  AL_MUX u6429 (
    .i0(Bomiu6),
    .i1(vis_r7_o[12]),
    .sel(Rdkiu6),
    .o(B7qhu6));  // ../RTL/cortexm0ds_logic.v(6979)
  buf u643 (vis_psp_o[14], Cfwpw6);  // ../RTL/cortexm0ds_logic.v(2085)
  AL_MUX u6430 (
    .i0(Bomiu6),
    .i1(vis_r6_o[12]),
    .sel(Kdkiu6),
    .o(U6qhu6));  // ../RTL/cortexm0ds_logic.v(6980)
  AL_MUX u6431 (
    .i0(Bomiu6),
    .i1(vis_r5_o[12]),
    .sel(Ddkiu6),
    .o(N6qhu6));  // ../RTL/cortexm0ds_logic.v(6981)
  AL_MUX u6432 (
    .i0(Bomiu6),
    .i1(vis_r4_o[12]),
    .sel(Wckiu6),
    .o(G6qhu6));  // ../RTL/cortexm0ds_logic.v(6982)
  AL_MUX u6433 (
    .i0(Bomiu6),
    .i1(vis_r11_o[12]),
    .sel(Afkiu6),
    .o(Z5qhu6));  // ../RTL/cortexm0ds_logic.v(6983)
  AL_MUX u6434 (
    .i0(Bomiu6),
    .i1(vis_r10_o[12]),
    .sel(Hfkiu6),
    .o(S5qhu6));  // ../RTL/cortexm0ds_logic.v(6984)
  AL_MUX u6435 (
    .i0(Bomiu6),
    .i1(vis_r9_o[12]),
    .sel(Ofkiu6),
    .o(L5qhu6));  // ../RTL/cortexm0ds_logic.v(6985)
  AL_MUX u6436 (
    .i0(Bomiu6),
    .i1(vis_r8_o[12]),
    .sel(Vfkiu6),
    .o(E5qhu6));  // ../RTL/cortexm0ds_logic.v(6986)
  AL_MUX u6437 (
    .i0(Bomiu6),
    .i1(vis_r3_o[12]),
    .sel(Pckiu6),
    .o(X4qhu6));  // ../RTL/cortexm0ds_logic.v(6987)
  AL_MUX u6438 (
    .i0(Bomiu6),
    .i1(vis_r2_o[12]),
    .sel(Ickiu6),
    .o(Q4qhu6));  // ../RTL/cortexm0ds_logic.v(6988)
  AL_MUX u6439 (
    .i0(Bomiu6),
    .i1(vis_r1_o[12]),
    .sel(Mx8iu6),
    .o(J4qhu6));  // ../RTL/cortexm0ds_logic.v(6989)
  buf u644 (Gqgpw6[24], Qmdax6);  // ../RTL/cortexm0ds_logic.v(2377)
  AL_MUX u6440 (
    .i0(Bomiu6),
    .i1(vis_r0_o[12]),
    .sel(Lf8iu6),
    .o(C4qhu6));  // ../RTL/cortexm0ds_logic.v(6990)
  or u6441 (Bomiu6, Iomiu6, Pomiu6);  // ../RTL/cortexm0ds_logic.v(6991)
  and u6442 (n1517, Womiu6, Dpmiu6);  // ../RTL/cortexm0ds_logic.v(6992)
  not u6443 (V3qhu6, n1517);  // ../RTL/cortexm0ds_logic.v(6992)
  and u6444 (Dpmiu6, Kpmiu6, Rpmiu6);  // ../RTL/cortexm0ds_logic.v(6993)
  and u6445 (n1518, Jl8iu6, Tugpw6[9]);  // ../RTL/cortexm0ds_logic.v(6994)
  not u6446 (Rpmiu6, n1518);  // ../RTL/cortexm0ds_logic.v(6994)
  buf u6447 (vis_r7_o[7], N1wax6);  // ../RTL/cortexm0ds_logic.v(2654)
  buf u6448 (vis_r7_o[19], Ljwax6);  // ../RTL/cortexm0ds_logic.v(2654)
  and u6449 (n1519, N5fpw6[10], Sdaiu6);  // ../RTL/cortexm0ds_logic.v(6996)
  not u645 (Evdpw6, Sbyax6);  // ../RTL/cortexm0ds_logic.v(2700)
  not u6450 (Fqmiu6, n1519);  // ../RTL/cortexm0ds_logic.v(6996)
  and u6451 (Ypmiu6, Mqmiu6, Tqmiu6);  // ../RTL/cortexm0ds_logic.v(6997)
  or u6452 (Tqmiu6, T2iiu6, Sn0iu6);  // ../RTL/cortexm0ds_logic.v(6998)
  and u6453 (n1520, Eafpw6[11], A3iiu6);  // ../RTL/cortexm0ds_logic.v(6999)
  not u6454 (Mqmiu6, n1520);  // ../RTL/cortexm0ds_logic.v(6999)
  and u6455 (n1521, vis_pc_o[10], Ok8iu6);  // ../RTL/cortexm0ds_logic.v(7000)
  not u6456 (Kpmiu6, n1521);  // ../RTL/cortexm0ds_logic.v(7000)
  and u6457 (Womiu6, Armiu6, Hrmiu6);  // ../RTL/cortexm0ds_logic.v(7001)
  or u6458 (Hrmiu6, Lm8iu6, Ormiu6);  // ../RTL/cortexm0ds_logic.v(7002)
  and u6459 (n1522, Zm8iu6, Q44iu6);  // ../RTL/cortexm0ds_logic.v(7003)
  buf u646 (Ahghu6, Pdyax6);  // ../RTL/cortexm0ds_logic.v(2701)
  not u6460 (Armiu6, n1522);  // ../RTL/cortexm0ds_logic.v(7003)
  AL_MUX u6461 (
    .i0(vis_psp_o[9]),
    .i1(Vrmiu6),
    .sel(Ydkiu6),
    .o(O3qhu6));  // ../RTL/cortexm0ds_logic.v(7004)
  AL_MUX u6462 (
    .i0(vis_msp_o[9]),
    .i1(Vrmiu6),
    .sel(Fekiu6),
    .o(H3qhu6));  // ../RTL/cortexm0ds_logic.v(7005)
  AL_MUX u6463 (
    .i0(Vrmiu6),
    .i1(vis_r14_o[11]),
    .sel(Mekiu6),
    .o(A3qhu6));  // ../RTL/cortexm0ds_logic.v(7006)
  AL_MUX u6464 (
    .i0(Vrmiu6),
    .i1(vis_r12_o[11]),
    .sel(Tekiu6),
    .o(T2qhu6));  // ../RTL/cortexm0ds_logic.v(7007)
  not u6465 (Tekiu6, Csmiu6);  // ../RTL/cortexm0ds_logic.v(7008)
  AL_MUX u6466 (
    .i0(Vrmiu6),
    .i1(vis_r7_o[11]),
    .sel(Rdkiu6),
    .o(M2qhu6));  // ../RTL/cortexm0ds_logic.v(7009)
  not u6467 (Rdkiu6, Jsmiu6);  // ../RTL/cortexm0ds_logic.v(7010)
  AL_MUX u6468 (
    .i0(Vrmiu6),
    .i1(vis_r6_o[11]),
    .sel(Kdkiu6),
    .o(F2qhu6));  // ../RTL/cortexm0ds_logic.v(7011)
  AL_MUX u6469 (
    .i0(Vrmiu6),
    .i1(vis_r5_o[11]),
    .sel(Ddkiu6),
    .o(Y1qhu6));  // ../RTL/cortexm0ds_logic.v(7012)
  buf u647 (Togpw6[11], F59bx6);  // ../RTL/cortexm0ds_logic.v(2378)
  not u6470 (Ddkiu6, Qsmiu6);  // ../RTL/cortexm0ds_logic.v(7013)
  AL_MUX u6471 (
    .i0(Vrmiu6),
    .i1(vis_r4_o[11]),
    .sel(Wckiu6),
    .o(R1qhu6));  // ../RTL/cortexm0ds_logic.v(7014)
  not u6472 (Wckiu6, Xsmiu6);  // ../RTL/cortexm0ds_logic.v(7015)
  AL_MUX u6473 (
    .i0(Vrmiu6),
    .i1(vis_r11_o[11]),
    .sel(Afkiu6),
    .o(K1qhu6));  // ../RTL/cortexm0ds_logic.v(7016)
  not u6474 (Afkiu6, Etmiu6);  // ../RTL/cortexm0ds_logic.v(7017)
  AL_MUX u6475 (
    .i0(Vrmiu6),
    .i1(vis_r10_o[11]),
    .sel(Hfkiu6),
    .o(D1qhu6));  // ../RTL/cortexm0ds_logic.v(7018)
  AL_MUX u6476 (
    .i0(Vrmiu6),
    .i1(vis_r9_o[11]),
    .sel(Ofkiu6),
    .o(W0qhu6));  // ../RTL/cortexm0ds_logic.v(7019)
  not u6477 (Ofkiu6, Ltmiu6);  // ../RTL/cortexm0ds_logic.v(7020)
  AL_MUX u6478 (
    .i0(Vrmiu6),
    .i1(vis_r8_o[11]),
    .sel(Vfkiu6),
    .o(P0qhu6));  // ../RTL/cortexm0ds_logic.v(7021)
  not u6479 (Vfkiu6, Stmiu6);  // ../RTL/cortexm0ds_logic.v(7022)
  buf u648 (Togpw6[10], C4dax6);  // ../RTL/cortexm0ds_logic.v(2378)
  AL_MUX u6480 (
    .i0(Vrmiu6),
    .i1(vis_r3_o[11]),
    .sel(Pckiu6),
    .o(I0qhu6));  // ../RTL/cortexm0ds_logic.v(7023)
  not u6481 (Pckiu6, Ztmiu6);  // ../RTL/cortexm0ds_logic.v(7024)
  AL_MUX u6482 (
    .i0(Vrmiu6),
    .i1(vis_r2_o[11]),
    .sel(Ickiu6),
    .o(B0qhu6));  // ../RTL/cortexm0ds_logic.v(7025)
  AL_MUX u6483 (
    .i0(Vrmiu6),
    .i1(vis_r1_o[11]),
    .sel(Mx8iu6),
    .o(Uzphu6));  // ../RTL/cortexm0ds_logic.v(7026)
  not u6484 (Mx8iu6, Gumiu6);  // ../RTL/cortexm0ds_logic.v(7027)
  AL_MUX u6485 (
    .i0(Vrmiu6),
    .i1(vis_r0_o[11]),
    .sel(Lf8iu6),
    .o(Nzphu6));  // ../RTL/cortexm0ds_logic.v(7028)
  not u6486 (Lf8iu6, Numiu6);  // ../RTL/cortexm0ds_logic.v(7029)
  or u6487 (Vrmiu6, Uumiu6, Bvmiu6);  // ../RTL/cortexm0ds_logic.v(7030)
  and u6488 (n1523, Ivmiu6, Pvmiu6);  // ../RTL/cortexm0ds_logic.v(7031)
  not u6489 (Gzphu6, n1523);  // ../RTL/cortexm0ds_logic.v(7031)
  buf u649 (Togpw6[9], Tcjbx6);  // ../RTL/cortexm0ds_logic.v(2378)
  and u6490 (Pvmiu6, Wvmiu6, Dwmiu6);  // ../RTL/cortexm0ds_logic.v(7032)
  and u6491 (n1524, Jl8iu6, Tugpw6[8]);  // ../RTL/cortexm0ds_logic.v(7033)
  not u6492 (Dwmiu6, n1524);  // ../RTL/cortexm0ds_logic.v(7033)
  buf u6493 (vis_r7_o[8], Lzwax6);  // ../RTL/cortexm0ds_logic.v(2654)
  buf u6494 (vis_r7_o[20], Lhwax6);  // ../RTL/cortexm0ds_logic.v(2654)
  and u6495 (n1525, N5fpw6[9], Sdaiu6);  // ../RTL/cortexm0ds_logic.v(7035)
  not u6496 (Rwmiu6, n1525);  // ../RTL/cortexm0ds_logic.v(7035)
  and u6497 (Kwmiu6, Ywmiu6, Fxmiu6);  // ../RTL/cortexm0ds_logic.v(7036)
  or u6498 (Fxmiu6, T2iiu6, Zn0iu6);  // ../RTL/cortexm0ds_logic.v(7037)
  and u6499 (n1526, Eafpw6[10], A3iiu6);  // ../RTL/cortexm0ds_logic.v(7038)
  buf u65 (Yenhu6, B7lpw6);  // ../RTL/cortexm0ds_logic.v(1831)
  buf u650 (Togpw6[7], U7dax6);  // ../RTL/cortexm0ds_logic.v(2378)
  not u6500 (Ywmiu6, n1526);  // ../RTL/cortexm0ds_logic.v(7038)
  and u6501 (n1527, vis_pc_o[9], Ok8iu6);  // ../RTL/cortexm0ds_logic.v(7039)
  not u6502 (Wvmiu6, n1527);  // ../RTL/cortexm0ds_logic.v(7039)
  and u6503 (Ivmiu6, Mxmiu6, Txmiu6);  // ../RTL/cortexm0ds_logic.v(7040)
  or u6504 (Txmiu6, Lm8iu6, Aymiu6);  // ../RTL/cortexm0ds_logic.v(7041)
  and u6505 (n1528, Zm8iu6, J44iu6);  // ../RTL/cortexm0ds_logic.v(7042)
  not u6506 (Mxmiu6, n1528);  // ../RTL/cortexm0ds_logic.v(7042)
  AL_MUX u6507 (
    .i0(vis_psp_o[8]),
    .i1(Hymiu6),
    .sel(Ydkiu6),
    .o(Zyphu6));  // ../RTL/cortexm0ds_logic.v(7043)
  AL_MUX u6508 (
    .i0(vis_msp_o[8]),
    .i1(Hymiu6),
    .sel(Fekiu6),
    .o(Syphu6));  // ../RTL/cortexm0ds_logic.v(7044)
  AL_MUX u6509 (
    .i0(Hymiu6),
    .i1(vis_r14_o[10]),
    .sel(Mekiu6),
    .o(Lyphu6));  // ../RTL/cortexm0ds_logic.v(7045)
  buf u651 (Togpw6[6], Zl9bx6);  // ../RTL/cortexm0ds_logic.v(2378)
  AL_MUX u6510 (
    .i0(vis_r12_o[10]),
    .i1(Hymiu6),
    .sel(Csmiu6),
    .o(Eyphu6));  // ../RTL/cortexm0ds_logic.v(7046)
  AL_MUX u6511 (
    .i0(vis_r7_o[10]),
    .i1(Hymiu6),
    .sel(Jsmiu6),
    .o(Xxphu6));  // ../RTL/cortexm0ds_logic.v(7047)
  AL_MUX u6512 (
    .i0(Hymiu6),
    .i1(vis_r6_o[10]),
    .sel(Kdkiu6),
    .o(Qxphu6));  // ../RTL/cortexm0ds_logic.v(7048)
  AL_MUX u6513 (
    .i0(vis_r5_o[10]),
    .i1(Hymiu6),
    .sel(Qsmiu6),
    .o(Jxphu6));  // ../RTL/cortexm0ds_logic.v(7049)
  AL_MUX u6514 (
    .i0(vis_r4_o[10]),
    .i1(Hymiu6),
    .sel(Xsmiu6),
    .o(Cxphu6));  // ../RTL/cortexm0ds_logic.v(7050)
  AL_MUX u6515 (
    .i0(vis_r11_o[10]),
    .i1(Hymiu6),
    .sel(Etmiu6),
    .o(Vwphu6));  // ../RTL/cortexm0ds_logic.v(7051)
  AL_MUX u6516 (
    .i0(Hymiu6),
    .i1(vis_r10_o[10]),
    .sel(Hfkiu6),
    .o(Owphu6));  // ../RTL/cortexm0ds_logic.v(7052)
  AL_MUX u6517 (
    .i0(vis_r9_o[10]),
    .i1(Hymiu6),
    .sel(Ltmiu6),
    .o(Hwphu6));  // ../RTL/cortexm0ds_logic.v(7053)
  AL_MUX u6518 (
    .i0(vis_r8_o[10]),
    .i1(Hymiu6),
    .sel(Stmiu6),
    .o(Awphu6));  // ../RTL/cortexm0ds_logic.v(7054)
  AL_MUX u6519 (
    .i0(vis_r3_o[10]),
    .i1(Hymiu6),
    .sel(Ztmiu6),
    .o(Tvphu6));  // ../RTL/cortexm0ds_logic.v(7055)
  buf u652 (Togpw6[5], Q9dax6);  // ../RTL/cortexm0ds_logic.v(2378)
  AL_MUX u6520 (
    .i0(Hymiu6),
    .i1(vis_r2_o[10]),
    .sel(Ickiu6),
    .o(Mvphu6));  // ../RTL/cortexm0ds_logic.v(7056)
  AL_MUX u6521 (
    .i0(vis_r1_o[10]),
    .i1(Hymiu6),
    .sel(Gumiu6),
    .o(Fvphu6));  // ../RTL/cortexm0ds_logic.v(7057)
  AL_MUX u6522 (
    .i0(vis_r0_o[10]),
    .i1(Hymiu6),
    .sel(Numiu6),
    .o(Yuphu6));  // ../RTL/cortexm0ds_logic.v(7058)
  or u6523 (Hymiu6, Oymiu6, Vymiu6);  // ../RTL/cortexm0ds_logic.v(7059)
  AL_MUX u6524 (
    .i0(L8ehu6),
    .i1(Czmiu6),
    .sel(Jzmiu6),
    .o(Ruphu6));  // ../RTL/cortexm0ds_logic.v(7060)
  and u6525 (Jzmiu6, Qzmiu6, HREADY);  // ../RTL/cortexm0ds_logic.v(7061)
  and u6526 (Qzmiu6, Xzmiu6, E0niu6);  // ../RTL/cortexm0ds_logic.v(7062)
  or u6527 (E0niu6, L0niu6, Bi0iu6);  // ../RTL/cortexm0ds_logic.v(7063)
  AL_MUX u6528 (
    .i0(S0niu6),
    .i1(Gh0iu6),
    .sel(Uzaiu6),
    .o(Czmiu6));  // ../RTL/cortexm0ds_logic.v(7064)
  and u6529 (n1529, Z0niu6, G1niu6);  // ../RTL/cortexm0ds_logic.v(7065)
  buf u653 (Jshpw6[8], Ke1qw6);  // ../RTL/cortexm0ds_logic.v(2372)
  not u6530 (Kuphu6, n1529);  // ../RTL/cortexm0ds_logic.v(7065)
  and u6531 (G1niu6, N1niu6, U1niu6);  // ../RTL/cortexm0ds_logic.v(7066)
  and u6532 (n1530, vis_pc_o[8], Ok8iu6);  // ../RTL/cortexm0ds_logic.v(7067)
  not u6533 (U1niu6, n1530);  // ../RTL/cortexm0ds_logic.v(7067)
  and u6534 (N1niu6, B2niu6, I2niu6);  // ../RTL/cortexm0ds_logic.v(7068)
  and u6535 (n1531, P2niu6, L8ehu6);  // ../RTL/cortexm0ds_logic.v(7069)
  not u6536 (I2niu6, n1531);  // ../RTL/cortexm0ds_logic.v(7069)
  and u6537 (P2niu6, Ql8iu6, Gc5iu6);  // ../RTL/cortexm0ds_logic.v(7070)
  and u6538 (n1532, Jl8iu6, Tugpw6[7]);  // ../RTL/cortexm0ds_logic.v(7071)
  not u6539 (B2niu6, n1532);  // ../RTL/cortexm0ds_logic.v(7071)
  buf u654 (Jshpw6[6], Vn9bx6);  // ../RTL/cortexm0ds_logic.v(2372)
  and u6540 (Z0niu6, W2niu6, D3niu6);  // ../RTL/cortexm0ds_logic.v(7072)
  and u6541 (n1533, W29iu6, Fkfpw6[9]);  // ../RTL/cortexm0ds_logic.v(7073)
  not u6542 (D3niu6, n1533);  // ../RTL/cortexm0ds_logic.v(7073)
  and u6543 (n1534, Zm8iu6, Ym4iu6);  // ../RTL/cortexm0ds_logic.v(7074)
  not u6544 (W2niu6, n1534);  // ../RTL/cortexm0ds_logic.v(7074)
  AL_MUX u6545 (
    .i0(vis_psp_o[7]),
    .i1(K3niu6),
    .sel(Ydkiu6),
    .o(Duphu6));  // ../RTL/cortexm0ds_logic.v(7075)
  AL_MUX u6546 (
    .i0(vis_msp_o[7]),
    .i1(K3niu6),
    .sel(Fekiu6),
    .o(Wtphu6));  // ../RTL/cortexm0ds_logic.v(7076)
  AL_MUX u6547 (
    .i0(K3niu6),
    .i1(vis_r14_o[9]),
    .sel(Mekiu6),
    .o(Ptphu6));  // ../RTL/cortexm0ds_logic.v(7077)
  AL_MUX u6548 (
    .i0(vis_r12_o[9]),
    .i1(K3niu6),
    .sel(Csmiu6),
    .o(Itphu6));  // ../RTL/cortexm0ds_logic.v(7078)
  AL_MUX u6549 (
    .i0(vis_r7_o[9]),
    .i1(K3niu6),
    .sel(Jsmiu6),
    .o(Btphu6));  // ../RTL/cortexm0ds_logic.v(7079)
  buf u655 (Jshpw6[5], Bf3qw6);  // ../RTL/cortexm0ds_logic.v(2372)
  AL_MUX u6550 (
    .i0(K3niu6),
    .i1(vis_r6_o[9]),
    .sel(Kdkiu6),
    .o(Usphu6));  // ../RTL/cortexm0ds_logic.v(7080)
  AL_MUX u6551 (
    .i0(vis_r5_o[9]),
    .i1(K3niu6),
    .sel(Qsmiu6),
    .o(Nsphu6));  // ../RTL/cortexm0ds_logic.v(7081)
  AL_MUX u6552 (
    .i0(vis_r4_o[9]),
    .i1(K3niu6),
    .sel(Xsmiu6),
    .o(Gsphu6));  // ../RTL/cortexm0ds_logic.v(7082)
  AL_MUX u6553 (
    .i0(vis_r11_o[9]),
    .i1(K3niu6),
    .sel(Etmiu6),
    .o(Zrphu6));  // ../RTL/cortexm0ds_logic.v(7083)
  AL_MUX u6554 (
    .i0(K3niu6),
    .i1(vis_r10_o[9]),
    .sel(Hfkiu6),
    .o(Srphu6));  // ../RTL/cortexm0ds_logic.v(7084)
  AL_MUX u6555 (
    .i0(vis_r9_o[9]),
    .i1(K3niu6),
    .sel(Ltmiu6),
    .o(Lrphu6));  // ../RTL/cortexm0ds_logic.v(7085)
  AL_MUX u6556 (
    .i0(vis_r8_o[9]),
    .i1(K3niu6),
    .sel(Stmiu6),
    .o(Erphu6));  // ../RTL/cortexm0ds_logic.v(7086)
  AL_MUX u6557 (
    .i0(vis_r3_o[9]),
    .i1(K3niu6),
    .sel(Ztmiu6),
    .o(Xqphu6));  // ../RTL/cortexm0ds_logic.v(7087)
  AL_MUX u6558 (
    .i0(K3niu6),
    .i1(vis_r2_o[9]),
    .sel(Ickiu6),
    .o(Qqphu6));  // ../RTL/cortexm0ds_logic.v(7088)
  AL_MUX u6559 (
    .i0(vis_r1_o[9]),
    .i1(K3niu6),
    .sel(Gumiu6),
    .o(Jqphu6));  // ../RTL/cortexm0ds_logic.v(7089)
  not u656 (Pkhpw6[1], n101[1]);  // ../RTL/cortexm0ds_logic.v(3356)
  AL_MUX u6560 (
    .i0(vis_r0_o[9]),
    .i1(K3niu6),
    .sel(Numiu6),
    .o(Cqphu6));  // ../RTL/cortexm0ds_logic.v(7090)
  or u6561 (K3niu6, S0niu6, R3niu6);  // ../RTL/cortexm0ds_logic.v(7091)
  and u6562 (n1535, Y3niu6, F4niu6);  // ../RTL/cortexm0ds_logic.v(7092)
  not u6563 (Vpphu6, n1535);  // ../RTL/cortexm0ds_logic.v(7092)
  and u6564 (F4niu6, M4niu6, T4niu6);  // ../RTL/cortexm0ds_logic.v(7093)
  and u6565 (n1536, Jl8iu6, Tugpw6[6]);  // ../RTL/cortexm0ds_logic.v(7094)
  not u6566 (T4niu6, n1536);  // ../RTL/cortexm0ds_logic.v(7094)
  buf u6567 (vis_r7_o[10], Lxwax6);  // ../RTL/cortexm0ds_logic.v(2654)
  buf u6568 (vis_r7_o[22], T9fbx6);  // ../RTL/cortexm0ds_logic.v(2654)
  and u6569 (n1537, N5fpw6[7], Sdaiu6);  // ../RTL/cortexm0ds_logic.v(7096)
  buf u657 (Qqdhu6, G0zax6);  // ../RTL/cortexm0ds_logic.v(2712)
  not u6570 (H5niu6, n1537);  // ../RTL/cortexm0ds_logic.v(7096)
  and u6571 (A5niu6, O5niu6, V5niu6);  // ../RTL/cortexm0ds_logic.v(7097)
  or u6572 (V5niu6, T2iiu6, Ve0iu6);  // ../RTL/cortexm0ds_logic.v(7098)
  and u6573 (n1538, Eafpw6[8], A3iiu6);  // ../RTL/cortexm0ds_logic.v(7099)
  not u6574 (O5niu6, n1538);  // ../RTL/cortexm0ds_logic.v(7099)
  and u6575 (n1539, vis_pc_o[7], Ok8iu6);  // ../RTL/cortexm0ds_logic.v(7100)
  not u6576 (M4niu6, n1539);  // ../RTL/cortexm0ds_logic.v(7100)
  and u6577 (Y3niu6, C6niu6, J6niu6);  // ../RTL/cortexm0ds_logic.v(7101)
  or u6578 (J6niu6, Lm8iu6, Q6niu6);  // ../RTL/cortexm0ds_logic.v(7102)
  and u6579 (n1540, Zm8iu6, Pl4iu6);  // ../RTL/cortexm0ds_logic.v(7103)
  buf u658 (Ndghu6, I2zax6);  // ../RTL/cortexm0ds_logic.v(2713)
  not u6580 (C6niu6, n1540);  // ../RTL/cortexm0ds_logic.v(7103)
  AL_MUX u6581 (
    .i0(vis_psp_o[6]),
    .i1(X6niu6),
    .sel(Ydkiu6),
    .o(Opphu6));  // ../RTL/cortexm0ds_logic.v(7104)
  AL_MUX u6582 (
    .i0(vis_msp_o[6]),
    .i1(X6niu6),
    .sel(Fekiu6),
    .o(Hpphu6));  // ../RTL/cortexm0ds_logic.v(7105)
  AL_MUX u6583 (
    .i0(X6niu6),
    .i1(vis_r14_o[8]),
    .sel(Mekiu6),
    .o(Apphu6));  // ../RTL/cortexm0ds_logic.v(7106)
  AL_MUX u6584 (
    .i0(vis_r12_o[8]),
    .i1(X6niu6),
    .sel(Csmiu6),
    .o(Tophu6));  // ../RTL/cortexm0ds_logic.v(7107)
  AL_MUX u6585 (
    .i0(vis_r7_o[8]),
    .i1(X6niu6),
    .sel(Jsmiu6),
    .o(Mophu6));  // ../RTL/cortexm0ds_logic.v(7108)
  AL_MUX u6586 (
    .i0(X6niu6),
    .i1(vis_r6_o[8]),
    .sel(Kdkiu6),
    .o(Fophu6));  // ../RTL/cortexm0ds_logic.v(7109)
  AL_MUX u6587 (
    .i0(vis_r5_o[8]),
    .i1(X6niu6),
    .sel(Qsmiu6),
    .o(Ynphu6));  // ../RTL/cortexm0ds_logic.v(7110)
  AL_MUX u6588 (
    .i0(vis_r4_o[8]),
    .i1(X6niu6),
    .sel(Xsmiu6),
    .o(Rnphu6));  // ../RTL/cortexm0ds_logic.v(7111)
  AL_MUX u6589 (
    .i0(vis_r11_o[8]),
    .i1(X6niu6),
    .sel(Etmiu6),
    .o(Knphu6));  // ../RTL/cortexm0ds_logic.v(7112)
  buf u659 (Togpw6[19], Uscax6);  // ../RTL/cortexm0ds_logic.v(2378)
  AL_MUX u6590 (
    .i0(X6niu6),
    .i1(vis_r10_o[8]),
    .sel(Hfkiu6),
    .o(Dnphu6));  // ../RTL/cortexm0ds_logic.v(7113)
  AL_MUX u6591 (
    .i0(vis_r9_o[8]),
    .i1(X6niu6),
    .sel(Ltmiu6),
    .o(Wmphu6));  // ../RTL/cortexm0ds_logic.v(7114)
  AL_MUX u6592 (
    .i0(vis_r8_o[8]),
    .i1(X6niu6),
    .sel(Stmiu6),
    .o(Pmphu6));  // ../RTL/cortexm0ds_logic.v(7115)
  AL_MUX u6593 (
    .i0(vis_r3_o[8]),
    .i1(X6niu6),
    .sel(Ztmiu6),
    .o(Imphu6));  // ../RTL/cortexm0ds_logic.v(7116)
  AL_MUX u6594 (
    .i0(X6niu6),
    .i1(vis_r2_o[8]),
    .sel(Ickiu6),
    .o(Bmphu6));  // ../RTL/cortexm0ds_logic.v(7117)
  AL_MUX u6595 (
    .i0(vis_r1_o[8]),
    .i1(X6niu6),
    .sel(Gumiu6),
    .o(Ulphu6));  // ../RTL/cortexm0ds_logic.v(7118)
  AL_MUX u6596 (
    .i0(vis_r0_o[8]),
    .i1(X6niu6),
    .sel(Numiu6),
    .o(Nlphu6));  // ../RTL/cortexm0ds_logic.v(7119)
  or u6597 (X6niu6, E7niu6, L7niu6);  // ../RTL/cortexm0ds_logic.v(7120)
  and u6598 (n1541, S7niu6, Z7niu6);  // ../RTL/cortexm0ds_logic.v(7121)
  not u6599 (Glphu6, n1541);  // ../RTL/cortexm0ds_logic.v(7121)
  buf u66 (Hknhu6, Y8lpw6);  // ../RTL/cortexm0ds_logic.v(1832)
  buf u660 (Togpw6[18], Rucax6);  // ../RTL/cortexm0ds_logic.v(2378)
  and u6600 (n1542, G8niu6, Ug8iu6);  // ../RTL/cortexm0ds_logic.v(7122)
  not u6601 (Z7niu6, n1542);  // ../RTL/cortexm0ds_logic.v(7122)
  AL_MUX u6602 (
    .i0(N8niu6),
    .i1(U8niu6),
    .sel(HREADY),
    .o(S7niu6));  // ../RTL/cortexm0ds_logic.v(7123)
  and u6603 (n1543, B9niu6, I9niu6);  // ../RTL/cortexm0ds_logic.v(7124)
  not u6604 (U8niu6, n1543);  // ../RTL/cortexm0ds_logic.v(7124)
  and u6605 (n1544, P9niu6, Ug8iu6);  // ../RTL/cortexm0ds_logic.v(7125)
  not u6606 (I9niu6, n1544);  // ../RTL/cortexm0ds_logic.v(7125)
  AL_MUX u6607 (
    .i0(W9niu6),
    .i1(Daniu6),
    .sel(Ug8iu6),
    .o(B9niu6));  // ../RTL/cortexm0ds_logic.v(7126)
  and u6608 (Daniu6, Kaniu6, Raniu6);  // ../RTL/cortexm0ds_logic.v(7127)
  and u6609 (n1545, Idfpw6[31], Eafpw6[31]);  // ../RTL/cortexm0ds_logic.v(7128)
  buf u661 (Togpw6[17], Btbbx6);  // ../RTL/cortexm0ds_logic.v(2378)
  not u6610 (Raniu6, n1545);  // ../RTL/cortexm0ds_logic.v(7128)
  AL_MUX u6611 (
    .i0(Eafpw6[31]),
    .i1(Idfpw6[31]),
    .sel(D5epw6),
    .o(Kaniu6));  // ../RTL/cortexm0ds_logic.v(7129)
  and u6612 (W9niu6, Yaniu6, Fbniu6);  // ../RTL/cortexm0ds_logic.v(7130)
  and u6613 (n1546, Mbniu6, Tbniu6);  // ../RTL/cortexm0ds_logic.v(7131)
  not u6614 (Fbniu6, n1546);  // ../RTL/cortexm0ds_logic.v(7131)
  or u6615 (Tbniu6, Cs8iu6, Acniu6);  // ../RTL/cortexm0ds_logic.v(7132)
  and u6616 (n1547, Acniu6, Hcniu6);  // ../RTL/cortexm0ds_logic.v(7133)
  not u6617 (Yaniu6, n1547);  // ../RTL/cortexm0ds_logic.v(7133)
  not u6618 (N8niu6, vis_apsr_o[0]);  // ../RTL/cortexm0ds_logic.v(7134)
  and u6619 (n1548, Ocniu6, Vcniu6);  // ../RTL/cortexm0ds_logic.v(7135)
  buf u662 (Togpw6[15], Lycax6);  // ../RTL/cortexm0ds_logic.v(2378)
  not u6620 (Zkphu6, n1548);  // ../RTL/cortexm0ds_logic.v(7135)
  and u6621 (Vcniu6, Cdniu6, Jdniu6);  // ../RTL/cortexm0ds_logic.v(7136)
  and u6622 (n1549, Ok8iu6, vis_pc_o[27]);  // ../RTL/cortexm0ds_logic.v(7137)
  not u6623 (Jdniu6, n1549);  // ../RTL/cortexm0ds_logic.v(7137)
  and u6624 (Cdniu6, Qdniu6, Xdniu6);  // ../RTL/cortexm0ds_logic.v(7138)
  and u6625 (n1550, Jl8iu6, V0epw6);  // ../RTL/cortexm0ds_logic.v(7139)
  not u6626 (Xdniu6, n1550);  // ../RTL/cortexm0ds_logic.v(7139)
  and u6627 (n1551, vis_apsr_o[0], Ql8iu6);  // ../RTL/cortexm0ds_logic.v(7140)
  not u6628 (Qdniu6, n1551);  // ../RTL/cortexm0ds_logic.v(7140)
  and u6629 (Ocniu6, Eeniu6, Leniu6);  // ../RTL/cortexm0ds_logic.v(7141)
  buf u663 (Togpw6[14], Buabx6);  // ../RTL/cortexm0ds_logic.v(2378)
  or u6630 (Leniu6, Lm8iu6, Seniu6);  // ../RTL/cortexm0ds_logic.v(7142)
  or u6631 (Eeniu6, Hx9iu6, Zeniu6);  // ../RTL/cortexm0ds_logic.v(7143)
  AL_MUX u6632 (
    .i0(vis_psp_o[26]),
    .i1(Gfniu6),
    .sel(Ydkiu6),
    .o(Skphu6));  // ../RTL/cortexm0ds_logic.v(7144)
  and u6633 (Ydkiu6, Nfniu6, Vrfhu6);  // ../RTL/cortexm0ds_logic.v(7145)
  AL_MUX u6634 (
    .i0(vis_msp_o[26]),
    .i1(Gfniu6),
    .sel(Fekiu6),
    .o(Lkphu6));  // ../RTL/cortexm0ds_logic.v(7147)
  or u6635 (n1552, Ufniu6, Vrfhu6);  // ../RTL/cortexm0ds_logic.v(7148)
  not u6636 (Fekiu6, n1552);  // ../RTL/cortexm0ds_logic.v(7148)
  and u6637 (Nfniu6, Bgniu6, Igniu6);  // ../RTL/cortexm0ds_logic.v(7149)
  not u6638 (Ufniu6, Nfniu6);  // ../RTL/cortexm0ds_logic.v(7149)
  or u6639 (n1553, Pgniu6, Wgniu6);  // ../RTL/cortexm0ds_logic.v(7150)
  buf u664 (Togpw6[13], I0dax6);  // ../RTL/cortexm0ds_logic.v(2378)
  not u6640 (Bgniu6, n1553);  // ../RTL/cortexm0ds_logic.v(7150)
  AL_MUX u6641 (
    .i0(Gfniu6),
    .i1(vis_r14_o[28]),
    .sel(Mekiu6),
    .o(Ekphu6));  // ../RTL/cortexm0ds_logic.v(7151)
  and u6642 (n1554, Dhniu6, Khniu6);  // ../RTL/cortexm0ds_logic.v(7152)
  not u6643 (Mekiu6, n1554);  // ../RTL/cortexm0ds_logic.v(7152)
  AL_MUX u6644 (
    .i0(vis_r12_o[28]),
    .i1(Gfniu6),
    .sel(Csmiu6),
    .o(Xjphu6));  // ../RTL/cortexm0ds_logic.v(7153)
  and u6645 (Csmiu6, Rhniu6, Khniu6);  // ../RTL/cortexm0ds_logic.v(7154)
  or u6646 (n1555, Yhniu6, Wgniu6);  // ../RTL/cortexm0ds_logic.v(7155)
  not u6647 (Rhniu6, n1555);  // ../RTL/cortexm0ds_logic.v(7155)
  AL_MUX u6648 (
    .i0(vis_r7_o[28]),
    .i1(Gfniu6),
    .sel(Jsmiu6),
    .o(Qjphu6));  // ../RTL/cortexm0ds_logic.v(7156)
  and u6649 (Jsmiu6, Finiu6, Miniu6);  // ../RTL/cortexm0ds_logic.v(7157)
  buf u665 (Jshpw6[12], Su8ax6);  // ../RTL/cortexm0ds_logic.v(2372)
  and u6650 (Finiu6, Tiniu6, Ajniu6);  // ../RTL/cortexm0ds_logic.v(7158)
  AL_MUX u6651 (
    .i0(Gfniu6),
    .i1(vis_r6_o[28]),
    .sel(Kdkiu6),
    .o(Jjphu6));  // ../RTL/cortexm0ds_logic.v(7159)
  and u6652 (n1556, Khniu6, Miniu6);  // ../RTL/cortexm0ds_logic.v(7160)
  not u6653 (Kdkiu6, n1556);  // ../RTL/cortexm0ds_logic.v(7160)
  AL_MUX u6654 (
    .i0(vis_r5_o[28]),
    .i1(Gfniu6),
    .sel(Qsmiu6),
    .o(Cjphu6));  // ../RTL/cortexm0ds_logic.v(7161)
  and u6655 (Qsmiu6, Hjniu6, Igniu6);  // ../RTL/cortexm0ds_logic.v(7162)
  or u6656 (n1557, Ojniu6, Pgniu6);  // ../RTL/cortexm0ds_logic.v(7163)
  not u6657 (Hjniu6, n1557);  // ../RTL/cortexm0ds_logic.v(7163)
  AL_MUX u6658 (
    .i0(vis_r4_o[28]),
    .i1(Gfniu6),
    .sel(Xsmiu6),
    .o(Viphu6));  // ../RTL/cortexm0ds_logic.v(7164)
  and u6659 (Xsmiu6, Vjniu6, Khniu6);  // ../RTL/cortexm0ds_logic.v(7165)
  buf u666 (Jshpw6[13], Kl8ax6);  // ../RTL/cortexm0ds_logic.v(2372)
  or u6660 (n1558, Ajniu6, Pgniu6);  // ../RTL/cortexm0ds_logic.v(7166)
  not u6661 (Khniu6, n1558);  // ../RTL/cortexm0ds_logic.v(7166)
  or u6662 (n1559, Yhniu6, Ojniu6);  // ../RTL/cortexm0ds_logic.v(7167)
  not u6663 (Vjniu6, n1559);  // ../RTL/cortexm0ds_logic.v(7167)
  AL_MUX u6664 (
    .i0(vis_r11_o[28]),
    .i1(Gfniu6),
    .sel(Etmiu6),
    .o(Oiphu6));  // ../RTL/cortexm0ds_logic.v(7168)
  and u6665 (Etmiu6, Ckniu6, Dhniu6);  // ../RTL/cortexm0ds_logic.v(7169)
  AL_MUX u6666 (
    .i0(Gfniu6),
    .i1(vis_r10_o[28]),
    .sel(Hfkiu6),
    .o(Hiphu6));  // ../RTL/cortexm0ds_logic.v(7170)
  and u6667 (n1560, Dhniu6, Jkniu6);  // ../RTL/cortexm0ds_logic.v(7171)
  not u6668 (Hfkiu6, n1560);  // ../RTL/cortexm0ds_logic.v(7171)
  or u6669 (n1561, Wgniu6, Qkniu6);  // ../RTL/cortexm0ds_logic.v(7172)
  buf u667 (Jshpw6[14], Yvabx6);  // ../RTL/cortexm0ds_logic.v(2372)
  not u6670 (Dhniu6, n1561);  // ../RTL/cortexm0ds_logic.v(7172)
  AL_MUX u6671 (
    .i0(vis_r9_o[28]),
    .i1(Gfniu6),
    .sel(Ltmiu6),
    .o(Aiphu6));  // ../RTL/cortexm0ds_logic.v(7173)
  and u6672 (Ltmiu6, Xkniu6, Igniu6);  // ../RTL/cortexm0ds_logic.v(7174)
  or u6673 (n1562, Tiniu6, Wgniu6);  // ../RTL/cortexm0ds_logic.v(7175)
  not u6674 (Xkniu6, n1562);  // ../RTL/cortexm0ds_logic.v(7175)
  AL_MUX u6675 (
    .i0(vis_r8_o[28]),
    .i1(Gfniu6),
    .sel(Stmiu6),
    .o(Thphu6));  // ../RTL/cortexm0ds_logic.v(7176)
  and u6676 (Stmiu6, Elniu6, Qkniu6);  // ../RTL/cortexm0ds_logic.v(7177)
  and u6677 (Elniu6, Jkniu6, Ojniu6);  // ../RTL/cortexm0ds_logic.v(7178)
  AL_MUX u6678 (
    .i0(vis_r3_o[28]),
    .i1(Gfniu6),
    .sel(Ztmiu6),
    .o(Mhphu6));  // ../RTL/cortexm0ds_logic.v(7179)
  and u6679 (Ztmiu6, Ckniu6, Miniu6);  // ../RTL/cortexm0ds_logic.v(7180)
  buf u668 (Jshpw6[16], Dpwpw6);  // ../RTL/cortexm0ds_logic.v(2372)
  and u6680 (Ckniu6, Pgniu6, Ajniu6);  // ../RTL/cortexm0ds_logic.v(7181)
  AL_MUX u6681 (
    .i0(Gfniu6),
    .i1(vis_r2_o[28]),
    .sel(Ickiu6),
    .o(Fhphu6));  // ../RTL/cortexm0ds_logic.v(7183)
  and u6682 (n1563, Miniu6, Jkniu6);  // ../RTL/cortexm0ds_logic.v(7184)
  not u6683 (Ickiu6, n1563);  // ../RTL/cortexm0ds_logic.v(7184)
  or u6684 (n1564, Ojniu6, Qkniu6);  // ../RTL/cortexm0ds_logic.v(7185)
  not u6685 (Miniu6, n1564);  // ../RTL/cortexm0ds_logic.v(7185)
  AL_MUX u6686 (
    .i0(vis_r1_o[28]),
    .i1(Gfniu6),
    .sel(Gumiu6),
    .o(Ygphu6));  // ../RTL/cortexm0ds_logic.v(7186)
  and u6687 (Gumiu6, Llniu6, Igniu6);  // ../RTL/cortexm0ds_logic.v(7187)
  and u6688 (Igniu6, Qkniu6, Ajniu6);  // ../RTL/cortexm0ds_logic.v(7188)
  or u6689 (n1565, Ojniu6, Tiniu6);  // ../RTL/cortexm0ds_logic.v(7189)
  buf u669 (Jshpw6[17], Yubbx6);  // ../RTL/cortexm0ds_logic.v(2372)
  not u6690 (Llniu6, n1565);  // ../RTL/cortexm0ds_logic.v(7189)
  AL_MUX u6691 (
    .i0(vis_r0_o[28]),
    .i1(Gfniu6),
    .sel(Numiu6),
    .o(Rgphu6));  // ../RTL/cortexm0ds_logic.v(7190)
  and u6692 (Numiu6, Slniu6, Qkniu6);  // ../RTL/cortexm0ds_logic.v(7191)
  not u6693 (Qkniu6, Yhniu6);  // ../RTL/cortexm0ds_logic.v(7192)
  or u6694 (Yhniu6, Zlniu6, Gmniu6);  // ../RTL/cortexm0ds_logic.v(7193)
  and u6695 (n1566, HREADY, Nmniu6);  // ../RTL/cortexm0ds_logic.v(7194)
  not u6696 (Zlniu6, n1566);  // ../RTL/cortexm0ds_logic.v(7194)
  and u6697 (Slniu6, Wgniu6, Jkniu6);  // ../RTL/cortexm0ds_logic.v(7195)
  or u6698 (n1567, Ajniu6, Tiniu6);  // ../RTL/cortexm0ds_logic.v(7196)
  not u6699 (Jkniu6, n1567);  // ../RTL/cortexm0ds_logic.v(7196)
  buf u67 (vis_r5_o[1], Plypw6);  // ../RTL/cortexm0ds_logic.v(1909)
  buf u670 (Jshpw6[18], Jl3qw6);  // ../RTL/cortexm0ds_logic.v(2372)
  and u6700 (Pgniu6, Umniu6, Bnniu6);  // ../RTL/cortexm0ds_logic.v(7197)
  not u6701 (Tiniu6, Pgniu6);  // ../RTL/cortexm0ds_logic.v(7197)
  and u6702 (Bnniu6, Inniu6, Pnniu6);  // ../RTL/cortexm0ds_logic.v(7198)
  and u6703 (n1568, S8fpw6[10], Wnniu6);  // ../RTL/cortexm0ds_logic.v(7199)
  not u6704 (Pnniu6, n1568);  // ../RTL/cortexm0ds_logic.v(7199)
  and u6705 (Inniu6, Doniu6, Koniu6);  // ../RTL/cortexm0ds_logic.v(7200)
  or u6706 (Koniu6, Roniu6, Yoniu6);  // ../RTL/cortexm0ds_logic.v(7201)
  or u6707 (Doniu6, Fpniu6, Mpniu6);  // ../RTL/cortexm0ds_logic.v(7202)
  and u6708 (n1569, Tpniu6, Aqniu6);  // ../RTL/cortexm0ds_logic.v(7203)
  not u6709 (Ajniu6, n1569);  // ../RTL/cortexm0ds_logic.v(7203)
  buf u671 (Bxghu6, Zszax6);  // ../RTL/cortexm0ds_logic.v(2726)
  and u6710 (Aqniu6, Hqniu6, Oqniu6);  // ../RTL/cortexm0ds_logic.v(7204)
  or u6711 (Oqniu6, Vqniu6, Mpniu6);  // ../RTL/cortexm0ds_logic.v(7205)
  and u6712 (n1570, S8fpw6[8], Wnniu6);  // ../RTL/cortexm0ds_logic.v(7206)
  not u6713 (Hqniu6, n1570);  // ../RTL/cortexm0ds_logic.v(7206)
  and u6714 (Tpniu6, Crniu6, Jrniu6);  // ../RTL/cortexm0ds_logic.v(7207)
  or u6715 (Jrniu6, Qrniu6, Yoniu6);  // ../RTL/cortexm0ds_logic.v(7208)
  and u6716 (Wgniu6, Umniu6, Xrniu6);  // ../RTL/cortexm0ds_logic.v(7210)
  not u6717 (Ojniu6, Wgniu6);  // ../RTL/cortexm0ds_logic.v(7210)
  and u6718 (Xrniu6, Esniu6, Lsniu6);  // ../RTL/cortexm0ds_logic.v(7211)
  or u6719 (Lsniu6, Ssniu6, Mpniu6);  // ../RTL/cortexm0ds_logic.v(7212)
  buf u672 (Dvghu6, Avzax6);  // ../RTL/cortexm0ds_logic.v(2727)
  and u6720 (Esniu6, Zsniu6, Gtniu6);  // ../RTL/cortexm0ds_logic.v(7213)
  and u6721 (n1571, S8fpw6[11], Wnniu6);  // ../RTL/cortexm0ds_logic.v(7214)
  not u6722 (Gtniu6, n1571);  // ../RTL/cortexm0ds_logic.v(7214)
  or u6723 (Zsniu6, Ntniu6, Yoniu6);  // ../RTL/cortexm0ds_logic.v(7215)
  and u6724 (Umniu6, Crniu6, Utniu6);  // ../RTL/cortexm0ds_logic.v(7216)
  and u6725 (Crniu6, Buniu6, HREADY);  // ../RTL/cortexm0ds_logic.v(7217)
  and u6726 (Buniu6, Nmniu6, Iuniu6);  // ../RTL/cortexm0ds_logic.v(7218)
  and u6727 (n1572, Puniu6, Wuniu6);  // ../RTL/cortexm0ds_logic.v(7219)
  not u6728 (Nmniu6, n1572);  // ../RTL/cortexm0ds_logic.v(7219)
  and u6729 (Wuniu6, Dvniu6, Kvniu6);  // ../RTL/cortexm0ds_logic.v(7220)
  not u673 (Tugpw6[8], n1272[8]);  // ../RTL/cortexm0ds_logic.v(16030)
  and u6730 (Kvniu6, Rvniu6, Yvniu6);  // ../RTL/cortexm0ds_logic.v(7221)
  and u6731 (n1573, Fwniu6, Toaiu6);  // ../RTL/cortexm0ds_logic.v(7222)
  not u6732 (Yvniu6, n1573);  // ../RTL/cortexm0ds_logic.v(7222)
  or u6733 (n1574, Knaiu6, Cyfpw6[4]);  // ../RTL/cortexm0ds_logic.v(7223)
  not u6734 (Fwniu6, n1574);  // ../RTL/cortexm0ds_logic.v(7223)
  and u6735 (Rvniu6, Mwniu6, Twniu6);  // ../RTL/cortexm0ds_logic.v(7224)
  and u6736 (Dvniu6, Axniu6, Hxniu6);  // ../RTL/cortexm0ds_logic.v(7225)
  and u6737 (n1575, Oxniu6, Vxniu6);  // ../RTL/cortexm0ds_logic.v(7226)
  not u6738 (Hxniu6, n1575);  // ../RTL/cortexm0ds_logic.v(7226)
  and u6739 (Axniu6, Cyniu6, Jyniu6);  // ../RTL/cortexm0ds_logic.v(7227)
  not u674 (Tugpw6[4], n1272[4]);  // ../RTL/cortexm0ds_logic.v(16030)
  and u6740 (n1576, Qyniu6, Xyniu6);  // ../RTL/cortexm0ds_logic.v(7228)
  not u6741 (Jyniu6, n1576);  // ../RTL/cortexm0ds_logic.v(7228)
  and u6742 (n1577, Ezniu6, Lzniu6);  // ../RTL/cortexm0ds_logic.v(7229)
  not u6743 (Xyniu6, n1577);  // ../RTL/cortexm0ds_logic.v(7229)
  or u6744 (Lzniu6, Szniu6, Nlaiu6);  // ../RTL/cortexm0ds_logic.v(7230)
  and u6745 (n1578, Zzniu6, Pugiu6);  // ../RTL/cortexm0ds_logic.v(7231)
  not u6746 (Cyniu6, n1578);  // ../RTL/cortexm0ds_logic.v(7231)
  and u6747 (Puniu6, G0oiu6, N0oiu6);  // ../RTL/cortexm0ds_logic.v(7232)
  and u6748 (N0oiu6, U0oiu6, B1oiu6);  // ../RTL/cortexm0ds_logic.v(7233)
  and u6749 (n1579, Y0jiu6, Wp0iu6);  // ../RTL/cortexm0ds_logic.v(7234)
  not u675 (Tugpw6[2], n1272[2]);  // ../RTL/cortexm0ds_logic.v(16030)
  not u6750 (B1oiu6, n1579);  // ../RTL/cortexm0ds_logic.v(7234)
  and u6751 (U0oiu6, I1oiu6, P1oiu6);  // ../RTL/cortexm0ds_logic.v(7235)
  and u6752 (n1580, W1oiu6, Geaiu6);  // ../RTL/cortexm0ds_logic.v(7236)
  not u6753 (P1oiu6, n1580);  // ../RTL/cortexm0ds_logic.v(7236)
  and u6754 (n1581, D2oiu6, K2oiu6);  // ../RTL/cortexm0ds_logic.v(7237)
  not u6755 (W1oiu6, n1581);  // ../RTL/cortexm0ds_logic.v(7237)
  and u6756 (n1582, R2oiu6, Fd0iu6);  // ../RTL/cortexm0ds_logic.v(7238)
  not u6757 (K2oiu6, n1582);  // ../RTL/cortexm0ds_logic.v(7238)
  or u6758 (n1583, Y2oiu6, Knaiu6);  // ../RTL/cortexm0ds_logic.v(7239)
  not u6759 (R2oiu6, n1583);  // ../RTL/cortexm0ds_logic.v(7239)
  not u676 (Tugpw6[1], n1272[1]);  // ../RTL/cortexm0ds_logic.v(16030)
  and u6760 (D2oiu6, F3oiu6, M3oiu6);  // ../RTL/cortexm0ds_logic.v(7240)
  and u6761 (n1584, T3oiu6, Md0iu6);  // ../RTL/cortexm0ds_logic.v(7241)
  not u6762 (M3oiu6, n1584);  // ../RTL/cortexm0ds_logic.v(7241)
  or u6763 (n1585, A4oiu6, Y7ghu6);  // ../RTL/cortexm0ds_logic.v(7242)
  not u6764 (T3oiu6, n1585);  // ../RTL/cortexm0ds_logic.v(7242)
  and u6765 (n1586, H4oiu6, O4oiu6);  // ../RTL/cortexm0ds_logic.v(7243)
  not u6766 (F3oiu6, n1586);  // ../RTL/cortexm0ds_logic.v(7243)
  and u6767 (n1587, Imaiu6, V4oiu6);  // ../RTL/cortexm0ds_logic.v(7244)
  not u6768 (I1oiu6, n1587);  // ../RTL/cortexm0ds_logic.v(7244)
  and u6769 (n1588, C5oiu6, J5oiu6);  // ../RTL/cortexm0ds_logic.v(7245)
  buf u677 (Gtgpw6[27], Cxcbx6);  // ../RTL/cortexm0ds_logic.v(2375)
  not u6770 (V4oiu6, n1588);  // ../RTL/cortexm0ds_logic.v(7245)
  and u6771 (J5oiu6, Q5oiu6, X5oiu6);  // ../RTL/cortexm0ds_logic.v(7246)
  and u6772 (n1589, E6oiu6, Cyfpw6[4]);  // ../RTL/cortexm0ds_logic.v(7247)
  not u6773 (Q5oiu6, n1589);  // ../RTL/cortexm0ds_logic.v(7247)
  and u6774 (C5oiu6, L6oiu6, S6oiu6);  // ../RTL/cortexm0ds_logic.v(7248)
  and u6775 (n1590, Pthiu6, Cyfpw6[7]);  // ../RTL/cortexm0ds_logic.v(7249)
  not u6776 (S6oiu6, n1590);  // ../RTL/cortexm0ds_logic.v(7249)
  AL_MUX u6777 (
    .i0(Z6oiu6),
    .i1(G7oiu6),
    .sel(Tr0iu6),
    .o(L6oiu6));  // ../RTL/cortexm0ds_logic.v(7250)
  and u6778 (G0oiu6, N7oiu6, U7oiu6);  // ../RTL/cortexm0ds_logic.v(7251)
  AL_MUX u6779 (
    .i0(B8oiu6),
    .i1(I8oiu6),
    .sel(Cyfpw6[6]),
    .o(U7oiu6));  // ../RTL/cortexm0ds_logic.v(7252)
  buf u678 (Gtgpw6[26], Zdcbx6);  // ../RTL/cortexm0ds_logic.v(2375)
  and u6780 (n1591, P8oiu6, Zraiu6);  // ../RTL/cortexm0ds_logic.v(7253)
  not u6781 (I8oiu6, n1591);  // ../RTL/cortexm0ds_logic.v(7253)
  or u6782 (B8oiu6, W8oiu6, D9oiu6);  // ../RTL/cortexm0ds_logic.v(7254)
  and u6783 (N7oiu6, K9oiu6, R9oiu6);  // ../RTL/cortexm0ds_logic.v(7255)
  and u6784 (n1592, Pthiu6, Mfjiu6);  // ../RTL/cortexm0ds_logic.v(7256)
  not u6785 (R9oiu6, n1592);  // ../RTL/cortexm0ds_logic.v(7256)
  AL_MUX u6786 (
    .i0(Y9oiu6),
    .i1(Faoiu6),
    .sel(H4ghu6),
    .o(K9oiu6));  // ../RTL/cortexm0ds_logic.v(7257)
  and u6787 (Faoiu6, Maoiu6, Taoiu6);  // ../RTL/cortexm0ds_logic.v(7258)
  and u6788 (n1593, Whfiu6, Pthiu6);  // ../RTL/cortexm0ds_logic.v(7259)
  not u6789 (Taoiu6, n1593);  // ../RTL/cortexm0ds_logic.v(7259)
  buf u679 (Gtgpw6[25], Htbax6);  // ../RTL/cortexm0ds_logic.v(2375)
  and u6790 (Maoiu6, Aboiu6, Hboiu6);  // ../RTL/cortexm0ds_logic.v(7260)
  and u6791 (n1594, Oboiu6, Vboiu6);  // ../RTL/cortexm0ds_logic.v(7261)
  not u6792 (Hboiu6, n1594);  // ../RTL/cortexm0ds_logic.v(7261)
  or u6793 (n1595, Ccoiu6, Qxaiu6);  // ../RTL/cortexm0ds_logic.v(7262)
  not u6794 (Oboiu6, n1595);  // ../RTL/cortexm0ds_logic.v(7262)
  and u6795 (n1596, Pugiu6, Jcoiu6);  // ../RTL/cortexm0ds_logic.v(7263)
  not u6796 (Aboiu6, n1596);  // ../RTL/cortexm0ds_logic.v(7263)
  and u6797 (n1597, Qcoiu6, Xcoiu6);  // ../RTL/cortexm0ds_logic.v(7264)
  not u6798 (Jcoiu6, n1597);  // ../RTL/cortexm0ds_logic.v(7264)
  and u6799 (n1598, Edoiu6, Ldoiu6);  // ../RTL/cortexm0ds_logic.v(7265)
  buf u68 (vis_r5_o[3], Nbppw6);  // ../RTL/cortexm0ds_logic.v(1909)
  buf u680 (Gtgpw6[24], Evbax6);  // ../RTL/cortexm0ds_logic.v(2375)
  not u6800 (Xcoiu6, n1598);  // ../RTL/cortexm0ds_logic.v(7265)
  or u6801 (n1599, Jcaiu6, Ii0iu6);  // ../RTL/cortexm0ds_logic.v(7266)
  not u6802 (Edoiu6, n1599);  // ../RTL/cortexm0ds_logic.v(7266)
  and u6803 (Y9oiu6, Sdoiu6, Zdoiu6);  // ../RTL/cortexm0ds_logic.v(7267)
  and u6804 (n1600, Geoiu6, Neoiu6);  // ../RTL/cortexm0ds_logic.v(7268)
  not u6805 (Zdoiu6, n1600);  // ../RTL/cortexm0ds_logic.v(7268)
  and u6806 (Sdoiu6, Ueoiu6, Bfoiu6);  // ../RTL/cortexm0ds_logic.v(7269)
  and u6807 (n1601, Ifoiu6, Pfoiu6);  // ../RTL/cortexm0ds_logic.v(7270)
  not u6808 (Bfoiu6, n1601);  // ../RTL/cortexm0ds_logic.v(7270)
  or u6809 (n1602, Wfoiu6, Y7ghu6);  // ../RTL/cortexm0ds_logic.v(7271)
  buf u681 (Gtgpw6[23], Tzgbx6);  // ../RTL/cortexm0ds_logic.v(2375)
  not u6810 (Ifoiu6, n1602);  // ../RTL/cortexm0ds_logic.v(7271)
  and u6811 (n1603, Dgoiu6, Fd0iu6);  // ../RTL/cortexm0ds_logic.v(7272)
  not u6812 (Ueoiu6, n1603);  // ../RTL/cortexm0ds_logic.v(7272)
  or u6813 (n1604, Ezniu6, Cyfpw6[4]);  // ../RTL/cortexm0ds_logic.v(7273)
  not u6814 (Dgoiu6, n1604);  // ../RTL/cortexm0ds_logic.v(7273)
  and u6815 (n1605, Acniu6, Kgoiu6);  // ../RTL/cortexm0ds_logic.v(7274)
  not u6816 (Gfniu6, n1605);  // ../RTL/cortexm0ds_logic.v(7274)
  AL_MUX u6817 (
    .i0(vis_apsr_o[3]),
    .i1(Rgoiu6),
    .sel(Y5liu6),
    .o(Kgphu6));  // ../RTL/cortexm0ds_logic.v(7275)
  and u6818 (Y5liu6, HREADY, Ygoiu6);  // ../RTL/cortexm0ds_logic.v(7276)
  and u6819 (n1606, Fhoiu6, Ug8iu6);  // ../RTL/cortexm0ds_logic.v(7277)
  buf u682 (Gtgpw6[22], Nnfbx6);  // ../RTL/cortexm0ds_logic.v(2375)
  not u6820 (Ygoiu6, n1606);  // ../RTL/cortexm0ds_logic.v(7277)
  and u6821 (n1607, Mhoiu6, Thoiu6);  // ../RTL/cortexm0ds_logic.v(7278)
  not u6822 (Rgoiu6, n1607);  // ../RTL/cortexm0ds_logic.v(7278)
  and u6823 (n1608, Ph8iu6, Aioiu6);  // ../RTL/cortexm0ds_logic.v(7279)
  not u6824 (Thoiu6, n1608);  // ../RTL/cortexm0ds_logic.v(7279)
  and u6825 (Mhoiu6, Hioiu6, Oioiu6);  // ../RTL/cortexm0ds_logic.v(7280)
  or u6826 (Oioiu6, O7liu6, Vioiu6);  // ../RTL/cortexm0ds_logic.v(7281)
  or u6827 (O7liu6, Ph8iu6, Yi8iu6);  // ../RTL/cortexm0ds_logic.v(7283)
  not u6828 (Ug8iu6, O7liu6);  // ../RTL/cortexm0ds_logic.v(7283)
  not u6829 (Yi8iu6, Cs8iu6);  // ../RTL/cortexm0ds_logic.v(7284)
  buf u683 (Gtgpw6[21], G8ebx6);  // ../RTL/cortexm0ds_logic.v(2375)
  not u6830 (Ph8iu6, Hcniu6);  // ../RTL/cortexm0ds_logic.v(7285)
  and u6831 (Hcniu6, Cjoiu6, Vr8iu6);  // ../RTL/cortexm0ds_logic.v(7286)
  and u6832 (n1609, Jjoiu6, Wofiu6);  // ../RTL/cortexm0ds_logic.v(7287)
  not u6833 (Vr8iu6, n1609);  // ../RTL/cortexm0ds_logic.v(7287)
  and u6834 (n1610, Jjoiu6, Qjoiu6);  // ../RTL/cortexm0ds_logic.v(7288)
  not u6835 (Cjoiu6, n1610);  // ../RTL/cortexm0ds_logic.v(7288)
  or u6836 (Hioiu6, Cs8iu6, Ualiu6);  // ../RTL/cortexm0ds_logic.v(7289)
  or u6837 (Cs8iu6, Mjfiu6, Uzaiu6);  // ../RTL/cortexm0ds_logic.v(7290)
  and u6838 (Uzaiu6, Xjoiu6, Ekoiu6);  // ../RTL/cortexm0ds_logic.v(7291)
  and u6839 (Ekoiu6, Lkoiu6, Skoiu6);  // ../RTL/cortexm0ds_logic.v(7292)
  buf u684 (Gtgpw6[20], Zodbx6);  // ../RTL/cortexm0ds_logic.v(2375)
  and u6840 (n1611, Zkoiu6, Gloiu6);  // ../RTL/cortexm0ds_logic.v(7293)
  not u6841 (Skoiu6, n1611);  // ../RTL/cortexm0ds_logic.v(7293)
  or u6842 (n1612, Nloiu6, Xe8iu6);  // ../RTL/cortexm0ds_logic.v(7294)
  not u6843 (Gloiu6, n1612);  // ../RTL/cortexm0ds_logic.v(7294)
  or u6844 (n1613, G7oiu6, Zraiu6);  // ../RTL/cortexm0ds_logic.v(7295)
  not u6845 (Zkoiu6, n1613);  // ../RTL/cortexm0ds_logic.v(7295)
  and u6846 (Lkoiu6, Twniu6, Uloiu6);  // ../RTL/cortexm0ds_logic.v(7296)
  and u6847 (Xjoiu6, Bmoiu6, Imoiu6);  // ../RTL/cortexm0ds_logic.v(7297)
  and u6848 (n1614, L0niu6, Tfjiu6);  // ../RTL/cortexm0ds_logic.v(7298)
  not u6849 (Bmoiu6, n1614);  // ../RTL/cortexm0ds_logic.v(7298)
  buf u685 (Gtgpw6[19], Bxbax6);  // ../RTL/cortexm0ds_logic.v(2375)
  and u6850 (n1615, Pmoiu6, Wmoiu6);  // ../RTL/cortexm0ds_logic.v(7299)
  not u6851 (Dgphu6, n1615);  // ../RTL/cortexm0ds_logic.v(7299)
  and u6852 (Wmoiu6, Dnoiu6, Knoiu6);  // ../RTL/cortexm0ds_logic.v(7300)
  and u6853 (n1616, Ok8iu6, vis_pc_o[30]);  // ../RTL/cortexm0ds_logic.v(7301)
  not u6854 (Knoiu6, n1616);  // ../RTL/cortexm0ds_logic.v(7301)
  and u6855 (Ok8iu6, Rnoiu6, W8aiu6);  // ../RTL/cortexm0ds_logic.v(7302)
  and u6856 (Rnoiu6, Ynoiu6, Lm8iu6);  // ../RTL/cortexm0ds_logic.v(7303)
  and u6857 (n1617, Fooiu6, Lraiu6);  // ../RTL/cortexm0ds_logic.v(7304)
  not u6858 (Ynoiu6, n1617);  // ../RTL/cortexm0ds_logic.v(7304)
  and u6859 (Fooiu6, Mooiu6, Tr0iu6);  // ../RTL/cortexm0ds_logic.v(7305)
  buf u686 (Gtgpw6[18], Yybax6);  // ../RTL/cortexm0ds_logic.v(2375)
  or u6860 (Mooiu6, Ttciu6, D7fpw6[3]);  // ../RTL/cortexm0ds_logic.v(7306)
  and u6861 (Dnoiu6, Tooiu6, Apoiu6);  // ../RTL/cortexm0ds_logic.v(7307)
  and u6862 (n1618, Jl8iu6, Ef1iu6);  // ../RTL/cortexm0ds_logic.v(7308)
  not u6863 (Apoiu6, n1618);  // ../RTL/cortexm0ds_logic.v(7308)
  and u6864 (Jl8iu6, Hpoiu6, Lm8iu6);  // ../RTL/cortexm0ds_logic.v(7309)
  and u6865 (n1619, Y7ghu6, Opoiu6);  // ../RTL/cortexm0ds_logic.v(7310)
  not u6866 (Hpoiu6, n1619);  // ../RTL/cortexm0ds_logic.v(7310)
  or u6867 (Opoiu6, Jojiu6, Cyfpw6[1]);  // ../RTL/cortexm0ds_logic.v(7311)
  and u6868 (n1620, vis_apsr_o[3], Ql8iu6);  // ../RTL/cortexm0ds_logic.v(7312)
  not u6869 (Tooiu6, n1620);  // ../RTL/cortexm0ds_logic.v(7312)
  buf u687 (Gtgpw6[17], Knbbx6);  // ../RTL/cortexm0ds_logic.v(2375)
  and u6870 (Ql8iu6, Vpoiu6, U19iu6);  // ../RTL/cortexm0ds_logic.v(7313)
  and u6871 (U19iu6, Cqoiu6, Jqoiu6);  // ../RTL/cortexm0ds_logic.v(7314)
  and u6872 (n1621, Qqoiu6, Xqoiu6);  // ../RTL/cortexm0ds_logic.v(7315)
  not u6873 (Jqoiu6, n1621);  // ../RTL/cortexm0ds_logic.v(7315)
  or u6874 (n1622, V4aiu6, R2aiu6);  // ../RTL/cortexm0ds_logic.v(7316)
  not u6875 (Xqoiu6, n1622);  // ../RTL/cortexm0ds_logic.v(7316)
  or u6876 (n1623, Q5aiu6, Prjiu6);  // ../RTL/cortexm0ds_logic.v(7317)
  not u6877 (Qqoiu6, n1623);  // ../RTL/cortexm0ds_logic.v(7317)
  and u6878 (Cqoiu6, Eroiu6, Lroiu6);  // ../RTL/cortexm0ds_logic.v(7318)
  and u6879 (n1624, Sroiu6, Zroiu6);  // ../RTL/cortexm0ds_logic.v(7319)
  buf u688 (Gtgpw6[16], V0cax6);  // ../RTL/cortexm0ds_logic.v(2375)
  not u6880 (Eroiu6, n1624);  // ../RTL/cortexm0ds_logic.v(7319)
  and u6881 (Sroiu6, D7fpw6[8], Nbkiu6);  // ../RTL/cortexm0ds_logic.v(7320)
  and u6882 (Vpoiu6, Frliu6, Lm8iu6);  // ../RTL/cortexm0ds_logic.v(7321)
  and u6883 (n1625, Twniu6, Gsoiu6);  // ../RTL/cortexm0ds_logic.v(7322)
  not u6884 (Frliu6, n1625);  // ../RTL/cortexm0ds_logic.v(7322)
  and u6885 (n1626, Nsoiu6, Usoiu6);  // ../RTL/cortexm0ds_logic.v(7323)
  not u6886 (Gsoiu6, n1626);  // ../RTL/cortexm0ds_logic.v(7323)
  and u6887 (Usoiu6, Btoiu6, D7fpw6[3]);  // ../RTL/cortexm0ds_logic.v(7324)
  or u6888 (n1627, Q5aiu6, Ttciu6);  // ../RTL/cortexm0ds_logic.v(7325)
  not u6889 (Nsoiu6, n1627);  // ../RTL/cortexm0ds_logic.v(7325)
  buf u689 (Gtgpw6[14], Koabx6);  // ../RTL/cortexm0ds_logic.v(2375)
  and u6890 (Pmoiu6, Itoiu6, Ptoiu6);  // ../RTL/cortexm0ds_logic.v(7326)
  or u6891 (Ptoiu6, Lm8iu6, Wtoiu6);  // ../RTL/cortexm0ds_logic.v(7327)
  not u6892 (Lm8iu6, W29iu6);  // ../RTL/cortexm0ds_logic.v(7328)
  and u6893 (W29iu6, Duoiu6, Hx9iu6);  // ../RTL/cortexm0ds_logic.v(7329)
  and u6894 (n1628, HREADY, Kuoiu6);  // ../RTL/cortexm0ds_logic.v(7330)
  not u6895 (Duoiu6, n1628);  // ../RTL/cortexm0ds_logic.v(7330)
  and u6896 (n1629, Ruoiu6, Yuoiu6);  // ../RTL/cortexm0ds_logic.v(7331)
  not u6897 (Kuoiu6, n1629);  // ../RTL/cortexm0ds_logic.v(7331)
  and u6898 (Yuoiu6, Fvoiu6, Mvoiu6);  // ../RTL/cortexm0ds_logic.v(7332)
  and u6899 (Mvoiu6, Tvoiu6, Awoiu6);  // ../RTL/cortexm0ds_logic.v(7333)
  buf u69 (vis_r5_o[2], Wjtpw6);  // ../RTL/cortexm0ds_logic.v(1909)
  buf u690 (Gtgpw6[12], M6cax6);  // ../RTL/cortexm0ds_logic.v(2375)
  and u6900 (n1630, Hwoiu6, Ia8iu6);  // ../RTL/cortexm0ds_logic.v(7334)
  not u6901 (Awoiu6, n1630);  // ../RTL/cortexm0ds_logic.v(7334)
  and u6902 (Hwoiu6, Vviiu6, D7fpw6[12]);  // ../RTL/cortexm0ds_logic.v(7335)
  and u6903 (n1631, Y0jiu6, Owoiu6);  // ../RTL/cortexm0ds_logic.v(7336)
  not u6904 (Tvoiu6, n1631);  // ../RTL/cortexm0ds_logic.v(7336)
  and u6905 (Fvoiu6, Vwoiu6, Cxoiu6);  // ../RTL/cortexm0ds_logic.v(7337)
  or u6906 (Cxoiu6, Jxoiu6, Qxoiu6);  // ../RTL/cortexm0ds_logic.v(7338)
  and u6907 (n1632, Xxoiu6, Zraiu6);  // ../RTL/cortexm0ds_logic.v(7339)
  not u6908 (Vwoiu6, n1632);  // ../RTL/cortexm0ds_logic.v(7339)
  and u6909 (n1633, Eyoiu6, Lyoiu6);  // ../RTL/cortexm0ds_logic.v(7340)
  buf u691 (Gtgpw6[10], J8cax6);  // ../RTL/cortexm0ds_logic.v(2375)
  not u6910 (Xxoiu6, n1633);  // ../RTL/cortexm0ds_logic.v(7340)
  and u6911 (Lyoiu6, Syoiu6, Td0iu6);  // ../RTL/cortexm0ds_logic.v(7341)
  and u6912 (n1634, Zyoiu6, Gzoiu6);  // ../RTL/cortexm0ds_logic.v(7342)
  not u6913 (Syoiu6, n1634);  // ../RTL/cortexm0ds_logic.v(7342)
  or u6914 (n1635, Lraiu6, Nzoiu6);  // ../RTL/cortexm0ds_logic.v(7343)
  not u6915 (Gzoiu6, n1635);  // ../RTL/cortexm0ds_logic.v(7343)
  and u6916 (Zyoiu6, Wliiu6, Dmiiu6);  // ../RTL/cortexm0ds_logic.v(7344)
  and u6917 (Eyoiu6, Uzoiu6, B0piu6);  // ../RTL/cortexm0ds_logic.v(7345)
  and u6918 (n1636, I0piu6, P0piu6);  // ../RTL/cortexm0ds_logic.v(7346)
  not u6919 (B0piu6, n1636);  // ../RTL/cortexm0ds_logic.v(7346)
  buf u692 (Gtgpw6[7], Bccax6);  // ../RTL/cortexm0ds_logic.v(2375)
  and u6920 (I0piu6, W0piu6, D7fpw6[13]);  // ../RTL/cortexm0ds_logic.v(7347)
  and u6921 (n1637, Vxniu6, D1piu6);  // ../RTL/cortexm0ds_logic.v(7348)
  not u6922 (Uzoiu6, n1637);  // ../RTL/cortexm0ds_logic.v(7348)
  and u6923 (Ruoiu6, K1piu6, R1piu6);  // ../RTL/cortexm0ds_logic.v(7349)
  and u6924 (R1piu6, Y1piu6, F2piu6);  // ../RTL/cortexm0ds_logic.v(7350)
  and u6925 (n1638, L0niu6, M2piu6);  // ../RTL/cortexm0ds_logic.v(7351)
  not u6926 (F2piu6, n1638);  // ../RTL/cortexm0ds_logic.v(7351)
  and u6927 (L0niu6, T2piu6, Md0iu6);  // ../RTL/cortexm0ds_logic.v(7352)
  or u6928 (n1639, A4oiu6, Mr0iu6);  // ../RTL/cortexm0ds_logic.v(7353)
  not u6929 (T2piu6, n1639);  // ../RTL/cortexm0ds_logic.v(7353)
  not u693 (Xudpw6, S11bx6);  // ../RTL/cortexm0ds_logic.v(2748)
  and u6930 (n1640, Geoiu6, Qe8iu6);  // ../RTL/cortexm0ds_logic.v(7354)
  not u6931 (Y1piu6, n1640);  // ../RTL/cortexm0ds_logic.v(7354)
  and u6932 (K1piu6, A3piu6, F85iu6);  // ../RTL/cortexm0ds_logic.v(7355)
  AL_MUX u6933 (
    .i0(H3piu6),
    .i1(O3piu6),
    .sel(Cyfpw6[3]),
    .o(A3piu6));  // ../RTL/cortexm0ds_logic.v(7356)
  and u6934 (n1641, V3piu6, W8aiu6);  // ../RTL/cortexm0ds_logic.v(7357)
  not u6935 (O3piu6, n1641);  // ../RTL/cortexm0ds_logic.v(7357)
  and u6936 (V3piu6, C4piu6, Nlaiu6);  // ../RTL/cortexm0ds_logic.v(7358)
  and u6937 (n1642, Lraiu6, J4piu6);  // ../RTL/cortexm0ds_logic.v(7359)
  not u6938 (C4piu6, n1642);  // ../RTL/cortexm0ds_logic.v(7359)
  and u6939 (n1643, Q4piu6, T0hhu6);  // ../RTL/cortexm0ds_logic.v(7360)
  buf u694 (Gtgpw6[6], Lg9bx6);  // ../RTL/cortexm0ds_logic.v(2375)
  not u6940 (J4piu6, n1643);  // ../RTL/cortexm0ds_logic.v(7360)
  and u6941 (Q4piu6, X4piu6, Ftjiu6);  // ../RTL/cortexm0ds_logic.v(7361)
  or u6942 (X4piu6, V4aiu6, R9aiu6);  // ../RTL/cortexm0ds_logic.v(7362)
  and u6943 (n1644, Zm8iu6, Lm1iu6);  // ../RTL/cortexm0ds_logic.v(7363)
  not u6944 (Itoiu6, n1644);  // ../RTL/cortexm0ds_logic.v(7363)
  and u6945 (Zm8iu6, E5piu6, HALTED);  // ../RTL/cortexm0ds_logic.v(7365)
  not u6946 (Hx9iu6, Zm8iu6);  // ../RTL/cortexm0ds_logic.v(7365)
  and u6947 (E5piu6, Ar1iu6, Npdhu6);  // ../RTL/cortexm0ds_logic.v(7366)
  or u6948 (Wfphu6, L5piu6, Ln7iu6);  // ../RTL/cortexm0ds_logic.v(7367)
  AL_MUX u6949 (
    .i0(Ppfpw6[16]),
    .i1(T15iu6),
    .sel(Zn7iu6),
    .o(L5piu6));  // ../RTL/cortexm0ds_logic.v(7368)
  not u695 (Qudpw6, W51bx6);  // ../RTL/cortexm0ds_logic.v(2750)
  and u6950 (Cpbiu6, A2ciu6, S5piu6);  // ../RTL/cortexm0ds_logic.v(7369)
  not u6951 (Zn7iu6, Cpbiu6);  // ../RTL/cortexm0ds_logic.v(7369)
  and u6952 (n1645, Z5piu6, G6piu6);  // ../RTL/cortexm0ds_logic.v(7370)
  not u6953 (S5piu6, n1645);  // ../RTL/cortexm0ds_logic.v(7370)
  or u6954 (n1646, N6piu6, C0ehu6);  // ../RTL/cortexm0ds_logic.v(7371)
  not u6955 (G6piu6, n1646);  // ../RTL/cortexm0ds_logic.v(7371)
  or u6956 (n1647, Qqhiu6, Juzhu6);  // ../RTL/cortexm0ds_logic.v(7372)
  not u6957 (Z5piu6, n1647);  // ../RTL/cortexm0ds_logic.v(7372)
  not u6958 (A2ciu6, Ln7iu6);  // ../RTL/cortexm0ds_logic.v(7373)
  or u6959 (Ln7iu6, H2ciu6, Ivfhu6);  // ../RTL/cortexm0ds_logic.v(7374)
  buf u696 (Trgpw6[20], Wqdbx6);  // ../RTL/cortexm0ds_logic.v(2376)
  not u6960 (H2ciu6, Jm7iu6);  // ../RTL/cortexm0ds_logic.v(7375)
  or u6961 (Jm7iu6, Wofiu6, U6piu6);  // ../RTL/cortexm0ds_logic.v(7376)
  and u6962 (Go7iu6, Svdpw6, Vobiu6);  // ../RTL/cortexm0ds_logic.v(7377)
  not u6963 (T15iu6, Go7iu6);  // ../RTL/cortexm0ds_logic.v(7377)
  or u6964 (Pfphu6, Ex4iu6, B7piu6);  // ../RTL/cortexm0ds_logic.v(7378)
  and u6965 (B7piu6, Dhgpw6[0], I7piu6);  // ../RTL/cortexm0ds_logic.v(7379)
  and u6966 (n1648, Scbiu6, T24iu6);  // ../RTL/cortexm0ds_logic.v(7380)
  not u6967 (I7piu6, n1648);  // ../RTL/cortexm0ds_logic.v(7380)
  and u6968 (n1649, P7piu6, W7piu6);  // ../RTL/cortexm0ds_logic.v(7381)
  not u6969 (Ex4iu6, n1649);  // ../RTL/cortexm0ds_logic.v(7381)
  not u697 (Judpw6, Ca1bx6);  // ../RTL/cortexm0ds_logic.v(2752)
  and u6970 (n1650, D8piu6, Tu4iu6);  // ../RTL/cortexm0ds_logic.v(7382)
  not u6971 (W7piu6, n1650);  // ../RTL/cortexm0ds_logic.v(7382)
  and u6972 (Tu4iu6, K8piu6, R8piu6);  // ../RTL/cortexm0ds_logic.v(7383)
  and u6973 (R8piu6, Y8piu6, F9piu6);  // ../RTL/cortexm0ds_logic.v(7384)
  and u6974 (F9piu6, M9piu6, T9piu6);  // ../RTL/cortexm0ds_logic.v(7385)
  and u6975 (T9piu6, Aapiu6, Asliu6);  // ../RTL/cortexm0ds_logic.v(7386)
  or u6976 (n1651, W74iu6, I74iu6);  // ../RTL/cortexm0ds_logic.v(7387)
  not u6977 (Aapiu6, n1651);  // ../RTL/cortexm0ds_logic.v(7387)
  or u6978 (n1652, Y84iu6, R84iu6);  // ../RTL/cortexm0ds_logic.v(7388)
  not u6979 (M9piu6, n1652);  // ../RTL/cortexm0ds_logic.v(7388)
  buf u698 (Trgpw6[22], Kpfbx6);  // ../RTL/cortexm0ds_logic.v(2376)
  and u6980 (Y8piu6, Hapiu6, Oapiu6);  // ../RTL/cortexm0ds_logic.v(7389)
  or u6981 (n1653, T94iu6, F94iu6);  // ../RTL/cortexm0ds_logic.v(7390)
  not u6982 (Oapiu6, n1653);  // ../RTL/cortexm0ds_logic.v(7390)
  and u6983 (Hapiu6, Lm1iu6, Rykiu6);  // ../RTL/cortexm0ds_logic.v(7391)
  and u6984 (K8piu6, Vapiu6, Cbpiu6);  // ../RTL/cortexm0ds_logic.v(7392)
  and u6985 (Cbpiu6, Jbpiu6, Qbpiu6);  // ../RTL/cortexm0ds_logic.v(7393)
  and u6986 (Qbpiu6, Xbpiu6, P74iu6);  // ../RTL/cortexm0ds_logic.v(7394)
  and u6987 (Xbpiu6, M94iu6, Z54iu6);  // ../RTL/cortexm0ds_logic.v(7395)
  and u6988 (Jbpiu6, U64iu6, B74iu6);  // ../RTL/cortexm0ds_logic.v(7396)
  and u6989 (Vapiu6, Ecpiu6, Lcpiu6);  // ../RTL/cortexm0ds_logic.v(7397)
  not u699 (Cudpw6, Ie1bx6);  // ../RTL/cortexm0ds_logic.v(2754)
  and u6990 (Lcpiu6, G64iu6, N64iu6);  // ../RTL/cortexm0ds_logic.v(7398)
  or u6991 (n1654, Duhiu6, Ps4iu6);  // ../RTL/cortexm0ds_logic.v(7399)
  not u6992 (Ecpiu6, n1654);  // ../RTL/cortexm0ds_logic.v(7399)
  and u6993 (D8piu6, T24iu6, O34iu6);  // ../RTL/cortexm0ds_logic.v(7400)
  and u6994 (n1655, Scpiu6, Zcpiu6);  // ../RTL/cortexm0ds_logic.v(7401)
  not u6995 (P7piu6, n1655);  // ../RTL/cortexm0ds_logic.v(7401)
  and u6996 (Zcpiu6, Gdpiu6, Jehhu6);  // ../RTL/cortexm0ds_logic.v(7402)
  and u6997 (Gdpiu6, Ndpiu6, Udpiu6);  // ../RTL/cortexm0ds_logic.v(7403)
  and u6998 (n1656, Bepiu6, Zrhiu6);  // ../RTL/cortexm0ds_logic.v(7404)
  not u6999 (Ndpiu6, n1656);  // ../RTL/cortexm0ds_logic.v(7404)
  buf u7 (HTRANS[0], 1'b0);  // ../RTL/cortexm0ds_logic.v(1730)
  buf u70 (vis_r8_o[31], Qmrax6);  // ../RTL/cortexm0ds_logic.v(2579)
  buf u700 (Trgpw6[21], Daebx6);  // ../RTL/cortexm0ds_logic.v(2376)
  or u7000 (n1657, LOCKUP, C0ehu6);  // ../RTL/cortexm0ds_logic.v(7405)
  not u7001 (Zrhiu6, n1657);  // ../RTL/cortexm0ds_logic.v(7405)
  and u7002 (Bepiu6, Uc5iu6, Sb5iu6);  // ../RTL/cortexm0ds_logic.v(7406)
  and u7003 (n1658, Iepiu6, K2aiu6);  // ../RTL/cortexm0ds_logic.v(7407)
  not u7004 (Uc5iu6, n1658);  // ../RTL/cortexm0ds_logic.v(7407)
  and u7005 (Scpiu6, Hbhhu6, HREADY);  // ../RTL/cortexm0ds_logic.v(7408)
  and u7006 (n1659, Pepiu6, Wepiu6);  // ../RTL/cortexm0ds_logic.v(7409)
  not u7007 (Ifphu6, n1659);  // ../RTL/cortexm0ds_logic.v(7409)
  and u7008 (n1660, Dfpiu6, Lx4iu6);  // ../RTL/cortexm0ds_logic.v(7410)
  not u7009 (Wepiu6, n1660);  // ../RTL/cortexm0ds_logic.v(7410)
  not u701 (Vtdpw6, Oi1bx6);  // ../RTL/cortexm0ds_logic.v(2756)
  or u7010 (Lx4iu6, Kfpiu6, Rfpiu6);  // ../RTL/cortexm0ds_logic.v(7411)
  and u7011 (n1661, Eh6iu6, Yfpiu6);  // ../RTL/cortexm0ds_logic.v(7412)
  not u7012 (Dfpiu6, n1661);  // ../RTL/cortexm0ds_logic.v(7412)
  and u7013 (n1662, Dhgpw6[2], Yfpiu6);  // ../RTL/cortexm0ds_logic.v(7413)
  not u7014 (Pepiu6, n1662);  // ../RTL/cortexm0ds_logic.v(7413)
  and u7015 (n1663, Scbiu6, Ud4iu6);  // ../RTL/cortexm0ds_logic.v(7414)
  not u7016 (Yfpiu6, n1663);  // ../RTL/cortexm0ds_logic.v(7414)
  and u7017 (Scbiu6, Fgpiu6, A2nhu6);  // ../RTL/cortexm0ds_logic.v(7415)
  and u7018 (n1664, Mgpiu6, Tgpiu6);  // ../RTL/cortexm0ds_logic.v(7416)
  not u7019 (Bfphu6, n1664);  // ../RTL/cortexm0ds_logic.v(7416)
  buf u702 (Trgpw6[19], Gkeax6);  // ../RTL/cortexm0ds_logic.v(2376)
  and u7020 (n1665, Rfpiu6, Ahpiu6);  // ../RTL/cortexm0ds_logic.v(7417)
  not u7021 (Tgpiu6, n1665);  // ../RTL/cortexm0ds_logic.v(7417)
  and u7022 (n1666, Eh6iu6, Hhpiu6);  // ../RTL/cortexm0ds_logic.v(7418)
  not u7023 (Ahpiu6, n1666);  // ../RTL/cortexm0ds_logic.v(7418)
  and u7024 (Rfpiu6, Ohpiu6, Yuhhu6);  // ../RTL/cortexm0ds_logic.v(7419)
  or u7025 (n1667, E81iu6, Vhpiu6);  // ../RTL/cortexm0ds_logic.v(7420)
  not u7026 (Ohpiu6, n1667);  // ../RTL/cortexm0ds_logic.v(7420)
  and u7027 (Vhpiu6, Cipiu6, Jipiu6);  // ../RTL/cortexm0ds_logic.v(7421)
  and u7028 (n1668, Qipiu6, Xipiu6);  // ../RTL/cortexm0ds_logic.v(7422)
  not u7029 (Jipiu6, n1668);  // ../RTL/cortexm0ds_logic.v(7422)
  not u703 (Otdpw6, Um1bx6);  // ../RTL/cortexm0ds_logic.v(2758)
  AL_MUX u7030 (
    .i0(Lwgpw6[1]),
    .i1(Lwgpw6[0]),
    .sel(Ejpiu6),
    .o(Qipiu6));  // ../RTL/cortexm0ds_logic.v(7423)
  or u7031 (Cipiu6, Ljpiu6, Ty0iu6);  // ../RTL/cortexm0ds_logic.v(7424)
  or u7032 (Ty0iu6, Lwgpw6[0], Lwgpw6[1]);  // ../RTL/cortexm0ds_logic.v(7425)
  and u7033 (n1669, Sjpiu6, Lwgpw6[2]);  // ../RTL/cortexm0ds_logic.v(7426)
  not u7034 (E81iu6, n1669);  // ../RTL/cortexm0ds_logic.v(7426)
  and u7035 (n1670, Hwmhu6, Hhpiu6);  // ../RTL/cortexm0ds_logic.v(7427)
  not u7036 (Mgpiu6, n1670);  // ../RTL/cortexm0ds_logic.v(7427)
  and u7037 (n1671, Ws4iu6, Ps4iu6);  // ../RTL/cortexm0ds_logic.v(7428)
  not u7038 (Hhpiu6, n1671);  // ../RTL/cortexm0ds_logic.v(7428)
  and u7039 (n1672, Zjpiu6, Gkpiu6);  // ../RTL/cortexm0ds_logic.v(7429)
  buf u704 (Trgpw6[18], Dmeax6);  // ../RTL/cortexm0ds_logic.v(2376)
  not u7040 (Uephu6, n1672);  // ../RTL/cortexm0ds_logic.v(7429)
  and u7041 (n1673, Kfpiu6, Nkpiu6);  // ../RTL/cortexm0ds_logic.v(7430)
  not u7042 (Gkpiu6, n1673);  // ../RTL/cortexm0ds_logic.v(7430)
  and u7043 (n1674, Eh6iu6, Ukpiu6);  // ../RTL/cortexm0ds_logic.v(7431)
  not u7044 (Nkpiu6, n1674);  // ../RTL/cortexm0ds_logic.v(7431)
  and u7045 (Kfpiu6, Blpiu6, Mekhu6);  // ../RTL/cortexm0ds_logic.v(7432)
  or u7046 (n1675, Yx0iu6, Ilpiu6);  // ../RTL/cortexm0ds_logic.v(7433)
  not u7047 (Blpiu6, n1675);  // ../RTL/cortexm0ds_logic.v(7433)
  and u7048 (Ilpiu6, Plpiu6, Wlpiu6);  // ../RTL/cortexm0ds_logic.v(7434)
  and u7049 (n1676, Dmpiu6, Xipiu6);  // ../RTL/cortexm0ds_logic.v(7435)
  not u705 (Htdpw6, Ar1bx6);  // ../RTL/cortexm0ds_logic.v(2760)
  not u7050 (Wlpiu6, n1676);  // ../RTL/cortexm0ds_logic.v(7435)
  and u7051 (Xipiu6, Kmpiu6, Rmpiu6);  // ../RTL/cortexm0ds_logic.v(7436)
  or u7052 (Rmpiu6, Z18iu6, Ympiu6);  // ../RTL/cortexm0ds_logic.v(7437)
  or u7053 (n1677, HMASTER, L18iu6);  // ../RTL/cortexm0ds_logic.v(7438)
  not u7054 (Kmpiu6, n1677);  // ../RTL/cortexm0ds_logic.v(7438)
  AL_MUX u7055 (
    .i0(R2hpw6[0]),
    .i1(R2hpw6[1]),
    .sel(Fnpiu6),
    .o(Dmpiu6));  // ../RTL/cortexm0ds_logic.v(7439)
  or u7056 (Plpiu6, Ljpiu6, Nv0iu6);  // ../RTL/cortexm0ds_logic.v(7440)
  or u7057 (Nv0iu6, R2hpw6[0], R2hpw6[1]);  // ../RTL/cortexm0ds_logic.v(7441)
  and u7058 (n1678, Mnpiu6, Sufpw6[1]);  // ../RTL/cortexm0ds_logic.v(7442)
  not u7059 (Ljpiu6, n1678);  // ../RTL/cortexm0ds_logic.v(7442)
  buf u706 (Trgpw6[15], Xpeax6);  // ../RTL/cortexm0ds_logic.v(2376)
  and u7060 (Mnpiu6, Sufpw6[0], K9aiu6);  // ../RTL/cortexm0ds_logic.v(7443)
  and u7061 (n1679, Sjpiu6, R2hpw6[2]);  // ../RTL/cortexm0ds_logic.v(7444)
  not u7062 (Yx0iu6, n1679);  // ../RTL/cortexm0ds_logic.v(7444)
  and u7063 (Sjpiu6, E5hhu6, Jehhu6);  // ../RTL/cortexm0ds_logic.v(7445)
  and u7064 (n1680, Vxmhu6, Ukpiu6);  // ../RTL/cortexm0ds_logic.v(7446)
  not u7065 (Zjpiu6, n1680);  // ../RTL/cortexm0ds_logic.v(7446)
  and u7066 (n1681, Eg7iu6, Ps4iu6);  // ../RTL/cortexm0ds_logic.v(7447)
  not u7067 (Ukpiu6, n1681);  // ../RTL/cortexm0ds_logic.v(7447)
  not u7068 (Ps4iu6, A2nhu6);  // ../RTL/cortexm0ds_logic.v(7448)
  and u7069 (n1682, Tnpiu6, Aopiu6);  // ../RTL/cortexm0ds_logic.v(7449)
  not u707 (Atdpw6, Gv1bx6);  // ../RTL/cortexm0ds_logic.v(2762)
  not u7070 (Nephu6, n1682);  // ../RTL/cortexm0ds_logic.v(7449)
  and u7071 (Aopiu6, Hopiu6, Oopiu6);  // ../RTL/cortexm0ds_logic.v(7450)
  and u7072 (n1683, Tnhpw6[1], Bo1iu6);  // ../RTL/cortexm0ds_logic.v(7451)
  not u7073 (Oopiu6, n1683);  // ../RTL/cortexm0ds_logic.v(7451)
  and u7074 (Hopiu6, Vopiu6, Po1iu6);  // ../RTL/cortexm0ds_logic.v(7452)
  and u7075 (n1684, Wo1iu6, Cppiu6);  // ../RTL/cortexm0ds_logic.v(7453)
  not u7076 (Vopiu6, n1684);  // ../RTL/cortexm0ds_logic.v(7453)
  and u7077 (n1685, Jppiu6, Qppiu6);  // ../RTL/cortexm0ds_logic.v(7454)
  not u7078 (Cppiu6, n1685);  // ../RTL/cortexm0ds_logic.v(7454)
  and u7079 (Qppiu6, Xppiu6, Eqpiu6);  // ../RTL/cortexm0ds_logic.v(7455)
  buf u708 (Trgpw6[16], Aoeax6);  // ../RTL/cortexm0ds_logic.v(2376)
  and u7080 (Eqpiu6, Lqpiu6, Sqpiu6);  // ../RTL/cortexm0ds_logic.v(7456)
  and u7081 (Sqpiu6, Zqpiu6, Grpiu6);  // ../RTL/cortexm0ds_logic.v(7457)
  and u7082 (n1686, R2hpw6[1], Eg7iu6);  // ../RTL/cortexm0ds_logic.v(7458)
  not u7083 (Grpiu6, n1686);  // ../RTL/cortexm0ds_logic.v(7458)
  and u7084 (n1687, Dhgpw6[1], Fgpiu6);  // ../RTL/cortexm0ds_logic.v(7459)
  not u7085 (Zqpiu6, n1687);  // ../RTL/cortexm0ds_logic.v(7459)
  and u7086 (Lqpiu6, Nrpiu6, Urpiu6);  // ../RTL/cortexm0ds_logic.v(7460)
  and u7087 (n1688, G4hpw6[1], Sg7iu6);  // ../RTL/cortexm0ds_logic.v(7461)
  not u7088 (Urpiu6, n1688);  // ../RTL/cortexm0ds_logic.v(7461)
  and u7089 (n1689, Aygpw6[1], Jf7iu6);  // ../RTL/cortexm0ds_logic.v(7462)
  not u709 (Tsdpw6, Mz1bx6);  // ../RTL/cortexm0ds_logic.v(2764)
  not u7090 (Nrpiu6, n1689);  // ../RTL/cortexm0ds_logic.v(7462)
  and u7091 (Xppiu6, Bspiu6, Ispiu6);  // ../RTL/cortexm0ds_logic.v(7463)
  and u7092 (n1690, Ar1iu6, Fkfpw6[1]);  // ../RTL/cortexm0ds_logic.v(7464)
  not u7093 (Ispiu6, n1690);  // ../RTL/cortexm0ds_logic.v(7464)
  and u7094 (Bspiu6, Pspiu6, Wspiu6);  // ../RTL/cortexm0ds_logic.v(7465)
  or u7095 (Wspiu6, Duhiu6, Udpiu6);  // ../RTL/cortexm0ds_logic.v(7466)
  and u7096 (n1691, Lwgpw6[1], Ws4iu6);  // ../RTL/cortexm0ds_logic.v(7467)
  not u7097 (Pspiu6, n1691);  // ../RTL/cortexm0ds_logic.v(7467)
  and u7098 (Jppiu6, Dtpiu6, Ktpiu6);  // ../RTL/cortexm0ds_logic.v(7468)
  and u7099 (Ktpiu6, Rtpiu6, Ytpiu6);  // ../RTL/cortexm0ds_logic.v(7469)
  buf u71 (Fnnhu6, Ahlpw6);  // ../RTL/cortexm0ds_logic.v(1837)
  buf u710 (Trgpw6[14], Hqabx6);  // ../RTL/cortexm0ds_logic.v(2376)
  and u7100 (Ytpiu6, Fupiu6, Mupiu6);  // ../RTL/cortexm0ds_logic.v(7470)
  and u7101 (n1692, HRDATA[1], St1iu6);  // ../RTL/cortexm0ds_logic.v(7471)
  not u7102 (Mupiu6, n1692);  // ../RTL/cortexm0ds_logic.v(7471)
  and u7103 (n1693, Zt1iu6, Pzgpw6[1]);  // ../RTL/cortexm0ds_logic.v(7472)
  not u7104 (Fupiu6, n1693);  // ../RTL/cortexm0ds_logic.v(7472)
  and u7105 (Rtpiu6, Tupiu6, Avpiu6);  // ../RTL/cortexm0ds_logic.v(7473)
  and u7106 (n1694, Kw1iu6, V5hpw6[1]);  // ../RTL/cortexm0ds_logic.v(7474)
  not u7107 (Avpiu6, n1694);  // ../RTL/cortexm0ds_logic.v(7474)
  and u7108 (n1695, Iv1iu6, vis_pc_o[0]);  // ../RTL/cortexm0ds_logic.v(7475)
  not u7109 (Tupiu6, n1695);  // ../RTL/cortexm0ds_logic.v(7475)
  not u711 (Msdpw6, S32bx6);  // ../RTL/cortexm0ds_logic.v(2766)
  and u7110 (Dtpiu6, Hvpiu6, Ovpiu6);  // ../RTL/cortexm0ds_logic.v(7476)
  and u7111 (Hvpiu6, Vvpiu6, Yw1iu6);  // ../RTL/cortexm0ds_logic.v(7477)
  and u7112 (Tnpiu6, Cwpiu6, Jwpiu6);  // ../RTL/cortexm0ds_logic.v(7478)
  and u7113 (n1696, Qwpiu6, Aphpw6[2]);  // ../RTL/cortexm0ds_logic.v(7479)
  not u7114 (Jwpiu6, n1696);  // ../RTL/cortexm0ds_logic.v(7479)
  and u7115 (n1697, Uthpw6[1], Sf1iu6);  // ../RTL/cortexm0ds_logic.v(7480)
  not u7116 (Cwpiu6, n1697);  // ../RTL/cortexm0ds_logic.v(7480)
  and u7117 (n1698, Xwpiu6, Expiu6);  // ../RTL/cortexm0ds_logic.v(7481)
  not u7118 (Gephu6, n1698);  // ../RTL/cortexm0ds_logic.v(7481)
  and u7119 (n1699, Uthpw6[2], Sf1iu6);  // ../RTL/cortexm0ds_logic.v(7482)
  buf u712 (Trgpw6[13], Ureax6);  // ../RTL/cortexm0ds_logic.v(2376)
  not u7120 (Expiu6, n1699);  // ../RTL/cortexm0ds_logic.v(7482)
  and u7121 (Xwpiu6, Lxpiu6, Sxpiu6);  // ../RTL/cortexm0ds_logic.v(7483)
  and u7122 (n1700, Wo1iu6, Zxpiu6);  // ../RTL/cortexm0ds_logic.v(7484)
  not u7123 (Sxpiu6, n1700);  // ../RTL/cortexm0ds_logic.v(7484)
  and u7124 (n1701, Gypiu6, Nypiu6);  // ../RTL/cortexm0ds_logic.v(7485)
  not u7125 (Zxpiu6, n1701);  // ../RTL/cortexm0ds_logic.v(7485)
  and u7126 (Nypiu6, Uypiu6, Bzpiu6);  // ../RTL/cortexm0ds_logic.v(7486)
  and u7127 (Bzpiu6, Izpiu6, Pzpiu6);  // ../RTL/cortexm0ds_logic.v(7487)
  and u7128 (Pzpiu6, Wzpiu6, D0qiu6);  // ../RTL/cortexm0ds_logic.v(7488)
  and u7129 (n1702, K0qiu6, Hbhhu6);  // ../RTL/cortexm0ds_logic.v(7489)
  not u713 (Fsdpw6, Y72bx6);  // ../RTL/cortexm0ds_logic.v(2768)
  not u7130 (D0qiu6, n1702);  // ../RTL/cortexm0ds_logic.v(7489)
  or u7131 (Grwiu6, Duhiu6, Zwciu6);  // ../RTL/cortexm0ds_logic.v(7490)
  not u7132 (K0qiu6, Grwiu6);  // ../RTL/cortexm0ds_logic.v(7490)
  and u7133 (Izpiu6, R0qiu6, Y0qiu6);  // ../RTL/cortexm0ds_logic.v(7491)
  and u7134 (n1703, Eg7iu6, R2hpw6[2]);  // ../RTL/cortexm0ds_logic.v(7492)
  not u7135 (Y0qiu6, n1703);  // ../RTL/cortexm0ds_logic.v(7492)
  and u7136 (R0qiu6, F1qiu6, M1qiu6);  // ../RTL/cortexm0ds_logic.v(7493)
  and u7137 (n1704, T1qiu6, A2qiu6);  // ../RTL/cortexm0ds_logic.v(7494)
  not u7138 (M1qiu6, n1704);  // ../RTL/cortexm0ds_logic.v(7494)
  AL_MUX u7139 (
    .i0(H2qiu6),
    .i1(O2qiu6),
    .sel(X8hpw6[5]),
    .o(T1qiu6));  // ../RTL/cortexm0ds_logic.v(7495)
  buf u714 (Gtgpw6[5], Xdcax6);  // ../RTL/cortexm0ds_logic.v(2375)
  or u7140 (O2qiu6, V2qiu6, C3qiu6);  // ../RTL/cortexm0ds_logic.v(7496)
  and u7141 (V2qiu6, Dr6iu6, Vm6iu6);  // ../RTL/cortexm0ds_logic.v(7497)
  or u7142 (n1705, J3qiu6, Dr6iu6);  // ../RTL/cortexm0ds_logic.v(7498)
  not u7143 (H2qiu6, n1705);  // ../RTL/cortexm0ds_logic.v(7498)
  and u7144 (n1706, Q3qiu6, Fl6iu6);  // ../RTL/cortexm0ds_logic.v(7499)
  not u7145 (F1qiu6, n1706);  // ../RTL/cortexm0ds_logic.v(7499)
  and u7146 (Uypiu6, X3qiu6, E4qiu6);  // ../RTL/cortexm0ds_logic.v(7500)
  and u7147 (E4qiu6, L4qiu6, S4qiu6);  // ../RTL/cortexm0ds_logic.v(7501)
  and u7148 (n1707, Aygpw6[2], Jf7iu6);  // ../RTL/cortexm0ds_logic.v(7502)
  not u7149 (S4qiu6, n1707);  // ../RTL/cortexm0ds_logic.v(7502)
  not u715 (Yrdpw6, Cc2bx6);  // ../RTL/cortexm0ds_logic.v(2770)
  and u7150 (L4qiu6, Z4qiu6, G5qiu6);  // ../RTL/cortexm0ds_logic.v(7503)
  and u7151 (n1708, Dhgpw6[2], Fgpiu6);  // ../RTL/cortexm0ds_logic.v(7504)
  not u7152 (G5qiu6, n1708);  // ../RTL/cortexm0ds_logic.v(7504)
  and u7153 (n1709, G4hpw6[2], Sg7iu6);  // ../RTL/cortexm0ds_logic.v(7505)
  not u7154 (Z4qiu6, n1709);  // ../RTL/cortexm0ds_logic.v(7505)
  and u7155 (X3qiu6, N5qiu6, U5qiu6);  // ../RTL/cortexm0ds_logic.v(7506)
  and u7156 (n1710, Togpw6[2], Vr1iu6);  // ../RTL/cortexm0ds_logic.v(7507)
  not u7157 (U5qiu6, n1710);  // ../RTL/cortexm0ds_logic.v(7507)
  and u7158 (n1711, Ws4iu6, Lwgpw6[2]);  // ../RTL/cortexm0ds_logic.v(7508)
  not u7159 (N5qiu6, n1711);  // ../RTL/cortexm0ds_logic.v(7508)
  buf u716 (Trgpw6[12], Rteax6);  // ../RTL/cortexm0ds_logic.v(2376)
  and u7160 (Gypiu6, B6qiu6, I6qiu6);  // ../RTL/cortexm0ds_logic.v(7509)
  and u7161 (I6qiu6, P6qiu6, W6qiu6);  // ../RTL/cortexm0ds_logic.v(7510)
  and u7162 (W6qiu6, D7qiu6, K7qiu6);  // ../RTL/cortexm0ds_logic.v(7511)
  and u7163 (n1712, HRDATA[2], St1iu6);  // ../RTL/cortexm0ds_logic.v(7512)
  not u7164 (K7qiu6, n1712);  // ../RTL/cortexm0ds_logic.v(7512)
  and u7165 (D7qiu6, R7qiu6, Y7qiu6);  // ../RTL/cortexm0ds_logic.v(7513)
  and u7166 (n1713, Gtgpw6[2], Cs1iu6);  // ../RTL/cortexm0ds_logic.v(7514)
  not u7167 (Y7qiu6, n1713);  // ../RTL/cortexm0ds_logic.v(7514)
  and u7168 (n1714, Ar1iu6, Fkfpw6[2]);  // ../RTL/cortexm0ds_logic.v(7515)
  not u7169 (R7qiu6, n1714);  // ../RTL/cortexm0ds_logic.v(7515)
  not u717 (Rrdpw6, Ig2bx6);  // ../RTL/cortexm0ds_logic.v(2772)
  and u7170 (P6qiu6, F8qiu6, M8qiu6);  // ../RTL/cortexm0ds_logic.v(7516)
  and u7171 (n1715, E1hpw6[2], Zt1iu6);  // ../RTL/cortexm0ds_logic.v(7517)
  not u7172 (M8qiu6, n1715);  // ../RTL/cortexm0ds_logic.v(7517)
  and u7173 (n1716, Gqgpw6[2], Xs1iu6);  // ../RTL/cortexm0ds_logic.v(7518)
  not u7174 (F8qiu6, n1716);  // ../RTL/cortexm0ds_logic.v(7518)
  and u7175 (B6qiu6, T8qiu6, A9qiu6);  // ../RTL/cortexm0ds_logic.v(7519)
  and u7176 (A9qiu6, H9qiu6, O9qiu6);  // ../RTL/cortexm0ds_logic.v(7520)
  and u7177 (n1717, Iv1iu6, vis_pc_o[1]);  // ../RTL/cortexm0ds_logic.v(7521)
  not u7178 (O9qiu6, n1717);  // ../RTL/cortexm0ds_logic.v(7521)
  and u7179 (H9qiu6, V9qiu6, Caqiu6);  // ../RTL/cortexm0ds_logic.v(7522)
  buf u718 (Trgpw6[11], N19bx6);  // ../RTL/cortexm0ds_logic.v(2376)
  and u7180 (n1718, Trgpw6[2], Dw1iu6);  // ../RTL/cortexm0ds_logic.v(7523)
  not u7181 (Caqiu6, n1718);  // ../RTL/cortexm0ds_logic.v(7523)
  and u7182 (n1719, K7hpw6[2], Kw1iu6);  // ../RTL/cortexm0ds_logic.v(7524)
  not u7183 (V9qiu6, n1719);  // ../RTL/cortexm0ds_logic.v(7524)
  and u7184 (T8qiu6, Jaqiu6, Qaqiu6);  // ../RTL/cortexm0ds_logic.v(7525)
  and u7185 (n1720, Tnhpw6[2], Bo1iu6);  // ../RTL/cortexm0ds_logic.v(7526)
  not u7186 (Lxpiu6, n1720);  // ../RTL/cortexm0ds_logic.v(7526)
  and u7187 (n1721, Xaqiu6, Ebqiu6);  // ../RTL/cortexm0ds_logic.v(7527)
  not u7188 (Zdphu6, n1721);  // ../RTL/cortexm0ds_logic.v(7527)
  and u7189 (n1722, Uthpw6[3], Sf1iu6);  // ../RTL/cortexm0ds_logic.v(7528)
  not u719 (Krdpw6, Ok2bx6);  // ../RTL/cortexm0ds_logic.v(2774)
  not u7190 (Ebqiu6, n1722);  // ../RTL/cortexm0ds_logic.v(7528)
  and u7191 (Xaqiu6, Lbqiu6, Sbqiu6);  // ../RTL/cortexm0ds_logic.v(7529)
  and u7192 (n1723, Wo1iu6, Zbqiu6);  // ../RTL/cortexm0ds_logic.v(7530)
  not u7193 (Sbqiu6, n1723);  // ../RTL/cortexm0ds_logic.v(7530)
  and u7194 (n1724, Gcqiu6, Ncqiu6);  // ../RTL/cortexm0ds_logic.v(7531)
  not u7195 (Zbqiu6, n1724);  // ../RTL/cortexm0ds_logic.v(7531)
  and u7196 (Ncqiu6, Ucqiu6, Bdqiu6);  // ../RTL/cortexm0ds_logic.v(7532)
  and u7197 (Bdqiu6, Idqiu6, Pdqiu6);  // ../RTL/cortexm0ds_logic.v(7533)
  and u7198 (Pdqiu6, Wdqiu6, Deqiu6);  // ../RTL/cortexm0ds_logic.v(7534)
  and u7199 (n1725, Dhgpw6[3], Fgpiu6);  // ../RTL/cortexm0ds_logic.v(7535)
  buf u72 (H2fpw6[0], Shopw6);  // ../RTL/cortexm0ds_logic.v(2444)
  buf u720 (Trgpw6[7], Gzeax6);  // ../RTL/cortexm0ds_logic.v(2376)
  not u7200 (Deqiu6, n1725);  // ../RTL/cortexm0ds_logic.v(7535)
  and u7201 (Wdqiu6, Keqiu6, Reqiu6);  // ../RTL/cortexm0ds_logic.v(7536)
  and u7202 (n1726, Yeqiu6, Ffqiu6);  // ../RTL/cortexm0ds_logic.v(7537)
  not u7203 (Keqiu6, n1726);  // ../RTL/cortexm0ds_logic.v(7537)
  or u7204 (n1727, Mfqiu6, X8hpw6[0]);  // ../RTL/cortexm0ds_logic.v(7538)
  not u7205 (Yeqiu6, n1727);  // ../RTL/cortexm0ds_logic.v(7538)
  and u7206 (Idqiu6, Tfqiu6, Agqiu6);  // ../RTL/cortexm0ds_logic.v(7539)
  and u7207 (n1728, G4hpw6[3], Sg7iu6);  // ../RTL/cortexm0ds_logic.v(7540)
  not u7208 (Agqiu6, n1728);  // ../RTL/cortexm0ds_logic.v(7540)
  and u7209 (n1729, Aygpw6[3], Jf7iu6);  // ../RTL/cortexm0ds_logic.v(7541)
  not u721 (Drdpw6, Uo2bx6);  // ../RTL/cortexm0ds_logic.v(2776)
  not u7210 (Tfqiu6, n1729);  // ../RTL/cortexm0ds_logic.v(7541)
  and u7211 (Ucqiu6, Hgqiu6, Ogqiu6);  // ../RTL/cortexm0ds_logic.v(7542)
  and u7212 (Ogqiu6, Vgqiu6, Chqiu6);  // ../RTL/cortexm0ds_logic.v(7543)
  and u7213 (n1730, Togpw6[3], Vr1iu6);  // ../RTL/cortexm0ds_logic.v(7544)
  not u7214 (Chqiu6, n1730);  // ../RTL/cortexm0ds_logic.v(7544)
  or u7215 (Vgqiu6, Jhqiu6, Duhiu6);  // ../RTL/cortexm0ds_logic.v(7545)
  and u7216 (Hgqiu6, Qhqiu6, Xhqiu6);  // ../RTL/cortexm0ds_logic.v(7546)
  and u7217 (n1731, Gtgpw6[3], Cs1iu6);  // ../RTL/cortexm0ds_logic.v(7547)
  not u7218 (Xhqiu6, n1731);  // ../RTL/cortexm0ds_logic.v(7547)
  and u7219 (n1732, Ar1iu6, Fkfpw6[3]);  // ../RTL/cortexm0ds_logic.v(7548)
  buf u722 (Trgpw6[9], B9jbx6);  // ../RTL/cortexm0ds_logic.v(2376)
  not u7220 (Qhqiu6, n1732);  // ../RTL/cortexm0ds_logic.v(7548)
  and u7221 (Gcqiu6, Eiqiu6, Liqiu6);  // ../RTL/cortexm0ds_logic.v(7549)
  and u7222 (Liqiu6, Siqiu6, Ziqiu6);  // ../RTL/cortexm0ds_logic.v(7550)
  and u7223 (Ziqiu6, Gjqiu6, Njqiu6);  // ../RTL/cortexm0ds_logic.v(7551)
  and u7224 (n1733, Gqgpw6[3], Xs1iu6);  // ../RTL/cortexm0ds_logic.v(7552)
  not u7225 (Njqiu6, n1733);  // ../RTL/cortexm0ds_logic.v(7552)
  and u7226 (Gjqiu6, Ujqiu6, Bkqiu6);  // ../RTL/cortexm0ds_logic.v(7553)
  and u7227 (n1734, HRDATA[3], St1iu6);  // ../RTL/cortexm0ds_logic.v(7554)
  not u7228 (Bkqiu6, n1734);  // ../RTL/cortexm0ds_logic.v(7554)
  and u7229 (n1735, E1hpw6[3], Zt1iu6);  // ../RTL/cortexm0ds_logic.v(7555)
  not u723 (Wqdpw6, At2bx6);  // ../RTL/cortexm0ds_logic.v(2778)
  not u7230 (Ujqiu6, n1735);  // ../RTL/cortexm0ds_logic.v(7555)
  and u7231 (Siqiu6, Ikqiu6, Pkqiu6);  // ../RTL/cortexm0ds_logic.v(7556)
  and u7232 (n1736, Trgpw6[3], Dw1iu6);  // ../RTL/cortexm0ds_logic.v(7557)
  not u7233 (Pkqiu6, n1736);  // ../RTL/cortexm0ds_logic.v(7557)
  and u7234 (n1737, K7hpw6[3], Kw1iu6);  // ../RTL/cortexm0ds_logic.v(7558)
  not u7235 (Ikqiu6, n1737);  // ../RTL/cortexm0ds_logic.v(7558)
  and u7236 (Eiqiu6, Wkqiu6, Dlqiu6);  // ../RTL/cortexm0ds_logic.v(7559)
  and u7237 (Dlqiu6, Vvpiu6, Klqiu6);  // ../RTL/cortexm0ds_logic.v(7560)
  and u7238 (n1738, Iv1iu6, vis_pc_o[2]);  // ../RTL/cortexm0ds_logic.v(7561)
  not u7239 (Klqiu6, n1738);  // ../RTL/cortexm0ds_logic.v(7561)
  buf u724 (Trgpw6[8], Kxeax6);  // ../RTL/cortexm0ds_logic.v(2376)
  or u7240 (n1739, Rlqiu6, Ylqiu6);  // ../RTL/cortexm0ds_logic.v(7562)
  not u7241 (Vvpiu6, n1739);  // ../RTL/cortexm0ds_logic.v(7562)
  AL_MUX u7242 (
    .i0(Fmqiu6),
    .i1(Q3qiu6),
    .sel(X8hpw6[4]),
    .o(Rlqiu6));  // ../RTL/cortexm0ds_logic.v(7563)
  and u7243 (Fmqiu6, Mmqiu6, X8hpw6[1]);  // ../RTL/cortexm0ds_logic.v(7564)
  and u7244 (Wkqiu6, Tmqiu6, Anqiu6);  // ../RTL/cortexm0ds_logic.v(7565)
  and u7245 (n1740, Tnhpw6[3], Bo1iu6);  // ../RTL/cortexm0ds_logic.v(7566)
  not u7246 (Lbqiu6, n1740);  // ../RTL/cortexm0ds_logic.v(7566)
  and u7247 (n1741, Hnqiu6, Onqiu6);  // ../RTL/cortexm0ds_logic.v(7567)
  not u7248 (Sdphu6, n1741);  // ../RTL/cortexm0ds_logic.v(7567)
  and u7249 (Onqiu6, Vnqiu6, Coqiu6);  // ../RTL/cortexm0ds_logic.v(7568)
  not u725 (Pqdpw6, Gx2bx6);  // ../RTL/cortexm0ds_logic.v(2780)
  and u7250 (n1742, Wo1iu6, Joqiu6);  // ../RTL/cortexm0ds_logic.v(7569)
  not u7251 (Coqiu6, n1742);  // ../RTL/cortexm0ds_logic.v(7569)
  and u7252 (n1743, Qoqiu6, Xoqiu6);  // ../RTL/cortexm0ds_logic.v(7570)
  not u7253 (Joqiu6, n1743);  // ../RTL/cortexm0ds_logic.v(7570)
  and u7254 (Xoqiu6, Epqiu6, Lpqiu6);  // ../RTL/cortexm0ds_logic.v(7571)
  and u7255 (Lpqiu6, Spqiu6, Zpqiu6);  // ../RTL/cortexm0ds_logic.v(7572)
  and u7256 (Zpqiu6, Gqqiu6, Nqqiu6);  // ../RTL/cortexm0ds_logic.v(7573)
  and u7257 (n1744, ECOREVNUM[16], Uqqiu6);  // ../RTL/cortexm0ds_logic.v(7574)
  not u7258 (Nqqiu6, n1744);  // ../RTL/cortexm0ds_logic.v(7574)
  and u7259 (Gqqiu6, Brqiu6, Irqiu6);  // ../RTL/cortexm0ds_logic.v(7575)
  buf u726 (Trgpw6[6], Hi9bx6);  // ../RTL/cortexm0ds_logic.v(2376)
  and u7260 (n1745, ECOREVNUM[12], Prqiu6);  // ../RTL/cortexm0ds_logic.v(7576)
  not u7261 (Brqiu6, n1745);  // ../RTL/cortexm0ds_logic.v(7576)
  and u7262 (Spqiu6, Wrqiu6, Dsqiu6);  // ../RTL/cortexm0ds_logic.v(7577)
  and u7263 (n1746, ECOREVNUM[4], Ksqiu6);  // ../RTL/cortexm0ds_logic.v(7578)
  not u7264 (Dsqiu6, n1746);  // ../RTL/cortexm0ds_logic.v(7578)
  and u7265 (n1747, ECOREVNUM[8], Rsqiu6);  // ../RTL/cortexm0ds_logic.v(7579)
  not u7266 (Wrqiu6, n1747);  // ../RTL/cortexm0ds_logic.v(7579)
  and u7267 (Epqiu6, Ysqiu6, Ftqiu6);  // ../RTL/cortexm0ds_logic.v(7580)
  and u7268 (Ftqiu6, Mtqiu6, Ttqiu6);  // ../RTL/cortexm0ds_logic.v(7581)
  and u7269 (n1748, Aygpw6[4], Jf7iu6);  // ../RTL/cortexm0ds_logic.v(7582)
  not u727 (Iqdpw6, M13bx6);  // ../RTL/cortexm0ds_logic.v(2782)
  not u7270 (Ttqiu6, n1748);  // ../RTL/cortexm0ds_logic.v(7582)
  and u7271 (Mtqiu6, Auqiu6, Huqiu6);  // ../RTL/cortexm0ds_logic.v(7583)
  and u7272 (n1749, Dhgpw6[4], Fgpiu6);  // ../RTL/cortexm0ds_logic.v(7584)
  not u7273 (Huqiu6, n1749);  // ../RTL/cortexm0ds_logic.v(7584)
  and u7274 (n1750, G4hpw6[4], Sg7iu6);  // ../RTL/cortexm0ds_logic.v(7585)
  not u7275 (Auqiu6, n1750);  // ../RTL/cortexm0ds_logic.v(7585)
  and u7276 (Ysqiu6, Ouqiu6, Vuqiu6);  // ../RTL/cortexm0ds_logic.v(7586)
  and u7277 (n1751, Togpw6[4], Vr1iu6);  // ../RTL/cortexm0ds_logic.v(7587)
  not u7278 (Vuqiu6, n1751);  // ../RTL/cortexm0ds_logic.v(7587)
  and u7279 (n1752, Gtgpw6[4], Cs1iu6);  // ../RTL/cortexm0ds_logic.v(7588)
  buf u728 (Trgpw6[5], C1fax6);  // ../RTL/cortexm0ds_logic.v(2376)
  not u7280 (Ouqiu6, n1752);  // ../RTL/cortexm0ds_logic.v(7588)
  and u7281 (Qoqiu6, Cvqiu6, Jvqiu6);  // ../RTL/cortexm0ds_logic.v(7589)
  and u7282 (Jvqiu6, Qvqiu6, Xvqiu6);  // ../RTL/cortexm0ds_logic.v(7590)
  and u7283 (Xvqiu6, Ewqiu6, Lwqiu6);  // ../RTL/cortexm0ds_logic.v(7591)
  and u7284 (n1753, E1hpw6[4], Zt1iu6);  // ../RTL/cortexm0ds_logic.v(7592)
  not u7285 (Lwqiu6, n1753);  // ../RTL/cortexm0ds_logic.v(7592)
  and u7286 (Ewqiu6, Swqiu6, Zwqiu6);  // ../RTL/cortexm0ds_logic.v(7593)
  and u7287 (n1754, Ar1iu6, Fkfpw6[4]);  // ../RTL/cortexm0ds_logic.v(7594)
  not u7288 (Zwqiu6, n1754);  // ../RTL/cortexm0ds_logic.v(7594)
  and u7289 (n1755, HRDATA[4], St1iu6);  // ../RTL/cortexm0ds_logic.v(7595)
  not u729 (Bqdpw6, S53bx6);  // ../RTL/cortexm0ds_logic.v(2784)
  not u7290 (Swqiu6, n1755);  // ../RTL/cortexm0ds_logic.v(7595)
  and u7291 (Qvqiu6, Gxqiu6, Nxqiu6);  // ../RTL/cortexm0ds_logic.v(7596)
  and u7292 (n1756, Gqgpw6[4], Xs1iu6);  // ../RTL/cortexm0ds_logic.v(7597)
  not u7293 (Nxqiu6, n1756);  // ../RTL/cortexm0ds_logic.v(7597)
  and u7294 (n1757, Trgpw6[4], Dw1iu6);  // ../RTL/cortexm0ds_logic.v(7598)
  not u7295 (Gxqiu6, n1757);  // ../RTL/cortexm0ds_logic.v(7598)
  and u7296 (Cvqiu6, Uxqiu6, Byqiu6);  // ../RTL/cortexm0ds_logic.v(7599)
  and u7297 (Byqiu6, Iyqiu6, Pyqiu6);  // ../RTL/cortexm0ds_logic.v(7600)
  and u7298 (n1758, Wyqiu6, Dzqiu6);  // ../RTL/cortexm0ds_logic.v(7601)
  not u7299 (Pyqiu6, n1758);  // ../RTL/cortexm0ds_logic.v(7601)
  buf u73 (vis_r8_o[30], Qkrax6);  // ../RTL/cortexm0ds_logic.v(2579)
  buf u730 (Trgpw6[4], Y2fax6);  // ../RTL/cortexm0ds_logic.v(2376)
  and u7300 (Iyqiu6, Kzqiu6, Rzqiu6);  // ../RTL/cortexm0ds_logic.v(7602)
  and u7301 (n1759, K7hpw6[4], Kw1iu6);  // ../RTL/cortexm0ds_logic.v(7603)
  not u7302 (Rzqiu6, n1759);  // ../RTL/cortexm0ds_logic.v(7603)
  and u7303 (n1760, vis_pc_o[3], Iv1iu6);  // ../RTL/cortexm0ds_logic.v(7604)
  not u7304 (Kzqiu6, n1760);  // ../RTL/cortexm0ds_logic.v(7604)
  and u7305 (Uxqiu6, Yzqiu6, F0riu6);  // ../RTL/cortexm0ds_logic.v(7605)
  and u7306 (n1761, Jshpw6[4], Bo1iu6);  // ../RTL/cortexm0ds_logic.v(7606)
  not u7307 (Vnqiu6, n1761);  // ../RTL/cortexm0ds_logic.v(7606)
  and u7308 (Hnqiu6, M0riu6, T0riu6);  // ../RTL/cortexm0ds_logic.v(7607)
  and u7309 (n1762, Qwpiu6, Cynhu6);  // ../RTL/cortexm0ds_logic.v(7608)
  not u731 (Updpw6, Y93bx6);  // ../RTL/cortexm0ds_logic.v(2786)
  not u7310 (T0riu6, n1762);  // ../RTL/cortexm0ds_logic.v(7608)
  and u7311 (n1763, Uthpw6[4], Sf1iu6);  // ../RTL/cortexm0ds_logic.v(7609)
  not u7312 (M0riu6, n1763);  // ../RTL/cortexm0ds_logic.v(7609)
  and u7313 (n1764, A1riu6, H1riu6);  // ../RTL/cortexm0ds_logic.v(7610)
  not u7314 (Ldphu6, n1764);  // ../RTL/cortexm0ds_logic.v(7610)
  and u7315 (H1riu6, O1riu6, V1riu6);  // ../RTL/cortexm0ds_logic.v(7611)
  and u7316 (n1765, Wo1iu6, C2riu6);  // ../RTL/cortexm0ds_logic.v(7612)
  not u7317 (O1riu6, n1765);  // ../RTL/cortexm0ds_logic.v(7612)
  and u7318 (n1766, J2riu6, Q2riu6);  // ../RTL/cortexm0ds_logic.v(7613)
  not u7319 (C2riu6, n1766);  // ../RTL/cortexm0ds_logic.v(7613)
  buf u732 (Trgpw6[3], U4fax6);  // ../RTL/cortexm0ds_logic.v(2376)
  and u7320 (Q2riu6, X2riu6, E3riu6);  // ../RTL/cortexm0ds_logic.v(7614)
  and u7321 (E3riu6, L3riu6, S3riu6);  // ../RTL/cortexm0ds_logic.v(7615)
  and u7322 (S3riu6, Z3riu6, G4riu6);  // ../RTL/cortexm0ds_logic.v(7616)
  and u7323 (n1767, ECOREVNUM[17], Uqqiu6);  // ../RTL/cortexm0ds_logic.v(7617)
  not u7324 (G4riu6, n1767);  // ../RTL/cortexm0ds_logic.v(7617)
  and u7325 (Z3riu6, N4riu6, Irqiu6);  // ../RTL/cortexm0ds_logic.v(7618)
  not u7326 (Irqiu6, U4riu6);  // ../RTL/cortexm0ds_logic.v(7619)
  and u7327 (n1768, ECOREVNUM[13], Prqiu6);  // ../RTL/cortexm0ds_logic.v(7620)
  not u7328 (N4riu6, n1768);  // ../RTL/cortexm0ds_logic.v(7620)
  and u7329 (L3riu6, B5riu6, I5riu6);  // ../RTL/cortexm0ds_logic.v(7621)
  not u733 (Npdpw6, Ee3bx6);  // ../RTL/cortexm0ds_logic.v(2788)
  and u7330 (n1769, ECOREVNUM[5], Ksqiu6);  // ../RTL/cortexm0ds_logic.v(7622)
  not u7331 (I5riu6, n1769);  // ../RTL/cortexm0ds_logic.v(7622)
  and u7332 (n1770, ECOREVNUM[9], Rsqiu6);  // ../RTL/cortexm0ds_logic.v(7623)
  not u7333 (B5riu6, n1770);  // ../RTL/cortexm0ds_logic.v(7623)
  and u7334 (X2riu6, P5riu6, W5riu6);  // ../RTL/cortexm0ds_logic.v(7624)
  and u7335 (W5riu6, D6riu6, K6riu6);  // ../RTL/cortexm0ds_logic.v(7625)
  and u7336 (n1771, Togpw6[5], Vr1iu6);  // ../RTL/cortexm0ds_logic.v(7626)
  not u7337 (K6riu6, n1771);  // ../RTL/cortexm0ds_logic.v(7626)
  and u7338 (n1772, Gtgpw6[5], Cs1iu6);  // ../RTL/cortexm0ds_logic.v(7627)
  not u7339 (D6riu6, n1772);  // ../RTL/cortexm0ds_logic.v(7627)
  buf u734 (vis_r4_o[0], Bauax6);  // ../RTL/cortexm0ds_logic.v(2626)
  and u7340 (P5riu6, R6riu6, Y6riu6);  // ../RTL/cortexm0ds_logic.v(7628)
  and u7341 (n1773, Ar1iu6, Fkfpw6[5]);  // ../RTL/cortexm0ds_logic.v(7629)
  not u7342 (Y6riu6, n1773);  // ../RTL/cortexm0ds_logic.v(7629)
  and u7343 (n1774, HRDATA[5], St1iu6);  // ../RTL/cortexm0ds_logic.v(7630)
  not u7344 (R6riu6, n1774);  // ../RTL/cortexm0ds_logic.v(7630)
  and u7345 (J2riu6, F7riu6, M7riu6);  // ../RTL/cortexm0ds_logic.v(7631)
  and u7346 (M7riu6, T7riu6, A8riu6);  // ../RTL/cortexm0ds_logic.v(7632)
  and u7347 (A8riu6, H8riu6, O8riu6);  // ../RTL/cortexm0ds_logic.v(7633)
  and u7348 (n1775, E1hpw6[5], Zt1iu6);  // ../RTL/cortexm0ds_logic.v(7634)
  not u7349 (O8riu6, n1775);  // ../RTL/cortexm0ds_logic.v(7634)
  not u735 (Gpdpw6, Ki3bx6);  // ../RTL/cortexm0ds_logic.v(2790)
  and u7350 (n1776, Gqgpw6[5], Xs1iu6);  // ../RTL/cortexm0ds_logic.v(7635)
  not u7351 (H8riu6, n1776);  // ../RTL/cortexm0ds_logic.v(7635)
  and u7352 (T7riu6, V8riu6, C9riu6);  // ../RTL/cortexm0ds_logic.v(7636)
  and u7353 (n1777, Trgpw6[5], Dw1iu6);  // ../RTL/cortexm0ds_logic.v(7637)
  not u7354 (C9riu6, n1777);  // ../RTL/cortexm0ds_logic.v(7637)
  and u7355 (n1778, K7hpw6[5], Kw1iu6);  // ../RTL/cortexm0ds_logic.v(7638)
  not u7356 (V8riu6, n1778);  // ../RTL/cortexm0ds_logic.v(7638)
  and u7357 (F7riu6, J9riu6, Q9riu6);  // ../RTL/cortexm0ds_logic.v(7639)
  and u7358 (Q9riu6, F0riu6, X9riu6);  // ../RTL/cortexm0ds_logic.v(7640)
  and u7359 (n1779, vis_pc_o[4], Iv1iu6);  // ../RTL/cortexm0ds_logic.v(7641)
  buf u736 (Trgpw6[27], Zycbx6);  // ../RTL/cortexm0ds_logic.v(2376)
  not u7360 (X9riu6, n1779);  // ../RTL/cortexm0ds_logic.v(7641)
  and u7361 (J9riu6, Eariu6, Lariu6);  // ../RTL/cortexm0ds_logic.v(7642)
  and u7362 (A1riu6, Sariu6, Zariu6);  // ../RTL/cortexm0ds_logic.v(7643)
  and u7363 (n1780, Jshpw6[5], Bo1iu6);  // ../RTL/cortexm0ds_logic.v(7644)
  not u7364 (Zariu6, n1780);  // ../RTL/cortexm0ds_logic.v(7644)
  and u7365 (n1781, Uthpw6[5], Sf1iu6);  // ../RTL/cortexm0ds_logic.v(7645)
  not u7366 (Sariu6, n1781);  // ../RTL/cortexm0ds_logic.v(7645)
  and u7367 (n1782, Gbriu6, Nbriu6);  // ../RTL/cortexm0ds_logic.v(7646)
  not u7368 (Edphu6, n1782);  // ../RTL/cortexm0ds_logic.v(7646)
  and u7369 (Nbriu6, Ubriu6, Bcriu6);  // ../RTL/cortexm0ds_logic.v(7647)
  not u737 (Zodpw6, Om3bx6);  // ../RTL/cortexm0ds_logic.v(2792)
  and u7370 (n1783, Wo1iu6, Icriu6);  // ../RTL/cortexm0ds_logic.v(7648)
  not u7371 (Ubriu6, n1783);  // ../RTL/cortexm0ds_logic.v(7648)
  and u7372 (n1784, Pcriu6, Wcriu6);  // ../RTL/cortexm0ds_logic.v(7649)
  not u7373 (Icriu6, n1784);  // ../RTL/cortexm0ds_logic.v(7649)
  and u7374 (Wcriu6, Ddriu6, Kdriu6);  // ../RTL/cortexm0ds_logic.v(7650)
  and u7375 (Kdriu6, Rdriu6, Ydriu6);  // ../RTL/cortexm0ds_logic.v(7651)
  and u7376 (Ydriu6, Feriu6, Reqiu6);  // ../RTL/cortexm0ds_logic.v(7652)
  or u7377 (n1785, U4riu6, Ve7iu6);  // ../RTL/cortexm0ds_logic.v(7653)
  not u7378 (Feriu6, n1785);  // ../RTL/cortexm0ds_logic.v(7653)
  and u7379 (Rdriu6, Meriu6, Teriu6);  // ../RTL/cortexm0ds_logic.v(7654)
  buf u738 (Trgpw6[25], Mgeax6);  // ../RTL/cortexm0ds_logic.v(2376)
  and u7380 (n1786, ECOREVNUM[14], Prqiu6);  // ../RTL/cortexm0ds_logic.v(7655)
  not u7381 (Teriu6, n1786);  // ../RTL/cortexm0ds_logic.v(7655)
  and u7382 (n1787, ECOREVNUM[18], Uqqiu6);  // ../RTL/cortexm0ds_logic.v(7656)
  not u7383 (Meriu6, n1787);  // ../RTL/cortexm0ds_logic.v(7656)
  and u7384 (Ddriu6, Afriu6, Hfriu6);  // ../RTL/cortexm0ds_logic.v(7657)
  and u7385 (Hfriu6, Ofriu6, Vfriu6);  // ../RTL/cortexm0ds_logic.v(7658)
  and u7386 (n1788, ECOREVNUM[6], Ksqiu6);  // ../RTL/cortexm0ds_logic.v(7659)
  not u7387 (Vfriu6, n1788);  // ../RTL/cortexm0ds_logic.v(7659)
  and u7388 (n1789, ECOREVNUM[10], Rsqiu6);  // ../RTL/cortexm0ds_logic.v(7660)
  not u7389 (Ofriu6, n1789);  // ../RTL/cortexm0ds_logic.v(7660)
  not u739 (Sodpw6, Sq3bx6);  // ../RTL/cortexm0ds_logic.v(2794)
  and u7390 (Afriu6, Cgriu6, Jgriu6);  // ../RTL/cortexm0ds_logic.v(7661)
  and u7391 (n1790, Togpw6[6], Vr1iu6);  // ../RTL/cortexm0ds_logic.v(7662)
  not u7392 (Jgriu6, n1790);  // ../RTL/cortexm0ds_logic.v(7662)
  and u7393 (n1791, Gtgpw6[6], Cs1iu6);  // ../RTL/cortexm0ds_logic.v(7663)
  not u7394 (Cgriu6, n1791);  // ../RTL/cortexm0ds_logic.v(7663)
  and u7395 (Pcriu6, Qgriu6, Xgriu6);  // ../RTL/cortexm0ds_logic.v(7664)
  and u7396 (Xgriu6, Ehriu6, Lhriu6);  // ../RTL/cortexm0ds_logic.v(7665)
  and u7397 (Lhriu6, Shriu6, Zhriu6);  // ../RTL/cortexm0ds_logic.v(7666)
  and u7398 (n1792, E1hpw6[6], Zt1iu6);  // ../RTL/cortexm0ds_logic.v(7667)
  not u7399 (Zhriu6, n1792);  // ../RTL/cortexm0ds_logic.v(7667)
  not u74 (Zehpw6[0], n7[0]);  // ../RTL/cortexm0ds_logic.v(3185)
  buf u740 (Trgpw6[24], Jieax6);  // ../RTL/cortexm0ds_logic.v(2376)
  and u7400 (Shriu6, Giriu6, Niriu6);  // ../RTL/cortexm0ds_logic.v(7668)
  and u7401 (n1793, Ar1iu6, Fkfpw6[6]);  // ../RTL/cortexm0ds_logic.v(7669)
  not u7402 (Niriu6, n1793);  // ../RTL/cortexm0ds_logic.v(7669)
  and u7403 (n1794, HRDATA[6], St1iu6);  // ../RTL/cortexm0ds_logic.v(7670)
  not u7404 (Giriu6, n1794);  // ../RTL/cortexm0ds_logic.v(7670)
  and u7405 (Ehriu6, Uiriu6, Bjriu6);  // ../RTL/cortexm0ds_logic.v(7671)
  and u7406 (n1795, Gqgpw6[6], Xs1iu6);  // ../RTL/cortexm0ds_logic.v(7672)
  not u7407 (Bjriu6, n1795);  // ../RTL/cortexm0ds_logic.v(7672)
  and u7408 (n1796, Trgpw6[6], Dw1iu6);  // ../RTL/cortexm0ds_logic.v(7673)
  not u7409 (Uiriu6, n1796);  // ../RTL/cortexm0ds_logic.v(7673)
  buf u741 (Togpw6[3], Iddax6);  // ../RTL/cortexm0ds_logic.v(2378)
  and u7410 (Qgriu6, Ijriu6, Pjriu6);  // ../RTL/cortexm0ds_logic.v(7674)
  and u7411 (Pjriu6, Wjriu6, Dkriu6);  // ../RTL/cortexm0ds_logic.v(7675)
  and u7412 (n1797, K7hpw6[6], Kw1iu6);  // ../RTL/cortexm0ds_logic.v(7676)
  not u7413 (Dkriu6, n1797);  // ../RTL/cortexm0ds_logic.v(7676)
  and u7414 (n1798, vis_pc_o[5], Iv1iu6);  // ../RTL/cortexm0ds_logic.v(7677)
  not u7415 (Wjriu6, n1798);  // ../RTL/cortexm0ds_logic.v(7677)
  and u7416 (Ijriu6, Kkriu6, Lariu6);  // ../RTL/cortexm0ds_logic.v(7678)
  and u7417 (Gbriu6, Rkriu6, Ykriu6);  // ../RTL/cortexm0ds_logic.v(7679)
  and u7418 (n1799, Jshpw6[6], Bo1iu6);  // ../RTL/cortexm0ds_logic.v(7680)
  not u7419 (Ykriu6, n1799);  // ../RTL/cortexm0ds_logic.v(7680)
  buf u742 (Engpw6[28], K6gax6);  // ../RTL/cortexm0ds_logic.v(2368)
  and u7420 (n1800, Uthpw6[6], Sf1iu6);  // ../RTL/cortexm0ds_logic.v(7681)
  not u7421 (Rkriu6, n1800);  // ../RTL/cortexm0ds_logic.v(7681)
  and u7422 (n1801, Flriu6, Mlriu6);  // ../RTL/cortexm0ds_logic.v(7682)
  not u7423 (Xcphu6, n1801);  // ../RTL/cortexm0ds_logic.v(7682)
  and u7424 (n1802, Uthpw6[7], Sf1iu6);  // ../RTL/cortexm0ds_logic.v(7683)
  not u7425 (Mlriu6, n1802);  // ../RTL/cortexm0ds_logic.v(7683)
  and u7426 (Flriu6, Tlriu6, Amriu6);  // ../RTL/cortexm0ds_logic.v(7684)
  and u7427 (n1803, Wo1iu6, Hmriu6);  // ../RTL/cortexm0ds_logic.v(7685)
  not u7428 (Amriu6, n1803);  // ../RTL/cortexm0ds_logic.v(7685)
  and u7429 (n1804, Omriu6, Vmriu6);  // ../RTL/cortexm0ds_logic.v(7686)
  buf u743 (Plgpw6[28], H8gax6);  // ../RTL/cortexm0ds_logic.v(2369)
  not u7430 (Hmriu6, n1804);  // ../RTL/cortexm0ds_logic.v(7686)
  and u7431 (Vmriu6, Cnriu6, Jnriu6);  // ../RTL/cortexm0ds_logic.v(7687)
  and u7432 (Jnriu6, Qnriu6, Xnriu6);  // ../RTL/cortexm0ds_logic.v(7688)
  and u7433 (Xnriu6, Eoriu6, Loriu6);  // ../RTL/cortexm0ds_logic.v(7689)
  and u7434 (n1805, ECOREVNUM[15], Prqiu6);  // ../RTL/cortexm0ds_logic.v(7690)
  not u7435 (Loriu6, n1805);  // ../RTL/cortexm0ds_logic.v(7690)
  and u7436 (Prqiu6, Soriu6, A2qiu6);  // ../RTL/cortexm0ds_logic.v(7691)
  and u7437 (Soriu6, Dzqiu6, Cvciu6);  // ../RTL/cortexm0ds_logic.v(7692)
  and u7438 (n1806, ECOREVNUM[19], Uqqiu6);  // ../RTL/cortexm0ds_logic.v(7693)
  not u7439 (Eoriu6, n1806);  // ../RTL/cortexm0ds_logic.v(7693)
  buf u744 (Uthpw6[31], Uunpw6);  // ../RTL/cortexm0ds_logic.v(1882)
  and u7440 (Uqqiu6, Zoriu6, Wyqiu6);  // ../RTL/cortexm0ds_logic.v(7694)
  or u7441 (n1807, Fl6iu6, Mfqiu6);  // ../RTL/cortexm0ds_logic.v(7695)
  not u7442 (Zoriu6, n1807);  // ../RTL/cortexm0ds_logic.v(7695)
  and u7443 (Qnriu6, Gpriu6, Npriu6);  // ../RTL/cortexm0ds_logic.v(7696)
  and u7444 (n1808, ECOREVNUM[7], Ksqiu6);  // ../RTL/cortexm0ds_logic.v(7697)
  not u7445 (Npriu6, n1808);  // ../RTL/cortexm0ds_logic.v(7697)
  and u7446 (Ksqiu6, Upriu6, A2qiu6);  // ../RTL/cortexm0ds_logic.v(7698)
  and u7447 (Upriu6, Bqriu6, Cvciu6);  // ../RTL/cortexm0ds_logic.v(7699)
  and u7448 (n1809, ECOREVNUM[11], Rsqiu6);  // ../RTL/cortexm0ds_logic.v(7700)
  not u7449 (Gpriu6, n1809);  // ../RTL/cortexm0ds_logic.v(7700)
  buf u745 (Uthpw6[30], X42qw6);  // ../RTL/cortexm0ds_logic.v(1882)
  and u7450 (Rsqiu6, Iqriu6, X8hpw6[4]);  // ../RTL/cortexm0ds_logic.v(7701)
  and u7451 (Cnriu6, Pqriu6, Wqriu6);  // ../RTL/cortexm0ds_logic.v(7702)
  and u7452 (Wqriu6, Drriu6, Krriu6);  // ../RTL/cortexm0ds_logic.v(7703)
  and u7453 (n1810, Togpw6[7], Vr1iu6);  // ../RTL/cortexm0ds_logic.v(7704)
  not u7454 (Krriu6, n1810);  // ../RTL/cortexm0ds_logic.v(7704)
  and u7455 (n1811, Gtgpw6[7], Cs1iu6);  // ../RTL/cortexm0ds_logic.v(7705)
  not u7456 (Drriu6, n1811);  // ../RTL/cortexm0ds_logic.v(7705)
  and u7457 (Pqriu6, Rrriu6, Yrriu6);  // ../RTL/cortexm0ds_logic.v(7706)
  and u7458 (n1812, Ar1iu6, Fkfpw6[7]);  // ../RTL/cortexm0ds_logic.v(7707)
  not u7459 (Yrriu6, n1812);  // ../RTL/cortexm0ds_logic.v(7707)
  buf u746 (Uthpw6[29], Rr3qw6);  // ../RTL/cortexm0ds_logic.v(1882)
  and u7460 (n1813, HRDATA[7], St1iu6);  // ../RTL/cortexm0ds_logic.v(7708)
  not u7461 (Rrriu6, n1813);  // ../RTL/cortexm0ds_logic.v(7708)
  and u7462 (Omriu6, Fsriu6, Msriu6);  // ../RTL/cortexm0ds_logic.v(7709)
  and u7463 (Msriu6, Tsriu6, Atriu6);  // ../RTL/cortexm0ds_logic.v(7710)
  and u7464 (Atriu6, Htriu6, Otriu6);  // ../RTL/cortexm0ds_logic.v(7711)
  and u7465 (n1814, E1hpw6[7], Zt1iu6);  // ../RTL/cortexm0ds_logic.v(7712)
  not u7466 (Otriu6, n1814);  // ../RTL/cortexm0ds_logic.v(7712)
  and u7467 (n1815, Gqgpw6[7], Xs1iu6);  // ../RTL/cortexm0ds_logic.v(7713)
  not u7468 (Htriu6, n1815);  // ../RTL/cortexm0ds_logic.v(7713)
  and u7469 (Tsriu6, Vtriu6, Curiu6);  // ../RTL/cortexm0ds_logic.v(7714)
  buf u747 (X8hpw6[5], Zm8ax6);  // ../RTL/cortexm0ds_logic.v(2046)
  and u7470 (n1816, Trgpw6[7], Dw1iu6);  // ../RTL/cortexm0ds_logic.v(7715)
  not u7471 (Curiu6, n1816);  // ../RTL/cortexm0ds_logic.v(7715)
  and u7472 (n1817, K7hpw6[7], Kw1iu6);  // ../RTL/cortexm0ds_logic.v(7716)
  not u7473 (Vtriu6, n1817);  // ../RTL/cortexm0ds_logic.v(7716)
  and u7474 (Fsriu6, Juriu6, Quriu6);  // ../RTL/cortexm0ds_logic.v(7717)
  and u7475 (Quriu6, F0riu6, Xuriu6);  // ../RTL/cortexm0ds_logic.v(7718)
  and u7476 (n1818, vis_pc_o[6], Iv1iu6);  // ../RTL/cortexm0ds_logic.v(7719)
  not u7477 (Xuriu6, n1818);  // ../RTL/cortexm0ds_logic.v(7719)
  and u7478 (F0riu6, Evriu6, Lvriu6);  // ../RTL/cortexm0ds_logic.v(7720)
  and u7479 (Lvriu6, Wzpiu6, Svriu6);  // ../RTL/cortexm0ds_logic.v(7721)
  buf u748 (X8hpw6[4], Di3qw6);  // ../RTL/cortexm0ds_logic.v(2046)
  and u7480 (Wzpiu6, Zvriu6, Reqiu6);  // ../RTL/cortexm0ds_logic.v(7722)
  and u7481 (n1819, Gwriu6, Wyqiu6);  // ../RTL/cortexm0ds_logic.v(7723)
  not u7482 (Zvriu6, n1819);  // ../RTL/cortexm0ds_logic.v(7723)
  or u7483 (n1820, Nwriu6, X8hpw6[4]);  // ../RTL/cortexm0ds_logic.v(7724)
  not u7484 (Gwriu6, n1820);  // ../RTL/cortexm0ds_logic.v(7724)
  and u7485 (Evriu6, Uwriu6, Bxriu6);  // ../RTL/cortexm0ds_logic.v(7725)
  and u7486 (n1821, Ixriu6, Fl6iu6);  // ../RTL/cortexm0ds_logic.v(7726)
  not u7487 (Bxriu6, n1821);  // ../RTL/cortexm0ds_logic.v(7726)
  and u7488 (Juriu6, Pxriu6, Lariu6);  // ../RTL/cortexm0ds_logic.v(7727)
  and u7489 (Lariu6, Wxriu6, Dyriu6);  // ../RTL/cortexm0ds_logic.v(7728)
  buf u749 (X8hpw6[3], D43qw6);  // ../RTL/cortexm0ds_logic.v(2046)
  and u7490 (n1822, Kyriu6, Ixriu6);  // ../RTL/cortexm0ds_logic.v(7729)
  not u7491 (Dyriu6, n1822);  // ../RTL/cortexm0ds_logic.v(7729)
  or u7492 (n1823, Fl6iu6, Vm6iu6);  // ../RTL/cortexm0ds_logic.v(7730)
  not u7493 (Kyriu6, n1823);  // ../RTL/cortexm0ds_logic.v(7730)
  and u7494 (n1824, Ryriu6, Cvciu6);  // ../RTL/cortexm0ds_logic.v(7731)
  not u7495 (Wxriu6, n1824);  // ../RTL/cortexm0ds_logic.v(7731)
  and u7496 (n1825, Jshpw6[7], Bo1iu6);  // ../RTL/cortexm0ds_logic.v(7732)
  not u7497 (Tlriu6, n1825);  // ../RTL/cortexm0ds_logic.v(7732)
  and u7498 (n1826, Yyriu6, Fzriu6);  // ../RTL/cortexm0ds_logic.v(7733)
  not u7499 (Qcphu6, n1826);  // ../RTL/cortexm0ds_logic.v(7733)
  buf u75 (vis_r5_o[16], Cdwpw6);  // ../RTL/cortexm0ds_logic.v(1909)
  buf u750 (X8hpw6[1], Le2qw6);  // ../RTL/cortexm0ds_logic.v(2046)
  and u7500 (n1827, Uthpw6[8], Sf1iu6);  // ../RTL/cortexm0ds_logic.v(7734)
  not u7501 (Fzriu6, n1827);  // ../RTL/cortexm0ds_logic.v(7734)
  and u7502 (Yyriu6, Mzriu6, Tzriu6);  // ../RTL/cortexm0ds_logic.v(7735)
  and u7503 (n1828, Wo1iu6, A0siu6);  // ../RTL/cortexm0ds_logic.v(7736)
  not u7504 (Tzriu6, n1828);  // ../RTL/cortexm0ds_logic.v(7736)
  and u7505 (n1829, H0siu6, O0siu6);  // ../RTL/cortexm0ds_logic.v(7737)
  not u7506 (A0siu6, n1829);  // ../RTL/cortexm0ds_logic.v(7737)
  and u7507 (O0siu6, V0siu6, C1siu6);  // ../RTL/cortexm0ds_logic.v(7738)
  and u7508 (C1siu6, J1siu6, Q1siu6);  // ../RTL/cortexm0ds_logic.v(7739)
  and u7509 (n1830, Gtgpw6[8], Cs1iu6);  // ../RTL/cortexm0ds_logic.v(7740)
  buf u751 (R2hpw6[2], P0bax6);  // ../RTL/cortexm0ds_logic.v(2268)
  not u7510 (Q1siu6, n1830);  // ../RTL/cortexm0ds_logic.v(7740)
  and u7511 (J1siu6, X1siu6, Reqiu6);  // ../RTL/cortexm0ds_logic.v(7741)
  and u7512 (n1831, Togpw6[8], Vr1iu6);  // ../RTL/cortexm0ds_logic.v(7742)
  not u7513 (X1siu6, n1831);  // ../RTL/cortexm0ds_logic.v(7742)
  and u7514 (V0siu6, E2siu6, L2siu6);  // ../RTL/cortexm0ds_logic.v(7743)
  and u7515 (n1832, E1hpw6[8], Zt1iu6);  // ../RTL/cortexm0ds_logic.v(7744)
  not u7516 (L2siu6, n1832);  // ../RTL/cortexm0ds_logic.v(7744)
  and u7517 (E2siu6, S2siu6, Z2siu6);  // ../RTL/cortexm0ds_logic.v(7745)
  and u7518 (n1833, Ar1iu6, Fkfpw6[8]);  // ../RTL/cortexm0ds_logic.v(7746)
  not u7519 (Z2siu6, n1833);  // ../RTL/cortexm0ds_logic.v(7746)
  buf u752 (R2hpw6[1], L2bax6);  // ../RTL/cortexm0ds_logic.v(2268)
  and u7520 (n1834, HRDATA[8], St1iu6);  // ../RTL/cortexm0ds_logic.v(7747)
  not u7521 (S2siu6, n1834);  // ../RTL/cortexm0ds_logic.v(7747)
  and u7522 (H0siu6, G3siu6, N3siu6);  // ../RTL/cortexm0ds_logic.v(7748)
  and u7523 (N3siu6, U3siu6, B4siu6);  // ../RTL/cortexm0ds_logic.v(7749)
  and u7524 (n1835, K7hpw6[8], Kw1iu6);  // ../RTL/cortexm0ds_logic.v(7750)
  not u7525 (B4siu6, n1835);  // ../RTL/cortexm0ds_logic.v(7750)
  and u7526 (U3siu6, I4siu6, P4siu6);  // ../RTL/cortexm0ds_logic.v(7751)
  and u7527 (n1836, Gqgpw6[8], Xs1iu6);  // ../RTL/cortexm0ds_logic.v(7752)
  not u7528 (P4siu6, n1836);  // ../RTL/cortexm0ds_logic.v(7752)
  and u7529 (n1837, Trgpw6[8], Dw1iu6);  // ../RTL/cortexm0ds_logic.v(7753)
  buf u753 (Jfgpw6[0], Yzspw6);  // ../RTL/cortexm0ds_logic.v(2010)
  not u7530 (I4siu6, n1837);  // ../RTL/cortexm0ds_logic.v(7753)
  and u7531 (G3siu6, W4siu6, D5siu6);  // ../RTL/cortexm0ds_logic.v(7754)
  and u7532 (n1838, vis_pc_o[7], Iv1iu6);  // ../RTL/cortexm0ds_logic.v(7755)
  not u7533 (D5siu6, n1838);  // ../RTL/cortexm0ds_logic.v(7755)
  and u7534 (n1839, Jshpw6[8], Bo1iu6);  // ../RTL/cortexm0ds_logic.v(7756)
  not u7535 (Mzriu6, n1839);  // ../RTL/cortexm0ds_logic.v(7756)
  and u7536 (n1840, K5siu6, R5siu6);  // ../RTL/cortexm0ds_logic.v(7757)
  not u7537 (Jcphu6, n1840);  // ../RTL/cortexm0ds_logic.v(7757)
  and u7538 (n1841, Uthpw6[9], Sf1iu6);  // ../RTL/cortexm0ds_logic.v(7758)
  not u7539 (R5siu6, n1841);  // ../RTL/cortexm0ds_logic.v(7758)
  buf u754 (Jshpw6[20], Nwdbx6);  // ../RTL/cortexm0ds_logic.v(2372)
  and u7540 (K5siu6, Y5siu6, F6siu6);  // ../RTL/cortexm0ds_logic.v(7759)
  and u7541 (n1842, Wo1iu6, M6siu6);  // ../RTL/cortexm0ds_logic.v(7760)
  not u7542 (F6siu6, n1842);  // ../RTL/cortexm0ds_logic.v(7760)
  and u7543 (n1843, T6siu6, A7siu6);  // ../RTL/cortexm0ds_logic.v(7761)
  not u7544 (M6siu6, n1843);  // ../RTL/cortexm0ds_logic.v(7761)
  and u7545 (A7siu6, H7siu6, O7siu6);  // ../RTL/cortexm0ds_logic.v(7762)
  and u7546 (O7siu6, V7siu6, C8siu6);  // ../RTL/cortexm0ds_logic.v(7763)
  and u7547 (n1844, Gtgpw6[9], Cs1iu6);  // ../RTL/cortexm0ds_logic.v(7764)
  not u7548 (C8siu6, n1844);  // ../RTL/cortexm0ds_logic.v(7764)
  and u7549 (V7siu6, J8siu6, Reqiu6);  // ../RTL/cortexm0ds_logic.v(7765)
  buf u755 (Uthpw6[27], N0cbx6);  // ../RTL/cortexm0ds_logic.v(1882)
  and u7550 (n1845, Togpw6[9], Vr1iu6);  // ../RTL/cortexm0ds_logic.v(7766)
  not u7551 (J8siu6, n1845);  // ../RTL/cortexm0ds_logic.v(7766)
  and u7552 (H7siu6, Q8siu6, X8siu6);  // ../RTL/cortexm0ds_logic.v(7767)
  and u7553 (n1846, E1hpw6[9], Zt1iu6);  // ../RTL/cortexm0ds_logic.v(7768)
  not u7554 (X8siu6, n1846);  // ../RTL/cortexm0ds_logic.v(7768)
  and u7555 (Q8siu6, E9siu6, L9siu6);  // ../RTL/cortexm0ds_logic.v(7769)
  and u7556 (n1847, Ar1iu6, Fkfpw6[9]);  // ../RTL/cortexm0ds_logic.v(7770)
  not u7557 (L9siu6, n1847);  // ../RTL/cortexm0ds_logic.v(7770)
  and u7558 (n1848, HRDATA[9], St1iu6);  // ../RTL/cortexm0ds_logic.v(7771)
  not u7559 (E9siu6, n1848);  // ../RTL/cortexm0ds_logic.v(7771)
  buf u756 (Uthpw6[26], Cncbx6);  // ../RTL/cortexm0ds_logic.v(1882)
  and u7560 (T6siu6, S9siu6, Z9siu6);  // ../RTL/cortexm0ds_logic.v(7772)
  and u7561 (Z9siu6, Gasiu6, Nasiu6);  // ../RTL/cortexm0ds_logic.v(7773)
  and u7562 (n1849, K7hpw6[9], Kw1iu6);  // ../RTL/cortexm0ds_logic.v(7774)
  not u7563 (Nasiu6, n1849);  // ../RTL/cortexm0ds_logic.v(7774)
  and u7564 (Gasiu6, Uasiu6, Bbsiu6);  // ../RTL/cortexm0ds_logic.v(7775)
  and u7565 (n1850, Gqgpw6[9], Xs1iu6);  // ../RTL/cortexm0ds_logic.v(7776)
  not u7566 (Bbsiu6, n1850);  // ../RTL/cortexm0ds_logic.v(7776)
  and u7567 (n1851, Trgpw6[9], Dw1iu6);  // ../RTL/cortexm0ds_logic.v(7777)
  not u7568 (Uasiu6, n1851);  // ../RTL/cortexm0ds_logic.v(7777)
  and u7569 (S9siu6, Ibsiu6, Pbsiu6);  // ../RTL/cortexm0ds_logic.v(7778)
  buf u757 (Uthpw6[25], Fl2qw6);  // ../RTL/cortexm0ds_logic.v(1882)
  and u7570 (n1852, vis_pc_o[8], Iv1iu6);  // ../RTL/cortexm0ds_logic.v(7779)
  not u7571 (Pbsiu6, n1852);  // ../RTL/cortexm0ds_logic.v(7779)
  and u7572 (n1853, Jshpw6[9], Bo1iu6);  // ../RTL/cortexm0ds_logic.v(7780)
  not u7573 (Y5siu6, n1853);  // ../RTL/cortexm0ds_logic.v(7780)
  and u7574 (n1854, Wbsiu6, Dcsiu6);  // ../RTL/cortexm0ds_logic.v(7781)
  not u7575 (Ccphu6, n1854);  // ../RTL/cortexm0ds_logic.v(7781)
  and u7576 (n1855, Uthpw6[10], Sf1iu6);  // ../RTL/cortexm0ds_logic.v(7782)
  not u7577 (Dcsiu6, n1855);  // ../RTL/cortexm0ds_logic.v(7782)
  and u7578 (Wbsiu6, Kcsiu6, Rcsiu6);  // ../RTL/cortexm0ds_logic.v(7783)
  and u7579 (n1856, Wo1iu6, Ycsiu6);  // ../RTL/cortexm0ds_logic.v(7784)
  buf u758 (Uthpw6[23], F8dbx6);  // ../RTL/cortexm0ds_logic.v(1882)
  not u7580 (Rcsiu6, n1856);  // ../RTL/cortexm0ds_logic.v(7784)
  and u7581 (n1857, Fdsiu6, Mdsiu6);  // ../RTL/cortexm0ds_logic.v(7785)
  not u7582 (Ycsiu6, n1857);  // ../RTL/cortexm0ds_logic.v(7785)
  and u7583 (Mdsiu6, Tdsiu6, Aesiu6);  // ../RTL/cortexm0ds_logic.v(7786)
  and u7584 (Aesiu6, Hesiu6, Oesiu6);  // ../RTL/cortexm0ds_logic.v(7787)
  and u7585 (n1858, Togpw6[10], Vr1iu6);  // ../RTL/cortexm0ds_logic.v(7788)
  not u7586 (Oesiu6, n1858);  // ../RTL/cortexm0ds_logic.v(7788)
  and u7587 (Hesiu6, Vesiu6, Reqiu6);  // ../RTL/cortexm0ds_logic.v(7789)
  and u7588 (n1859, Yc7iu6, S3hhu6);  // ../RTL/cortexm0ds_logic.v(7790)
  not u7589 (Vesiu6, n1859);  // ../RTL/cortexm0ds_logic.v(7790)
  buf u759 (Uthpw6[22], Qwfbx6);  // ../RTL/cortexm0ds_logic.v(1882)
  and u7590 (Tdsiu6, Cfsiu6, Jfsiu6);  // ../RTL/cortexm0ds_logic.v(7791)
  and u7591 (n1860, HRDATA[10], St1iu6);  // ../RTL/cortexm0ds_logic.v(7792)
  not u7592 (Jfsiu6, n1860);  // ../RTL/cortexm0ds_logic.v(7792)
  and u7593 (Cfsiu6, Qfsiu6, Xfsiu6);  // ../RTL/cortexm0ds_logic.v(7793)
  and u7594 (n1861, Gtgpw6[10], Cs1iu6);  // ../RTL/cortexm0ds_logic.v(7794)
  not u7595 (Xfsiu6, n1861);  // ../RTL/cortexm0ds_logic.v(7794)
  and u7596 (n1862, Ar1iu6, Fkfpw6[10]);  // ../RTL/cortexm0ds_logic.v(7795)
  not u7597 (Qfsiu6, n1862);  // ../RTL/cortexm0ds_logic.v(7795)
  and u7598 (Fdsiu6, Egsiu6, Lgsiu6);  // ../RTL/cortexm0ds_logic.v(7796)
  and u7599 (Lgsiu6, Sgsiu6, Zgsiu6);  // ../RTL/cortexm0ds_logic.v(7797)
  buf u76 (vis_r5_o[17], Yfupw6);  // ../RTL/cortexm0ds_logic.v(1909)
  buf u760 (R4gpw6[0], Nv9bx6);  // ../RTL/cortexm0ds_logic.v(2815)
  and u7600 (n1863, Trgpw6[10], Dw1iu6);  // ../RTL/cortexm0ds_logic.v(7798)
  not u7601 (Zgsiu6, n1863);  // ../RTL/cortexm0ds_logic.v(7798)
  and u7602 (Sgsiu6, Ghsiu6, Nhsiu6);  // ../RTL/cortexm0ds_logic.v(7799)
  and u7603 (n1864, E1hpw6[10], Zt1iu6);  // ../RTL/cortexm0ds_logic.v(7800)
  not u7604 (Nhsiu6, n1864);  // ../RTL/cortexm0ds_logic.v(7800)
  and u7605 (n1865, Gqgpw6[10], Xs1iu6);  // ../RTL/cortexm0ds_logic.v(7801)
  not u7606 (Ghsiu6, n1865);  // ../RTL/cortexm0ds_logic.v(7801)
  and u7607 (Egsiu6, Uhsiu6, Bisiu6);  // ../RTL/cortexm0ds_logic.v(7802)
  and u7608 (Uhsiu6, Iisiu6, Pisiu6);  // ../RTL/cortexm0ds_logic.v(7803)
  and u7609 (n1866, K7hpw6[10], Kw1iu6);  // ../RTL/cortexm0ds_logic.v(7804)
  buf u761 (Togpw6[27], T2dbx6);  // ../RTL/cortexm0ds_logic.v(2378)
  not u7610 (Pisiu6, n1866);  // ../RTL/cortexm0ds_logic.v(7804)
  and u7611 (n1867, vis_pc_o[9], Iv1iu6);  // ../RTL/cortexm0ds_logic.v(7805)
  not u7612 (Iisiu6, n1867);  // ../RTL/cortexm0ds_logic.v(7805)
  and u7613 (n1868, Jshpw6[10], Bo1iu6);  // ../RTL/cortexm0ds_logic.v(7806)
  not u7614 (Kcsiu6, n1868);  // ../RTL/cortexm0ds_logic.v(7806)
  and u7615 (n1869, Wisiu6, Djsiu6);  // ../RTL/cortexm0ds_logic.v(7807)
  not u7616 (Vbphu6, n1869);  // ../RTL/cortexm0ds_logic.v(7807)
  and u7617 (n1870, Uthpw6[11], Sf1iu6);  // ../RTL/cortexm0ds_logic.v(7808)
  not u7618 (Djsiu6, n1870);  // ../RTL/cortexm0ds_logic.v(7808)
  and u7619 (Wisiu6, Kjsiu6, Rjsiu6);  // ../RTL/cortexm0ds_logic.v(7809)
  buf u762 (Togpw6[26], Qjcbx6);  // ../RTL/cortexm0ds_logic.v(2378)
  and u7620 (n1871, Wo1iu6, Yjsiu6);  // ../RTL/cortexm0ds_logic.v(7810)
  not u7621 (Rjsiu6, n1871);  // ../RTL/cortexm0ds_logic.v(7810)
  and u7622 (n1872, Fksiu6, Mksiu6);  // ../RTL/cortexm0ds_logic.v(7811)
  not u7623 (Yjsiu6, n1872);  // ../RTL/cortexm0ds_logic.v(7811)
  and u7624 (Mksiu6, Tksiu6, Alsiu6);  // ../RTL/cortexm0ds_logic.v(7812)
  and u7625 (Alsiu6, Hlsiu6, Olsiu6);  // ../RTL/cortexm0ds_logic.v(7813)
  and u7626 (n1873, Gtgpw6[11], Cs1iu6);  // ../RTL/cortexm0ds_logic.v(7814)
  not u7627 (Olsiu6, n1873);  // ../RTL/cortexm0ds_logic.v(7814)
  and u7628 (Hlsiu6, Vlsiu6, Reqiu6);  // ../RTL/cortexm0ds_logic.v(7815)
  and u7629 (n1874, Togpw6[11], Vr1iu6);  // ../RTL/cortexm0ds_logic.v(7816)
  buf u763 (Togpw6[25], Apcax6);  // ../RTL/cortexm0ds_logic.v(2378)
  not u7630 (Vlsiu6, n1874);  // ../RTL/cortexm0ds_logic.v(7816)
  and u7631 (Tksiu6, Cmsiu6, Jmsiu6);  // ../RTL/cortexm0ds_logic.v(7817)
  and u7632 (n1875, E1hpw6[11], Zt1iu6);  // ../RTL/cortexm0ds_logic.v(7818)
  not u7633 (Jmsiu6, n1875);  // ../RTL/cortexm0ds_logic.v(7818)
  and u7634 (Cmsiu6, Qmsiu6, Xmsiu6);  // ../RTL/cortexm0ds_logic.v(7819)
  and u7635 (n1876, Ar1iu6, Fkfpw6[11]);  // ../RTL/cortexm0ds_logic.v(7820)
  not u7636 (Xmsiu6, n1876);  // ../RTL/cortexm0ds_logic.v(7820)
  and u7637 (n1877, HRDATA[11], St1iu6);  // ../RTL/cortexm0ds_logic.v(7821)
  not u7638 (Qmsiu6, n1877);  // ../RTL/cortexm0ds_logic.v(7821)
  and u7639 (Fksiu6, Ensiu6, Lnsiu6);  // ../RTL/cortexm0ds_logic.v(7822)
  buf u764 (Togpw6[23], K5hbx6);  // ../RTL/cortexm0ds_logic.v(2378)
  and u7640 (Lnsiu6, Snsiu6, Znsiu6);  // ../RTL/cortexm0ds_logic.v(7823)
  and u7641 (n1878, K7hpw6[11], Kw1iu6);  // ../RTL/cortexm0ds_logic.v(7824)
  not u7642 (Znsiu6, n1878);  // ../RTL/cortexm0ds_logic.v(7824)
  and u7643 (Snsiu6, Gosiu6, Nosiu6);  // ../RTL/cortexm0ds_logic.v(7825)
  and u7644 (n1879, Gqgpw6[11], Xs1iu6);  // ../RTL/cortexm0ds_logic.v(7826)
  not u7645 (Nosiu6, n1879);  // ../RTL/cortexm0ds_logic.v(7826)
  and u7646 (n1880, Trgpw6[11], Dw1iu6);  // ../RTL/cortexm0ds_logic.v(7827)
  not u7647 (Gosiu6, n1880);  // ../RTL/cortexm0ds_logic.v(7827)
  and u7648 (Ensiu6, Uosiu6, Bpsiu6);  // ../RTL/cortexm0ds_logic.v(7828)
  and u7649 (n1881, vis_pc_o[10], Iv1iu6);  // ../RTL/cortexm0ds_logic.v(7829)
  buf u765 (Togpw6[22], Etfbx6);  // ../RTL/cortexm0ds_logic.v(2378)
  not u7650 (Bpsiu6, n1881);  // ../RTL/cortexm0ds_logic.v(7829)
  and u7651 (n1882, Jshpw6[11], Bo1iu6);  // ../RTL/cortexm0ds_logic.v(7830)
  not u7652 (Kjsiu6, n1882);  // ../RTL/cortexm0ds_logic.v(7830)
  and u7653 (n1883, Ipsiu6, Ppsiu6);  // ../RTL/cortexm0ds_logic.v(7831)
  not u7654 (Obphu6, n1883);  // ../RTL/cortexm0ds_logic.v(7831)
  and u7655 (Ppsiu6, Wpsiu6, Po1iu6);  // ../RTL/cortexm0ds_logic.v(7832)
  and u7656 (n1884, Wo1iu6, Dqsiu6);  // ../RTL/cortexm0ds_logic.v(7833)
  not u7657 (Wpsiu6, n1884);  // ../RTL/cortexm0ds_logic.v(7833)
  and u7658 (n1885, Kqsiu6, Rqsiu6);  // ../RTL/cortexm0ds_logic.v(7834)
  not u7659 (Dqsiu6, n1885);  // ../RTL/cortexm0ds_logic.v(7834)
  buf u766 (Togpw6[21], Xdebx6);  // ../RTL/cortexm0ds_logic.v(2378)
  and u7660 (Rqsiu6, Yqsiu6, Frsiu6);  // ../RTL/cortexm0ds_logic.v(7835)
  and u7661 (Frsiu6, Mrsiu6, Trsiu6);  // ../RTL/cortexm0ds_logic.v(7836)
  and u7662 (n1886, Gtgpw6[12], Cs1iu6);  // ../RTL/cortexm0ds_logic.v(7837)
  not u7663 (Trsiu6, n1886);  // ../RTL/cortexm0ds_logic.v(7837)
  and u7664 (Mrsiu6, Assiu6, Hssiu6);  // ../RTL/cortexm0ds_logic.v(7838)
  and u7665 (n1887, Togpw6[12], Vr1iu6);  // ../RTL/cortexm0ds_logic.v(7839)
  not u7666 (Assiu6, n1887);  // ../RTL/cortexm0ds_logic.v(7839)
  and u7667 (Yqsiu6, Ossiu6, Vssiu6);  // ../RTL/cortexm0ds_logic.v(7840)
  and u7668 (n1888, E1hpw6[12], Zt1iu6);  // ../RTL/cortexm0ds_logic.v(7841)
  not u7669 (Vssiu6, n1888);  // ../RTL/cortexm0ds_logic.v(7841)
  buf u767 (vis_psp_o[12], S98ax6);  // ../RTL/cortexm0ds_logic.v(2085)
  and u7670 (Ossiu6, Ctsiu6, Jtsiu6);  // ../RTL/cortexm0ds_logic.v(7842)
  and u7671 (n1889, Ar1iu6, Fkfpw6[12]);  // ../RTL/cortexm0ds_logic.v(7843)
  not u7672 (Jtsiu6, n1889);  // ../RTL/cortexm0ds_logic.v(7843)
  and u7673 (n1890, HRDATA[12], St1iu6);  // ../RTL/cortexm0ds_logic.v(7844)
  not u7674 (Ctsiu6, n1890);  // ../RTL/cortexm0ds_logic.v(7844)
  and u7675 (Kqsiu6, Qtsiu6, Xtsiu6);  // ../RTL/cortexm0ds_logic.v(7845)
  and u7676 (Xtsiu6, Eusiu6, Lusiu6);  // ../RTL/cortexm0ds_logic.v(7846)
  and u7677 (n1891, K7hpw6[12], Kw1iu6);  // ../RTL/cortexm0ds_logic.v(7847)
  not u7678 (Lusiu6, n1891);  // ../RTL/cortexm0ds_logic.v(7847)
  and u7679 (Eusiu6, Susiu6, Zusiu6);  // ../RTL/cortexm0ds_logic.v(7848)
  buf u768 (H8gpw6[0], Wgipw6);  // ../RTL/cortexm0ds_logic.v(1877)
  and u7680 (n1892, Gqgpw6[12], Xs1iu6);  // ../RTL/cortexm0ds_logic.v(7849)
  not u7681 (Zusiu6, n1892);  // ../RTL/cortexm0ds_logic.v(7849)
  and u7682 (n1893, Trgpw6[12], Dw1iu6);  // ../RTL/cortexm0ds_logic.v(7850)
  not u7683 (Susiu6, n1893);  // ../RTL/cortexm0ds_logic.v(7850)
  and u7684 (Qtsiu6, Gvsiu6, Nvsiu6);  // ../RTL/cortexm0ds_logic.v(7851)
  and u7685 (Gvsiu6, Uvsiu6, Bwsiu6);  // ../RTL/cortexm0ds_logic.v(7852)
  and u7686 (n1894, vis_pc_o[11], Iv1iu6);  // ../RTL/cortexm0ds_logic.v(7853)
  not u7687 (Bwsiu6, n1894);  // ../RTL/cortexm0ds_logic.v(7853)
  and u7688 (Ipsiu6, Iwsiu6, Pwsiu6);  // ../RTL/cortexm0ds_logic.v(7854)
  and u7689 (n1895, Jshpw6[12], Bo1iu6);  // ../RTL/cortexm0ds_logic.v(7855)
  buf u769 (vis_psp_o[16], Pcxpw6);  // ../RTL/cortexm0ds_logic.v(2085)
  not u7690 (Pwsiu6, n1895);  // ../RTL/cortexm0ds_logic.v(7855)
  and u7691 (n1896, Uthpw6[12], Sf1iu6);  // ../RTL/cortexm0ds_logic.v(7856)
  not u7692 (Iwsiu6, n1896);  // ../RTL/cortexm0ds_logic.v(7856)
  and u7693 (n1897, Wwsiu6, Dxsiu6);  // ../RTL/cortexm0ds_logic.v(7857)
  not u7694 (Hbphu6, n1897);  // ../RTL/cortexm0ds_logic.v(7857)
  and u7695 (Dxsiu6, Kxsiu6, Po1iu6);  // ../RTL/cortexm0ds_logic.v(7858)
  and u7696 (n1898, Wo1iu6, Rxsiu6);  // ../RTL/cortexm0ds_logic.v(7859)
  not u7697 (Kxsiu6, n1898);  // ../RTL/cortexm0ds_logic.v(7859)
  and u7698 (n1899, Yxsiu6, Fysiu6);  // ../RTL/cortexm0ds_logic.v(7860)
  not u7699 (Rxsiu6, n1899);  // ../RTL/cortexm0ds_logic.v(7860)
  buf u77 (vis_r5_o[18], Paxpw6);  // ../RTL/cortexm0ds_logic.v(1909)
  buf u770 (vis_r12_o[2], Misax6);  // ../RTL/cortexm0ds_logic.v(2599)
  and u7700 (Fysiu6, Mysiu6, Tysiu6);  // ../RTL/cortexm0ds_logic.v(7861)
  and u7701 (Tysiu6, Azsiu6, Hzsiu6);  // ../RTL/cortexm0ds_logic.v(7862)
  and u7702 (n1900, Ar1iu6, Fkfpw6[13]);  // ../RTL/cortexm0ds_logic.v(7863)
  not u7703 (Hzsiu6, n1900);  // ../RTL/cortexm0ds_logic.v(7863)
  and u7704 (Azsiu6, Ozsiu6, Vzsiu6);  // ../RTL/cortexm0ds_logic.v(7864)
  and u7705 (n1901, Togpw6[13], Vr1iu6);  // ../RTL/cortexm0ds_logic.v(7865)
  not u7706 (Vzsiu6, n1901);  // ../RTL/cortexm0ds_logic.v(7865)
  and u7707 (n1902, Gtgpw6[13], Cs1iu6);  // ../RTL/cortexm0ds_logic.v(7866)
  not u7708 (Ozsiu6, n1902);  // ../RTL/cortexm0ds_logic.v(7866)
  and u7709 (Mysiu6, C0tiu6, J0tiu6);  // ../RTL/cortexm0ds_logic.v(7867)
  buf u771 (vis_r12_o[4], Lksax6);  // ../RTL/cortexm0ds_logic.v(2599)
  and u7710 (n1903, Gqgpw6[13], Xs1iu6);  // ../RTL/cortexm0ds_logic.v(7868)
  not u7711 (J0tiu6, n1903);  // ../RTL/cortexm0ds_logic.v(7868)
  and u7712 (C0tiu6, Q0tiu6, X0tiu6);  // ../RTL/cortexm0ds_logic.v(7869)
  and u7713 (n1904, HRDATA[13], St1iu6);  // ../RTL/cortexm0ds_logic.v(7870)
  not u7714 (X0tiu6, n1904);  // ../RTL/cortexm0ds_logic.v(7870)
  and u7715 (n1905, E1hpw6[13], Zt1iu6);  // ../RTL/cortexm0ds_logic.v(7871)
  not u7716 (Q0tiu6, n1905);  // ../RTL/cortexm0ds_logic.v(7871)
  and u7717 (Yxsiu6, E1tiu6, L1tiu6);  // ../RTL/cortexm0ds_logic.v(7872)
  and u7718 (L1tiu6, S1tiu6, Z1tiu6);  // ../RTL/cortexm0ds_logic.v(7873)
  and u7719 (n1906, vis_pc_o[12], Iv1iu6);  // ../RTL/cortexm0ds_logic.v(7874)
  buf u772 (L8ehu6, F26bx6);  // ../RTL/cortexm0ds_logic.v(2835)
  not u7720 (Z1tiu6, n1906);  // ../RTL/cortexm0ds_logic.v(7874)
  and u7721 (S1tiu6, G2tiu6, N2tiu6);  // ../RTL/cortexm0ds_logic.v(7875)
  and u7722 (n1907, Trgpw6[13], Dw1iu6);  // ../RTL/cortexm0ds_logic.v(7876)
  not u7723 (N2tiu6, n1907);  // ../RTL/cortexm0ds_logic.v(7876)
  and u7724 (n1908, K7hpw6[13], Kw1iu6);  // ../RTL/cortexm0ds_logic.v(7877)
  not u7725 (G2tiu6, n1908);  // ../RTL/cortexm0ds_logic.v(7877)
  and u7726 (E1tiu6, U2tiu6, Yw1iu6);  // ../RTL/cortexm0ds_logic.v(7878)
  and u7727 (Wwsiu6, B3tiu6, I3tiu6);  // ../RTL/cortexm0ds_logic.v(7879)
  and u7728 (n1909, Jshpw6[13], Bo1iu6);  // ../RTL/cortexm0ds_logic.v(7880)
  not u7729 (I3tiu6, n1909);  // ../RTL/cortexm0ds_logic.v(7880)
  buf u773 (vis_psp_o[5], A7zpw6);  // ../RTL/cortexm0ds_logic.v(2085)
  and u7730 (n1910, Uthpw6[13], Sf1iu6);  // ../RTL/cortexm0ds_logic.v(7881)
  not u7731 (B3tiu6, n1910);  // ../RTL/cortexm0ds_logic.v(7881)
  and u7732 (n1911, P3tiu6, W3tiu6);  // ../RTL/cortexm0ds_logic.v(7882)
  not u7733 (Abphu6, n1911);  // ../RTL/cortexm0ds_logic.v(7882)
  and u7734 (W3tiu6, D4tiu6, Po1iu6);  // ../RTL/cortexm0ds_logic.v(7883)
  and u7735 (n1912, Wo1iu6, K4tiu6);  // ../RTL/cortexm0ds_logic.v(7884)
  not u7736 (D4tiu6, n1912);  // ../RTL/cortexm0ds_logic.v(7884)
  and u7737 (n1913, R4tiu6, Y4tiu6);  // ../RTL/cortexm0ds_logic.v(7885)
  not u7738 (K4tiu6, n1913);  // ../RTL/cortexm0ds_logic.v(7885)
  and u7739 (Y4tiu6, F5tiu6, M5tiu6);  // ../RTL/cortexm0ds_logic.v(7886)
  buf u774 (vis_r4_o[12], Vbvax6);  // ../RTL/cortexm0ds_logic.v(2626)
  and u7740 (M5tiu6, T5tiu6, A6tiu6);  // ../RTL/cortexm0ds_logic.v(7887)
  and u7741 (n1914, Ar1iu6, Fkfpw6[14]);  // ../RTL/cortexm0ds_logic.v(7888)
  not u7742 (A6tiu6, n1914);  // ../RTL/cortexm0ds_logic.v(7888)
  and u7743 (T5tiu6, H6tiu6, O6tiu6);  // ../RTL/cortexm0ds_logic.v(7889)
  and u7744 (n1915, Togpw6[14], Vr1iu6);  // ../RTL/cortexm0ds_logic.v(7890)
  not u7745 (O6tiu6, n1915);  // ../RTL/cortexm0ds_logic.v(7890)
  and u7746 (n1916, Gtgpw6[14], Cs1iu6);  // ../RTL/cortexm0ds_logic.v(7891)
  not u7747 (H6tiu6, n1916);  // ../RTL/cortexm0ds_logic.v(7891)
  and u7748 (F5tiu6, V6tiu6, C7tiu6);  // ../RTL/cortexm0ds_logic.v(7892)
  and u7749 (n1917, Gqgpw6[14], Xs1iu6);  // ../RTL/cortexm0ds_logic.v(7893)
  buf u775 (vis_r14_o[9], Qxibx6);  // ../RTL/cortexm0ds_logic.v(2497)
  not u7750 (C7tiu6, n1917);  // ../RTL/cortexm0ds_logic.v(7893)
  and u7751 (V6tiu6, J7tiu6, Q7tiu6);  // ../RTL/cortexm0ds_logic.v(7894)
  and u7752 (n1918, HRDATA[14], St1iu6);  // ../RTL/cortexm0ds_logic.v(7895)
  not u7753 (Q7tiu6, n1918);  // ../RTL/cortexm0ds_logic.v(7895)
  and u7754 (n1919, E1hpw6[14], Zt1iu6);  // ../RTL/cortexm0ds_logic.v(7896)
  not u7755 (J7tiu6, n1919);  // ../RTL/cortexm0ds_logic.v(7896)
  and u7756 (R4tiu6, X7tiu6, E8tiu6);  // ../RTL/cortexm0ds_logic.v(7897)
  and u7757 (E8tiu6, L8tiu6, S8tiu6);  // ../RTL/cortexm0ds_logic.v(7898)
  and u7758 (n1920, vis_pc_o[13], Iv1iu6);  // ../RTL/cortexm0ds_logic.v(7899)
  not u7759 (S8tiu6, n1920);  // ../RTL/cortexm0ds_logic.v(7899)
  buf u776 (vis_r8_o[18], O0sax6);  // ../RTL/cortexm0ds_logic.v(2579)
  and u7760 (L8tiu6, Z8tiu6, G9tiu6);  // ../RTL/cortexm0ds_logic.v(7900)
  and u7761 (n1921, Trgpw6[14], Dw1iu6);  // ../RTL/cortexm0ds_logic.v(7901)
  not u7762 (G9tiu6, n1921);  // ../RTL/cortexm0ds_logic.v(7901)
  and u7763 (n1922, K7hpw6[14], Kw1iu6);  // ../RTL/cortexm0ds_logic.v(7902)
  not u7764 (Z8tiu6, n1922);  // ../RTL/cortexm0ds_logic.v(7902)
  and u7765 (X7tiu6, N9tiu6, Uvsiu6);  // ../RTL/cortexm0ds_logic.v(7903)
  and u7766 (P3tiu6, U9tiu6, Batiu6);  // ../RTL/cortexm0ds_logic.v(7904)
  and u7767 (n1923, Jshpw6[14], Bo1iu6);  // ../RTL/cortexm0ds_logic.v(7905)
  not u7768 (Batiu6, n1923);  // ../RTL/cortexm0ds_logic.v(7905)
  and u7769 (n1924, Uthpw6[14], Sf1iu6);  // ../RTL/cortexm0ds_logic.v(7906)
  buf u777 (vis_psp_o[6], O41qw6);  // ../RTL/cortexm0ds_logic.v(2085)
  not u7770 (U9tiu6, n1924);  // ../RTL/cortexm0ds_logic.v(7906)
  and u7771 (n1925, Iatiu6, Patiu6);  // ../RTL/cortexm0ds_logic.v(7907)
  not u7772 (Taphu6, n1925);  // ../RTL/cortexm0ds_logic.v(7907)
  and u7773 (Patiu6, Watiu6, Po1iu6);  // ../RTL/cortexm0ds_logic.v(7908)
  and u7774 (n1926, Wo1iu6, Dbtiu6);  // ../RTL/cortexm0ds_logic.v(7909)
  not u7775 (Watiu6, n1926);  // ../RTL/cortexm0ds_logic.v(7909)
  and u7776 (n1927, Kbtiu6, Rbtiu6);  // ../RTL/cortexm0ds_logic.v(7910)
  not u7777 (Dbtiu6, n1927);  // ../RTL/cortexm0ds_logic.v(7910)
  and u7778 (Rbtiu6, Ybtiu6, Fctiu6);  // ../RTL/cortexm0ds_logic.v(7911)
  and u7779 (Fctiu6, Mctiu6, Tctiu6);  // ../RTL/cortexm0ds_logic.v(7912)
  buf u778 (vis_r1_o[29], Izppw6);  // ../RTL/cortexm0ds_logic.v(1876)
  and u7780 (n1928, Ar1iu6, Fkfpw6[15]);  // ../RTL/cortexm0ds_logic.v(7913)
  not u7781 (Tctiu6, n1928);  // ../RTL/cortexm0ds_logic.v(7913)
  and u7782 (Mctiu6, Adtiu6, Hdtiu6);  // ../RTL/cortexm0ds_logic.v(7914)
  and u7783 (n1929, Togpw6[15], Vr1iu6);  // ../RTL/cortexm0ds_logic.v(7915)
  not u7784 (Hdtiu6, n1929);  // ../RTL/cortexm0ds_logic.v(7915)
  and u7785 (n1930, Gtgpw6[15], Cs1iu6);  // ../RTL/cortexm0ds_logic.v(7916)
  not u7786 (Adtiu6, n1930);  // ../RTL/cortexm0ds_logic.v(7916)
  and u7787 (Ybtiu6, Odtiu6, Vdtiu6);  // ../RTL/cortexm0ds_logic.v(7917)
  and u7788 (n1931, Gqgpw6[15], Xs1iu6);  // ../RTL/cortexm0ds_logic.v(7918)
  not u7789 (Vdtiu6, n1931);  // ../RTL/cortexm0ds_logic.v(7918)
  buf u779 (vis_r0_o[8], Tu0qw6);  // ../RTL/cortexm0ds_logic.v(1875)
  and u7790 (Odtiu6, Cetiu6, Jetiu6);  // ../RTL/cortexm0ds_logic.v(7919)
  and u7791 (n1932, HRDATA[15], St1iu6);  // ../RTL/cortexm0ds_logic.v(7920)
  not u7792 (Jetiu6, n1932);  // ../RTL/cortexm0ds_logic.v(7920)
  and u7793 (n1933, E1hpw6[15], Zt1iu6);  // ../RTL/cortexm0ds_logic.v(7921)
  not u7794 (Cetiu6, n1933);  // ../RTL/cortexm0ds_logic.v(7921)
  and u7795 (Kbtiu6, Qetiu6, Xetiu6);  // ../RTL/cortexm0ds_logic.v(7922)
  and u7796 (Xetiu6, Eftiu6, Lftiu6);  // ../RTL/cortexm0ds_logic.v(7923)
  and u7797 (n1934, vis_pc_o[14], Iv1iu6);  // ../RTL/cortexm0ds_logic.v(7924)
  not u7798 (Lftiu6, n1934);  // ../RTL/cortexm0ds_logic.v(7924)
  and u7799 (Eftiu6, Sftiu6, Zftiu6);  // ../RTL/cortexm0ds_logic.v(7925)
  buf u78 (Ulnhu6, Zslpw6);  // ../RTL/cortexm0ds_logic.v(1844)
  buf u780 (Tzfpw6[15], Nbxax6);  // ../RTL/cortexm0ds_logic.v(2007)
  and u7800 (n1935, Trgpw6[15], Dw1iu6);  // ../RTL/cortexm0ds_logic.v(7926)
  not u7801 (Zftiu6, n1935);  // ../RTL/cortexm0ds_logic.v(7926)
  and u7802 (n1936, K7hpw6[15], Kw1iu6);  // ../RTL/cortexm0ds_logic.v(7927)
  not u7803 (Sftiu6, n1936);  // ../RTL/cortexm0ds_logic.v(7927)
  and u7804 (Qetiu6, Ggtiu6, Uvsiu6);  // ../RTL/cortexm0ds_logic.v(7928)
  and u7805 (Iatiu6, Ngtiu6, Ugtiu6);  // ../RTL/cortexm0ds_logic.v(7929)
  and u7806 (n1937, Jshpw6[15], Bo1iu6);  // ../RTL/cortexm0ds_logic.v(7930)
  not u7807 (Ugtiu6, n1937);  // ../RTL/cortexm0ds_logic.v(7930)
  and u7808 (n1938, Uthpw6[15], Sf1iu6);  // ../RTL/cortexm0ds_logic.v(7931)
  not u7809 (Ngtiu6, n1938);  // ../RTL/cortexm0ds_logic.v(7931)
  buf u781 (Shhpw6[26], A6cbx6);  // ../RTL/cortexm0ds_logic.v(1941)
  and u7810 (n1939, Bhtiu6, Ihtiu6);  // ../RTL/cortexm0ds_logic.v(7932)
  not u7811 (Maphu6, n1939);  // ../RTL/cortexm0ds_logic.v(7932)
  and u7812 (Ihtiu6, Phtiu6, Whtiu6);  // ../RTL/cortexm0ds_logic.v(7933)
  and u7813 (n1940, Wo1iu6, Ditiu6);  // ../RTL/cortexm0ds_logic.v(7934)
  not u7814 (Whtiu6, n1940);  // ../RTL/cortexm0ds_logic.v(7934)
  and u7815 (n1941, Kitiu6, Ritiu6);  // ../RTL/cortexm0ds_logic.v(7935)
  not u7816 (Ditiu6, n1941);  // ../RTL/cortexm0ds_logic.v(7935)
  and u7817 (Ritiu6, Yitiu6, Fjtiu6);  // ../RTL/cortexm0ds_logic.v(7936)
  and u7818 (Fjtiu6, Mjtiu6, Tjtiu6);  // ../RTL/cortexm0ds_logic.v(7937)
  and u7819 (n1942, Ar1iu6, Fkfpw6[16]);  // ../RTL/cortexm0ds_logic.v(7938)
  buf u782 (vis_r12_o[28], Rpibx6);  // ../RTL/cortexm0ds_logic.v(2599)
  not u7820 (Tjtiu6, n1942);  // ../RTL/cortexm0ds_logic.v(7938)
  and u7821 (Mjtiu6, Aktiu6, Hktiu6);  // ../RTL/cortexm0ds_logic.v(7939)
  and u7822 (n1943, Togpw6[16], Vr1iu6);  // ../RTL/cortexm0ds_logic.v(7940)
  not u7823 (Hktiu6, n1943);  // ../RTL/cortexm0ds_logic.v(7940)
  and u7824 (n1944, Gtgpw6[16], Cs1iu6);  // ../RTL/cortexm0ds_logic.v(7941)
  not u7825 (Aktiu6, n1944);  // ../RTL/cortexm0ds_logic.v(7941)
  and u7826 (Yitiu6, Oktiu6, Vktiu6);  // ../RTL/cortexm0ds_logic.v(7942)
  and u7827 (n1945, Gqgpw6[16], Xs1iu6);  // ../RTL/cortexm0ds_logic.v(7943)
  not u7828 (Vktiu6, n1945);  // ../RTL/cortexm0ds_logic.v(7943)
  and u7829 (Oktiu6, Cltiu6, Jltiu6);  // ../RTL/cortexm0ds_logic.v(7944)
  buf u783 (vis_r0_o[12], Ebnpw6);  // ../RTL/cortexm0ds_logic.v(1875)
  and u7830 (n1946, HRDATA[16], St1iu6);  // ../RTL/cortexm0ds_logic.v(7945)
  not u7831 (Jltiu6, n1946);  // ../RTL/cortexm0ds_logic.v(7945)
  and u7832 (n1947, E1hpw6[16], Zt1iu6);  // ../RTL/cortexm0ds_logic.v(7946)
  not u7833 (Cltiu6, n1947);  // ../RTL/cortexm0ds_logic.v(7946)
  and u7834 (Kitiu6, Qltiu6, Xltiu6);  // ../RTL/cortexm0ds_logic.v(7947)
  and u7835 (Xltiu6, Emtiu6, Lmtiu6);  // ../RTL/cortexm0ds_logic.v(7948)
  and u7836 (n1948, vis_pc_o[15], Iv1iu6);  // ../RTL/cortexm0ds_logic.v(7949)
  not u7837 (Lmtiu6, n1948);  // ../RTL/cortexm0ds_logic.v(7949)
  and u7838 (Emtiu6, Smtiu6, Zmtiu6);  // ../RTL/cortexm0ds_logic.v(7950)
  and u7839 (n1949, Trgpw6[16], Dw1iu6);  // ../RTL/cortexm0ds_logic.v(7951)
  buf u784 (Tzfpw6[19], Nr7ax6);  // ../RTL/cortexm0ds_logic.v(2007)
  not u7840 (Zmtiu6, n1949);  // ../RTL/cortexm0ds_logic.v(7951)
  and u7841 (n1950, K7hpw6[16], Kw1iu6);  // ../RTL/cortexm0ds_logic.v(7952)
  not u7842 (Smtiu6, n1950);  // ../RTL/cortexm0ds_logic.v(7952)
  and u7843 (Qltiu6, Gntiu6, Nntiu6);  // ../RTL/cortexm0ds_logic.v(7953)
  and u7844 (n1951, Jshpw6[16], Bo1iu6);  // ../RTL/cortexm0ds_logic.v(7954)
  not u7845 (Phtiu6, n1951);  // ../RTL/cortexm0ds_logic.v(7954)
  and u7846 (Bhtiu6, Untiu6, Botiu6);  // ../RTL/cortexm0ds_logic.v(7955)
  and u7847 (n1952, Uthpw6[16], Sf1iu6);  // ../RTL/cortexm0ds_logic.v(7956)
  not u7848 (Botiu6, n1952);  // ../RTL/cortexm0ds_logic.v(7956)
  and u7849 (n1953, Iotiu6, Potiu6);  // ../RTL/cortexm0ds_logic.v(7957)
  buf u785 (Shhpw6[30], Ra2qw6);  // ../RTL/cortexm0ds_logic.v(1941)
  not u7850 (Faphu6, n1953);  // ../RTL/cortexm0ds_logic.v(7957)
  and u7851 (Potiu6, Wotiu6, Dptiu6);  // ../RTL/cortexm0ds_logic.v(7958)
  and u7852 (n1954, Wo1iu6, Kptiu6);  // ../RTL/cortexm0ds_logic.v(7959)
  not u7853 (Dptiu6, n1954);  // ../RTL/cortexm0ds_logic.v(7959)
  and u7854 (n1955, Rptiu6, Yptiu6);  // ../RTL/cortexm0ds_logic.v(7960)
  not u7855 (Kptiu6, n1955);  // ../RTL/cortexm0ds_logic.v(7960)
  and u7856 (Yptiu6, Fqtiu6, Mqtiu6);  // ../RTL/cortexm0ds_logic.v(7961)
  and u7857 (Mqtiu6, Tqtiu6, Artiu6);  // ../RTL/cortexm0ds_logic.v(7962)
  and u7858 (n1956, Ar1iu6, Fkfpw6[17]);  // ../RTL/cortexm0ds_logic.v(7963)
  not u7859 (Artiu6, n1956);  // ../RTL/cortexm0ds_logic.v(7963)
  buf u786 (Shhpw6[1], M8ipw6);  // ../RTL/cortexm0ds_logic.v(1941)
  and u7860 (Tqtiu6, Hrtiu6, Ortiu6);  // ../RTL/cortexm0ds_logic.v(7964)
  and u7861 (n1957, Togpw6[17], Vr1iu6);  // ../RTL/cortexm0ds_logic.v(7965)
  not u7862 (Ortiu6, n1957);  // ../RTL/cortexm0ds_logic.v(7965)
  and u7863 (n1958, Gtgpw6[17], Cs1iu6);  // ../RTL/cortexm0ds_logic.v(7966)
  not u7864 (Hrtiu6, n1958);  // ../RTL/cortexm0ds_logic.v(7966)
  and u7865 (Fqtiu6, Vrtiu6, Cstiu6);  // ../RTL/cortexm0ds_logic.v(7967)
  and u7866 (n1959, Gqgpw6[17], Xs1iu6);  // ../RTL/cortexm0ds_logic.v(7968)
  not u7867 (Cstiu6, n1959);  // ../RTL/cortexm0ds_logic.v(7968)
  and u7868 (Vrtiu6, Jstiu6, Qstiu6);  // ../RTL/cortexm0ds_logic.v(7969)
  and u7869 (n1960, HRDATA[17], St1iu6);  // ../RTL/cortexm0ds_logic.v(7970)
  buf u787 (vis_r9_o[14], S18ax6);  // ../RTL/cortexm0ds_logic.v(1898)
  not u7870 (Qstiu6, n1960);  // ../RTL/cortexm0ds_logic.v(7970)
  and u7871 (n1961, E1hpw6[17], Zt1iu6);  // ../RTL/cortexm0ds_logic.v(7971)
  not u7872 (Jstiu6, n1961);  // ../RTL/cortexm0ds_logic.v(7971)
  and u7873 (Rptiu6, Xstiu6, Ettiu6);  // ../RTL/cortexm0ds_logic.v(7972)
  and u7874 (Ettiu6, Lttiu6, Sttiu6);  // ../RTL/cortexm0ds_logic.v(7973)
  and u7875 (n1962, vis_pc_o[16], Iv1iu6);  // ../RTL/cortexm0ds_logic.v(7974)
  not u7876 (Sttiu6, n1962);  // ../RTL/cortexm0ds_logic.v(7974)
  and u7877 (Lttiu6, Zttiu6, Gutiu6);  // ../RTL/cortexm0ds_logic.v(7975)
  and u7878 (n1963, Trgpw6[17], Dw1iu6);  // ../RTL/cortexm0ds_logic.v(7976)
  not u7879 (Gutiu6, n1963);  // ../RTL/cortexm0ds_logic.v(7976)
  buf u788 (vis_r3_o[19], D86bx6);  // ../RTL/cortexm0ds_logic.v(2694)
  and u7880 (n1964, K7hpw6[17], Kw1iu6);  // ../RTL/cortexm0ds_logic.v(7977)
  not u7881 (Zttiu6, n1964);  // ../RTL/cortexm0ds_logic.v(7977)
  and u7882 (Xstiu6, Nutiu6, Nntiu6);  // ../RTL/cortexm0ds_logic.v(7978)
  and u7883 (Nntiu6, Reqiu6, Uutiu6);  // ../RTL/cortexm0ds_logic.v(7979)
  and u7884 (n1965, HALTED, Bvtiu6);  // ../RTL/cortexm0ds_logic.v(7980)
  not u7885 (Uutiu6, n1965);  // ../RTL/cortexm0ds_logic.v(7980)
  and u7886 (n1966, Jshpw6[17], Bo1iu6);  // ../RTL/cortexm0ds_logic.v(7981)
  not u7887 (Wotiu6, n1966);  // ../RTL/cortexm0ds_logic.v(7981)
  and u7888 (Iotiu6, Untiu6, Ivtiu6);  // ../RTL/cortexm0ds_logic.v(7982)
  and u7889 (n1967, Uthpw6[17], Sf1iu6);  // ../RTL/cortexm0ds_logic.v(7983)
  buf u789 (vis_msp_o[14], Tg0qw6);  // ../RTL/cortexm0ds_logic.v(2097)
  not u7890 (Ivtiu6, n1967);  // ../RTL/cortexm0ds_logic.v(7983)
  and u7891 (n1968, Pvtiu6, Wvtiu6);  // ../RTL/cortexm0ds_logic.v(7984)
  not u7892 (Y9phu6, n1968);  // ../RTL/cortexm0ds_logic.v(7984)
  and u7893 (Wvtiu6, Dwtiu6, Kwtiu6);  // ../RTL/cortexm0ds_logic.v(7985)
  and u7894 (n1969, Wo1iu6, Rwtiu6);  // ../RTL/cortexm0ds_logic.v(7986)
  not u7895 (Kwtiu6, n1969);  // ../RTL/cortexm0ds_logic.v(7986)
  and u7896 (n1970, Ywtiu6, Fxtiu6);  // ../RTL/cortexm0ds_logic.v(7987)
  not u7897 (Rwtiu6, n1970);  // ../RTL/cortexm0ds_logic.v(7987)
  and u7898 (Fxtiu6, Mxtiu6, Txtiu6);  // ../RTL/cortexm0ds_logic.v(7988)
  and u7899 (Txtiu6, Aytiu6, Hytiu6);  // ../RTL/cortexm0ds_logic.v(7989)
  buf u79 (Pinhu6, Oulpw6);  // ../RTL/cortexm0ds_logic.v(1845)
  buf u790 (vis_r11_o[11], Cg7bx6);  // ../RTL/cortexm0ds_logic.v(1874)
  or u7900 (Hytiu6, Duhiu6, Qa5iu6);  // ../RTL/cortexm0ds_logic.v(7990)
  and u7901 (Aytiu6, Oytiu6, Reqiu6);  // ../RTL/cortexm0ds_logic.v(7991)
  and u7902 (n1971, Togpw6[18], Vr1iu6);  // ../RTL/cortexm0ds_logic.v(7992)
  not u7903 (Oytiu6, n1971);  // ../RTL/cortexm0ds_logic.v(7992)
  and u7904 (Mxtiu6, Vytiu6, Cztiu6);  // ../RTL/cortexm0ds_logic.v(7993)
  and u7905 (n1972, HRDATA[18], St1iu6);  // ../RTL/cortexm0ds_logic.v(7994)
  not u7906 (Cztiu6, n1972);  // ../RTL/cortexm0ds_logic.v(7994)
  and u7907 (Vytiu6, Jztiu6, Qztiu6);  // ../RTL/cortexm0ds_logic.v(7995)
  and u7908 (n1973, Gtgpw6[18], Cs1iu6);  // ../RTL/cortexm0ds_logic.v(7996)
  not u7909 (Qztiu6, n1973);  // ../RTL/cortexm0ds_logic.v(7996)
  buf u791 (Hrfpw6[6], L8kax6);  // ../RTL/cortexm0ds_logic.v(2428)
  and u7910 (n1974, Ar1iu6, Fkfpw6[18]);  // ../RTL/cortexm0ds_logic.v(7997)
  not u7911 (Jztiu6, n1974);  // ../RTL/cortexm0ds_logic.v(7997)
  and u7912 (Ywtiu6, Xztiu6, E0uiu6);  // ../RTL/cortexm0ds_logic.v(7998)
  and u7913 (E0uiu6, L0uiu6, S0uiu6);  // ../RTL/cortexm0ds_logic.v(7999)
  and u7914 (n1975, Trgpw6[18], Dw1iu6);  // ../RTL/cortexm0ds_logic.v(8000)
  not u7915 (S0uiu6, n1975);  // ../RTL/cortexm0ds_logic.v(8000)
  and u7916 (L0uiu6, Z0uiu6, G1uiu6);  // ../RTL/cortexm0ds_logic.v(8001)
  and u7917 (n1976, E1hpw6[18], Zt1iu6);  // ../RTL/cortexm0ds_logic.v(8002)
  not u7918 (G1uiu6, n1976);  // ../RTL/cortexm0ds_logic.v(8002)
  and u7919 (n1977, Gqgpw6[18], Xs1iu6);  // ../RTL/cortexm0ds_logic.v(8003)
  buf u792 (Gqgpw6[6], Dk9bx6);  // ../RTL/cortexm0ds_logic.v(2377)
  not u7920 (Z0uiu6, n1977);  // ../RTL/cortexm0ds_logic.v(8003)
  and u7921 (Xztiu6, N1uiu6, U1uiu6);  // ../RTL/cortexm0ds_logic.v(8004)
  and u7922 (N1uiu6, B2uiu6, I2uiu6);  // ../RTL/cortexm0ds_logic.v(8005)
  and u7923 (n1978, K7hpw6[18], Kw1iu6);  // ../RTL/cortexm0ds_logic.v(8006)
  not u7924 (I2uiu6, n1978);  // ../RTL/cortexm0ds_logic.v(8006)
  and u7925 (n1979, vis_pc_o[17], Iv1iu6);  // ../RTL/cortexm0ds_logic.v(8007)
  not u7926 (B2uiu6, n1979);  // ../RTL/cortexm0ds_logic.v(8007)
  and u7927 (n1980, Jshpw6[18], Bo1iu6);  // ../RTL/cortexm0ds_logic.v(8008)
  not u7928 (Dwtiu6, n1980);  // ../RTL/cortexm0ds_logic.v(8008)
  and u7929 (Pvtiu6, Untiu6, P2uiu6);  // ../RTL/cortexm0ds_logic.v(8009)
  buf u793 (Vbgpw6[12], E90bx6);  // ../RTL/cortexm0ds_logic.v(3092)
  and u7930 (n1981, Uthpw6[18], Sf1iu6);  // ../RTL/cortexm0ds_logic.v(8010)
  not u7931 (P2uiu6, n1981);  // ../RTL/cortexm0ds_logic.v(8010)
  and u7932 (n1982, W2uiu6, D3uiu6);  // ../RTL/cortexm0ds_logic.v(8011)
  not u7933 (R9phu6, n1982);  // ../RTL/cortexm0ds_logic.v(8011)
  and u7934 (D3uiu6, K3uiu6, Po1iu6);  // ../RTL/cortexm0ds_logic.v(8012)
  and u7935 (n1983, Wo1iu6, R3uiu6);  // ../RTL/cortexm0ds_logic.v(8013)
  not u7936 (K3uiu6, n1983);  // ../RTL/cortexm0ds_logic.v(8013)
  and u7937 (n1984, Y3uiu6, F4uiu6);  // ../RTL/cortexm0ds_logic.v(8014)
  not u7938 (R3uiu6, n1984);  // ../RTL/cortexm0ds_logic.v(8014)
  and u7939 (F4uiu6, M4uiu6, T4uiu6);  // ../RTL/cortexm0ds_logic.v(8015)
  buf u794 (vis_r8_o[23], Qirax6);  // ../RTL/cortexm0ds_logic.v(2579)
  and u7940 (T4uiu6, A5uiu6, H5uiu6);  // ../RTL/cortexm0ds_logic.v(8016)
  or u7941 (H5uiu6, Duhiu6, Dp8iu6);  // ../RTL/cortexm0ds_logic.v(8017)
  and u7942 (A5uiu6, O5uiu6, Reqiu6);  // ../RTL/cortexm0ds_logic.v(8018)
  and u7943 (n1985, Togpw6[19], Vr1iu6);  // ../RTL/cortexm0ds_logic.v(8019)
  not u7944 (O5uiu6, n1985);  // ../RTL/cortexm0ds_logic.v(8019)
  and u7945 (M4uiu6, V5uiu6, C6uiu6);  // ../RTL/cortexm0ds_logic.v(8020)
  and u7946 (n1986, HRDATA[19], St1iu6);  // ../RTL/cortexm0ds_logic.v(8021)
  not u7947 (C6uiu6, n1986);  // ../RTL/cortexm0ds_logic.v(8021)
  and u7948 (V5uiu6, J6uiu6, Q6uiu6);  // ../RTL/cortexm0ds_logic.v(8022)
  and u7949 (n1987, Gtgpw6[19], Cs1iu6);  // ../RTL/cortexm0ds_logic.v(8023)
  buf u795 (vis_psp_o[11], Vnkpw6);  // ../RTL/cortexm0ds_logic.v(2085)
  not u7950 (Q6uiu6, n1987);  // ../RTL/cortexm0ds_logic.v(8023)
  and u7951 (n1988, Ar1iu6, Fkfpw6[19]);  // ../RTL/cortexm0ds_logic.v(8024)
  not u7952 (J6uiu6, n1988);  // ../RTL/cortexm0ds_logic.v(8024)
  and u7953 (Y3uiu6, X6uiu6, E7uiu6);  // ../RTL/cortexm0ds_logic.v(8025)
  and u7954 (E7uiu6, L7uiu6, S7uiu6);  // ../RTL/cortexm0ds_logic.v(8026)
  and u7955 (n1989, Trgpw6[19], Dw1iu6);  // ../RTL/cortexm0ds_logic.v(8027)
  not u7956 (S7uiu6, n1989);  // ../RTL/cortexm0ds_logic.v(8027)
  and u7957 (L7uiu6, Z7uiu6, G8uiu6);  // ../RTL/cortexm0ds_logic.v(8028)
  and u7958 (n1990, E1hpw6[19], Zt1iu6);  // ../RTL/cortexm0ds_logic.v(8029)
  not u7959 (G8uiu6, n1990);  // ../RTL/cortexm0ds_logic.v(8029)
  buf u796 (vis_r9_o[19], Jnvpw6);  // ../RTL/cortexm0ds_logic.v(1898)
  and u7960 (n1991, Gqgpw6[19], Xs1iu6);  // ../RTL/cortexm0ds_logic.v(8030)
  not u7961 (Z7uiu6, n1991);  // ../RTL/cortexm0ds_logic.v(8030)
  and u7962 (X6uiu6, N8uiu6, U8uiu6);  // ../RTL/cortexm0ds_logic.v(8031)
  and u7963 (N8uiu6, B9uiu6, I9uiu6);  // ../RTL/cortexm0ds_logic.v(8032)
  and u7964 (n1992, K7hpw6[19], Kw1iu6);  // ../RTL/cortexm0ds_logic.v(8033)
  not u7965 (I9uiu6, n1992);  // ../RTL/cortexm0ds_logic.v(8033)
  and u7966 (n1993, vis_pc_o[18], Iv1iu6);  // ../RTL/cortexm0ds_logic.v(8034)
  not u7967 (B9uiu6, n1993);  // ../RTL/cortexm0ds_logic.v(8034)
  and u7968 (W2uiu6, P9uiu6, W9uiu6);  // ../RTL/cortexm0ds_logic.v(8035)
  and u7969 (n1994, Jshpw6[19], Bo1iu6);  // ../RTL/cortexm0ds_logic.v(8036)
  buf u797 (vis_r3_o[24], Ni5bx6);  // ../RTL/cortexm0ds_logic.v(2694)
  not u7970 (W9uiu6, n1994);  // ../RTL/cortexm0ds_logic.v(8036)
  and u7971 (n1995, Uthpw6[19], Sf1iu6);  // ../RTL/cortexm0ds_logic.v(8037)
  not u7972 (P9uiu6, n1995);  // ../RTL/cortexm0ds_logic.v(8037)
  and u7973 (n1996, Dauiu6, Kauiu6);  // ../RTL/cortexm0ds_logic.v(8038)
  not u7974 (K9phu6, n1996);  // ../RTL/cortexm0ds_logic.v(8038)
  and u7975 (Kauiu6, Rauiu6, V1riu6);  // ../RTL/cortexm0ds_logic.v(8039)
  and u7976 (n1997, Wo1iu6, Yauiu6);  // ../RTL/cortexm0ds_logic.v(8040)
  not u7977 (Rauiu6, n1997);  // ../RTL/cortexm0ds_logic.v(8040)
  and u7978 (n1998, Fbuiu6, Mbuiu6);  // ../RTL/cortexm0ds_logic.v(8041)
  not u7979 (Yauiu6, n1998);  // ../RTL/cortexm0ds_logic.v(8041)
  buf u798 (vis_msp_o[19], T60qw6);  // ../RTL/cortexm0ds_logic.v(2097)
  and u7980 (Mbuiu6, Tbuiu6, Acuiu6);  // ../RTL/cortexm0ds_logic.v(8042)
  and u7981 (Acuiu6, Hcuiu6, Ocuiu6);  // ../RTL/cortexm0ds_logic.v(8043)
  and u7982 (n1999, Ar1iu6, Fkfpw6[20]);  // ../RTL/cortexm0ds_logic.v(8044)
  not u7983 (Ocuiu6, n1999);  // ../RTL/cortexm0ds_logic.v(8044)
  and u7984 (Hcuiu6, Vcuiu6, Cduiu6);  // ../RTL/cortexm0ds_logic.v(8045)
  and u7985 (n2000, Togpw6[20], Vr1iu6);  // ../RTL/cortexm0ds_logic.v(8046)
  not u7986 (Cduiu6, n2000);  // ../RTL/cortexm0ds_logic.v(8046)
  and u7987 (n2001, Gtgpw6[20], Cs1iu6);  // ../RTL/cortexm0ds_logic.v(8047)
  not u7988 (Vcuiu6, n2001);  // ../RTL/cortexm0ds_logic.v(8047)
  and u7989 (Tbuiu6, Jduiu6, Qduiu6);  // ../RTL/cortexm0ds_logic.v(8048)
  buf u799 (vis_r11_o[16], Cbwpw6);  // ../RTL/cortexm0ds_logic.v(1874)
  and u7990 (n2002, Gqgpw6[20], Xs1iu6);  // ../RTL/cortexm0ds_logic.v(8049)
  not u7991 (Qduiu6, n2002);  // ../RTL/cortexm0ds_logic.v(8049)
  and u7992 (Jduiu6, Xduiu6, Eeuiu6);  // ../RTL/cortexm0ds_logic.v(8050)
  and u7993 (n2003, HRDATA[20], St1iu6);  // ../RTL/cortexm0ds_logic.v(8051)
  not u7994 (Eeuiu6, n2003);  // ../RTL/cortexm0ds_logic.v(8051)
  and u7995 (n2004, E1hpw6[20], Zt1iu6);  // ../RTL/cortexm0ds_logic.v(8052)
  not u7996 (Xduiu6, n2004);  // ../RTL/cortexm0ds_logic.v(8052)
  and u7997 (Fbuiu6, Leuiu6, Seuiu6);  // ../RTL/cortexm0ds_logic.v(8053)
  and u7998 (Seuiu6, Zeuiu6, Gfuiu6);  // ../RTL/cortexm0ds_logic.v(8054)
  and u7999 (n2005, vis_pc_o[19], Iv1iu6);  // ../RTL/cortexm0ds_logic.v(8055)
  buf u8 (nTDOEN, 1'b0);  // ../RTL/cortexm0ds_logic.v(1731)
  buf u80 (B7nhu6, Kwlpw6);  // ../RTL/cortexm0ds_logic.v(1846)
  buf u800 (Hrfpw6[11], Smjax6);  // ../RTL/cortexm0ds_logic.v(2428)
  not u8000 (Gfuiu6, n2005);  // ../RTL/cortexm0ds_logic.v(8055)
  and u8001 (Zeuiu6, Nfuiu6, Ufuiu6);  // ../RTL/cortexm0ds_logic.v(8056)
  and u8002 (n2006, Trgpw6[20], Dw1iu6);  // ../RTL/cortexm0ds_logic.v(8057)
  not u8003 (Ufuiu6, n2006);  // ../RTL/cortexm0ds_logic.v(8057)
  and u8004 (n2007, K7hpw6[20], Kw1iu6);  // ../RTL/cortexm0ds_logic.v(8058)
  not u8005 (Nfuiu6, n2007);  // ../RTL/cortexm0ds_logic.v(8058)
  and u8006 (Leuiu6, Bguiu6, Yw1iu6);  // ../RTL/cortexm0ds_logic.v(8059)
  and u8007 (Dauiu6, Iguiu6, Pguiu6);  // ../RTL/cortexm0ds_logic.v(8060)
  and u8008 (n2008, Jshpw6[20], Bo1iu6);  // ../RTL/cortexm0ds_logic.v(8061)
  not u8009 (Pguiu6, n2008);  // ../RTL/cortexm0ds_logic.v(8061)
  buf u801 (Gqgpw6[11], J39bx6);  // ../RTL/cortexm0ds_logic.v(2377)
  and u8010 (n2009, Uthpw6[20], Sf1iu6);  // ../RTL/cortexm0ds_logic.v(8062)
  not u8011 (Iguiu6, n2009);  // ../RTL/cortexm0ds_logic.v(8062)
  and u8012 (n2010, Wguiu6, Dhuiu6);  // ../RTL/cortexm0ds_logic.v(8063)
  not u8013 (D9phu6, n2010);  // ../RTL/cortexm0ds_logic.v(8063)
  and u8014 (Dhuiu6, Khuiu6, V1riu6);  // ../RTL/cortexm0ds_logic.v(8064)
  and u8015 (n2011, Wo1iu6, Rhuiu6);  // ../RTL/cortexm0ds_logic.v(8065)
  not u8016 (Khuiu6, n2011);  // ../RTL/cortexm0ds_logic.v(8065)
  and u8017 (n2012, Yhuiu6, Fiuiu6);  // ../RTL/cortexm0ds_logic.v(8066)
  not u8018 (Rhuiu6, n2012);  // ../RTL/cortexm0ds_logic.v(8066)
  and u8019 (Fiuiu6, Miuiu6, Tiuiu6);  // ../RTL/cortexm0ds_logic.v(8067)
  buf u802 (Vbgpw6[17], Jj0bx6);  // ../RTL/cortexm0ds_logic.v(3092)
  and u8020 (Tiuiu6, Ajuiu6, Hjuiu6);  // ../RTL/cortexm0ds_logic.v(8068)
  and u8021 (n2013, Ar1iu6, Fkfpw6[21]);  // ../RTL/cortexm0ds_logic.v(8069)
  not u8022 (Hjuiu6, n2013);  // ../RTL/cortexm0ds_logic.v(8069)
  and u8023 (Ajuiu6, Ojuiu6, Vjuiu6);  // ../RTL/cortexm0ds_logic.v(8070)
  and u8024 (n2014, Togpw6[21], Vr1iu6);  // ../RTL/cortexm0ds_logic.v(8071)
  not u8025 (Vjuiu6, n2014);  // ../RTL/cortexm0ds_logic.v(8071)
  and u8026 (n2015, Gtgpw6[21], Cs1iu6);  // ../RTL/cortexm0ds_logic.v(8072)
  not u8027 (Ojuiu6, n2015);  // ../RTL/cortexm0ds_logic.v(8072)
  and u8028 (Miuiu6, Ckuiu6, Jkuiu6);  // ../RTL/cortexm0ds_logic.v(8073)
  and u8029 (n2016, Gqgpw6[21], Xs1iu6);  // ../RTL/cortexm0ds_logic.v(8074)
  not u803 (Lodpw6, Jp9bx6);  // ../RTL/cortexm0ds_logic.v(2902)
  not u8030 (Jkuiu6, n2016);  // ../RTL/cortexm0ds_logic.v(8074)
  and u8031 (Ckuiu6, Qkuiu6, Xkuiu6);  // ../RTL/cortexm0ds_logic.v(8075)
  and u8032 (n2017, HRDATA[21], St1iu6);  // ../RTL/cortexm0ds_logic.v(8076)
  not u8033 (Xkuiu6, n2017);  // ../RTL/cortexm0ds_logic.v(8076)
  and u8034 (n2018, E1hpw6[21], Zt1iu6);  // ../RTL/cortexm0ds_logic.v(8077)
  not u8035 (Qkuiu6, n2018);  // ../RTL/cortexm0ds_logic.v(8077)
  and u8036 (Yhuiu6, Eluiu6, Lluiu6);  // ../RTL/cortexm0ds_logic.v(8078)
  and u8037 (Lluiu6, Sluiu6, Zluiu6);  // ../RTL/cortexm0ds_logic.v(8079)
  and u8038 (n2019, vis_pc_o[20], Iv1iu6);  // ../RTL/cortexm0ds_logic.v(8080)
  not u8039 (Zluiu6, n2019);  // ../RTL/cortexm0ds_logic.v(8080)
  buf u804 (Trgpw6[26], Wfcbx6);  // ../RTL/cortexm0ds_logic.v(2376)
  and u8040 (Sluiu6, Gmuiu6, Nmuiu6);  // ../RTL/cortexm0ds_logic.v(8081)
  and u8041 (n2020, Trgpw6[21], Dw1iu6);  // ../RTL/cortexm0ds_logic.v(8082)
  not u8042 (Nmuiu6, n2020);  // ../RTL/cortexm0ds_logic.v(8082)
  and u8043 (n2021, K7hpw6[21], Kw1iu6);  // ../RTL/cortexm0ds_logic.v(8083)
  not u8044 (Gmuiu6, n2021);  // ../RTL/cortexm0ds_logic.v(8083)
  and u8045 (Eluiu6, Umuiu6, Yw1iu6);  // ../RTL/cortexm0ds_logic.v(8084)
  and u8046 (Wguiu6, Bnuiu6, Inuiu6);  // ../RTL/cortexm0ds_logic.v(8085)
  and u8047 (n2022, Jshpw6[21], Bo1iu6);  // ../RTL/cortexm0ds_logic.v(8086)
  not u8048 (Inuiu6, n2022);  // ../RTL/cortexm0ds_logic.v(8086)
  and u8049 (n2023, Uthpw6[21], Sf1iu6);  // ../RTL/cortexm0ds_logic.v(8087)
  not u805 (Tugpw6[3], n1272[3]);  // ../RTL/cortexm0ds_logic.v(16030)
  not u8050 (Bnuiu6, n2023);  // ../RTL/cortexm0ds_logic.v(8087)
  and u8051 (n2024, Pnuiu6, Wnuiu6);  // ../RTL/cortexm0ds_logic.v(8088)
  not u8052 (W8phu6, n2024);  // ../RTL/cortexm0ds_logic.v(8088)
  and u8053 (Wnuiu6, Douiu6, V1riu6);  // ../RTL/cortexm0ds_logic.v(8089)
  and u8054 (n2025, Wo1iu6, Kouiu6);  // ../RTL/cortexm0ds_logic.v(8090)
  not u8055 (Douiu6, n2025);  // ../RTL/cortexm0ds_logic.v(8090)
  and u8056 (n2026, Rouiu6, Youiu6);  // ../RTL/cortexm0ds_logic.v(8091)
  not u8057 (Kouiu6, n2026);  // ../RTL/cortexm0ds_logic.v(8091)
  and u8058 (Youiu6, Fpuiu6, Mpuiu6);  // ../RTL/cortexm0ds_logic.v(8092)
  and u8059 (Mpuiu6, Tpuiu6, Aquiu6);  // ../RTL/cortexm0ds_logic.v(8093)
  buf u806 (Jshpw6[19], Ym3qw6);  // ../RTL/cortexm0ds_logic.v(2372)
  and u8060 (n2027, Ar1iu6, Fkfpw6[22]);  // ../RTL/cortexm0ds_logic.v(8094)
  not u8061 (Aquiu6, n2027);  // ../RTL/cortexm0ds_logic.v(8094)
  and u8062 (Tpuiu6, Hquiu6, Oquiu6);  // ../RTL/cortexm0ds_logic.v(8095)
  and u8063 (n2028, Togpw6[22], Vr1iu6);  // ../RTL/cortexm0ds_logic.v(8096)
  not u8064 (Oquiu6, n2028);  // ../RTL/cortexm0ds_logic.v(8096)
  and u8065 (n2029, Gtgpw6[22], Cs1iu6);  // ../RTL/cortexm0ds_logic.v(8097)
  not u8066 (Hquiu6, n2029);  // ../RTL/cortexm0ds_logic.v(8097)
  and u8067 (Fpuiu6, Vquiu6, Cruiu6);  // ../RTL/cortexm0ds_logic.v(8098)
  and u8068 (n2030, Gqgpw6[22], Xs1iu6);  // ../RTL/cortexm0ds_logic.v(8099)
  not u8069 (Cruiu6, n2030);  // ../RTL/cortexm0ds_logic.v(8099)
  buf u807 (Uthpw6[14], Sd8ax6);  // ../RTL/cortexm0ds_logic.v(1882)
  and u8070 (Vquiu6, Jruiu6, Qruiu6);  // ../RTL/cortexm0ds_logic.v(8100)
  and u8071 (n2031, HRDATA[22], St1iu6);  // ../RTL/cortexm0ds_logic.v(8101)
  not u8072 (Qruiu6, n2031);  // ../RTL/cortexm0ds_logic.v(8101)
  and u8073 (n2032, E1hpw6[22], Zt1iu6);  // ../RTL/cortexm0ds_logic.v(8102)
  not u8074 (Jruiu6, n2032);  // ../RTL/cortexm0ds_logic.v(8102)
  and u8075 (Rouiu6, Xruiu6, Esuiu6);  // ../RTL/cortexm0ds_logic.v(8103)
  and u8076 (Esuiu6, Lsuiu6, Ssuiu6);  // ../RTL/cortexm0ds_logic.v(8104)
  and u8077 (n2033, vis_pc_o[21], Iv1iu6);  // ../RTL/cortexm0ds_logic.v(8105)
  not u8078 (Ssuiu6, n2033);  // ../RTL/cortexm0ds_logic.v(8105)
  and u8079 (Lsuiu6, Zsuiu6, Gtuiu6);  // ../RTL/cortexm0ds_logic.v(8106)
  buf u808 (Uthpw6[28], Idqpw6);  // ../RTL/cortexm0ds_logic.v(1882)
  and u8080 (n2034, Trgpw6[22], Dw1iu6);  // ../RTL/cortexm0ds_logic.v(8107)
  not u8081 (Gtuiu6, n2034);  // ../RTL/cortexm0ds_logic.v(8107)
  and u8082 (n2035, K7hpw6[22], Kw1iu6);  // ../RTL/cortexm0ds_logic.v(8108)
  not u8083 (Zsuiu6, n2035);  // ../RTL/cortexm0ds_logic.v(8108)
  and u8084 (Xruiu6, Ntuiu6, Yw1iu6);  // ../RTL/cortexm0ds_logic.v(8109)
  and u8085 (Pnuiu6, Utuiu6, Buuiu6);  // ../RTL/cortexm0ds_logic.v(8110)
  and u8086 (n2036, Jshpw6[22], Bo1iu6);  // ../RTL/cortexm0ds_logic.v(8111)
  not u8087 (Buuiu6, n2036);  // ../RTL/cortexm0ds_logic.v(8111)
  and u8088 (n2037, Uthpw6[22], Sf1iu6);  // ../RTL/cortexm0ds_logic.v(8112)
  not u8089 (Utuiu6, n2037);  // ../RTL/cortexm0ds_logic.v(8112)
  buf u809 (Togpw6[4], Mbdax6);  // ../RTL/cortexm0ds_logic.v(2378)
  and u8090 (n2038, Iuuiu6, Puuiu6);  // ../RTL/cortexm0ds_logic.v(8113)
  not u8091 (P8phu6, n2038);  // ../RTL/cortexm0ds_logic.v(8113)
  and u8092 (n2039, Uthpw6[23], Sf1iu6);  // ../RTL/cortexm0ds_logic.v(8114)
  not u8093 (Puuiu6, n2039);  // ../RTL/cortexm0ds_logic.v(8114)
  and u8094 (Iuuiu6, Wuuiu6, Dvuiu6);  // ../RTL/cortexm0ds_logic.v(8115)
  and u8095 (n2040, Wo1iu6, Kvuiu6);  // ../RTL/cortexm0ds_logic.v(8116)
  not u8096 (Dvuiu6, n2040);  // ../RTL/cortexm0ds_logic.v(8116)
  and u8097 (n2041, Rvuiu6, Yvuiu6);  // ../RTL/cortexm0ds_logic.v(8117)
  not u8098 (Kvuiu6, n2041);  // ../RTL/cortexm0ds_logic.v(8117)
  and u8099 (Yvuiu6, Fwuiu6, Mwuiu6);  // ../RTL/cortexm0ds_logic.v(8118)
  buf u81 (Ubnhu6, Gylpw6);  // ../RTL/cortexm0ds_logic.v(1847)
  buf u810 (Togpw6[12], F2dax6);  // ../RTL/cortexm0ds_logic.v(2378)
  and u8100 (Mwuiu6, Twuiu6, Axuiu6);  // ../RTL/cortexm0ds_logic.v(8119)
  and u8101 (n2042, Ar1iu6, Fkfpw6[23]);  // ../RTL/cortexm0ds_logic.v(8120)
  not u8102 (Axuiu6, n2042);  // ../RTL/cortexm0ds_logic.v(8120)
  and u8103 (Twuiu6, Hxuiu6, Oxuiu6);  // ../RTL/cortexm0ds_logic.v(8121)
  and u8104 (n2043, Togpw6[23], Vr1iu6);  // ../RTL/cortexm0ds_logic.v(8122)
  not u8105 (Oxuiu6, n2043);  // ../RTL/cortexm0ds_logic.v(8122)
  and u8106 (n2044, Gtgpw6[23], Cs1iu6);  // ../RTL/cortexm0ds_logic.v(8123)
  not u8107 (Hxuiu6, n2044);  // ../RTL/cortexm0ds_logic.v(8123)
  and u8108 (Fwuiu6, Vxuiu6, Cyuiu6);  // ../RTL/cortexm0ds_logic.v(8124)
  and u8109 (n2045, Gqgpw6[23], Xs1iu6);  // ../RTL/cortexm0ds_logic.v(8125)
  buf u811 (Togpw6[20], Qudbx6);  // ../RTL/cortexm0ds_logic.v(2378)
  not u8110 (Cyuiu6, n2045);  // ../RTL/cortexm0ds_logic.v(8125)
  and u8111 (Vxuiu6, Jyuiu6, Qyuiu6);  // ../RTL/cortexm0ds_logic.v(8126)
  and u8112 (n2046, HRDATA[23], St1iu6);  // ../RTL/cortexm0ds_logic.v(8127)
  not u8113 (Qyuiu6, n2046);  // ../RTL/cortexm0ds_logic.v(8127)
  and u8114 (n2047, E1hpw6[23], Zt1iu6);  // ../RTL/cortexm0ds_logic.v(8128)
  not u8115 (Jyuiu6, n2047);  // ../RTL/cortexm0ds_logic.v(8128)
  and u8116 (Rvuiu6, Xyuiu6, Ezuiu6);  // ../RTL/cortexm0ds_logic.v(8129)
  and u8117 (Ezuiu6, Lzuiu6, Szuiu6);  // ../RTL/cortexm0ds_logic.v(8130)
  and u8118 (n2048, vis_pc_o[22], Iv1iu6);  // ../RTL/cortexm0ds_logic.v(8131)
  not u8119 (Szuiu6, n2048);  // ../RTL/cortexm0ds_logic.v(8131)
  buf u812 (Togpw6[28], Yogax6);  // ../RTL/cortexm0ds_logic.v(2378)
  and u8120 (Lzuiu6, Zzuiu6, G0viu6);  // ../RTL/cortexm0ds_logic.v(8132)
  and u8121 (n2049, Trgpw6[23], Dw1iu6);  // ../RTL/cortexm0ds_logic.v(8133)
  not u8122 (G0viu6, n2049);  // ../RTL/cortexm0ds_logic.v(8133)
  and u8123 (n2050, K7hpw6[23], Kw1iu6);  // ../RTL/cortexm0ds_logic.v(8134)
  not u8124 (Zzuiu6, n2050);  // ../RTL/cortexm0ds_logic.v(8134)
  and u8125 (Xyuiu6, N0viu6, Yw1iu6);  // ../RTL/cortexm0ds_logic.v(8135)
  and u8126 (n2051, Jshpw6[23], Bo1iu6);  // ../RTL/cortexm0ds_logic.v(8136)
  not u8127 (Wuuiu6, n2051);  // ../RTL/cortexm0ds_logic.v(8136)
  and u8128 (n2052, U0viu6, B1viu6);  // ../RTL/cortexm0ds_logic.v(8137)
  not u8129 (I8phu6, n2052);  // ../RTL/cortexm0ds_logic.v(8137)
  buf u813 (X8hpw6[6], Sqwpw6);  // ../RTL/cortexm0ds_logic.v(2046)
  and u8130 (B1viu6, I1viu6, Bcriu6);  // ../RTL/cortexm0ds_logic.v(8138)
  and u8131 (n2053, Wo1iu6, P1viu6);  // ../RTL/cortexm0ds_logic.v(8139)
  not u8132 (I1viu6, n2053);  // ../RTL/cortexm0ds_logic.v(8139)
  and u8133 (n2054, W1viu6, D2viu6);  // ../RTL/cortexm0ds_logic.v(8140)
  not u8134 (P1viu6, n2054);  // ../RTL/cortexm0ds_logic.v(8140)
  and u8135 (D2viu6, K2viu6, R2viu6);  // ../RTL/cortexm0ds_logic.v(8141)
  and u8136 (R2viu6, Y2viu6, F3viu6);  // ../RTL/cortexm0ds_logic.v(8142)
  and u8137 (F3viu6, M3viu6, T3viu6);  // ../RTL/cortexm0ds_logic.v(8143)
  and u8138 (n2055, Vxmhu6, Eg7iu6);  // ../RTL/cortexm0ds_logic.v(8144)
  not u8139 (T3viu6, n2055);  // ../RTL/cortexm0ds_logic.v(8144)
  buf u814 (Jshpw6[11], B79bx6);  // ../RTL/cortexm0ds_logic.v(2372)
  and u8140 (n2056, Yc7iu6, E5hhu6);  // ../RTL/cortexm0ds_logic.v(8145)
  not u8141 (M3viu6, n2056);  // ../RTL/cortexm0ds_logic.v(8145)
  and u8142 (Y2viu6, A4viu6, H4viu6);  // ../RTL/cortexm0ds_logic.v(8146)
  and u8143 (n2057, Togpw6[24], Vr1iu6);  // ../RTL/cortexm0ds_logic.v(8147)
  not u8144 (H4viu6, n2057);  // ../RTL/cortexm0ds_logic.v(8147)
  and u8145 (n2058, R6hhu6, Bvtiu6);  // ../RTL/cortexm0ds_logic.v(8148)
  not u8146 (A4viu6, n2058);  // ../RTL/cortexm0ds_logic.v(8148)
  and u8147 (K2viu6, O4viu6, V4viu6);  // ../RTL/cortexm0ds_logic.v(8149)
  and u8148 (V4viu6, C5viu6, J5viu6);  // ../RTL/cortexm0ds_logic.v(8150)
  and u8149 (n2059, Hwmhu6, Ws4iu6);  // ../RTL/cortexm0ds_logic.v(8151)
  buf u815 (vis_r4_o[18], V1vax6);  // ../RTL/cortexm0ds_logic.v(2626)
  not u8150 (J5viu6, n2059);  // ../RTL/cortexm0ds_logic.v(8151)
  and u8151 (n2060, Gtgpw6[24], Cs1iu6);  // ../RTL/cortexm0ds_logic.v(8152)
  not u8152 (C5viu6, n2060);  // ../RTL/cortexm0ds_logic.v(8152)
  and u8153 (O4viu6, Q5viu6, X5viu6);  // ../RTL/cortexm0ds_logic.v(8153)
  and u8154 (n2061, Ar1iu6, Fkfpw6[24]);  // ../RTL/cortexm0ds_logic.v(8154)
  not u8155 (X5viu6, n2061);  // ../RTL/cortexm0ds_logic.v(8154)
  and u8156 (n2062, HRDATA[24], St1iu6);  // ../RTL/cortexm0ds_logic.v(8155)
  not u8157 (Q5viu6, n2062);  // ../RTL/cortexm0ds_logic.v(8155)
  and u8158 (W1viu6, E6viu6, L6viu6);  // ../RTL/cortexm0ds_logic.v(8156)
  and u8159 (L6viu6, S6viu6, Z6viu6);  // ../RTL/cortexm0ds_logic.v(8157)
  buf u816 (vis_r4_o[10], Vdvax6);  // ../RTL/cortexm0ds_logic.v(2626)
  and u8160 (Z6viu6, G7viu6, N7viu6);  // ../RTL/cortexm0ds_logic.v(8158)
  and u8161 (n2063, E1hpw6[24], Zt1iu6);  // ../RTL/cortexm0ds_logic.v(8159)
  not u8162 (N7viu6, n2063);  // ../RTL/cortexm0ds_logic.v(8159)
  and u8163 (n2064, Gqgpw6[24], Xs1iu6);  // ../RTL/cortexm0ds_logic.v(8160)
  not u8164 (G7viu6, n2064);  // ../RTL/cortexm0ds_logic.v(8160)
  and u8165 (S6viu6, U7viu6, B8viu6);  // ../RTL/cortexm0ds_logic.v(8161)
  and u8166 (n2065, Trgpw6[24], Dw1iu6);  // ../RTL/cortexm0ds_logic.v(8162)
  not u8167 (B8viu6, n2065);  // ../RTL/cortexm0ds_logic.v(8162)
  and u8168 (n2066, K7hpw6[24], Kw1iu6);  // ../RTL/cortexm0ds_logic.v(8163)
  not u8169 (U7viu6, n2066);  // ../RTL/cortexm0ds_logic.v(8163)
  buf u817 (vis_r8_o[15], Zz7bx6);  // ../RTL/cortexm0ds_logic.v(2579)
  and u8170 (E6viu6, I8viu6, P8viu6);  // ../RTL/cortexm0ds_logic.v(8164)
  and u8171 (I8viu6, Yw1iu6, W8viu6);  // ../RTL/cortexm0ds_logic.v(8165)
  and u8172 (n2067, vis_pc_o[23], Iv1iu6);  // ../RTL/cortexm0ds_logic.v(8166)
  not u8173 (W8viu6, n2067);  // ../RTL/cortexm0ds_logic.v(8166)
  and u8174 (U0viu6, D9viu6, K9viu6);  // ../RTL/cortexm0ds_logic.v(8167)
  and u8175 (n2068, Jshpw6[24], Bo1iu6);  // ../RTL/cortexm0ds_logic.v(8168)
  not u8176 (K9viu6, n2068);  // ../RTL/cortexm0ds_logic.v(8168)
  and u8177 (n2069, Uthpw6[24], Sf1iu6);  // ../RTL/cortexm0ds_logic.v(8169)
  not u8178 (D9viu6, n2069);  // ../RTL/cortexm0ds_logic.v(8169)
  and u8179 (n2070, R9viu6, Y9viu6);  // ../RTL/cortexm0ds_logic.v(8170)
  buf u818 (vis_r9_o[11], Cc7bx6);  // ../RTL/cortexm0ds_logic.v(1898)
  not u8180 (B8phu6, n2070);  // ../RTL/cortexm0ds_logic.v(8170)
  and u8181 (Y9viu6, Faviu6, Bcriu6);  // ../RTL/cortexm0ds_logic.v(8171)
  and u8182 (n2071, Wo1iu6, Maviu6);  // ../RTL/cortexm0ds_logic.v(8173)
  not u8183 (Faviu6, n2071);  // ../RTL/cortexm0ds_logic.v(8173)
  and u8184 (n2072, Taviu6, Abviu6);  // ../RTL/cortexm0ds_logic.v(8174)
  not u8185 (Maviu6, n2072);  // ../RTL/cortexm0ds_logic.v(8174)
  and u8186 (Abviu6, Hbviu6, Obviu6);  // ../RTL/cortexm0ds_logic.v(8175)
  and u8187 (Obviu6, Vbviu6, Ccviu6);  // ../RTL/cortexm0ds_logic.v(8176)
  and u8188 (n2073, Gtgpw6[25], Cs1iu6);  // ../RTL/cortexm0ds_logic.v(8177)
  not u8189 (Ccviu6, n2073);  // ../RTL/cortexm0ds_logic.v(8177)
  buf u819 (vis_r3_o[16], De6bx6);  // ../RTL/cortexm0ds_logic.v(2694)
  and u8190 (Vbviu6, Jcviu6, Qcviu6);  // ../RTL/cortexm0ds_logic.v(8178)
  and u8191 (n2074, Togpw6[25], Vr1iu6);  // ../RTL/cortexm0ds_logic.v(8179)
  not u8192 (Qcviu6, n2074);  // ../RTL/cortexm0ds_logic.v(8179)
  and u8193 (n2075, D8hhu6, Bvtiu6);  // ../RTL/cortexm0ds_logic.v(8180)
  not u8194 (Jcviu6, n2075);  // ../RTL/cortexm0ds_logic.v(8180)
  and u8195 (Hbviu6, Xcviu6, Edviu6);  // ../RTL/cortexm0ds_logic.v(8181)
  and u8196 (n2076, E1hpw6[25], Zt1iu6);  // ../RTL/cortexm0ds_logic.v(8182)
  not u8197 (Edviu6, n2076);  // ../RTL/cortexm0ds_logic.v(8182)
  and u8198 (Xcviu6, Ldviu6, Sdviu6);  // ../RTL/cortexm0ds_logic.v(8183)
  and u8199 (n2077, Ar1iu6, Fkfpw6[25]);  // ../RTL/cortexm0ds_logic.v(8184)
  buf u82 (vis_r14_o[13], N3oax6);  // ../RTL/cortexm0ds_logic.v(2497)
  buf u820 (vis_msp_o[11], Ti0qw6);  // ../RTL/cortexm0ds_logic.v(2097)
  not u8200 (Sdviu6, n2077);  // ../RTL/cortexm0ds_logic.v(8184)
  and u8201 (n2078, HRDATA[25], St1iu6);  // ../RTL/cortexm0ds_logic.v(8185)
  not u8202 (Ldviu6, n2078);  // ../RTL/cortexm0ds_logic.v(8185)
  and u8203 (Taviu6, Zdviu6, Geviu6);  // ../RTL/cortexm0ds_logic.v(8186)
  and u8204 (Geviu6, Neviu6, Ueviu6);  // ../RTL/cortexm0ds_logic.v(8187)
  and u8205 (n2079, K7hpw6[25], Kw1iu6);  // ../RTL/cortexm0ds_logic.v(8188)
  not u8206 (Ueviu6, n2079);  // ../RTL/cortexm0ds_logic.v(8188)
  and u8207 (Neviu6, Bfviu6, Ifviu6);  // ../RTL/cortexm0ds_logic.v(8189)
  and u8208 (n2080, Gqgpw6[25], Xs1iu6);  // ../RTL/cortexm0ds_logic.v(8190)
  not u8209 (Ifviu6, n2080);  // ../RTL/cortexm0ds_logic.v(8190)
  buf u821 (vis_r11_o[8], Q01qw6);  // ../RTL/cortexm0ds_logic.v(1874)
  and u8210 (n2081, Trgpw6[25], Dw1iu6);  // ../RTL/cortexm0ds_logic.v(8191)
  not u8211 (Bfviu6, n2081);  // ../RTL/cortexm0ds_logic.v(8191)
  and u8212 (Zdviu6, Pfviu6, Wfviu6);  // ../RTL/cortexm0ds_logic.v(8192)
  and u8213 (Pfviu6, Yw1iu6, Dgviu6);  // ../RTL/cortexm0ds_logic.v(8193)
  and u8214 (n2082, vis_pc_o[24], Iv1iu6);  // ../RTL/cortexm0ds_logic.v(8194)
  not u8215 (Dgviu6, n2082);  // ../RTL/cortexm0ds_logic.v(8194)
  and u8216 (R9viu6, Kgviu6, Rgviu6);  // ../RTL/cortexm0ds_logic.v(8195)
  and u8217 (n2083, Jshpw6[25], Bo1iu6);  // ../RTL/cortexm0ds_logic.v(8196)
  not u8218 (Rgviu6, n2083);  // ../RTL/cortexm0ds_logic.v(8196)
  and u8219 (n2084, Uthpw6[25], Sf1iu6);  // ../RTL/cortexm0ds_logic.v(8197)
  buf u822 (Hrfpw6[3], Vqjbx6);  // ../RTL/cortexm0ds_logic.v(2428)
  not u8220 (Kgviu6, n2084);  // ../RTL/cortexm0ds_logic.v(8197)
  and u8221 (n2085, Ygviu6, Fhviu6);  // ../RTL/cortexm0ds_logic.v(8198)
  not u8222 (U7phu6, n2085);  // ../RTL/cortexm0ds_logic.v(8198)
  and u8223 (Fhviu6, Mhviu6, V1riu6);  // ../RTL/cortexm0ds_logic.v(8199)
  and u8224 (n2086, Wo1iu6, Thviu6);  // ../RTL/cortexm0ds_logic.v(8200)
  not u8225 (Mhviu6, n2086);  // ../RTL/cortexm0ds_logic.v(8200)
  and u8226 (n2087, Aiviu6, Hiviu6);  // ../RTL/cortexm0ds_logic.v(8201)
  not u8227 (Thviu6, n2087);  // ../RTL/cortexm0ds_logic.v(8201)
  and u8228 (Hiviu6, Oiviu6, Viviu6);  // ../RTL/cortexm0ds_logic.v(8202)
  and u8229 (Viviu6, Cjviu6, Jjviu6);  // ../RTL/cortexm0ds_logic.v(8203)
  buf u823 (Gqgpw6[3], B9eax6);  // ../RTL/cortexm0ds_logic.v(2377)
  and u8230 (n2088, Ar1iu6, Fkfpw6[26]);  // ../RTL/cortexm0ds_logic.v(8204)
  not u8231 (Jjviu6, n2088);  // ../RTL/cortexm0ds_logic.v(8204)
  and u8232 (Cjviu6, Qjviu6, Xjviu6);  // ../RTL/cortexm0ds_logic.v(8205)
  and u8233 (n2089, Togpw6[26], Vr1iu6);  // ../RTL/cortexm0ds_logic.v(8206)
  not u8234 (Xjviu6, n2089);  // ../RTL/cortexm0ds_logic.v(8206)
  and u8235 (n2090, Gtgpw6[26], Cs1iu6);  // ../RTL/cortexm0ds_logic.v(8207)
  not u8236 (Qjviu6, n2090);  // ../RTL/cortexm0ds_logic.v(8207)
  and u8237 (Oiviu6, Ekviu6, Lkviu6);  // ../RTL/cortexm0ds_logic.v(8208)
  and u8238 (n2091, Gqgpw6[26], Xs1iu6);  // ../RTL/cortexm0ds_logic.v(8209)
  not u8239 (Lkviu6, n2091);  // ../RTL/cortexm0ds_logic.v(8209)
  buf u824 (Vbgpw6[9], Tkjbx6);  // ../RTL/cortexm0ds_logic.v(3092)
  and u8240 (Ekviu6, Skviu6, Zkviu6);  // ../RTL/cortexm0ds_logic.v(8210)
  and u8241 (n2092, HRDATA[26], St1iu6);  // ../RTL/cortexm0ds_logic.v(8211)
  not u8242 (Zkviu6, n2092);  // ../RTL/cortexm0ds_logic.v(8211)
  and u8243 (n2093, E1hpw6[26], Zt1iu6);  // ../RTL/cortexm0ds_logic.v(8212)
  not u8244 (Skviu6, n2093);  // ../RTL/cortexm0ds_logic.v(8212)
  and u8245 (Aiviu6, Glviu6, Nlviu6);  // ../RTL/cortexm0ds_logic.v(8213)
  and u8246 (Nlviu6, Ulviu6, Bmviu6);  // ../RTL/cortexm0ds_logic.v(8214)
  and u8247 (n2094, vis_pc_o[25], Iv1iu6);  // ../RTL/cortexm0ds_logic.v(8215)
  not u8248 (Bmviu6, n2094);  // ../RTL/cortexm0ds_logic.v(8215)
  and u8249 (Ulviu6, Imviu6, Pmviu6);  // ../RTL/cortexm0ds_logic.v(8216)
  buf u825 (vis_r1_o[22], Tpebx6);  // ../RTL/cortexm0ds_logic.v(1876)
  and u8250 (n2095, Trgpw6[26], Dw1iu6);  // ../RTL/cortexm0ds_logic.v(8217)
  not u8251 (Pmviu6, n2095);  // ../RTL/cortexm0ds_logic.v(8217)
  and u8252 (n2096, K7hpw6[26], Kw1iu6);  // ../RTL/cortexm0ds_logic.v(8218)
  not u8253 (Imviu6, n2096);  // ../RTL/cortexm0ds_logic.v(8218)
  and u8254 (Glviu6, Wmviu6, Yw1iu6);  // ../RTL/cortexm0ds_logic.v(8219)
  and u8255 (Ygviu6, Dnviu6, Knviu6);  // ../RTL/cortexm0ds_logic.v(8220)
  and u8256 (n2097, Jshpw6[26], Bo1iu6);  // ../RTL/cortexm0ds_logic.v(8221)
  not u8257 (Knviu6, n2097);  // ../RTL/cortexm0ds_logic.v(8221)
  and u8258 (n2098, Uthpw6[26], Sf1iu6);  // ../RTL/cortexm0ds_logic.v(8222)
  not u8259 (Dnviu6, n2098);  // ../RTL/cortexm0ds_logic.v(8222)
  buf u826 (E1hpw6[6], Pe9bx6);  // ../RTL/cortexm0ds_logic.v(2367)
  and u8260 (n2099, Rnviu6, Ynviu6);  // ../RTL/cortexm0ds_logic.v(8223)
  not u8261 (N7phu6, n2099);  // ../RTL/cortexm0ds_logic.v(8223)
  and u8262 (n2100, Uthpw6[27], Sf1iu6);  // ../RTL/cortexm0ds_logic.v(8224)
  not u8263 (Ynviu6, n2100);  // ../RTL/cortexm0ds_logic.v(8224)
  and u8264 (Rnviu6, Foviu6, Moviu6);  // ../RTL/cortexm0ds_logic.v(8225)
  and u8265 (n2101, Wo1iu6, Toviu6);  // ../RTL/cortexm0ds_logic.v(8226)
  not u8266 (Moviu6, n2101);  // ../RTL/cortexm0ds_logic.v(8226)
  and u8267 (n2102, Apviu6, Hpviu6);  // ../RTL/cortexm0ds_logic.v(8227)
  not u8268 (Toviu6, n2102);  // ../RTL/cortexm0ds_logic.v(8227)
  and u8269 (Hpviu6, Opviu6, Vpviu6);  // ../RTL/cortexm0ds_logic.v(8228)
  not u827 (Tugpw6[7], n1272[7]);  // ../RTL/cortexm0ds_logic.v(16030)
  and u8270 (Vpviu6, Cqviu6, Jqviu6);  // ../RTL/cortexm0ds_logic.v(8229)
  and u8271 (n2103, Ar1iu6, Fkfpw6[27]);  // ../RTL/cortexm0ds_logic.v(8230)
  not u8272 (Jqviu6, n2103);  // ../RTL/cortexm0ds_logic.v(8230)
  and u8273 (Cqviu6, Qqviu6, Xqviu6);  // ../RTL/cortexm0ds_logic.v(8231)
  and u8274 (n2104, Togpw6[27], Vr1iu6);  // ../RTL/cortexm0ds_logic.v(8232)
  not u8275 (Xqviu6, n2104);  // ../RTL/cortexm0ds_logic.v(8232)
  and u8276 (n2105, Gtgpw6[27], Cs1iu6);  // ../RTL/cortexm0ds_logic.v(8233)
  not u8277 (Qqviu6, n2105);  // ../RTL/cortexm0ds_logic.v(8233)
  and u8278 (Opviu6, Erviu6, Lrviu6);  // ../RTL/cortexm0ds_logic.v(8234)
  and u8279 (n2106, Gqgpw6[27], Xs1iu6);  // ../RTL/cortexm0ds_logic.v(8235)
  not u828 (Eodpw6, L3bbx6);  // ../RTL/cortexm0ds_logic.v(2927)
  not u8280 (Lrviu6, n2106);  // ../RTL/cortexm0ds_logic.v(8235)
  and u8281 (Erviu6, Srviu6, Zrviu6);  // ../RTL/cortexm0ds_logic.v(8236)
  and u8282 (n2107, HRDATA[27], St1iu6);  // ../RTL/cortexm0ds_logic.v(8237)
  not u8283 (Zrviu6, n2107);  // ../RTL/cortexm0ds_logic.v(8237)
  and u8284 (n2108, E1hpw6[27], Zt1iu6);  // ../RTL/cortexm0ds_logic.v(8238)
  not u8285 (Srviu6, n2108);  // ../RTL/cortexm0ds_logic.v(8238)
  and u8286 (Apviu6, Gsviu6, Nsviu6);  // ../RTL/cortexm0ds_logic.v(8239)
  and u8287 (Nsviu6, Usviu6, Btviu6);  // ../RTL/cortexm0ds_logic.v(8240)
  and u8288 (n2109, vis_pc_o[26], Iv1iu6);  // ../RTL/cortexm0ds_logic.v(8241)
  not u8289 (Btviu6, n2109);  // ../RTL/cortexm0ds_logic.v(8241)
  buf u829 (Gtgpw6[4], Tfcax6);  // ../RTL/cortexm0ds_logic.v(2375)
  and u8290 (Usviu6, Itviu6, Ptviu6);  // ../RTL/cortexm0ds_logic.v(8242)
  and u8291 (n2110, Trgpw6[27], Dw1iu6);  // ../RTL/cortexm0ds_logic.v(8243)
  not u8292 (Ptviu6, n2110);  // ../RTL/cortexm0ds_logic.v(8243)
  and u8293 (n2111, K7hpw6[27], Kw1iu6);  // ../RTL/cortexm0ds_logic.v(8244)
  not u8294 (Itviu6, n2111);  // ../RTL/cortexm0ds_logic.v(8244)
  and u8295 (Gsviu6, Wtviu6, Yw1iu6);  // ../RTL/cortexm0ds_logic.v(8245)
  and u8296 (n2112, Jshpw6[27], Bo1iu6);  // ../RTL/cortexm0ds_logic.v(8246)
  not u8297 (Foviu6, n2112);  // ../RTL/cortexm0ds_logic.v(8246)
  and u8298 (n2113, Duviu6, Kuviu6);  // ../RTL/cortexm0ds_logic.v(8247)
  not u8299 (G7phu6, n2113);  // ../RTL/cortexm0ds_logic.v(8247)
  buf u83 (vis_r8_o[22], Tvebx6);  // ../RTL/cortexm0ds_logic.v(2579)
  buf u830 (vis_r12_o[3], Jusax6);  // ../RTL/cortexm0ds_logic.v(2599)
  and u8300 (Kuviu6, Ruviu6, Yuviu6);  // ../RTL/cortexm0ds_logic.v(8248)
  and u8301 (n2114, Wo1iu6, Fvviu6);  // ../RTL/cortexm0ds_logic.v(8249)
  not u8302 (Yuviu6, n2114);  // ../RTL/cortexm0ds_logic.v(8249)
  and u8303 (n2115, Mvviu6, Tvviu6);  // ../RTL/cortexm0ds_logic.v(8250)
  not u8304 (Fvviu6, n2115);  // ../RTL/cortexm0ds_logic.v(8250)
  and u8305 (Tvviu6, Awviu6, Hwviu6);  // ../RTL/cortexm0ds_logic.v(8251)
  and u8306 (Hwviu6, Owviu6, Vwviu6);  // ../RTL/cortexm0ds_logic.v(8252)
  and u8307 (n2116, Ar1iu6, Fkfpw6[28]);  // ../RTL/cortexm0ds_logic.v(8253)
  not u8308 (Vwviu6, n2116);  // ../RTL/cortexm0ds_logic.v(8253)
  and u8309 (Owviu6, Cxviu6, Jxviu6);  // ../RTL/cortexm0ds_logic.v(8254)
  buf u831 (vis_r4_o[22], T3fbx6);  // ../RTL/cortexm0ds_logic.v(2626)
  and u8310 (n2117, Togpw6[28], Vr1iu6);  // ../RTL/cortexm0ds_logic.v(8255)
  not u8311 (Jxviu6, n2117);  // ../RTL/cortexm0ds_logic.v(8255)
  and u8312 (n2118, Gtgpw6[28], Cs1iu6);  // ../RTL/cortexm0ds_logic.v(8256)
  not u8313 (Cxviu6, n2118);  // ../RTL/cortexm0ds_logic.v(8256)
  and u8314 (Awviu6, Qxviu6, Xxviu6);  // ../RTL/cortexm0ds_logic.v(8257)
  and u8315 (n2119, Gqgpw6[28], Xs1iu6);  // ../RTL/cortexm0ds_logic.v(8258)
  not u8316 (Xxviu6, n2119);  // ../RTL/cortexm0ds_logic.v(8258)
  and u8317 (Qxviu6, Eyviu6, Lyviu6);  // ../RTL/cortexm0ds_logic.v(8259)
  and u8318 (n2120, HRDATA[28], St1iu6);  // ../RTL/cortexm0ds_logic.v(8260)
  not u8319 (Lyviu6, n2120);  // ../RTL/cortexm0ds_logic.v(8260)
  buf u832 (Mdhpw6[3], Rilpw6);  // ../RTL/cortexm0ds_logic.v(1838)
  and u8320 (n2121, E1hpw6[28], Zt1iu6);  // ../RTL/cortexm0ds_logic.v(8261)
  not u8321 (Eyviu6, n2121);  // ../RTL/cortexm0ds_logic.v(8261)
  and u8322 (Mvviu6, Syviu6, Zyviu6);  // ../RTL/cortexm0ds_logic.v(8262)
  and u8323 (Zyviu6, Gzviu6, Nzviu6);  // ../RTL/cortexm0ds_logic.v(8263)
  and u8324 (n2122, Iv1iu6, vis_pc_o[27]);  // ../RTL/cortexm0ds_logic.v(8264)
  not u8325 (Nzviu6, n2122);  // ../RTL/cortexm0ds_logic.v(8264)
  and u8326 (Gzviu6, Uzviu6, B0wiu6);  // ../RTL/cortexm0ds_logic.v(8265)
  and u8327 (n2123, Trgpw6[28], Dw1iu6);  // ../RTL/cortexm0ds_logic.v(8266)
  not u8328 (B0wiu6, n2123);  // ../RTL/cortexm0ds_logic.v(8266)
  and u8329 (n2124, K7hpw6[28], Kw1iu6);  // ../RTL/cortexm0ds_logic.v(8267)
  buf u833 (vis_r4_o[6], Yfuax6);  // ../RTL/cortexm0ds_logic.v(2626)
  not u8330 (Uzviu6, n2124);  // ../RTL/cortexm0ds_logic.v(8267)
  and u8331 (Syviu6, I0wiu6, Yw1iu6);  // ../RTL/cortexm0ds_logic.v(8268)
  and u8332 (n2125, Jshpw6[28], Bo1iu6);  // ../RTL/cortexm0ds_logic.v(8269)
  not u8333 (Ruviu6, n2125);  // ../RTL/cortexm0ds_logic.v(8269)
  and u8334 (Duviu6, P0wiu6, W0wiu6);  // ../RTL/cortexm0ds_logic.v(8270)
  and u8335 (n2126, ECOREVNUM[20], Tx1iu6);  // ../RTL/cortexm0ds_logic.v(8271)
  not u8336 (W0wiu6, n2126);  // ../RTL/cortexm0ds_logic.v(8271)
  and u8337 (n2127, Uthpw6[28], Sf1iu6);  // ../RTL/cortexm0ds_logic.v(8272)
  not u8338 (P0wiu6, n2127);  // ../RTL/cortexm0ds_logic.v(8272)
  and u8339 (n2128, D1wiu6, K1wiu6);  // ../RTL/cortexm0ds_logic.v(8273)
  buf u834 (vis_r14_o[3], R7nax6);  // ../RTL/cortexm0ds_logic.v(2497)
  not u8340 (Z6phu6, n2128);  // ../RTL/cortexm0ds_logic.v(8273)
  and u8341 (K1wiu6, R1wiu6, Y1wiu6);  // ../RTL/cortexm0ds_logic.v(8274)
  and u8342 (n2129, Jshpw6[29], Bo1iu6);  // ../RTL/cortexm0ds_logic.v(8275)
  not u8343 (Y1wiu6, n2129);  // ../RTL/cortexm0ds_logic.v(8275)
  and u8344 (R1wiu6, F2wiu6, Po1iu6);  // ../RTL/cortexm0ds_logic.v(8276)
  and u8345 (n2130, Wo1iu6, M2wiu6);  // ../RTL/cortexm0ds_logic.v(8277)
  not u8346 (F2wiu6, n2130);  // ../RTL/cortexm0ds_logic.v(8277)
  and u8347 (n2131, T2wiu6, A3wiu6);  // ../RTL/cortexm0ds_logic.v(8278)
  not u8348 (M2wiu6, n2131);  // ../RTL/cortexm0ds_logic.v(8278)
  and u8349 (A3wiu6, H3wiu6, O3wiu6);  // ../RTL/cortexm0ds_logic.v(8279)
  buf u835 (vis_r8_o[12], Oasax6);  // ../RTL/cortexm0ds_logic.v(2579)
  and u8350 (O3wiu6, V3wiu6, C4wiu6);  // ../RTL/cortexm0ds_logic.v(8280)
  and u8351 (n2132, J4wiu6, C3qiu6);  // ../RTL/cortexm0ds_logic.v(8281)
  not u8352 (C4wiu6, n2132);  // ../RTL/cortexm0ds_logic.v(8281)
  and u8353 (J4wiu6, Q4wiu6, X4wiu6);  // ../RTL/cortexm0ds_logic.v(8282)
  and u8354 (n2133, Ar1iu6, Fkfpw6[29]);  // ../RTL/cortexm0ds_logic.v(8283)
  not u8355 (V3wiu6, n2133);  // ../RTL/cortexm0ds_logic.v(8283)
  and u8356 (H3wiu6, E5wiu6, L5wiu6);  // ../RTL/cortexm0ds_logic.v(8284)
  and u8357 (n2134, HRDATA[29], St1iu6);  // ../RTL/cortexm0ds_logic.v(8285)
  not u8358 (L5wiu6, n2134);  // ../RTL/cortexm0ds_logic.v(8285)
  and u8359 (n2135, E1hpw6[29], Zt1iu6);  // ../RTL/cortexm0ds_logic.v(8286)
  buf u836 (vis_r9_o[8], Ry0qw6);  // ../RTL/cortexm0ds_logic.v(1898)
  not u8360 (E5wiu6, n2135);  // ../RTL/cortexm0ds_logic.v(8286)
  and u8361 (T2wiu6, S5wiu6, Z5wiu6);  // ../RTL/cortexm0ds_logic.v(8287)
  and u8362 (Z5wiu6, G6wiu6, N6wiu6);  // ../RTL/cortexm0ds_logic.v(8288)
  and u8363 (n2136, K7hpw6[29], Kw1iu6);  // ../RTL/cortexm0ds_logic.v(8289)
  not u8364 (N6wiu6, n2136);  // ../RTL/cortexm0ds_logic.v(8289)
  and u8365 (n2137, Iv1iu6, vis_pc_o[28]);  // ../RTL/cortexm0ds_logic.v(8290)
  not u8366 (G6wiu6, n2137);  // ../RTL/cortexm0ds_logic.v(8290)
  and u8367 (S5wiu6, U6wiu6, Yw1iu6);  // ../RTL/cortexm0ds_logic.v(8291)
  and u8368 (D1wiu6, B7wiu6, I7wiu6);  // ../RTL/cortexm0ds_logic.v(8292)
  and u8369 (n2138, ECOREVNUM[21], Tx1iu6);  // ../RTL/cortexm0ds_logic.v(8293)
  buf u837 (vis_r3_o[13], Di6bx6);  // ../RTL/cortexm0ds_logic.v(2694)
  not u8370 (I7wiu6, n2138);  // ../RTL/cortexm0ds_logic.v(8293)
  and u8371 (n2139, Uthpw6[29], Sf1iu6);  // ../RTL/cortexm0ds_logic.v(8294)
  not u8372 (B7wiu6, n2139);  // ../RTL/cortexm0ds_logic.v(8294)
  and u8373 (n2140, P7wiu6, W7wiu6);  // ../RTL/cortexm0ds_logic.v(8295)
  not u8374 (S6phu6, n2140);  // ../RTL/cortexm0ds_logic.v(8295)
  and u8375 (W7wiu6, D8wiu6, K8wiu6);  // ../RTL/cortexm0ds_logic.v(8296)
  and u8376 (n2141, Jshpw6[30], Bo1iu6);  // ../RTL/cortexm0ds_logic.v(8297)
  not u8377 (K8wiu6, n2141);  // ../RTL/cortexm0ds_logic.v(8297)
  and u8378 (D8wiu6, R8wiu6, Po1iu6);  // ../RTL/cortexm0ds_logic.v(8298)
  and u8379 (n2142, Wo1iu6, Y8wiu6);  // ../RTL/cortexm0ds_logic.v(8299)
  buf u838 (vis_msp_o[8], Tm0qw6);  // ../RTL/cortexm0ds_logic.v(2097)
  not u8380 (R8wiu6, n2142);  // ../RTL/cortexm0ds_logic.v(8299)
  and u8381 (n2143, F9wiu6, M9wiu6);  // ../RTL/cortexm0ds_logic.v(8300)
  not u8382 (Y8wiu6, n2143);  // ../RTL/cortexm0ds_logic.v(8300)
  and u8383 (M9wiu6, T9wiu6, Aawiu6);  // ../RTL/cortexm0ds_logic.v(8301)
  and u8384 (Aawiu6, Hawiu6, Oawiu6);  // ../RTL/cortexm0ds_logic.v(8302)
  and u8385 (n2144, Ar1iu6, Fkfpw6[30]);  // ../RTL/cortexm0ds_logic.v(8303)
  not u8386 (Oawiu6, n2144);  // ../RTL/cortexm0ds_logic.v(8303)
  and u8387 (Hawiu6, Vawiu6, Cbwiu6);  // ../RTL/cortexm0ds_logic.v(8304)
  and u8388 (n2145, Ligpw6[27], Vr1iu6);  // ../RTL/cortexm0ds_logic.v(8305)
  not u8389 (Cbwiu6, n2145);  // ../RTL/cortexm0ds_logic.v(8305)
  buf u839 (vis_r11_o[5], T3kpw6);  // ../RTL/cortexm0ds_logic.v(1874)
  and u8390 (n2146, Engpw6[27], Cs1iu6);  // ../RTL/cortexm0ds_logic.v(8306)
  not u8391 (Vawiu6, n2146);  // ../RTL/cortexm0ds_logic.v(8306)
  and u8392 (T9wiu6, Jbwiu6, Qbwiu6);  // ../RTL/cortexm0ds_logic.v(8307)
  and u8393 (n2147, Akgpw6[27], Xs1iu6);  // ../RTL/cortexm0ds_logic.v(8308)
  not u8394 (Qbwiu6, n2147);  // ../RTL/cortexm0ds_logic.v(8308)
  and u8395 (Jbwiu6, Xbwiu6, Ecwiu6);  // ../RTL/cortexm0ds_logic.v(8309)
  and u8396 (n2148, HRDATA[30], St1iu6);  // ../RTL/cortexm0ds_logic.v(8310)
  not u8397 (Ecwiu6, n2148);  // ../RTL/cortexm0ds_logic.v(8310)
  and u8398 (n2149, E1hpw6[30], Zt1iu6);  // ../RTL/cortexm0ds_logic.v(8311)
  not u8399 (Xbwiu6, n2149);  // ../RTL/cortexm0ds_logic.v(8311)
  buf u84 (Jshpw6[10], H4ypw6);  // ../RTL/cortexm0ds_logic.v(2372)
  buf u840 (vis_r11_o[31], Efnpw6);  // ../RTL/cortexm0ds_logic.v(1874)
  and u8400 (F9wiu6, Lcwiu6, Scwiu6);  // ../RTL/cortexm0ds_logic.v(8312)
  and u8401 (Scwiu6, Zcwiu6, Gdwiu6);  // ../RTL/cortexm0ds_logic.v(8313)
  and u8402 (n2150, Iv1iu6, vis_pc_o[29]);  // ../RTL/cortexm0ds_logic.v(8314)
  not u8403 (Gdwiu6, n2150);  // ../RTL/cortexm0ds_logic.v(8314)
  and u8404 (Zcwiu6, Ndwiu6, Udwiu6);  // ../RTL/cortexm0ds_logic.v(8315)
  and u8405 (n2151, Plgpw6[27], Dw1iu6);  // ../RTL/cortexm0ds_logic.v(8316)
  not u8406 (Udwiu6, n2151);  // ../RTL/cortexm0ds_logic.v(8316)
  and u8407 (n2152, K7hpw6[30], Kw1iu6);  // ../RTL/cortexm0ds_logic.v(8317)
  not u8408 (Ndwiu6, n2152);  // ../RTL/cortexm0ds_logic.v(8317)
  and u8409 (Lcwiu6, Bewiu6, Yw1iu6);  // ../RTL/cortexm0ds_logic.v(8318)
  buf u841 (Sufpw6[1], J0iax6);  // ../RTL/cortexm0ds_logic.v(2404)
  and u8410 (P7wiu6, Iewiu6, Pewiu6);  // ../RTL/cortexm0ds_logic.v(8319)
  and u8411 (n2153, ECOREVNUM[22], Tx1iu6);  // ../RTL/cortexm0ds_logic.v(8320)
  not u8412 (Pewiu6, n2153);  // ../RTL/cortexm0ds_logic.v(8320)
  and u8413 (n2154, Uthpw6[30], Sf1iu6);  // ../RTL/cortexm0ds_logic.v(8321)
  not u8414 (Iewiu6, n2154);  // ../RTL/cortexm0ds_logic.v(8321)
  and u8415 (n2155, Wewiu6, Dfwiu6);  // ../RTL/cortexm0ds_logic.v(8322)
  not u8416 (L6phu6, n2155);  // ../RTL/cortexm0ds_logic.v(8322)
  and u8417 (Dfwiu6, Kfwiu6, Rfwiu6);  // ../RTL/cortexm0ds_logic.v(8323)
  and u8418 (n2156, Qwpiu6, Aphpw6[1]);  // ../RTL/cortexm0ds_logic.v(8324)
  not u8419 (Rfwiu6, n2156);  // ../RTL/cortexm0ds_logic.v(8324)
  buf u842 (Vbgpw6[6], Nt9bx6);  // ../RTL/cortexm0ds_logic.v(3092)
  or u8420 (Bcriu6, Yfwiu6, Vo4iu6);  // ../RTL/cortexm0ds_logic.v(8325)
  not u8421 (Qwpiu6, Bcriu6);  // ../RTL/cortexm0ds_logic.v(8325)
  and u8422 (Kfwiu6, Fgwiu6, Mgwiu6);  // ../RTL/cortexm0ds_logic.v(8326)
  and u8423 (n2157, Tnhpw6[0], Bo1iu6);  // ../RTL/cortexm0ds_logic.v(8327)
  not u8424 (Mgwiu6, n2157);  // ../RTL/cortexm0ds_logic.v(8327)
  and u8425 (Bo1iu6, Tgwiu6, Vo4iu6);  // ../RTL/cortexm0ds_logic.v(8328)
  and u8426 (Tgwiu6, Ahwiu6, Hhwiu6);  // ../RTL/cortexm0ds_logic.v(8330)
  not u8427 (Yfwiu6, Tgwiu6);  // ../RTL/cortexm0ds_logic.v(8330)
  or u8428 (n2158, Wu9iu6, Ho4iu6);  // ../RTL/cortexm0ds_logic.v(8331)
  not u8429 (Hhwiu6, n2158);  // ../RTL/cortexm0ds_logic.v(8331)
  buf u843 (Aygpw6[1], Hdbax6);  // ../RTL/cortexm0ds_logic.v(2278)
  or u8430 (n2159, Ohwiu6, Sf1iu6);  // ../RTL/cortexm0ds_logic.v(8332)
  not u8431 (Ahwiu6, n2159);  // ../RTL/cortexm0ds_logic.v(8332)
  and u8432 (n2160, Wo1iu6, Vhwiu6);  // ../RTL/cortexm0ds_logic.v(8333)
  not u8433 (Fgwiu6, n2160);  // ../RTL/cortexm0ds_logic.v(8333)
  and u8434 (n2161, Ciwiu6, Jiwiu6);  // ../RTL/cortexm0ds_logic.v(8334)
  not u8435 (Vhwiu6, n2161);  // ../RTL/cortexm0ds_logic.v(8334)
  and u8436 (Jiwiu6, Qiwiu6, Xiwiu6);  // ../RTL/cortexm0ds_logic.v(8335)
  and u8437 (Xiwiu6, Ejwiu6, Ljwiu6);  // ../RTL/cortexm0ds_logic.v(8336)
  and u8438 (Ljwiu6, Sjwiu6, Zjwiu6);  // ../RTL/cortexm0ds_logic.v(8337)
  and u8439 (n2162, Gkwiu6, A2qiu6);  // ../RTL/cortexm0ds_logic.v(8338)
  buf u844 (K7hpw6[30], J59ax6);  // ../RTL/cortexm0ds_logic.v(2366)
  not u8440 (Zjwiu6, n2162);  // ../RTL/cortexm0ds_logic.v(8338)
  and u8441 (Gkwiu6, Nkwiu6, Ukwiu6);  // ../RTL/cortexm0ds_logic.v(8339)
  or u8442 (n2163, Q3qiu6, U4riu6);  // ../RTL/cortexm0ds_logic.v(8340)
  not u8443 (Sjwiu6, n2163);  // ../RTL/cortexm0ds_logic.v(8340)
  and u8444 (U4riu6, Ffqiu6, C3qiu6);  // ../RTL/cortexm0ds_logic.v(8341)
  and u8445 (Q3qiu6, Blwiu6, X8hpw6[1]);  // ../RTL/cortexm0ds_logic.v(8342)
  and u8446 (Blwiu6, Nkwiu6, Ilwiu6);  // ../RTL/cortexm0ds_logic.v(8343)
  and u8447 (Ejwiu6, Plwiu6, Wlwiu6);  // ../RTL/cortexm0ds_logic.v(8344)
  and u8448 (n2164, G4hpw6[0], Sg7iu6);  // ../RTL/cortexm0ds_logic.v(8345)
  not u8449 (Wlwiu6, n2164);  // ../RTL/cortexm0ds_logic.v(8345)
  buf u845 (R4gpw6[63], Cy4bx6);  // ../RTL/cortexm0ds_logic.v(2815)
  and u8450 (Sg7iu6, Dmwiu6, Q4wiu6);  // ../RTL/cortexm0ds_logic.v(8346)
  and u8451 (Plwiu6, Kmwiu6, Rmwiu6);  // ../RTL/cortexm0ds_logic.v(8347)
  and u8452 (n2165, R2hpw6[0], Eg7iu6);  // ../RTL/cortexm0ds_logic.v(8348)
  not u8453 (Rmwiu6, n2165);  // ../RTL/cortexm0ds_logic.v(8348)
  and u8454 (Eg7iu6, Vuciu6, Nkwiu6);  // ../RTL/cortexm0ds_logic.v(8349)
  and u8455 (n2166, Dhgpw6[0], Fgpiu6);  // ../RTL/cortexm0ds_logic.v(8350)
  not u8456 (Kmwiu6, n2166);  // ../RTL/cortexm0ds_logic.v(8350)
  and u8457 (Fgpiu6, Ymwiu6, Fnwiu6);  // ../RTL/cortexm0ds_logic.v(8351)
  and u8458 (Ymwiu6, Mnwiu6, Ilwiu6);  // ../RTL/cortexm0ds_logic.v(8352)
  and u8459 (Qiwiu6, Tnwiu6, Aowiu6);  // ../RTL/cortexm0ds_logic.v(8353)
  buf u846 (vis_r5_o[24], Yvspw6);  // ../RTL/cortexm0ds_logic.v(1909)
  and u8460 (Aowiu6, Howiu6, Oowiu6);  // ../RTL/cortexm0ds_logic.v(8354)
  and u8461 (n2167, Kohhu6, Ve7iu6);  // ../RTL/cortexm0ds_logic.v(8355)
  not u8462 (Oowiu6, n2167);  // ../RTL/cortexm0ds_logic.v(8355)
  and u8463 (Ve7iu6, Vowiu6, Cpwiu6);  // ../RTL/cortexm0ds_logic.v(8356)
  and u8464 (Howiu6, Jpwiu6, Qpwiu6);  // ../RTL/cortexm0ds_logic.v(8357)
  and u8465 (n2168, Yc7iu6, H2hhu6);  // ../RTL/cortexm0ds_logic.v(8358)
  not u8466 (Qpwiu6, n2168);  // ../RTL/cortexm0ds_logic.v(8358)
  and u8467 (Yc7iu6, Xpwiu6, Dzqiu6);  // ../RTL/cortexm0ds_logic.v(8359)
  and u8468 (Xpwiu6, Q4wiu6, Cvciu6);  // ../RTL/cortexm0ds_logic.v(8360)
  and u8469 (n2169, Aygpw6[0], Jf7iu6);  // ../RTL/cortexm0ds_logic.v(8361)
  buf u847 (vis_r5_o[25], Z9tpw6);  // ../RTL/cortexm0ds_logic.v(1909)
  not u8470 (Jpwiu6, n2169);  // ../RTL/cortexm0ds_logic.v(8361)
  and u8471 (Jf7iu6, Dmwiu6, Mnwiu6);  // ../RTL/cortexm0ds_logic.v(8362)
  and u8472 (Dmwiu6, Eqwiu6, C3qiu6);  // ../RTL/cortexm0ds_logic.v(8363)
  and u8473 (Tnwiu6, Lqwiu6, Sqwiu6);  // ../RTL/cortexm0ds_logic.v(8364)
  and u8474 (n2170, Lwgpw6[0], Ws4iu6);  // ../RTL/cortexm0ds_logic.v(8365)
  not u8475 (Sqwiu6, n2170);  // ../RTL/cortexm0ds_logic.v(8365)
  or u8476 (Is4iu6, Zqwiu6, Mfqiu6);  // ../RTL/cortexm0ds_logic.v(8366)
  not u8477 (Ws4iu6, Is4iu6);  // ../RTL/cortexm0ds_logic.v(8366)
  and u8478 (Lqwiu6, Grwiu6, Nrwiu6);  // ../RTL/cortexm0ds_logic.v(8367)
  and u8479 (n2171, Qhhhu6, Vr1iu6);  // ../RTL/cortexm0ds_logic.v(8368)
  buf u848 (vis_r8_o[3], Pdmpw6);  // ../RTL/cortexm0ds_logic.v(2579)
  not u8480 (Nrwiu6, n2171);  // ../RTL/cortexm0ds_logic.v(8368)
  and u8481 (Vr1iu6, Vuciu6, Urwiu6);  // ../RTL/cortexm0ds_logic.v(8369)
  buf u8482 (Osehu6, Ozkbx6[22]);  // ../RTL/cortexm0ds_logic.v(3176)
  not u8483 (Duhiu6, Bvtiu6);  // ../RTL/cortexm0ds_logic.v(8371)
  and u8484 (Bvtiu6, Fnwiu6, Vuciu6);  // ../RTL/cortexm0ds_logic.v(8372)
  and u8485 (Fnwiu6, Bswiu6, Dr6iu6);  // ../RTL/cortexm0ds_logic.v(8373)
  and u8486 (Ciwiu6, Iswiu6, Pswiu6);  // ../RTL/cortexm0ds_logic.v(8374)
  and u8487 (Pswiu6, Wswiu6, Dtwiu6);  // ../RTL/cortexm0ds_logic.v(8375)
  and u8488 (Dtwiu6, Ktwiu6, Rtwiu6);  // ../RTL/cortexm0ds_logic.v(8376)
  and u8489 (n2172, HRDATA[0], St1iu6);  // ../RTL/cortexm0ds_logic.v(8377)
  buf u849 (K7hpw6[31], Q2gax6);  // ../RTL/cortexm0ds_logic.v(2366)
  not u8490 (Rtwiu6, n2172);  // ../RTL/cortexm0ds_logic.v(8377)
  and u8491 (St1iu6, Ytwiu6, Ur4iu6);  // ../RTL/cortexm0ds_logic.v(8378)
  and u8492 (Ur4iu6, Fuwiu6, Q4wiu6);  // ../RTL/cortexm0ds_logic.v(8379)
  and u8493 (Fuwiu6, Cvciu6, Ukwiu6);  // ../RTL/cortexm0ds_logic.v(8380)
  and u8494 (Ktwiu6, Muwiu6, Tuwiu6);  // ../RTL/cortexm0ds_logic.v(8381)
  and u8495 (n2173, Smhhu6, Cs1iu6);  // ../RTL/cortexm0ds_logic.v(8382)
  not u8496 (Tuwiu6, n2173);  // ../RTL/cortexm0ds_logic.v(8382)
  and u8497 (Cs1iu6, Cpwiu6, Avwiu6);  // ../RTL/cortexm0ds_logic.v(8383)
  and u8498 (n2174, Ar1iu6, Fkfpw6[0]);  // ../RTL/cortexm0ds_logic.v(8384)
  not u8499 (Muwiu6, n2174);  // ../RTL/cortexm0ds_logic.v(8384)
  buf u85 (K7hpw6[18], Xc9ax6);  // ../RTL/cortexm0ds_logic.v(2366)
  buf u850 (vis_r14_o[30], S1nax6);  // ../RTL/cortexm0ds_logic.v(2497)
  and u8500 (Ar1iu6, Rzciu6, D5eiu6);  // ../RTL/cortexm0ds_logic.v(8385)
  and u8501 (Wswiu6, Hvwiu6, Ovwiu6);  // ../RTL/cortexm0ds_logic.v(8386)
  and u8502 (n2175, Alhhu6, Dw1iu6);  // ../RTL/cortexm0ds_logic.v(8387)
  not u8503 (Ovwiu6, n2175);  // ../RTL/cortexm0ds_logic.v(8387)
  and u8504 (Dw1iu6, Avwiu6, Urwiu6);  // ../RTL/cortexm0ds_logic.v(8388)
  and u8505 (Urwiu6, Vvwiu6, X8hpw6[6]);  // ../RTL/cortexm0ds_logic.v(8389)
  or u8506 (n2176, X8hpw6[0], X8hpw6[5]);  // ../RTL/cortexm0ds_logic.v(8390)
  not u8507 (Vvwiu6, n2176);  // ../RTL/cortexm0ds_logic.v(8390)
  and u8508 (Hvwiu6, Cwwiu6, Jwwiu6);  // ../RTL/cortexm0ds_logic.v(8391)
  and u8509 (n2177, Zt1iu6, Pzgpw6[0]);  // ../RTL/cortexm0ds_logic.v(8392)
  buf u851 (vis_r3_o[4], J3xax6);  // ../RTL/cortexm0ds_logic.v(2694)
  not u8510 (Jwwiu6, n2177);  // ../RTL/cortexm0ds_logic.v(8392)
  and u8511 (Zt1iu6, Avwiu6, Nkwiu6);  // ../RTL/cortexm0ds_logic.v(8393)
  and u8512 (Avwiu6, Dzqiu6, Mnwiu6);  // ../RTL/cortexm0ds_logic.v(8394)
  and u8513 (n2178, Ijhhu6, Xs1iu6);  // ../RTL/cortexm0ds_logic.v(8395)
  not u8514 (Cwwiu6, n2178);  // ../RTL/cortexm0ds_logic.v(8395)
  and u8515 (Xs1iu6, Cpwiu6, Vuciu6);  // ../RTL/cortexm0ds_logic.v(8396)
  and u8516 (Vuciu6, Mnwiu6, Ukwiu6);  // ../RTL/cortexm0ds_logic.v(8397)
  and u8517 (Iswiu6, Qwwiu6, Xwwiu6);  // ../RTL/cortexm0ds_logic.v(8398)
  or u8518 (n2179, Exwiu6, Ylqiu6);  // ../RTL/cortexm0ds_logic.v(8399)
  not u8519 (Xwwiu6, n2179);  // ../RTL/cortexm0ds_logic.v(8399)
  buf u852 (vis_r7_o[30], Rpvax6);  // ../RTL/cortexm0ds_logic.v(2654)
  and u8520 (n2180, Lxwiu6, Sxwiu6);  // ../RTL/cortexm0ds_logic.v(8400)
  not u8521 (Ylqiu6, n2180);  // ../RTL/cortexm0ds_logic.v(8400)
  and u8522 (n2181, Zxwiu6, Ffqiu6);  // ../RTL/cortexm0ds_logic.v(8401)
  not u8523 (Sxwiu6, n2181);  // ../RTL/cortexm0ds_logic.v(8401)
  and u8524 (Zxwiu6, Ilwiu6, Dr6iu6);  // ../RTL/cortexm0ds_logic.v(8402)
  and u8525 (n2182, Gywiu6, A2qiu6);  // ../RTL/cortexm0ds_logic.v(8403)
  not u8526 (Lxwiu6, n2182);  // ../RTL/cortexm0ds_logic.v(8403)
  and u8527 (Gywiu6, Bswiu6, Nywiu6);  // ../RTL/cortexm0ds_logic.v(8404)
  and u8528 (n2183, Yw1iu6, Uywiu6);  // ../RTL/cortexm0ds_logic.v(8405)
  not u8529 (Exwiu6, n2183);  // ../RTL/cortexm0ds_logic.v(8405)
  buf u853 (vis_msp_o[25], T00qw6);  // ../RTL/cortexm0ds_logic.v(2097)
  and u8530 (n2184, Kw1iu6, V5hpw6[0]);  // ../RTL/cortexm0ds_logic.v(8406)
  not u8531 (Uywiu6, n2184);  // ../RTL/cortexm0ds_logic.v(8406)
  or u8532 (n2185, Nwriu6, Zqwiu6);  // ../RTL/cortexm0ds_logic.v(8407)
  not u8533 (Kw1iu6, n2185);  // ../RTL/cortexm0ds_logic.v(8407)
  not u8534 (Nwriu6, Dzqiu6);  // ../RTL/cortexm0ds_logic.v(8408)
  and u8535 (Yw1iu6, Bzwiu6, Uvsiu6);  // ../RTL/cortexm0ds_logic.v(8409)
  and u8536 (Uvsiu6, Izwiu6, Reqiu6);  // ../RTL/cortexm0ds_logic.v(8410)
  and u8537 (n2186, Iv1iu6, Pzwiu6);  // ../RTL/cortexm0ds_logic.v(8411)
  not u8538 (Reqiu6, n2186);  // ../RTL/cortexm0ds_logic.v(8411)
  and u8539 (Iv1iu6, Wzwiu6, Vowiu6);  // ../RTL/cortexm0ds_logic.v(8412)
  buf u854 (vis_r11_o[22], T1fbx6);  // ../RTL/cortexm0ds_logic.v(1874)
  and u8540 (Vowiu6, Q4wiu6, Ukwiu6);  // ../RTL/cortexm0ds_logic.v(8413)
  and u8541 (Wzwiu6, X8hpw6[0], Bswiu6);  // ../RTL/cortexm0ds_logic.v(8414)
  and u8542 (n2187, D0xiu6, K0xiu6);  // ../RTL/cortexm0ds_logic.v(8415)
  not u8543 (Izwiu6, n2187);  // ../RTL/cortexm0ds_logic.v(8415)
  and u8544 (D0xiu6, Bqriu6, Q4wiu6);  // ../RTL/cortexm0ds_logic.v(8416)
  and u8545 (Bzwiu6, R0xiu6, Hssiu6);  // ../RTL/cortexm0ds_logic.v(8417)
  and u8546 (n2188, Y0xiu6, Mnwiu6);  // ../RTL/cortexm0ds_logic.v(8418)
  not u8547 (Hssiu6, n2188);  // ../RTL/cortexm0ds_logic.v(8418)
  or u8548 (n2189, Fl6iu6, X8hpw6[1]);  // ../RTL/cortexm0ds_logic.v(8419)
  not u8549 (Mnwiu6, n2189);  // ../RTL/cortexm0ds_logic.v(8419)
  or u855 (Qbfpw6[25], Vj8ju6, M75ju6);  // ../RTL/cortexm0ds_logic.v(9482)
  and u8550 (Y0xiu6, Ilwiu6, K0xiu6);  // ../RTL/cortexm0ds_logic.v(8420)
  or u8551 (R0xiu6, Zqwiu6, J3qiu6);  // ../RTL/cortexm0ds_logic.v(8421)
  not u8552 (J3qiu6, Bqriu6);  // ../RTL/cortexm0ds_logic.v(8422)
  and u8553 (n2190, Nkwiu6, Q4wiu6);  // ../RTL/cortexm0ds_logic.v(8423)
  not u8554 (Zqwiu6, n2190);  // ../RTL/cortexm0ds_logic.v(8423)
  and u8555 (Qwwiu6, F1xiu6, M1xiu6);  // ../RTL/cortexm0ds_logic.v(8424)
  and u8556 (F1xiu6, Uwriu6, Qaqiu6);  // ../RTL/cortexm0ds_logic.v(8425)
  and u8557 (Qaqiu6, Anqiu6, T1xiu6);  // ../RTL/cortexm0ds_logic.v(8426)
  and u8558 (n2191, Ffqiu6, Nywiu6);  // ../RTL/cortexm0ds_logic.v(8427)
  not u8559 (T1xiu6, n2191);  // ../RTL/cortexm0ds_logic.v(8427)
  buf u856 (vis_r4_o[28], Rhibx6);  // ../RTL/cortexm0ds_logic.v(2626)
  not u8560 (Nywiu6, A2xiu6);  // ../RTL/cortexm0ds_logic.v(8428)
  AL_MUX u8561 (
    .i0(H2xiu6),
    .i1(Mfqiu6),
    .sel(X8hpw6[0]),
    .o(A2xiu6));  // ../RTL/cortexm0ds_logic.v(8429)
  not u8562 (Mfqiu6, Ukwiu6);  // ../RTL/cortexm0ds_logic.v(8430)
  and u8563 (Ffqiu6, O2xiu6, X8hpw6[1]);  // ../RTL/cortexm0ds_logic.v(8431)
  and u8564 (O2xiu6, Bswiu6, Fl6iu6);  // ../RTL/cortexm0ds_logic.v(8432)
  and u8565 (Anqiu6, V2xiu6, C3xiu6);  // ../RTL/cortexm0ds_logic.v(8433)
  and u8566 (n2192, Mmqiu6, A2qiu6);  // ../RTL/cortexm0ds_logic.v(8434)
  not u8567 (C3xiu6, n2192);  // ../RTL/cortexm0ds_logic.v(8434)
  and u8568 (Mmqiu6, Nkwiu6, Bqriu6);  // ../RTL/cortexm0ds_logic.v(8435)
  and u8569 (Nkwiu6, J3xiu6, X8hpw6[0]);  // ../RTL/cortexm0ds_logic.v(8436)
  buf u857 (Jfgpw6[1], I5xax6);  // ../RTL/cortexm0ds_logic.v(2010)
  or u8570 (n2193, Zh6iu6, X8hpw6[5]);  // ../RTL/cortexm0ds_logic.v(8437)
  not u8571 (J3xiu6, n2193);  // ../RTL/cortexm0ds_logic.v(8437)
  and u8572 (n2194, Bswiu6, Q3xiu6);  // ../RTL/cortexm0ds_logic.v(8438)
  not u8573 (V2xiu6, n2194);  // ../RTL/cortexm0ds_logic.v(8438)
  and u8574 (n2195, X3xiu6, E4xiu6);  // ../RTL/cortexm0ds_logic.v(8439)
  not u8575 (Q3xiu6, n2195);  // ../RTL/cortexm0ds_logic.v(8439)
  and u8576 (n2196, Ryriu6, Dr6iu6);  // ../RTL/cortexm0ds_logic.v(8440)
  not u8577 (E4xiu6, n2196);  // ../RTL/cortexm0ds_logic.v(8440)
  and u8578 (Ryriu6, A2qiu6, L4xiu6);  // ../RTL/cortexm0ds_logic.v(8441)
  or u8579 (L4xiu6, Ilwiu6, Ukwiu6);  // ../RTL/cortexm0ds_logic.v(8442)
  buf u858 (vis_r5_o[20], Llppw6);  // ../RTL/cortexm0ds_logic.v(1909)
  and u8580 (n2197, A2qiu6, C3qiu6);  // ../RTL/cortexm0ds_logic.v(8443)
  not u8581 (X3xiu6, n2197);  // ../RTL/cortexm0ds_logic.v(8443)
  and u8582 (C3qiu6, Dzqiu6, X8hpw6[0]);  // ../RTL/cortexm0ds_logic.v(8444)
  and u8583 (A2qiu6, X8hpw6[1], X8hpw6[4]);  // ../RTL/cortexm0ds_logic.v(8445)
  or u8584 (n2198, Zh6iu6, Wj6iu6);  // ../RTL/cortexm0ds_logic.v(8446)
  not u8585 (Bswiu6, n2198);  // ../RTL/cortexm0ds_logic.v(8446)
  not u8586 (Zh6iu6, X8hpw6[6]);  // ../RTL/cortexm0ds_logic.v(8447)
  and u8587 (Uwriu6, S4xiu6, Z4xiu6);  // ../RTL/cortexm0ds_logic.v(8448)
  and u8588 (n2199, Fl6iu6, G5xiu6);  // ../RTL/cortexm0ds_logic.v(8449)
  not u8589 (Z4xiu6, n2199);  // ../RTL/cortexm0ds_logic.v(8449)
  buf u859 (vis_r8_o[2], Serax6);  // ../RTL/cortexm0ds_logic.v(2579)
  or u8590 (G5xiu6, N5xiu6, Iqriu6);  // ../RTL/cortexm0ds_logic.v(8450)
  and u8591 (Iqriu6, Ixriu6, Vm6iu6);  // ../RTL/cortexm0ds_logic.v(8451)
  and u8592 (Ixriu6, U5xiu6, X8hpw6[1]);  // ../RTL/cortexm0ds_logic.v(8452)
  and u8593 (U5xiu6, K0xiu6, X8hpw6[2]);  // ../RTL/cortexm0ds_logic.v(8453)
  and u8594 (K0xiu6, Eqwiu6, X8hpw6[0]);  // ../RTL/cortexm0ds_logic.v(8454)
  or u8595 (n2200, Wj6iu6, X8hpw6[6]);  // ../RTL/cortexm0ds_logic.v(8455)
  not u8596 (Eqwiu6, n2200);  // ../RTL/cortexm0ds_logic.v(8455)
  not u8597 (Wj6iu6, X8hpw6[5]);  // ../RTL/cortexm0ds_logic.v(8456)
  and u8598 (N5xiu6, Wyqiu6, Ukwiu6);  // ../RTL/cortexm0ds_logic.v(8457)
  and u8599 (Ukwiu6, Eo6iu6, Vm6iu6);  // ../RTL/cortexm0ds_logic.v(8458)
  buf u86 (vis_r2_o[29], Vkqax6);  // ../RTL/cortexm0ds_logic.v(2551)
  buf u860 (vis_r14_o[29], Nlnax6);  // ../RTL/cortexm0ds_logic.v(2497)
  and u8600 (Wyqiu6, B6xiu6, X8hpw6[1]);  // ../RTL/cortexm0ds_logic.v(8459)
  and u8601 (B6xiu6, X8hpw6[0], X4wiu6);  // ../RTL/cortexm0ds_logic.v(8460)
  or u8602 (S4xiu6, Svriu6, H2xiu6);  // ../RTL/cortexm0ds_logic.v(8461)
  or u8603 (n2201, Bqriu6, Dzqiu6);  // ../RTL/cortexm0ds_logic.v(8462)
  not u8604 (H2xiu6, n2201);  // ../RTL/cortexm0ds_logic.v(8462)
  and u8605 (Dzqiu6, X8hpw6[3], Eo6iu6);  // ../RTL/cortexm0ds_logic.v(8463)
  not u8606 (Eo6iu6, X8hpw6[2]);  // ../RTL/cortexm0ds_logic.v(8464)
  and u8607 (Bqriu6, X8hpw6[3], X8hpw6[2]);  // ../RTL/cortexm0ds_logic.v(8465)
  and u8608 (n2202, I6xiu6, X8hpw6[1]);  // ../RTL/cortexm0ds_logic.v(8466)
  not u8609 (Svriu6, n2202);  // ../RTL/cortexm0ds_logic.v(8466)
  buf u861 (vis_r3_o[3], U3yax6);  // ../RTL/cortexm0ds_logic.v(2694)
  and u8610 (I6xiu6, Cvciu6, Fl6iu6);  // ../RTL/cortexm0ds_logic.v(8467)
  not u8611 (Fl6iu6, X8hpw6[4]);  // ../RTL/cortexm0ds_logic.v(8468)
  and u8612 (Cvciu6, X4wiu6, Dr6iu6);  // ../RTL/cortexm0ds_logic.v(8469)
  not u8613 (Dr6iu6, X8hpw6[0]);  // ../RTL/cortexm0ds_logic.v(8470)
  or u8614 (n2203, X8hpw6[5], X8hpw6[6]);  // ../RTL/cortexm0ds_logic.v(8471)
  not u8615 (X4wiu6, n2203);  // ../RTL/cortexm0ds_logic.v(8471)
  and u8616 (Wo1iu6, P6xiu6, W6xiu6);  // ../RTL/cortexm0ds_logic.v(8472)
  and u8617 (P6xiu6, D7xiu6, K7xiu6);  // ../RTL/cortexm0ds_logic.v(8473)
  and u8618 (n2204, R7xiu6, Y7xiu6);  // ../RTL/cortexm0ds_logic.v(8474)
  not u8619 (K7xiu6, n2204);  // ../RTL/cortexm0ds_logic.v(8474)
  buf u862 (vis_r7_o[29], M9wax6);  // ../RTL/cortexm0ds_logic.v(2654)
  or u8620 (Y7xiu6, Xp4iu6, C44iu6);  // ../RTL/cortexm0ds_logic.v(8475)
  not u8621 (D7xiu6, Sf1iu6);  // ../RTL/cortexm0ds_logic.v(8476)
  and u8622 (Wewiu6, Untiu6, F8xiu6);  // ../RTL/cortexm0ds_logic.v(8477)
  and u8623 (n2205, Uthpw6[0], Sf1iu6);  // ../RTL/cortexm0ds_logic.v(8478)
  not u8624 (F8xiu6, n2205);  // ../RTL/cortexm0ds_logic.v(8478)
  and u8625 (Untiu6, V1riu6, Po1iu6);  // ../RTL/cortexm0ds_logic.v(8479)
  and u8626 (n2206, M8xiu6, C44iu6);  // ../RTL/cortexm0ds_logic.v(8480)
  not u8627 (Po1iu6, n2206);  // ../RTL/cortexm0ds_logic.v(8480)
  not u8628 (V1riu6, Tx1iu6);  // ../RTL/cortexm0ds_logic.v(8481)
  and u8629 (Tx1iu6, M8xiu6, Vo4iu6);  // ../RTL/cortexm0ds_logic.v(8482)
  buf u863 (vis_msp_o[24], Tyzpw6);  // ../RTL/cortexm0ds_logic.v(2097)
  and u8630 (M8xiu6, T8xiu6, A9xiu6);  // ../RTL/cortexm0ds_logic.v(8483)
  or u8631 (n2207, R7xiu6, W6xiu6);  // ../RTL/cortexm0ds_logic.v(8484)
  not u8632 (A9xiu6, n2207);  // ../RTL/cortexm0ds_logic.v(8484)
  and u8633 (W6xiu6, Sq4iu6, H9xiu6);  // ../RTL/cortexm0ds_logic.v(8486)
  not u8634 (Ohwiu6, W6xiu6);  // ../RTL/cortexm0ds_logic.v(8486)
  not u8635 (R7xiu6, Ho4iu6);  // ../RTL/cortexm0ds_logic.v(8487)
  or u8636 (n2208, Sf1iu6, Xp4iu6);  // ../RTL/cortexm0ds_logic.v(8488)
  not u8637 (T8xiu6, n2208);  // ../RTL/cortexm0ds_logic.v(8488)
  not u8638 (Xp4iu6, Wu9iu6);  // ../RTL/cortexm0ds_logic.v(8489)
  or u8639 (Sf1iu6, O9xiu6, Npzhu6);  // ../RTL/cortexm0ds_logic.v(8490)
  buf u864 (vis_r11_o[21], Rdkpw6);  // ../RTL/cortexm0ds_logic.v(1874)
  not u8640 (Npzhu6, Sqhpw6[1]);  // ../RTL/cortexm0ds_logic.v(8491)
  AL_MUX u8641 (
    .i0(Fszhu6),
    .i1(V9xiu6),
    .sel(Sqhpw6[0]),
    .o(O9xiu6));  // ../RTL/cortexm0ds_logic.v(8492)
  buf u8642 (Cuehu6, Ozkbx6[21]);  // ../RTL/cortexm0ds_logic.v(3176)
  and u8643 (Pqzhu6, Caxiu6, Wu9iu6);  // ../RTL/cortexm0ds_logic.v(8494)
  and u8644 (Wu9iu6, Cjhpw6[1], Iqzhu6);  // ../RTL/cortexm0ds_logic.v(8495)
  or u8645 (n2209, C44iu6, Eq4iu6);  // ../RTL/cortexm0ds_logic.v(8496)
  not u8646 (Caxiu6, n2209);  // ../RTL/cortexm0ds_logic.v(8496)
  not u8647 (C44iu6, Vo4iu6);  // ../RTL/cortexm0ds_logic.v(8497)
  and u8648 (Vo4iu6, Cjhpw6[0], Iqzhu6);  // ../RTL/cortexm0ds_logic.v(8498)
  not u8649 (Fszhu6, Drzhu6);  // ../RTL/cortexm0ds_logic.v(8499)
  buf u865 (Hrfpw6[16], Tajax6);  // ../RTL/cortexm0ds_logic.v(2428)
  and u8650 (Drzhu6, HREADY, Jaxiu6);  // ../RTL/cortexm0ds_logic.v(8500)
  and u8651 (n2210, Qaxiu6, Xaxiu6);  // ../RTL/cortexm0ds_logic.v(8501)
  not u8652 (Jaxiu6, n2210);  // ../RTL/cortexm0ds_logic.v(8501)
  and u8653 (Aj9pw6, HMASTER, Ebxiu6);  // ../RTL/cortexm0ds_logic.v(8502)
  not u8654 (Xaxiu6, Aj9pw6);  // ../RTL/cortexm0ds_logic.v(8502)
  and u8655 (J5phu6, Fk7iu6, Lbxiu6);  // ../RTL/cortexm0ds_logic.v(8503)
  and u8656 (n2211, Sbxiu6, Zbxiu6);  // ../RTL/cortexm0ds_logic.v(8504)
  not u8657 (Lbxiu6, n2211);  // ../RTL/cortexm0ds_logic.v(8504)
  and u8658 (n2212, Xudpw6, IRQ[0]);  // ../RTL/cortexm0ds_logic.v(8505)
  not u8659 (Zbxiu6, n2212);  // ../RTL/cortexm0ds_logic.v(8505)
  buf u866 (vis_r4_o[27], Wnuax6);  // ../RTL/cortexm0ds_logic.v(2626)
  and u8660 (Sbxiu6, Gcxiu6, Yj7iu6);  // ../RTL/cortexm0ds_logic.v(8506)
  and u8661 (n2213, Kwfiu6, HWDATA[0]);  // ../RTL/cortexm0ds_logic.v(8507)
  not u8662 (Yj7iu6, n2213);  // ../RTL/cortexm0ds_logic.v(8507)
  and u8663 (n2214, Odgpw6[0], Ncxiu6);  // ../RTL/cortexm0ds_logic.v(8508)
  not u8664 (Gcxiu6, n2214);  // ../RTL/cortexm0ds_logic.v(8508)
  and u8665 (n2215, K66iu6, HWDATA[0]);  // ../RTL/cortexm0ds_logic.v(8509)
  not u8666 (Ncxiu6, n2215);  // ../RTL/cortexm0ds_logic.v(8509)
  or u8667 (Fk7iu6, Sb5iu6, Ucxiu6);  // ../RTL/cortexm0ds_logic.v(8510)
  and u8668 (C5phu6, Dogiu6, Bdxiu6);  // ../RTL/cortexm0ds_logic.v(8511)
  and u8669 (n2216, Idxiu6, Pdxiu6);  // ../RTL/cortexm0ds_logic.v(8512)
  buf u867 (K7hpw6[27], Itcbx6);  // ../RTL/cortexm0ds_logic.v(2366)
  not u8670 (Bdxiu6, n2216);  // ../RTL/cortexm0ds_logic.v(8512)
  and u8671 (n2217, Fsdpw6, IRQ[1]);  // ../RTL/cortexm0ds_logic.v(8513)
  not u8672 (Pdxiu6, n2217);  // ../RTL/cortexm0ds_logic.v(8513)
  and u8673 (Idxiu6, Wdxiu6, Wngiu6);  // ../RTL/cortexm0ds_logic.v(8514)
  and u8674 (n2218, Kwfiu6, I4eiu6);  // ../RTL/cortexm0ds_logic.v(8515)
  not u8675 (Wngiu6, n2218);  // ../RTL/cortexm0ds_logic.v(8515)
  and u8676 (n2219, Odgpw6[1], Dexiu6);  // ../RTL/cortexm0ds_logic.v(8516)
  not u8677 (Wdxiu6, n2219);  // ../RTL/cortexm0ds_logic.v(8516)
  and u8678 (n2220, K66iu6, I4eiu6);  // ../RTL/cortexm0ds_logic.v(8517)
  not u8679 (Dexiu6, n2220);  // ../RTL/cortexm0ds_logic.v(8517)
  buf u868 (Jfgpw6[4], Ztupw6);  // ../RTL/cortexm0ds_logic.v(2010)
  and u8680 (I4eiu6, Npdhu6, HWDATA[1]);  // ../RTL/cortexm0ds_logic.v(8518)
  or u8681 (Dogiu6, Sb5iu6, Kexiu6);  // ../RTL/cortexm0ds_logic.v(8519)
  and u8682 (V4phu6, Zlgiu6, Rexiu6);  // ../RTL/cortexm0ds_logic.v(8521)
  and u8683 (n2221, Yexiu6, Ffxiu6);  // ../RTL/cortexm0ds_logic.v(8522)
  not u8684 (Rexiu6, n2221);  // ../RTL/cortexm0ds_logic.v(8522)
  and u8685 (n2222, Eodpw6, IRQ[2]);  // ../RTL/cortexm0ds_logic.v(8523)
  not u8686 (Ffxiu6, n2222);  // ../RTL/cortexm0ds_logic.v(8523)
  and u8687 (Yexiu6, Mfxiu6, Slgiu6);  // ../RTL/cortexm0ds_logic.v(8524)
  and u8688 (n2223, G3eiu6, Kwfiu6);  // ../RTL/cortexm0ds_logic.v(8525)
  not u8689 (Slgiu6, n2223);  // ../RTL/cortexm0ds_logic.v(8525)
  buf u869 (vis_r5_o[28], Rjibx6);  // ../RTL/cortexm0ds_logic.v(1909)
  and u8690 (n2224, Odgpw6[2], Tfxiu6);  // ../RTL/cortexm0ds_logic.v(8526)
  not u8691 (Mfxiu6, n2224);  // ../RTL/cortexm0ds_logic.v(8526)
  and u8692 (n2225, G3eiu6, K66iu6);  // ../RTL/cortexm0ds_logic.v(8527)
  not u8693 (Tfxiu6, n2225);  // ../RTL/cortexm0ds_logic.v(8527)
  or u8694 (Zlgiu6, Sb5iu6, Agxiu6);  // ../RTL/cortexm0ds_logic.v(8528)
  and u8695 (O4phu6, Xefiu6, Hgxiu6);  // ../RTL/cortexm0ds_logic.v(8529)
  and u8696 (n2226, Ogxiu6, Vgxiu6);  // ../RTL/cortexm0ds_logic.v(8530)
  not u8697 (Hgxiu6, n2226);  // ../RTL/cortexm0ds_logic.v(8530)
  and u8698 (n2227, Jndpw6, IRQ[3]);  // ../RTL/cortexm0ds_logic.v(8531)
  not u8699 (Vgxiu6, n2227);  // ../RTL/cortexm0ds_logic.v(8531)
  buf u87 (vis_r2_o[14], U2rax6);  // ../RTL/cortexm0ds_logic.v(2551)
  buf u870 (vis_r5_o[29], Lhppw6);  // ../RTL/cortexm0ds_logic.v(1909)
  and u8700 (Ogxiu6, Chxiu6, Qefiu6);  // ../RTL/cortexm0ds_logic.v(8532)
  and u8701 (n2228, Kwfiu6, HWDATA[3]);  // ../RTL/cortexm0ds_logic.v(8533)
  not u8702 (Qefiu6, n2228);  // ../RTL/cortexm0ds_logic.v(8533)
  and u8703 (n2229, Odgpw6[3], Jhxiu6);  // ../RTL/cortexm0ds_logic.v(8534)
  not u8704 (Chxiu6, n2229);  // ../RTL/cortexm0ds_logic.v(8534)
  and u8705 (n2230, K66iu6, HWDATA[3]);  // ../RTL/cortexm0ds_logic.v(8535)
  not u8706 (Jhxiu6, n2230);  // ../RTL/cortexm0ds_logic.v(8535)
  or u8707 (Xefiu6, Sb5iu6, Qhxiu6);  // ../RTL/cortexm0ds_logic.v(8536)
  and u8708 (H4phu6, Tcfiu6, Xhxiu6);  // ../RTL/cortexm0ds_logic.v(8537)
  and u8709 (n2231, Eixiu6, Lixiu6);  // ../RTL/cortexm0ds_logic.v(8538)
  buf u871 (vis_r5_o[30], N7ppw6);  // ../RTL/cortexm0ds_logic.v(1909)
  not u8710 (Xhxiu6, n2231);  // ../RTL/cortexm0ds_logic.v(8538)
  and u8711 (n2232, Qndpw6, IRQ[4]);  // ../RTL/cortexm0ds_logic.v(8539)
  not u8712 (Lixiu6, n2232);  // ../RTL/cortexm0ds_logic.v(8539)
  and u8713 (Eixiu6, Sixiu6, Mcfiu6);  // ../RTL/cortexm0ds_logic.v(8540)
  and u8714 (n2233, Kwfiu6, HWDATA[4]);  // ../RTL/cortexm0ds_logic.v(8541)
  not u8715 (Mcfiu6, n2233);  // ../RTL/cortexm0ds_logic.v(8541)
  and u8716 (n2234, Odgpw6[4], Zixiu6);  // ../RTL/cortexm0ds_logic.v(8542)
  not u8717 (Sixiu6, n2234);  // ../RTL/cortexm0ds_logic.v(8542)
  and u8718 (n2235, K66iu6, HWDATA[4]);  // ../RTL/cortexm0ds_logic.v(8543)
  not u8719 (Zixiu6, n2235);  // ../RTL/cortexm0ds_logic.v(8543)
  buf u872 (vis_r5_o[31], N9ppw6);  // ../RTL/cortexm0ds_logic.v(1909)
  or u8720 (Tcfiu6, Sb5iu6, Gjxiu6);  // ../RTL/cortexm0ds_logic.v(8544)
  and u8721 (A4phu6, Pafiu6, Njxiu6);  // ../RTL/cortexm0ds_logic.v(8546)
  and u8722 (n2236, Ujxiu6, Bkxiu6);  // ../RTL/cortexm0ds_logic.v(8547)
  not u8723 (Njxiu6, n2236);  // ../RTL/cortexm0ds_logic.v(8547)
  and u8724 (n2237, Gpdpw6, IRQ[5]);  // ../RTL/cortexm0ds_logic.v(8548)
  not u8725 (Bkxiu6, n2237);  // ../RTL/cortexm0ds_logic.v(8548)
  and u8726 (Ujxiu6, Ikxiu6, Iafiu6);  // ../RTL/cortexm0ds_logic.v(8549)
  and u8727 (n2238, Kwfiu6, HWDATA[5]);  // ../RTL/cortexm0ds_logic.v(8550)
  not u8728 (Iafiu6, n2238);  // ../RTL/cortexm0ds_logic.v(8550)
  and u8729 (n2239, Odgpw6[5], Pkxiu6);  // ../RTL/cortexm0ds_logic.v(8551)
  buf u873 (vis_r8_o[9], Oesax6);  // ../RTL/cortexm0ds_logic.v(2579)
  not u8730 (Ikxiu6, n2239);  // ../RTL/cortexm0ds_logic.v(8551)
  and u8731 (n2240, K66iu6, HWDATA[5]);  // ../RTL/cortexm0ds_logic.v(8552)
  not u8732 (Pkxiu6, n2240);  // ../RTL/cortexm0ds_logic.v(8552)
  or u8733 (Pafiu6, Sb5iu6, Wkxiu6);  // ../RTL/cortexm0ds_logic.v(8553)
  and u8734 (T3phu6, L8fiu6, Dlxiu6);  // ../RTL/cortexm0ds_logic.v(8554)
  and u8735 (n2241, Klxiu6, Rlxiu6);  // ../RTL/cortexm0ds_logic.v(8555)
  not u8736 (Dlxiu6, n2241);  // ../RTL/cortexm0ds_logic.v(8555)
  and u8737 (n2242, Lodpw6, IRQ[6]);  // ../RTL/cortexm0ds_logic.v(8556)
  not u8738 (Rlxiu6, n2242);  // ../RTL/cortexm0ds_logic.v(8556)
  and u8739 (Klxiu6, Ylxiu6, E8fiu6);  // ../RTL/cortexm0ds_logic.v(8557)
  buf u874 (Aphpw6[2], Dugax6);  // ../RTL/cortexm0ds_logic.v(2381)
  and u8740 (n2243, Kwfiu6, HWDATA[6]);  // ../RTL/cortexm0ds_logic.v(8558)
  not u8741 (E8fiu6, n2243);  // ../RTL/cortexm0ds_logic.v(8558)
  and u8742 (n2244, Odgpw6[6], Fmxiu6);  // ../RTL/cortexm0ds_logic.v(8559)
  not u8743 (Ylxiu6, n2244);  // ../RTL/cortexm0ds_logic.v(8559)
  and u8744 (n2245, K66iu6, HWDATA[6]);  // ../RTL/cortexm0ds_logic.v(8560)
  not u8745 (Fmxiu6, n2245);  // ../RTL/cortexm0ds_logic.v(8560)
  or u8746 (L8fiu6, Sb5iu6, Mmxiu6);  // ../RTL/cortexm0ds_logic.v(8561)
  and u8747 (M3phu6, H6fiu6, Tmxiu6);  // ../RTL/cortexm0ds_logic.v(8562)
  and u8748 (n2246, Anxiu6, Hnxiu6);  // ../RTL/cortexm0ds_logic.v(8563)
  not u8749 (Tmxiu6, n2246);  // ../RTL/cortexm0ds_logic.v(8563)
  buf u875 (vis_r9_o[5], Propw6);  // ../RTL/cortexm0ds_logic.v(1898)
  and u8750 (n2247, Zodpw6, IRQ[7]);  // ../RTL/cortexm0ds_logic.v(8564)
  not u8751 (Hnxiu6, n2247);  // ../RTL/cortexm0ds_logic.v(8564)
  and u8752 (Anxiu6, Onxiu6, A6fiu6);  // ../RTL/cortexm0ds_logic.v(8565)
  and u8753 (n2248, Kwfiu6, HWDATA[7]);  // ../RTL/cortexm0ds_logic.v(8566)
  not u8754 (A6fiu6, n2248);  // ../RTL/cortexm0ds_logic.v(8566)
  and u8755 (n2249, Odgpw6[7], Vnxiu6);  // ../RTL/cortexm0ds_logic.v(8567)
  not u8756 (Onxiu6, n2249);  // ../RTL/cortexm0ds_logic.v(8567)
  and u8757 (n2250, K66iu6, HWDATA[7]);  // ../RTL/cortexm0ds_logic.v(8568)
  not u8758 (Vnxiu6, n2250);  // ../RTL/cortexm0ds_logic.v(8568)
  or u8759 (H6fiu6, Sb5iu6, Coxiu6);  // ../RTL/cortexm0ds_logic.v(8569)
  buf u876 (vis_r3_o[10], Do6bx6);  // ../RTL/cortexm0ds_logic.v(2694)
  and u8760 (F3phu6, Mbgiu6, Joxiu6);  // ../RTL/cortexm0ds_logic.v(8570)
  and u8761 (n2251, Qoxiu6, Xoxiu6);  // ../RTL/cortexm0ds_logic.v(8571)
  not u8762 (Joxiu6, n2251);  // ../RTL/cortexm0ds_logic.v(8571)
  and u8763 (n2252, Judpw6, IRQ[10]);  // ../RTL/cortexm0ds_logic.v(8572)
  not u8764 (Xoxiu6, n2252);  // ../RTL/cortexm0ds_logic.v(8572)
  and u8765 (Qoxiu6, Epxiu6, Fbgiu6);  // ../RTL/cortexm0ds_logic.v(8573)
  and u8766 (n2253, Kwfiu6, HWDATA[10]);  // ../RTL/cortexm0ds_logic.v(8574)
  not u8767 (Fbgiu6, n2253);  // ../RTL/cortexm0ds_logic.v(8574)
  and u8768 (n2254, Odgpw6[10], Lpxiu6);  // ../RTL/cortexm0ds_logic.v(8575)
  not u8769 (Epxiu6, n2254);  // ../RTL/cortexm0ds_logic.v(8575)
  buf u877 (vis_msp_o[5], Uuzpw6);  // ../RTL/cortexm0ds_logic.v(2097)
  and u8770 (n2255, K66iu6, HWDATA[10]);  // ../RTL/cortexm0ds_logic.v(8576)
  not u8771 (Lpxiu6, n2255);  // ../RTL/cortexm0ds_logic.v(8576)
  or u8772 (Mbgiu6, Sb5iu6, Spxiu6);  // ../RTL/cortexm0ds_logic.v(8577)
  and u8773 (Y2phu6, I9giu6, Zpxiu6);  // ../RTL/cortexm0ds_logic.v(8578)
  and u8774 (n2256, Gqxiu6, Nqxiu6);  // ../RTL/cortexm0ds_logic.v(8579)
  not u8775 (Zpxiu6, n2256);  // ../RTL/cortexm0ds_logic.v(8579)
  and u8776 (n2257, Cudpw6, IRQ[11]);  // ../RTL/cortexm0ds_logic.v(8580)
  not u8777 (Nqxiu6, n2257);  // ../RTL/cortexm0ds_logic.v(8580)
  and u8778 (Gqxiu6, Uqxiu6, B9giu6);  // ../RTL/cortexm0ds_logic.v(8581)
  and u8779 (n2258, Kwfiu6, HWDATA[11]);  // ../RTL/cortexm0ds_logic.v(8582)
  buf u878 (vis_r11_o[2], Xhtpw6);  // ../RTL/cortexm0ds_logic.v(1874)
  not u8780 (B9giu6, n2258);  // ../RTL/cortexm0ds_logic.v(8582)
  and u8781 (n2259, Odgpw6[11], Brxiu6);  // ../RTL/cortexm0ds_logic.v(8583)
  not u8782 (Uqxiu6, n2259);  // ../RTL/cortexm0ds_logic.v(8583)
  and u8783 (n2260, K66iu6, HWDATA[11]);  // ../RTL/cortexm0ds_logic.v(8584)
  not u8784 (Brxiu6, n2260);  // ../RTL/cortexm0ds_logic.v(8584)
  or u8785 (I9giu6, Sb5iu6, Irxiu6);  // ../RTL/cortexm0ds_logic.v(8585)
  and u8786 (R2phu6, E7giu6, Prxiu6);  // ../RTL/cortexm0ds_logic.v(8586)
  and u8787 (n2261, Wrxiu6, Dsxiu6);  // ../RTL/cortexm0ds_logic.v(8587)
  not u8788 (Prxiu6, n2261);  // ../RTL/cortexm0ds_logic.v(8587)
  and u8789 (n2262, Qudpw6, IRQ[12]);  // ../RTL/cortexm0ds_logic.v(8588)
  buf u879 (vis_r11_o[28], Uqipw6);  // ../RTL/cortexm0ds_logic.v(1874)
  not u8790 (Dsxiu6, n2262);  // ../RTL/cortexm0ds_logic.v(8588)
  and u8791 (Wrxiu6, Ksxiu6, X6giu6);  // ../RTL/cortexm0ds_logic.v(8589)
  and u8792 (n2263, Kwfiu6, HWDATA[12]);  // ../RTL/cortexm0ds_logic.v(8590)
  not u8793 (X6giu6, n2263);  // ../RTL/cortexm0ds_logic.v(8590)
  and u8794 (n2264, Odgpw6[12], Rsxiu6);  // ../RTL/cortexm0ds_logic.v(8591)
  not u8795 (Ksxiu6, n2264);  // ../RTL/cortexm0ds_logic.v(8591)
  and u8796 (n2265, K66iu6, HWDATA[12]);  // ../RTL/cortexm0ds_logic.v(8592)
  not u8797 (Rsxiu6, n2265);  // ../RTL/cortexm0ds_logic.v(8592)
  or u8798 (E7giu6, Sb5iu6, Ysxiu6);  // ../RTL/cortexm0ds_logic.v(8593)
  and u8799 (K2phu6, A5giu6, Ftxiu6);  // ../RTL/cortexm0ds_logic.v(8594)
  buf u88 (Uthpw6[9], Mh1qw6);  // ../RTL/cortexm0ds_logic.v(1882)
  buf u880 (X3fpw6[1], Iixpw6);  // ../RTL/cortexm0ds_logic.v(1784)
  and u8800 (n2266, Mtxiu6, Ttxiu6);  // ../RTL/cortexm0ds_logic.v(8595)
  not u8801 (Ftxiu6, n2266);  // ../RTL/cortexm0ds_logic.v(8595)
  and u8802 (n2267, Vtdpw6, IRQ[13]);  // ../RTL/cortexm0ds_logic.v(8596)
  not u8803 (Ttxiu6, n2267);  // ../RTL/cortexm0ds_logic.v(8596)
  and u8804 (Mtxiu6, Auxiu6, T4giu6);  // ../RTL/cortexm0ds_logic.v(8597)
  and u8805 (n2268, Kwfiu6, HWDATA[13]);  // ../RTL/cortexm0ds_logic.v(8598)
  not u8806 (T4giu6, n2268);  // ../RTL/cortexm0ds_logic.v(8598)
  and u8807 (n2269, Odgpw6[13], Huxiu6);  // ../RTL/cortexm0ds_logic.v(8599)
  not u8808 (Auxiu6, n2269);  // ../RTL/cortexm0ds_logic.v(8599)
  and u8809 (n2270, K66iu6, HWDATA[13]);  // ../RTL/cortexm0ds_logic.v(8600)
  buf u881 (Vbgpw6[3], Owhbx6);  // ../RTL/cortexm0ds_logic.v(3092)
  not u8810 (Huxiu6, n2270);  // ../RTL/cortexm0ds_logic.v(8600)
  or u8811 (A5giu6, Sb5iu6, Ouxiu6);  // ../RTL/cortexm0ds_logic.v(8601)
  and u8812 (D2phu6, W2giu6, Vuxiu6);  // ../RTL/cortexm0ds_logic.v(8602)
  and u8813 (n2271, Cvxiu6, Jvxiu6);  // ../RTL/cortexm0ds_logic.v(8603)
  not u8814 (Vuxiu6, n2271);  // ../RTL/cortexm0ds_logic.v(8603)
  and u8815 (n2272, Otdpw6, IRQ[14]);  // ../RTL/cortexm0ds_logic.v(8604)
  not u8816 (Jvxiu6, n2272);  // ../RTL/cortexm0ds_logic.v(8604)
  and u8817 (Cvxiu6, Qvxiu6, P2giu6);  // ../RTL/cortexm0ds_logic.v(8605)
  and u8818 (n2273, Kwfiu6, HWDATA[14]);  // ../RTL/cortexm0ds_logic.v(8606)
  not u8819 (P2giu6, n2273);  // ../RTL/cortexm0ds_logic.v(8606)
  buf u882 (vis_r4_o[3], Acuax6);  // ../RTL/cortexm0ds_logic.v(2626)
  and u8820 (n2274, Odgpw6[14], Xvxiu6);  // ../RTL/cortexm0ds_logic.v(8607)
  not u8821 (Qvxiu6, n2274);  // ../RTL/cortexm0ds_logic.v(8607)
  and u8822 (n2275, K66iu6, HWDATA[14]);  // ../RTL/cortexm0ds_logic.v(8608)
  not u8823 (Xvxiu6, n2275);  // ../RTL/cortexm0ds_logic.v(8608)
  and u8824 (n2276, Clfiu6, R3giu6);  // ../RTL/cortexm0ds_logic.v(8609)
  not u8825 (W2giu6, n2276);  // ../RTL/cortexm0ds_logic.v(8609)
  and u8826 (W1phu6, S0giu6, Ewxiu6);  // ../RTL/cortexm0ds_logic.v(8610)
  and u8827 (n2277, Lwxiu6, Swxiu6);  // ../RTL/cortexm0ds_logic.v(8611)
  not u8828 (Ewxiu6, n2277);  // ../RTL/cortexm0ds_logic.v(8611)
  and u8829 (n2278, Lvdpw6, IRQ[15]);  // ../RTL/cortexm0ds_logic.v(8612)
  buf u883 (vis_r8_o[8], Ngsax6);  // ../RTL/cortexm0ds_logic.v(2579)
  not u8830 (Swxiu6, n2278);  // ../RTL/cortexm0ds_logic.v(8612)
  and u8831 (Lwxiu6, Zwxiu6, L0giu6);  // ../RTL/cortexm0ds_logic.v(8613)
  and u8832 (n2279, Fsdiu6, Kwfiu6);  // ../RTL/cortexm0ds_logic.v(8614)
  not u8833 (L0giu6, n2279);  // ../RTL/cortexm0ds_logic.v(8614)
  and u8834 (n2280, Odgpw6[15], Gxxiu6);  // ../RTL/cortexm0ds_logic.v(8615)
  not u8835 (Zwxiu6, n2280);  // ../RTL/cortexm0ds_logic.v(8615)
  and u8836 (n2281, Fsdiu6, K66iu6);  // ../RTL/cortexm0ds_logic.v(8616)
  not u8837 (Gxxiu6, n2281);  // ../RTL/cortexm0ds_logic.v(8616)
  and u8838 (Fsdiu6, Npdhu6, HWDATA[15]);  // ../RTL/cortexm0ds_logic.v(8617)
  or u8839 (S0giu6, Sb5iu6, Nxxiu6);  // ../RTL/cortexm0ds_logic.v(8618)
  buf u884 (B3gpw6[1], Uj4bx6);  // ../RTL/cortexm0ds_logic.v(2808)
  and u8840 (P1phu6, Mvhiu6, Uxxiu6);  // ../RTL/cortexm0ds_logic.v(8619)
  and u8841 (n2282, Byxiu6, Iyxiu6);  // ../RTL/cortexm0ds_logic.v(8620)
  not u8842 (Uxxiu6, n2282);  // ../RTL/cortexm0ds_logic.v(8620)
  and u8843 (n2283, Atdpw6, IRQ[16]);  // ../RTL/cortexm0ds_logic.v(8621)
  not u8844 (Iyxiu6, n2283);  // ../RTL/cortexm0ds_logic.v(8621)
  and u8845 (Byxiu6, Pyxiu6, Fvhiu6);  // ../RTL/cortexm0ds_logic.v(8622)
  and u8846 (n2284, Kwfiu6, HWDATA[16]);  // ../RTL/cortexm0ds_logic.v(8623)
  not u8847 (Fvhiu6, n2284);  // ../RTL/cortexm0ds_logic.v(8623)
  and u8848 (n2285, Odgpw6[16], Wyxiu6);  // ../RTL/cortexm0ds_logic.v(8624)
  not u8849 (Pyxiu6, n2285);  // ../RTL/cortexm0ds_logic.v(8624)
  buf u885 (vis_r9_o[4], Rjopw6);  // ../RTL/cortexm0ds_logic.v(1898)
  and u8850 (n2286, K66iu6, HWDATA[16]);  // ../RTL/cortexm0ds_logic.v(8625)
  not u8851 (Wyxiu6, n2286);  // ../RTL/cortexm0ds_logic.v(8625)
  and u8852 (n2287, Clfiu6, Hwhiu6);  // ../RTL/cortexm0ds_logic.v(8626)
  not u8853 (Mvhiu6, n2287);  // ../RTL/cortexm0ds_logic.v(8626)
  and u8854 (I1phu6, Npdiu6, Dzxiu6);  // ../RTL/cortexm0ds_logic.v(8627)
  and u8855 (n2288, Kzxiu6, Rzxiu6);  // ../RTL/cortexm0ds_logic.v(8628)
  not u8856 (Dzxiu6, n2288);  // ../RTL/cortexm0ds_logic.v(8628)
  and u8857 (n2289, Htdpw6, IRQ[17]);  // ../RTL/cortexm0ds_logic.v(8629)
  not u8858 (Rzxiu6, n2289);  // ../RTL/cortexm0ds_logic.v(8629)
  and u8859 (Kzxiu6, Yzxiu6, Gpdiu6);  // ../RTL/cortexm0ds_logic.v(8630)
  buf u886 (vis_r3_o[9], Dq6bx6);  // ../RTL/cortexm0ds_logic.v(2694)
  and u8860 (n2290, Kwfiu6, HWDATA[17]);  // ../RTL/cortexm0ds_logic.v(8631)
  not u8861 (Gpdiu6, n2290);  // ../RTL/cortexm0ds_logic.v(8631)
  and u8862 (n2291, Odgpw6[17], F0yiu6);  // ../RTL/cortexm0ds_logic.v(8632)
  not u8863 (Yzxiu6, n2291);  // ../RTL/cortexm0ds_logic.v(8632)
  and u8864 (n2292, K66iu6, HWDATA[17]);  // ../RTL/cortexm0ds_logic.v(8633)
  not u8865 (F0yiu6, n2292);  // ../RTL/cortexm0ds_logic.v(8633)
  or u8866 (Npdiu6, Sb5iu6, M0yiu6);  // ../RTL/cortexm0ds_logic.v(8634)
  and u8867 (B1phu6, Omdiu6, T0yiu6);  // ../RTL/cortexm0ds_logic.v(8635)
  and u8868 (n2293, A1yiu6, H1yiu6);  // ../RTL/cortexm0ds_logic.v(8636)
  not u8869 (T0yiu6, n2293);  // ../RTL/cortexm0ds_logic.v(8636)
  buf u887 (vis_msp_o[4], Vszpw6);  // ../RTL/cortexm0ds_logic.v(2097)
  and u8870 (n2294, Tsdpw6, IRQ[18]);  // ../RTL/cortexm0ds_logic.v(8637)
  not u8871 (H1yiu6, n2294);  // ../RTL/cortexm0ds_logic.v(8637)
  and u8872 (A1yiu6, O1yiu6, Hmdiu6);  // ../RTL/cortexm0ds_logic.v(8638)
  and u8873 (n2295, Kwfiu6, HWDATA[18]);  // ../RTL/cortexm0ds_logic.v(8639)
  not u8874 (Hmdiu6, n2295);  // ../RTL/cortexm0ds_logic.v(8639)
  and u8875 (n2296, Odgpw6[18], V1yiu6);  // ../RTL/cortexm0ds_logic.v(8640)
  not u8876 (O1yiu6, n2296);  // ../RTL/cortexm0ds_logic.v(8640)
  and u8877 (n2297, K66iu6, HWDATA[18]);  // ../RTL/cortexm0ds_logic.v(8641)
  not u8878 (V1yiu6, n2297);  // ../RTL/cortexm0ds_logic.v(8641)
  or u8879 (Omdiu6, Sb5iu6, C2yiu6);  // ../RTL/cortexm0ds_logic.v(8642)
  buf u888 (vis_r11_o[1], Qjypw6);  // ../RTL/cortexm0ds_logic.v(1874)
  and u8880 (U0phu6, Pjdiu6, J2yiu6);  // ../RTL/cortexm0ds_logic.v(8643)
  and u8881 (n2298, Q2yiu6, X2yiu6);  // ../RTL/cortexm0ds_logic.v(8644)
  not u8882 (J2yiu6, n2298);  // ../RTL/cortexm0ds_logic.v(8644)
  and u8883 (n2299, Msdpw6, IRQ[19]);  // ../RTL/cortexm0ds_logic.v(8645)
  not u8884 (X2yiu6, n2299);  // ../RTL/cortexm0ds_logic.v(8645)
  and u8885 (Q2yiu6, E3yiu6, Ijdiu6);  // ../RTL/cortexm0ds_logic.v(8646)
  and u8886 (n2300, Kwfiu6, HWDATA[19]);  // ../RTL/cortexm0ds_logic.v(8647)
  not u8887 (Ijdiu6, n2300);  // ../RTL/cortexm0ds_logic.v(8647)
  and u8888 (n2301, Odgpw6[19], L3yiu6);  // ../RTL/cortexm0ds_logic.v(8648)
  not u8889 (E3yiu6, n2301);  // ../RTL/cortexm0ds_logic.v(8648)
  buf u889 (vis_r11_o[27], Mjmpw6);  // ../RTL/cortexm0ds_logic.v(1874)
  and u8890 (n2302, K66iu6, HWDATA[19]);  // ../RTL/cortexm0ds_logic.v(8649)
  not u8891 (L3yiu6, n2302);  // ../RTL/cortexm0ds_logic.v(8649)
  or u8892 (Pjdiu6, Sb5iu6, S3yiu6);  // ../RTL/cortexm0ds_logic.v(8650)
  and u8893 (N0phu6, Qgdiu6, Z3yiu6);  // ../RTL/cortexm0ds_logic.v(8651)
  and u8894 (n2303, G4yiu6, N4yiu6);  // ../RTL/cortexm0ds_logic.v(8652)
  not u8895 (Z3yiu6, n2303);  // ../RTL/cortexm0ds_logic.v(8652)
  and u8896 (n2304, Yrdpw6, IRQ[20]);  // ../RTL/cortexm0ds_logic.v(8653)
  not u8897 (N4yiu6, n2304);  // ../RTL/cortexm0ds_logic.v(8653)
  and u8898 (G4yiu6, U4yiu6, Jgdiu6);  // ../RTL/cortexm0ds_logic.v(8654)
  and u8899 (n2305, Kwfiu6, HWDATA[20]);  // ../RTL/cortexm0ds_logic.v(8655)
  buf u89 (vis_r1_o[7], Dorpw6);  // ../RTL/cortexm0ds_logic.v(1876)
  or u890 (Qbfpw6[30], Dd5ju6, M75ju6);  // ../RTL/cortexm0ds_logic.v(9482)
  not u8900 (Jgdiu6, n2305);  // ../RTL/cortexm0ds_logic.v(8655)
  and u8901 (n2306, Odgpw6[20], B5yiu6);  // ../RTL/cortexm0ds_logic.v(8656)
  not u8902 (U4yiu6, n2306);  // ../RTL/cortexm0ds_logic.v(8656)
  and u8903 (n2307, K66iu6, HWDATA[20]);  // ../RTL/cortexm0ds_logic.v(8657)
  not u8904 (B5yiu6, n2307);  // ../RTL/cortexm0ds_logic.v(8657)
  or u8905 (Qgdiu6, Sb5iu6, I5yiu6);  // ../RTL/cortexm0ds_logic.v(8658)
  and u8906 (G0phu6, Rddiu6, P5yiu6);  // ../RTL/cortexm0ds_logic.v(8660)
  and u8907 (n2308, W5yiu6, D6yiu6);  // ../RTL/cortexm0ds_logic.v(8661)
  not u8908 (P5yiu6, n2308);  // ../RTL/cortexm0ds_logic.v(8661)
  and u8909 (n2309, Rrdpw6, IRQ[21]);  // ../RTL/cortexm0ds_logic.v(8662)
  buf u891 (Vbgpw6[2], L1bbx6);  // ../RTL/cortexm0ds_logic.v(3092)
  not u8910 (D6yiu6, n2309);  // ../RTL/cortexm0ds_logic.v(8662)
  and u8911 (W5yiu6, K6yiu6, Kddiu6);  // ../RTL/cortexm0ds_logic.v(8663)
  and u8912 (n2310, Kwfiu6, HWDATA[21]);  // ../RTL/cortexm0ds_logic.v(8664)
  not u8913 (Kddiu6, n2310);  // ../RTL/cortexm0ds_logic.v(8664)
  and u8914 (n2311, Odgpw6[21], R6yiu6);  // ../RTL/cortexm0ds_logic.v(8665)
  not u8915 (K6yiu6, n2311);  // ../RTL/cortexm0ds_logic.v(8665)
  and u8916 (n2312, K66iu6, HWDATA[21]);  // ../RTL/cortexm0ds_logic.v(8666)
  not u8917 (R6yiu6, n2312);  // ../RTL/cortexm0ds_logic.v(8666)
  or u8918 (Rddiu6, Sb5iu6, Y6yiu6);  // ../RTL/cortexm0ds_logic.v(8667)
  and u8919 (Zzohu6, Sadiu6, F7yiu6);  // ../RTL/cortexm0ds_logic.v(8668)
  buf u892 (vis_r4_o[2], D0uax6);  // ../RTL/cortexm0ds_logic.v(2626)
  and u8920 (n2313, M7yiu6, T7yiu6);  // ../RTL/cortexm0ds_logic.v(8669)
  not u8921 (F7yiu6, n2313);  // ../RTL/cortexm0ds_logic.v(8669)
  and u8922 (n2314, Xndpw6, IRQ[22]);  // ../RTL/cortexm0ds_logic.v(8670)
  not u8923 (T7yiu6, n2314);  // ../RTL/cortexm0ds_logic.v(8670)
  and u8924 (M7yiu6, A8yiu6, Ladiu6);  // ../RTL/cortexm0ds_logic.v(8671)
  and u8925 (n2315, Kwfiu6, HWDATA[22]);  // ../RTL/cortexm0ds_logic.v(8672)
  not u8926 (Ladiu6, n2315);  // ../RTL/cortexm0ds_logic.v(8672)
  and u8927 (n2316, Odgpw6[22], H8yiu6);  // ../RTL/cortexm0ds_logic.v(8673)
  not u8928 (A8yiu6, n2316);  // ../RTL/cortexm0ds_logic.v(8673)
  and u8929 (n2317, K66iu6, HWDATA[22]);  // ../RTL/cortexm0ds_logic.v(8674)
  buf u893 (vis_r8_o[7], Zvrpw6);  // ../RTL/cortexm0ds_logic.v(2579)
  not u8930 (H8yiu6, n2317);  // ../RTL/cortexm0ds_logic.v(8674)
  or u8931 (Sadiu6, Sb5iu6, O8yiu6);  // ../RTL/cortexm0ds_logic.v(8675)
  and u8932 (Szohu6, T7diu6, V8yiu6);  // ../RTL/cortexm0ds_logic.v(8676)
  and u8933 (n2318, C9yiu6, J9yiu6);  // ../RTL/cortexm0ds_logic.v(8677)
  not u8934 (V8yiu6, n2318);  // ../RTL/cortexm0ds_logic.v(8677)
  and u8935 (n2319, Drdpw6, IRQ[23]);  // ../RTL/cortexm0ds_logic.v(8678)
  not u8936 (J9yiu6, n2319);  // ../RTL/cortexm0ds_logic.v(8678)
  and u8937 (C9yiu6, Q9yiu6, M7diu6);  // ../RTL/cortexm0ds_logic.v(8679)
  and u8938 (n2320, Kwfiu6, HWDATA[23]);  // ../RTL/cortexm0ds_logic.v(8680)
  not u8939 (M7diu6, n2320);  // ../RTL/cortexm0ds_logic.v(8680)
  buf u894 (Aygpw6[4], Vibax6);  // ../RTL/cortexm0ds_logic.v(2278)
  and u8940 (n2321, Odgpw6[23], X9yiu6);  // ../RTL/cortexm0ds_logic.v(8681)
  not u8941 (Q9yiu6, n2321);  // ../RTL/cortexm0ds_logic.v(8681)
  and u8942 (n2322, K66iu6, HWDATA[23]);  // ../RTL/cortexm0ds_logic.v(8682)
  not u8943 (X9yiu6, n2322);  // ../RTL/cortexm0ds_logic.v(8682)
  or u8944 (T7diu6, Sb5iu6, Eayiu6);  // ../RTL/cortexm0ds_logic.v(8683)
  and u8945 (Lzohu6, Nufiu6, Layiu6);  // ../RTL/cortexm0ds_logic.v(8684)
  and u8946 (n2323, Sayiu6, Zayiu6);  // ../RTL/cortexm0ds_logic.v(8685)
  not u8947 (Layiu6, n2323);  // ../RTL/cortexm0ds_logic.v(8685)
  and u8948 (n2324, Pqdpw6, IRQ[26]);  // ../RTL/cortexm0ds_logic.v(8686)
  not u8949 (Zayiu6, n2324);  // ../RTL/cortexm0ds_logic.v(8686)
  not u895 (HPROT[3], n5200[1]);  // ../RTL/cortexm0ds_logic.v(15247)
  and u8950 (Sayiu6, Gbyiu6, Gufiu6);  // ../RTL/cortexm0ds_logic.v(8687)
  and u8951 (n2325, Kwfiu6, HWDATA[26]);  // ../RTL/cortexm0ds_logic.v(8688)
  not u8952 (Gufiu6, n2325);  // ../RTL/cortexm0ds_logic.v(8688)
  and u8953 (n2326, Odgpw6[26], Nbyiu6);  // ../RTL/cortexm0ds_logic.v(8689)
  not u8954 (Gbyiu6, n2326);  // ../RTL/cortexm0ds_logic.v(8689)
  and u8955 (n2327, K66iu6, HWDATA[26]);  // ../RTL/cortexm0ds_logic.v(8690)
  not u8956 (Nbyiu6, n2327);  // ../RTL/cortexm0ds_logic.v(8690)
  or u8957 (Nufiu6, Sb5iu6, Ubyiu6);  // ../RTL/cortexm0ds_logic.v(8691)
  and u8958 (Ezohu6, Jsfiu6, Bcyiu6);  // ../RTL/cortexm0ds_logic.v(8692)
  and u8959 (n2328, Icyiu6, Pcyiu6);  // ../RTL/cortexm0ds_logic.v(8693)
  buf u896 (vis_r0_o[1], Tdypw6);  // ../RTL/cortexm0ds_logic.v(1875)
  not u8960 (Bcyiu6, n2328);  // ../RTL/cortexm0ds_logic.v(8693)
  and u8961 (n2329, Iqdpw6, IRQ[27]);  // ../RTL/cortexm0ds_logic.v(8694)
  not u8962 (Pcyiu6, n2329);  // ../RTL/cortexm0ds_logic.v(8694)
  and u8963 (Icyiu6, Wcyiu6, Csfiu6);  // ../RTL/cortexm0ds_logic.v(8695)
  and u8964 (n2330, Kwfiu6, HWDATA[27]);  // ../RTL/cortexm0ds_logic.v(8696)
  not u8965 (Csfiu6, n2330);  // ../RTL/cortexm0ds_logic.v(8696)
  and u8966 (n2331, Odgpw6[27], Ddyiu6);  // ../RTL/cortexm0ds_logic.v(8697)
  not u8967 (Wcyiu6, n2331);  // ../RTL/cortexm0ds_logic.v(8697)
  and u8968 (n2332, K66iu6, HWDATA[27]);  // ../RTL/cortexm0ds_logic.v(8698)
  not u8969 (Ddyiu6, n2332);  // ../RTL/cortexm0ds_logic.v(8698)
  buf u897 (Tzfpw6[8], Ss0qw6);  // ../RTL/cortexm0ds_logic.v(2007)
  or u8970 (Jsfiu6, Sb5iu6, Kdyiu6);  // ../RTL/cortexm0ds_logic.v(8699)
  and u8971 (Xyohu6, Fqfiu6, Rdyiu6);  // ../RTL/cortexm0ds_logic.v(8700)
  and u8972 (n2333, Ydyiu6, Feyiu6);  // ../RTL/cortexm0ds_logic.v(8701)
  not u8973 (Rdyiu6, n2333);  // ../RTL/cortexm0ds_logic.v(8701)
  and u8974 (n2334, Bqdpw6, IRQ[28]);  // ../RTL/cortexm0ds_logic.v(8702)
  not u8975 (Feyiu6, n2334);  // ../RTL/cortexm0ds_logic.v(8702)
  and u8976 (Ydyiu6, Meyiu6, Ypfiu6);  // ../RTL/cortexm0ds_logic.v(8703)
  and u8977 (n2335, Kwfiu6, HWDATA[28]);  // ../RTL/cortexm0ds_logic.v(8704)
  not u8978 (Ypfiu6, n2335);  // ../RTL/cortexm0ds_logic.v(8704)
  and u8979 (n2336, Odgpw6[28], Teyiu6);  // ../RTL/cortexm0ds_logic.v(8705)
  buf u898 (Shhpw6[19], Cfvpw6);  // ../RTL/cortexm0ds_logic.v(1941)
  not u8980 (Meyiu6, n2336);  // ../RTL/cortexm0ds_logic.v(8705)
  and u8981 (n2337, K66iu6, HWDATA[28]);  // ../RTL/cortexm0ds_logic.v(8706)
  not u8982 (Teyiu6, n2337);  // ../RTL/cortexm0ds_logic.v(8706)
  or u8983 (Fqfiu6, Sb5iu6, Afyiu6);  // ../RTL/cortexm0ds_logic.v(8707)
  and u8984 (Qyohu6, Fgbiu6, Hfyiu6);  // ../RTL/cortexm0ds_logic.v(8708)
  and u8985 (n2338, Ofyiu6, Vfyiu6);  // ../RTL/cortexm0ds_logic.v(8709)
  not u8986 (Hfyiu6, n2338);  // ../RTL/cortexm0ds_logic.v(8709)
  and u8987 (n2339, Updpw6, IRQ[29]);  // ../RTL/cortexm0ds_logic.v(8710)
  not u8988 (Vfyiu6, n2339);  // ../RTL/cortexm0ds_logic.v(8710)
  and u8989 (Ofyiu6, Cgyiu6, Yfbiu6);  // ../RTL/cortexm0ds_logic.v(8711)
  buf u899 (vis_r12_o[21], Eetax6);  // ../RTL/cortexm0ds_logic.v(2599)
  and u8990 (n2340, Kwfiu6, HWDATA[29]);  // ../RTL/cortexm0ds_logic.v(8712)
  not u8991 (Yfbiu6, n2340);  // ../RTL/cortexm0ds_logic.v(8712)
  and u8992 (n2341, Odgpw6[29], Jgyiu6);  // ../RTL/cortexm0ds_logic.v(8713)
  not u8993 (Cgyiu6, n2341);  // ../RTL/cortexm0ds_logic.v(8713)
  and u8994 (n2342, K66iu6, HWDATA[29]);  // ../RTL/cortexm0ds_logic.v(8714)
  not u8995 (Jgyiu6, n2342);  // ../RTL/cortexm0ds_logic.v(8714)
  or u8996 (Fgbiu6, Sb5iu6, Qgyiu6);  // ../RTL/cortexm0ds_logic.v(8715)
  and u8997 (Jyohu6, Qxhiu6, Xgyiu6);  // ../RTL/cortexm0ds_logic.v(8716)
  and u8998 (n2343, Ehyiu6, Lhyiu6);  // ../RTL/cortexm0ds_logic.v(8717)
  not u8999 (Xgyiu6, n2343);  // ../RTL/cortexm0ds_logic.v(8717)
  buf u9 (WICENACK, 1'b0);  // ../RTL/cortexm0ds_logic.v(1732)
  buf u90 (vis_r0_o[27], E1npw6);  // ../RTL/cortexm0ds_logic.v(1875)
  buf u900 (vis_r9_o[3], Qpopw6);  // ../RTL/cortexm0ds_logic.v(1898)
  and u9000 (n2344, Zvdpw6, IRQ[30]);  // ../RTL/cortexm0ds_logic.v(8718)
  not u9001 (Lhyiu6, n2344);  // ../RTL/cortexm0ds_logic.v(8718)
  and u9002 (Ehyiu6, Shyiu6, Jxhiu6);  // ../RTL/cortexm0ds_logic.v(8719)
  and u9003 (n2345, Kwfiu6, HWDATA[30]);  // ../RTL/cortexm0ds_logic.v(8720)
  not u9004 (Jxhiu6, n2345);  // ../RTL/cortexm0ds_logic.v(8720)
  and u9005 (n2346, Odgpw6[30], Zhyiu6);  // ../RTL/cortexm0ds_logic.v(8721)
  not u9006 (Shyiu6, n2346);  // ../RTL/cortexm0ds_logic.v(8721)
  and u9007 (n2347, K66iu6, HWDATA[30]);  // ../RTL/cortexm0ds_logic.v(8722)
  not u9008 (Zhyiu6, n2347);  // ../RTL/cortexm0ds_logic.v(8722)
  or u9009 (Qxhiu6, Sb5iu6, Giyiu6);  // ../RTL/cortexm0ds_logic.v(8723)
  buf u901 (vis_r3_o[8], Cs6bx6);  // ../RTL/cortexm0ds_logic.v(2694)
  and u9010 (Cyohu6, Bebiu6, Niyiu6);  // ../RTL/cortexm0ds_logic.v(8724)
  and u9011 (n2348, Uiyiu6, Bjyiu6);  // ../RTL/cortexm0ds_logic.v(8725)
  not u9012 (Niyiu6, n2348);  // ../RTL/cortexm0ds_logic.v(8725)
  and u9013 (n2349, Npdpw6, IRQ[31]);  // ../RTL/cortexm0ds_logic.v(8726)
  not u9014 (Bjyiu6, n2349);  // ../RTL/cortexm0ds_logic.v(8726)
  and u9015 (Uiyiu6, Ijyiu6, Udbiu6);  // ../RTL/cortexm0ds_logic.v(8727)
  and u9016 (n2350, Kwfiu6, HWDATA[31]);  // ../RTL/cortexm0ds_logic.v(8728)
  not u9017 (Udbiu6, n2350);  // ../RTL/cortexm0ds_logic.v(8728)
  and u9018 (Kwfiu6, Pjyiu6, Yzciu6);  // ../RTL/cortexm0ds_logic.v(8729)
  and u9019 (Yzciu6, Wjyiu6, Npdhu6);  // ../RTL/cortexm0ds_logic.v(8730)
  buf u902 (vis_msp_o[3], Wqzpw6);  // ../RTL/cortexm0ds_logic.v(2097)
  and u9020 (n2351, Odgpw6[31], Dkyiu6);  // ../RTL/cortexm0ds_logic.v(8731)
  not u9021 (Ijyiu6, n2351);  // ../RTL/cortexm0ds_logic.v(8731)
  and u9022 (n2352, K66iu6, HWDATA[31]);  // ../RTL/cortexm0ds_logic.v(8732)
  not u9023 (Dkyiu6, n2352);  // ../RTL/cortexm0ds_logic.v(8732)
  and u9024 (K66iu6, Kkyiu6, D5eiu6);  // ../RTL/cortexm0ds_logic.v(8733)
  and u9025 (Kkyiu6, Pjyiu6, Npdhu6);  // ../RTL/cortexm0ds_logic.v(8734)
  and u9026 (n2353, Clfiu6, Webiu6);  // ../RTL/cortexm0ds_logic.v(8735)
  not u9027 (Bebiu6, n2353);  // ../RTL/cortexm0ds_logic.v(8735)
  and u9028 (Clfiu6, Rkyiu6, Ykyiu6);  // ../RTL/cortexm0ds_logic.v(8737)
  not u9029 (Sb5iu6, Clfiu6);  // ../RTL/cortexm0ds_logic.v(8737)
  buf u903 (vis_msp_o[29], Yizpw6);  // ../RTL/cortexm0ds_logic.v(2097)
  or u9030 (n2354, Xe8iu6, Ae0iu6);  // ../RTL/cortexm0ds_logic.v(8738)
  not u9031 (Ykyiu6, n2354);  // ../RTL/cortexm0ds_logic.v(8738)
  or u9032 (n2355, G7oiu6, Nloiu6);  // ../RTL/cortexm0ds_logic.v(8739)
  not u9033 (Rkyiu6, n2355);  // ../RTL/cortexm0ds_logic.v(8739)
  AL_MUX u9034 (
    .i0(Flyiu6),
    .i1(X3fpw6[3]),
    .sel(O25iu6),
    .o(Vxohu6));  // ../RTL/cortexm0ds_logic.v(8740)
  and u9035 (n2356, Mlyiu6, Tlyiu6);  // ../RTL/cortexm0ds_logic.v(8741)
  not u9036 (Flyiu6, n2356);  // ../RTL/cortexm0ds_logic.v(8741)
  and u9037 (Tlyiu6, Amyiu6, Hmyiu6);  // ../RTL/cortexm0ds_logic.v(8742)
  and u9038 (n2357, Omyiu6, S8fpw6[11]);  // ../RTL/cortexm0ds_logic.v(8743)
  not u9039 (Hmyiu6, n2357);  // ../RTL/cortexm0ds_logic.v(8743)
  buf u904 (vis_r11_o[26], Xztpw6);  // ../RTL/cortexm0ds_logic.v(1874)
  and u9040 (Amyiu6, Vmyiu6, Cnyiu6);  // ../RTL/cortexm0ds_logic.v(8744)
  and u9041 (n2358, Jnyiu6, D7fpw6[10]);  // ../RTL/cortexm0ds_logic.v(8745)
  not u9042 (Cnyiu6, n2358);  // ../RTL/cortexm0ds_logic.v(8745)
  and u9043 (Jnyiu6, D7fpw6[6], Qnyiu6);  // ../RTL/cortexm0ds_logic.v(8746)
  or u9044 (Qnyiu6, Xiiiu6, Mtjiu6);  // ../RTL/cortexm0ds_logic.v(8747)
  and u9045 (n2359, L45iu6, Xnyiu6);  // ../RTL/cortexm0ds_logic.v(8748)
  not u9046 (Vmyiu6, n2359);  // ../RTL/cortexm0ds_logic.v(8748)
  or u9047 (Xnyiu6, Eoyiu6, Loyiu6);  // ../RTL/cortexm0ds_logic.v(8749)
  and u9048 (Loyiu6, Soyiu6, N55iu6);  // ../RTL/cortexm0ds_logic.v(8750)
  or u9049 (n2360, K9aiu6, Zoyiu6);  // ../RTL/cortexm0ds_logic.v(8751)
  or u905 (Qbfpw6[29], N97ju6, M75ju6);  // ../RTL/cortexm0ds_logic.v(9482)
  not u9050 (Soyiu6, n2360);  // ../RTL/cortexm0ds_logic.v(8751)
  and u9051 (Mlyiu6, Gpyiu6, Npyiu6);  // ../RTL/cortexm0ds_logic.v(8752)
  and u9052 (n2361, A95iu6, D7fpw6[3]);  // ../RTL/cortexm0ds_logic.v(8753)
  not u9053 (Npyiu6, n2361);  // ../RTL/cortexm0ds_logic.v(8753)
  and u9054 (Oxohu6, Upyiu6, Bqyiu6);  // ../RTL/cortexm0ds_logic.v(8754)
  and u9055 (n2362, Iqyiu6, Pqyiu6);  // ../RTL/cortexm0ds_logic.v(8755)
  not u9056 (Bqyiu6, n2362);  // ../RTL/cortexm0ds_logic.v(8755)
  and u9057 (Pqyiu6, Wqyiu6, Dryiu6);  // ../RTL/cortexm0ds_logic.v(8756)
  and u9058 (Dryiu6, Kryiu6, Rryiu6);  // ../RTL/cortexm0ds_logic.v(8757)
  and u9059 (Rryiu6, Yryiu6, O4aiu6);  // ../RTL/cortexm0ds_logic.v(8758)
  buf u906 (Vbgpw6[1], Cxzax6);  // ../RTL/cortexm0ds_logic.v(3092)
  and u9060 (Kryiu6, Fsyiu6, Uloiu6);  // ../RTL/cortexm0ds_logic.v(8759)
  and u9061 (n2363, Msyiu6, Y0jiu6);  // ../RTL/cortexm0ds_logic.v(8760)
  not u9062 (Fsyiu6, n2363);  // ../RTL/cortexm0ds_logic.v(8760)
  or u9063 (n2364, Sijiu6, Cyfpw6[3]);  // ../RTL/cortexm0ds_logic.v(8761)
  not u9064 (Msyiu6, n2364);  // ../RTL/cortexm0ds_logic.v(8761)
  and u9065 (Wqyiu6, Tsyiu6, Atyiu6);  // ../RTL/cortexm0ds_logic.v(8762)
  and u9066 (n2365, Htyiu6, Otyiu6);  // ../RTL/cortexm0ds_logic.v(8763)
  not u9067 (Atyiu6, n2365);  // ../RTL/cortexm0ds_logic.v(8763)
  and u9068 (n2366, Vtyiu6, Cuyiu6);  // ../RTL/cortexm0ds_logic.v(8764)
  not u9069 (Otyiu6, n2366);  // ../RTL/cortexm0ds_logic.v(8764)
  buf u907 (vis_r4_o[1], Wruax6);  // ../RTL/cortexm0ds_logic.v(2626)
  and u9070 (n2367, Juyiu6, Quyiu6);  // ../RTL/cortexm0ds_logic.v(8765)
  not u9071 (Cuyiu6, n2367);  // ../RTL/cortexm0ds_logic.v(8765)
  and u9072 (Juyiu6, Xuyiu6, A95iu6);  // ../RTL/cortexm0ds_logic.v(8766)
  or u9073 (n2368, Evyiu6, P0piu6);  // ../RTL/cortexm0ds_logic.v(8767)
  not u9074 (Vtyiu6, n2368);  // ../RTL/cortexm0ds_logic.v(8767)
  and u9075 (Tsyiu6, Lvyiu6, Svyiu6);  // ../RTL/cortexm0ds_logic.v(8768)
  and u9076 (n2369, Zvyiu6, Ae0iu6);  // ../RTL/cortexm0ds_logic.v(8769)
  not u9077 (Svyiu6, n2369);  // ../RTL/cortexm0ds_logic.v(8769)
  and u9078 (Zvyiu6, D6kiu6, Gwyiu6);  // ../RTL/cortexm0ds_logic.v(8770)
  and u9079 (n2370, W8aiu6, Nwyiu6);  // ../RTL/cortexm0ds_logic.v(8771)
  not u908 (Xndpw6, Vyfbx6);  // ../RTL/cortexm0ds_logic.v(3018)
  not u9080 (Lvyiu6, n2370);  // ../RTL/cortexm0ds_logic.v(8771)
  and u9081 (n2371, Uwyiu6, Bxyiu6);  // ../RTL/cortexm0ds_logic.v(8772)
  not u9082 (Nwyiu6, n2371);  // ../RTL/cortexm0ds_logic.v(8772)
  and u9083 (n2372, Ixyiu6, Cyfpw6[7]);  // ../RTL/cortexm0ds_logic.v(8773)
  not u9084 (Bxyiu6, n2372);  // ../RTL/cortexm0ds_logic.v(8773)
  and u9085 (Ixyiu6, Cyfpw6[5], Pxyiu6);  // ../RTL/cortexm0ds_logic.v(8774)
  or u9086 (Uwyiu6, Lkaiu6, Wxyiu6);  // ../RTL/cortexm0ds_logic.v(8775)
  and u9087 (Iqyiu6, Dyyiu6, Kyyiu6);  // ../RTL/cortexm0ds_logic.v(8776)
  and u9088 (Kyyiu6, Ryyiu6, Yyyiu6);  // ../RTL/cortexm0ds_logic.v(8777)
  and u9089 (Yyyiu6, Fzyiu6, Mzyiu6);  // ../RTL/cortexm0ds_logic.v(8778)
  buf u909 (Trgpw6[10], Oveax6);  // ../RTL/cortexm0ds_logic.v(2376)
  and u9090 (n2373, Tzyiu6, Geaiu6);  // ../RTL/cortexm0ds_logic.v(8779)
  not u9091 (Mzyiu6, n2373);  // ../RTL/cortexm0ds_logic.v(8779)
  and u9092 (n2374, A0ziu6, H0ziu6);  // ../RTL/cortexm0ds_logic.v(8780)
  not u9093 (Tzyiu6, n2374);  // ../RTL/cortexm0ds_logic.v(8780)
  and u9094 (H0ziu6, O0ziu6, V0ziu6);  // ../RTL/cortexm0ds_logic.v(8781)
  and u9095 (n2375, C1ziu6, J1ziu6);  // ../RTL/cortexm0ds_logic.v(8782)
  not u9096 (V0ziu6, n2375);  // ../RTL/cortexm0ds_logic.v(8782)
  or u9097 (n2376, Q1ziu6, X1ziu6);  // ../RTL/cortexm0ds_logic.v(8783)
  not u9098 (C1ziu6, n2376);  // ../RTL/cortexm0ds_logic.v(8783)
  and u9099 (O0ziu6, E2ziu6, Gjjiu6);  // ../RTL/cortexm0ds_logic.v(8784)
  buf u91 (Ikghu6, Mnmpw6);  // ../RTL/cortexm0ds_logic.v(1860)
  buf u910 (Gtgpw6[15], S2cax6);  // ../RTL/cortexm0ds_logic.v(2375)
  and u9100 (n2377, L2ziu6, S2ziu6);  // ../RTL/cortexm0ds_logic.v(8785)
  not u9101 (Gjjiu6, n2377);  // ../RTL/cortexm0ds_logic.v(8785)
  and u9102 (L2ziu6, L45iu6, K9aiu6);  // ../RTL/cortexm0ds_logic.v(8786)
  and u9103 (A0ziu6, Z2ziu6, G3ziu6);  // ../RTL/cortexm0ds_logic.v(8787)
  and u9104 (n2378, U4kiu6, N3ziu6);  // ../RTL/cortexm0ds_logic.v(8788)
  not u9105 (G3ziu6, n2378);  // ../RTL/cortexm0ds_logic.v(8788)
  and u9106 (n2379, D1piu6, Xzmiu6);  // ../RTL/cortexm0ds_logic.v(8789)
  not u9107 (Z2ziu6, n2379);  // ../RTL/cortexm0ds_logic.v(8789)
  and u9108 (n2380, Imaiu6, U3ziu6);  // ../RTL/cortexm0ds_logic.v(8790)
  not u9109 (Fzyiu6, n2380);  // ../RTL/cortexm0ds_logic.v(8790)
  buf u911 (Jshpw6[15], Ad7ax6);  // ../RTL/cortexm0ds_logic.v(2372)
  and u9110 (n2381, B4ziu6, I4ziu6);  // ../RTL/cortexm0ds_logic.v(8791)
  not u9111 (U3ziu6, n2381);  // ../RTL/cortexm0ds_logic.v(8791)
  and u9112 (n2382, W0piu6, P4ziu6);  // ../RTL/cortexm0ds_logic.v(8792)
  not u9113 (I4ziu6, n2382);  // ../RTL/cortexm0ds_logic.v(8792)
  and u9114 (n2383, W4ziu6, D5ziu6);  // ../RTL/cortexm0ds_logic.v(8793)
  not u9115 (P4ziu6, n2383);  // ../RTL/cortexm0ds_logic.v(8793)
  and u9116 (n2384, K5ziu6, R5ziu6);  // ../RTL/cortexm0ds_logic.v(8794)
  not u9117 (D5ziu6, n2384);  // ../RTL/cortexm0ds_logic.v(8794)
  xor u9118 (n2385, Ndiiu6, Y5ziu6);  // ../RTL/cortexm0ds_logic.v(8795)
  not u9119 (R5ziu6, n2385);  // ../RTL/cortexm0ds_logic.v(8795)
  not u912 (Tugpw6[11], Iu9iu6);  // ../RTL/cortexm0ds_logic.v(16030)
  or u9120 (n2386, F6ziu6, D7fpw6[13]);  // ../RTL/cortexm0ds_logic.v(8796)
  not u9121 (K5ziu6, n2386);  // ../RTL/cortexm0ds_logic.v(8796)
  and u9122 (n2387, M6ziu6, X1ziu6);  // ../RTL/cortexm0ds_logic.v(8797)
  not u9123 (W4ziu6, n2387);  // ../RTL/cortexm0ds_logic.v(8797)
  and u9124 (n2388, T6ziu6, A7ziu6);  // ../RTL/cortexm0ds_logic.v(8798)
  not u9125 (M6ziu6, n2388);  // ../RTL/cortexm0ds_logic.v(8798)
  and u9126 (A7ziu6, H7ziu6, O7ziu6);  // ../RTL/cortexm0ds_logic.v(8799)
  and u9127 (n2389, V7ziu6, C8ziu6);  // ../RTL/cortexm0ds_logic.v(8800)
  not u9128 (H7ziu6, n2389);  // ../RTL/cortexm0ds_logic.v(8800)
  or u9129 (n2390, I6jiu6, D7fpw6[4]);  // ../RTL/cortexm0ds_logic.v(8801)
  buf u913 (Jshpw6[22], Bvfbx6);  // ../RTL/cortexm0ds_logic.v(2372)
  not u9130 (C8ziu6, n2390);  // ../RTL/cortexm0ds_logic.v(8801)
  and u9131 (V7ziu6, J8ziu6, D7fpw6[11]);  // ../RTL/cortexm0ds_logic.v(8802)
  and u9132 (T6ziu6, D7fpw6[13], Q8ziu6);  // ../RTL/cortexm0ds_logic.v(8803)
  and u9133 (n2391, X8ziu6, Tniiu6);  // ../RTL/cortexm0ds_logic.v(8804)
  not u9134 (Q8ziu6, n2391);  // ../RTL/cortexm0ds_logic.v(8804)
  and u9135 (n2392, E9ziu6, Q5aiu6);  // ../RTL/cortexm0ds_logic.v(8805)
  not u9136 (B4ziu6, n2392);  // ../RTL/cortexm0ds_logic.v(8805)
  and u9137 (n2393, L9ziu6, S9ziu6);  // ../RTL/cortexm0ds_logic.v(8806)
  not u9138 (E9ziu6, n2393);  // ../RTL/cortexm0ds_logic.v(8806)
  and u9139 (n2394, Jiiiu6, Z9ziu6);  // ../RTL/cortexm0ds_logic.v(8807)
  buf u914 (Uthpw6[24], Nrkpw6);  // ../RTL/cortexm0ds_logic.v(1882)
  not u9140 (S9ziu6, n2394);  // ../RTL/cortexm0ds_logic.v(8807)
  and u9141 (n2395, Gaziu6, Naziu6);  // ../RTL/cortexm0ds_logic.v(8808)
  not u9142 (Z9ziu6, n2395);  // ../RTL/cortexm0ds_logic.v(8808)
  or u9143 (Naziu6, Oviiu6, Gkiiu6);  // ../RTL/cortexm0ds_logic.v(8809)
  and u9144 (n2396, Dmiiu6, Uaziu6);  // ../RTL/cortexm0ds_logic.v(8810)
  not u9145 (L9ziu6, n2396);  // ../RTL/cortexm0ds_logic.v(8810)
  and u9146 (n2397, Bbziu6, Ibziu6);  // ../RTL/cortexm0ds_logic.v(8811)
  not u9147 (Uaziu6, n2397);  // ../RTL/cortexm0ds_logic.v(8811)
  or u9148 (n2398, D7fpw6[10], D7fpw6[12]);  // ../RTL/cortexm0ds_logic.v(8812)
  not u9149 (Ibziu6, n2398);  // ../RTL/cortexm0ds_logic.v(8812)
  buf u915 (Akgpw6[28], Eagax6);  // ../RTL/cortexm0ds_logic.v(2370)
  and u9150 (Bbziu6, Pbziu6, Wbziu6);  // ../RTL/cortexm0ds_logic.v(8813)
  xor u9151 (n2399, Dcziu6, D7fpw6[9]);  // ../RTL/cortexm0ds_logic.v(8814)
  not u9152 (Wbziu6, n2399);  // ../RTL/cortexm0ds_logic.v(8814)
  AL_MUX u9153 (
    .i0(Kcziu6),
    .i1(D7fpw6[7]),
    .sel(Ndiiu6),
    .o(Pbziu6));  // ../RTL/cortexm0ds_logic.v(8815)
  and u9154 (Ryyiu6, Rcziu6, Ycziu6);  // ../RTL/cortexm0ds_logic.v(8816)
  or u9155 (Ycziu6, E45iu6, Wthiu6);  // ../RTL/cortexm0ds_logic.v(8817)
  and u9156 (Dyyiu6, Fdziu6, Mdziu6);  // ../RTL/cortexm0ds_logic.v(8818)
  AL_MUX u9157 (
    .i0(Tdziu6),
    .i1(Aeziu6),
    .sel(D7fpw6[14]),
    .o(Mdziu6));  // ../RTL/cortexm0ds_logic.v(8819)
  and u9158 (n2400, Heziu6, Nriiu6);  // ../RTL/cortexm0ds_logic.v(8820)
  not u9159 (Aeziu6, n2400);  // ../RTL/cortexm0ds_logic.v(8820)
  buf u916 (Togpw6[8], Y5dax6);  // ../RTL/cortexm0ds_logic.v(2378)
  and u9160 (Heziu6, Aujiu6, K9aiu6);  // ../RTL/cortexm0ds_logic.v(8821)
  and u9161 (Fdziu6, Oeziu6, Veziu6);  // ../RTL/cortexm0ds_logic.v(8822)
  or u9162 (Upyiu6, H6ghu6, HREADY);  // ../RTL/cortexm0ds_logic.v(8823)
  and u9163 (n2401, Cfziu6, Jfziu6);  // ../RTL/cortexm0ds_logic.v(8824)
  not u9164 (Hxohu6, n2401);  // ../RTL/cortexm0ds_logic.v(8824)
  and u9165 (Jfziu6, Qfziu6, Xfziu6);  // ../RTL/cortexm0ds_logic.v(8825)
  and u9166 (n2402, Egziu6, Eafpw6[29]);  // ../RTL/cortexm0ds_logic.v(8826)
  not u9167 (Xfziu6, n2402);  // ../RTL/cortexm0ds_logic.v(8826)
  and u9168 (Qfziu6, Lgziu6, Sgziu6);  // ../RTL/cortexm0ds_logic.v(8827)
  and u9169 (n2403, Zgziu6, Fj8iu6);  // ../RTL/cortexm0ds_logic.v(8828)
  buf u917 (Togpw6[16], Owcax6);  // ../RTL/cortexm0ds_logic.v(2378)
  not u9170 (Lgziu6, n2403);  // ../RTL/cortexm0ds_logic.v(8828)
  and u9171 (n2404, Ghziu6, Nhziu6);  // ../RTL/cortexm0ds_logic.v(8829)
  not u9172 (Fj8iu6, n2404);  // ../RTL/cortexm0ds_logic.v(8829)
  and u9173 (Nhziu6, Uhziu6, Biziu6);  // ../RTL/cortexm0ds_logic.v(8830)
  or u9174 (Biziu6, Iiziu6, Piziu6);  // ../RTL/cortexm0ds_logic.v(8831)
  and u9175 (Uhziu6, Wiziu6, Djziu6);  // ../RTL/cortexm0ds_logic.v(8832)
  or u9176 (Wiziu6, Kjziu6, Rjziu6);  // ../RTL/cortexm0ds_logic.v(8833)
  and u9177 (Ghziu6, Yjziu6, Fkziu6);  // ../RTL/cortexm0ds_logic.v(8834)
  or u9178 (Fkziu6, Mkziu6, Tkziu6);  // ../RTL/cortexm0ds_logic.v(8835)
  or u9179 (Yjziu6, Alziu6, Hlziu6);  // ../RTL/cortexm0ds_logic.v(8836)
  buf u918 (Togpw6[24], Xqcax6);  // ../RTL/cortexm0ds_logic.v(2378)
  and u9180 (Cfziu6, Olziu6, Vlziu6);  // ../RTL/cortexm0ds_logic.v(8837)
  and u9181 (n2405, Zsfpw6[28], Cmziu6);  // ../RTL/cortexm0ds_logic.v(8838)
  not u9182 (Vlziu6, n2405);  // ../RTL/cortexm0ds_logic.v(8838)
  and u9183 (n2406, vis_pc_o[28], Jmziu6);  // ../RTL/cortexm0ds_logic.v(8839)
  not u9184 (Olziu6, n2406);  // ../RTL/cortexm0ds_logic.v(8839)
  not u9185 (Axohu6, Qmziu6);  // ../RTL/cortexm0ds_logic.v(8840)
  AL_MUX u9186 (
    .i0(Tfjiu6),
    .i1(Xmziu6),
    .sel(HREADY),
    .o(Qmziu6));  // ../RTL/cortexm0ds_logic.v(8841)
  and u9187 (Xmziu6, Enziu6, Lnziu6);  // ../RTL/cortexm0ds_logic.v(8842)
  and u9188 (Lnziu6, Snziu6, Znziu6);  // ../RTL/cortexm0ds_logic.v(8843)
  and u9189 (Znziu6, Goziu6, Noziu6);  // ../RTL/cortexm0ds_logic.v(8844)
  buf u919 (X8hpw6[2], Pe7ax6);  // ../RTL/cortexm0ds_logic.v(2046)
  or u9190 (n2407, Bi0iu6, Uoziu6);  // ../RTL/cortexm0ds_logic.v(8845)
  not u9191 (Noziu6, n2407);  // ../RTL/cortexm0ds_logic.v(8845)
  and u9192 (Goziu6, Bpziu6, Oaiiu6);  // ../RTL/cortexm0ds_logic.v(8846)
  and u9193 (n2408, Ipziu6, Qe8iu6);  // ../RTL/cortexm0ds_logic.v(8847)
  not u9194 (Bpziu6, n2408);  // ../RTL/cortexm0ds_logic.v(8847)
  and u9195 (Snziu6, Ppziu6, Wpziu6);  // ../RTL/cortexm0ds_logic.v(8848)
  and u9196 (n2409, Neoiu6, Dqziu6);  // ../RTL/cortexm0ds_logic.v(8849)
  not u9197 (Wpziu6, n2409);  // ../RTL/cortexm0ds_logic.v(8849)
  and u9198 (n2410, Kqziu6, Rqziu6);  // ../RTL/cortexm0ds_logic.v(8850)
  not u9199 (Dqziu6, n2410);  // ../RTL/cortexm0ds_logic.v(8850)
  buf u92 (K7hpw6[17], Qjbbx6);  // ../RTL/cortexm0ds_logic.v(2366)
  buf u920 (Jshpw6[7], Nd3qw6);  // ../RTL/cortexm0ds_logic.v(2372)
  and u9200 (n2411, Yqziu6, D1piu6);  // ../RTL/cortexm0ds_logic.v(8851)
  not u9201 (Rqziu6, n2411);  // ../RTL/cortexm0ds_logic.v(8851)
  and u9202 (Yqziu6, Frziu6, Cyfpw6[5]);  // ../RTL/cortexm0ds_logic.v(8852)
  and u9203 (Kqziu6, Ntgiu6, E4jiu6);  // ../RTL/cortexm0ds_logic.v(8853)
  and u9204 (Ppziu6, Mrziu6, Trziu6);  // ../RTL/cortexm0ds_logic.v(8854)
  and u9205 (n2412, Asziu6, Uriiu6);  // ../RTL/cortexm0ds_logic.v(8855)
  not u9206 (Trziu6, n2412);  // ../RTL/cortexm0ds_logic.v(8855)
  and u9207 (n2413, Hsziu6, Osziu6);  // ../RTL/cortexm0ds_logic.v(8856)
  not u9208 (Asziu6, n2413);  // ../RTL/cortexm0ds_logic.v(8856)
  and u9209 (n2414, Vsziu6, Ia8iu6);  // ../RTL/cortexm0ds_logic.v(8857)
  buf u921 (Jshpw6[21], Ufebx6);  // ../RTL/cortexm0ds_logic.v(2372)
  not u9210 (Osziu6, n2414);  // ../RTL/cortexm0ds_logic.v(8857)
  or u9211 (n2415, E4jiu6, Cyfpw6[3]);  // ../RTL/cortexm0ds_logic.v(8858)
  not u9212 (Vsziu6, n2415);  // ../RTL/cortexm0ds_logic.v(8858)
  or u9213 (Hsziu6, Ctziu6, Tfjiu6);  // ../RTL/cortexm0ds_logic.v(8859)
  or u9214 (Mrziu6, Ctziu6, As0iu6);  // ../RTL/cortexm0ds_logic.v(8860)
  and u9215 (Enziu6, Jtziu6, Qtziu6);  // ../RTL/cortexm0ds_logic.v(8861)
  and u9216 (Qtziu6, Xtziu6, Euziu6);  // ../RTL/cortexm0ds_logic.v(8862)
  and u9217 (Euziu6, Luziu6, Suziu6);  // ../RTL/cortexm0ds_logic.v(8863)
  and u9218 (n2416, Cyfpw6[7], Zuziu6);  // ../RTL/cortexm0ds_logic.v(8864)
  not u9219 (Suziu6, n2416);  // ../RTL/cortexm0ds_logic.v(8864)
  buf u922 (vis_r8_o[6], W9spw6);  // ../RTL/cortexm0ds_logic.v(2579)
  and u9220 (n2417, Gvziu6, Nvziu6);  // ../RTL/cortexm0ds_logic.v(8865)
  not u9221 (Zuziu6, n2417);  // ../RTL/cortexm0ds_logic.v(8865)
  or u9222 (Nvziu6, Q5aiu6, Uvziu6);  // ../RTL/cortexm0ds_logic.v(8866)
  and u9223 (Gvziu6, Bwziu6, Iwziu6);  // ../RTL/cortexm0ds_logic.v(8867)
  and u9224 (n2418, Pwziu6, Wwziu6);  // ../RTL/cortexm0ds_logic.v(8868)
  not u9225 (Iwziu6, n2418);  // ../RTL/cortexm0ds_logic.v(8868)
  or u9226 (n2419, Dxziu6, Cyfpw6[0]);  // ../RTL/cortexm0ds_logic.v(8869)
  not u9227 (Pwziu6, n2419);  // ../RTL/cortexm0ds_logic.v(8869)
  or u9228 (Bwziu6, Jojiu6, Ii0iu6);  // ../RTL/cortexm0ds_logic.v(8870)
  and u9229 (n2420, Kxziu6, Rxziu6);  // ../RTL/cortexm0ds_logic.v(8871)
  buf u923 (Aygpw6[3], Zgbax6);  // ../RTL/cortexm0ds_logic.v(2278)
  not u9230 (Luziu6, n2420);  // ../RTL/cortexm0ds_logic.v(8871)
  and u9231 (n2421, Yxziu6, Fyziu6);  // ../RTL/cortexm0ds_logic.v(8872)
  not u9232 (Rxziu6, n2421);  // ../RTL/cortexm0ds_logic.v(8872)
  and u9233 (Fyziu6, Myziu6, Tyziu6);  // ../RTL/cortexm0ds_logic.v(8873)
  and u9234 (n2422, Azziu6, Hzziu6);  // ../RTL/cortexm0ds_logic.v(8874)
  not u9235 (Tyziu6, n2422);  // ../RTL/cortexm0ds_logic.v(8874)
  or u9236 (n2423, Tfjiu6, D7fpw6[15]);  // ../RTL/cortexm0ds_logic.v(8875)
  not u9237 (Azziu6, n2423);  // ../RTL/cortexm0ds_logic.v(8875)
  or u9238 (n2424, P0piu6, Ozziu6);  // ../RTL/cortexm0ds_logic.v(8876)
  not u9239 (Myziu6, n2424);  // ../RTL/cortexm0ds_logic.v(8876)
  buf u924 (vis_r9_o[2], Yftpw6);  // ../RTL/cortexm0ds_logic.v(1898)
  and u9240 (Yxziu6, X3jiu6, Vzziu6);  // ../RTL/cortexm0ds_logic.v(8877)
  and u9241 (n2425, U0aiu6, D7fpw6[3]);  // ../RTL/cortexm0ds_logic.v(8878)
  not u9242 (Vzziu6, n2425);  // ../RTL/cortexm0ds_logic.v(8878)
  or u9243 (X3jiu6, Jjhiu6, Uriiu6);  // ../RTL/cortexm0ds_logic.v(8879)
  and u9244 (Xtziu6, Fniiu6, C00ju6);  // ../RTL/cortexm0ds_logic.v(8880)
  and u9245 (n2426, J00ju6, Zraiu6);  // ../RTL/cortexm0ds_logic.v(8881)
  not u9246 (C00ju6, n2426);  // ../RTL/cortexm0ds_logic.v(8881)
  and u9247 (n2427, Q00ju6, X00ju6);  // ../RTL/cortexm0ds_logic.v(8882)
  not u9248 (J00ju6, n2427);  // ../RTL/cortexm0ds_logic.v(8882)
  and u9249 (X00ju6, E10ju6, L10ju6);  // ../RTL/cortexm0ds_logic.v(8883)
  buf u925 (vis_r3_o[7], Og5bx6);  // ../RTL/cortexm0ds_logic.v(2694)
  and u9250 (L10ju6, S10ju6, Z10ju6);  // ../RTL/cortexm0ds_logic.v(8884)
  and u9251 (n2428, G20ju6, N20ju6);  // ../RTL/cortexm0ds_logic.v(8885)
  not u9252 (Z10ju6, n2428);  // ../RTL/cortexm0ds_logic.v(8885)
  or u9253 (n2429, Nsaiu6, Xe8iu6);  // ../RTL/cortexm0ds_logic.v(8886)
  not u9254 (G20ju6, n2429);  // ../RTL/cortexm0ds_logic.v(8886)
  and u9255 (S10ju6, U20ju6, W8oiu6);  // ../RTL/cortexm0ds_logic.v(8887)
  and u9256 (n2430, B30ju6, Mmjiu6);  // ../RTL/cortexm0ds_logic.v(8888)
  not u9257 (U20ju6, n2430);  // ../RTL/cortexm0ds_logic.v(8888)
  and u9258 (B30ju6, I30ju6, Gwyiu6);  // ../RTL/cortexm0ds_logic.v(8889)
  and u9259 (E10ju6, P30ju6, W30ju6);  // ../RTL/cortexm0ds_logic.v(8890)
  buf u926 (vis_msp_o[2], Ymzpw6);  // ../RTL/cortexm0ds_logic.v(2097)
  and u9260 (n2431, Hzziu6, D40ju6);  // ../RTL/cortexm0ds_logic.v(8891)
  not u9261 (W30ju6, n2431);  // ../RTL/cortexm0ds_logic.v(8891)
  and u9262 (n2432, K40ju6, R40ju6);  // ../RTL/cortexm0ds_logic.v(8892)
  not u9263 (D40ju6, n2432);  // ../RTL/cortexm0ds_logic.v(8892)
  and u9264 (n2433, Y40ju6, Ii0iu6);  // ../RTL/cortexm0ds_logic.v(8893)
  not u9265 (R40ju6, n2433);  // ../RTL/cortexm0ds_logic.v(8893)
  and u9266 (K40ju6, F50ju6, Xe8iu6);  // ../RTL/cortexm0ds_logic.v(8894)
  and u9267 (n2434, M50ju6, V9ghu6);  // ../RTL/cortexm0ds_logic.v(8895)
  not u9268 (F50ju6, n2434);  // ../RTL/cortexm0ds_logic.v(8895)
  or u9269 (n2435, P0biu6, Cyfpw6[6]);  // ../RTL/cortexm0ds_logic.v(8896)
  buf u927 (vis_msp_o[28], Ykzpw6);  // ../RTL/cortexm0ds_logic.v(2097)
  not u9270 (M50ju6, n2435);  // ../RTL/cortexm0ds_logic.v(8896)
  and u9271 (P30ju6, T50ju6, A60ju6);  // ../RTL/cortexm0ds_logic.v(8897)
  and u9272 (n2436, Omyiu6, H60ju6);  // ../RTL/cortexm0ds_logic.v(8898)
  not u9273 (A60ju6, n2436);  // ../RTL/cortexm0ds_logic.v(8898)
  and u9274 (n2437, O60ju6, V60ju6);  // ../RTL/cortexm0ds_logic.v(8899)
  not u9275 (H60ju6, n2437);  // ../RTL/cortexm0ds_logic.v(8899)
  and u9276 (n2438, Wp0iu6, Qyniu6);  // ../RTL/cortexm0ds_logic.v(8900)
  not u9277 (V60ju6, n2438);  // ../RTL/cortexm0ds_logic.v(8900)
  and u9278 (n2439, Yljiu6, C70ju6);  // ../RTL/cortexm0ds_logic.v(8901)
  not u9279 (T50ju6, n2439);  // ../RTL/cortexm0ds_logic.v(8901)
  buf u928 (vis_r11_o[25], Z7tpw6);  // ../RTL/cortexm0ds_logic.v(1874)
  and u9280 (n2440, Cyfpw6[7], J70ju6);  // ../RTL/cortexm0ds_logic.v(8902)
  not u9281 (C70ju6, n2440);  // ../RTL/cortexm0ds_logic.v(8902)
  or u9282 (J70ju6, As0iu6, Dxziu6);  // ../RTL/cortexm0ds_logic.v(8903)
  and u9283 (Q00ju6, Q70ju6, X70ju6);  // ../RTL/cortexm0ds_logic.v(8904)
  and u9284 (X70ju6, E80ju6, L80ju6);  // ../RTL/cortexm0ds_logic.v(8905)
  or u9285 (L80ju6, S80ju6, Ftjiu6);  // ../RTL/cortexm0ds_logic.v(8906)
  and u9286 (E80ju6, Z80ju6, G90ju6);  // ../RTL/cortexm0ds_logic.v(8907)
  and u9287 (n2441, N90ju6, Uriiu6);  // ../RTL/cortexm0ds_logic.v(8908)
  not u9288 (G90ju6, n2441);  // ../RTL/cortexm0ds_logic.v(8908)
  and u9289 (n2442, U90ju6, Ba0ju6);  // ../RTL/cortexm0ds_logic.v(8909)
  or u929 (Qbfpw6[28], Nn7ju6, M75ju6);  // ../RTL/cortexm0ds_logic.v(9482)
  not u9290 (N90ju6, n2442);  // ../RTL/cortexm0ds_logic.v(8909)
  and u9291 (Ba0ju6, Ia0ju6, Pa0ju6);  // ../RTL/cortexm0ds_logic.v(8910)
  and u9292 (n2443, Wa0ju6, Db0ju6);  // ../RTL/cortexm0ds_logic.v(8911)
  not u9293 (Pa0ju6, n2443);  // ../RTL/cortexm0ds_logic.v(8911)
  and u9294 (Wa0ju6, Nbkiu6, Oviiu6);  // ../RTL/cortexm0ds_logic.v(8912)
  and u9295 (Ia0ju6, Kb0ju6, Rb0ju6);  // ../RTL/cortexm0ds_logic.v(8913)
  and u9296 (U90ju6, Yb0ju6, Fc0ju6);  // ../RTL/cortexm0ds_logic.v(8914)
  and u9297 (n2444, P0piu6, Mc0ju6);  // ../RTL/cortexm0ds_logic.v(8915)
  not u9298 (Fc0ju6, n2444);  // ../RTL/cortexm0ds_logic.v(8915)
  and u9299 (n2445, Tc0ju6, Ad0ju6);  // ../RTL/cortexm0ds_logic.v(8916)
  buf u93 (vis_r2_o[28], R7ibx6);  // ../RTL/cortexm0ds_logic.v(2551)
  buf u930 (vis_r4_o[31], B8uax6);  // ../RTL/cortexm0ds_logic.v(2626)
  not u9300 (Mc0ju6, n2445);  // ../RTL/cortexm0ds_logic.v(8916)
  and u9301 (Ad0ju6, Hd0ju6, Od0ju6);  // ../RTL/cortexm0ds_logic.v(8917)
  and u9302 (n2446, D7fpw6[8], Vd0ju6);  // ../RTL/cortexm0ds_logic.v(8918)
  not u9303 (Hd0ju6, n2446);  // ../RTL/cortexm0ds_logic.v(8918)
  or u9304 (Vd0ju6, U5jiu6, Dcziu6);  // ../RTL/cortexm0ds_logic.v(8919)
  and u9305 (Tc0ju6, Ce0ju6, Je0ju6);  // ../RTL/cortexm0ds_logic.v(8920)
  AL_MUX u9306 (
    .i0(Qe0ju6),
    .i1(Kcziu6),
    .sel(I6jiu6),
    .o(Ce0ju6));  // ../RTL/cortexm0ds_logic.v(8921)
  or u9307 (Yb0ju6, Xe0ju6, H95iu6);  // ../RTL/cortexm0ds_logic.v(8922)
  and u9308 (n2447, J9kiu6, Ef0ju6);  // ../RTL/cortexm0ds_logic.v(8923)
  not u9309 (Z80ju6, n2447);  // ../RTL/cortexm0ds_logic.v(8923)
  buf u931 (K7hpw6[4], Tt9ax6);  // ../RTL/cortexm0ds_logic.v(2366)
  and u9310 (n2448, Lf0ju6, Sf0ju6);  // ../RTL/cortexm0ds_logic.v(8924)
  not u9311 (Ef0ju6, n2448);  // ../RTL/cortexm0ds_logic.v(8924)
  and u9312 (Sf0ju6, Zf0ju6, Gg0ju6);  // ../RTL/cortexm0ds_logic.v(8925)
  and u9313 (n2449, Ng0ju6, Oviiu6);  // ../RTL/cortexm0ds_logic.v(8926)
  not u9314 (Gg0ju6, n2449);  // ../RTL/cortexm0ds_logic.v(8926)
  and u9315 (n2450, I6jiu6, Je0ju6);  // ../RTL/cortexm0ds_logic.v(8927)
  not u9316 (Ng0ju6, n2450);  // ../RTL/cortexm0ds_logic.v(8927)
  or u9317 (Je0ju6, O95iu6, D7fpw6[9]);  // ../RTL/cortexm0ds_logic.v(8928)
  and u9318 (n2451, D7fpw6[13], Ug0ju6);  // ../RTL/cortexm0ds_logic.v(8929)
  not u9319 (Zf0ju6, n2451);  // ../RTL/cortexm0ds_logic.v(8929)
  buf u932 (vis_r14_o[27], Njnax6);  // ../RTL/cortexm0ds_logic.v(2497)
  and u9320 (n2452, Bh0ju6, Ih0ju6);  // ../RTL/cortexm0ds_logic.v(8930)
  not u9321 (Ug0ju6, n2452);  // ../RTL/cortexm0ds_logic.v(8930)
  or u9322 (Ih0ju6, Ph0ju6, D7fpw6[4]);  // ../RTL/cortexm0ds_logic.v(8931)
  or u9323 (Bh0ju6, Ndiiu6, Wh0ju6);  // ../RTL/cortexm0ds_logic.v(8932)
  and u9324 (Lf0ju6, Di0ju6, Ki0ju6);  // ../RTL/cortexm0ds_logic.v(8933)
  and u9325 (n2453, D7fpw6[12], Ri0ju6);  // ../RTL/cortexm0ds_logic.v(8934)
  not u9326 (Ki0ju6, n2453);  // ../RTL/cortexm0ds_logic.v(8934)
  and u9327 (n2454, Yi0ju6, Fj0ju6);  // ../RTL/cortexm0ds_logic.v(8935)
  not u9328 (Ri0ju6, n2454);  // ../RTL/cortexm0ds_logic.v(8935)
  and u9329 (Fj0ju6, Mj0ju6, Tj0ju6);  // ../RTL/cortexm0ds_logic.v(8936)
  buf u933 (vis_r3_o[1], Nq5bx6);  // ../RTL/cortexm0ds_logic.v(2694)
  and u9330 (n2455, Ak0ju6, Zwciu6);  // ../RTL/cortexm0ds_logic.v(8937)
  not u9331 (Tj0ju6, n2455);  // ../RTL/cortexm0ds_logic.v(8937)
  or u9332 (Mj0ju6, Hk0ju6, Oviiu6);  // ../RTL/cortexm0ds_logic.v(8938)
  and u9333 (Yi0ju6, Ok0ju6, Vk0ju6);  // ../RTL/cortexm0ds_logic.v(8939)
  or u9334 (Vk0ju6, Kcziu6, D7fpw6[10]);  // ../RTL/cortexm0ds_logic.v(8940)
  or u9335 (Ok0ju6, Ndiiu6, Qxoiu6);  // ../RTL/cortexm0ds_logic.v(8941)
  or u9336 (Di0ju6, Cl0ju6, D7fpw6[7]);  // ../RTL/cortexm0ds_logic.v(8942)
  not u9337 (Cl0ju6, Zroiu6);  // ../RTL/cortexm0ds_logic.v(8943)
  or u9338 (n2456, Jl0ju6, Ql0ju6);  // ../RTL/cortexm0ds_logic.v(8944)
  not u9339 (Q70ju6, n2456);  // ../RTL/cortexm0ds_logic.v(8944)
  buf u934 (Vbgpw6[24], Oxkpw6);  // ../RTL/cortexm0ds_logic.v(3092)
  or u9340 (n2457, Xl0ju6, D7fpw6[8]);  // ../RTL/cortexm0ds_logic.v(8945)
  not u9341 (Ql0ju6, n2457);  // ../RTL/cortexm0ds_logic.v(8945)
  AL_MUX u9342 (
    .i0(Em0ju6),
    .i1(Lraiu6),
    .sel(C0ehu6),
    .o(Jl0ju6));  // ../RTL/cortexm0ds_logic.v(8946)
  and u9343 (Em0ju6, Geoiu6, H4ghu6);  // ../RTL/cortexm0ds_logic.v(8947)
  or u9344 (Fniiu6, Hujiu6, D7fpw6[12]);  // ../RTL/cortexm0ds_logic.v(8948)
  and u9345 (Jtziu6, Lm0ju6, F85iu6);  // ../RTL/cortexm0ds_logic.v(8949)
  and u9346 (Lm0ju6, Sm0ju6, Zm0ju6);  // ../RTL/cortexm0ds_logic.v(8950)
  or u9347 (Zm0ju6, Wthiu6, Nloiu6);  // ../RTL/cortexm0ds_logic.v(8951)
  or u9348 (Sm0ju6, Taaiu6, Faaiu6);  // ../RTL/cortexm0ds_logic.v(8952)
  and u9349 (Twohu6, Gn0ju6, Nn0ju6);  // ../RTL/cortexm0ds_logic.v(8953)
  not u935 (Qndpw6, Eghbx6);  // ../RTL/cortexm0ds_logic.v(3045)
  and u9350 (n2458, Un0ju6, Bo0ju6);  // ../RTL/cortexm0ds_logic.v(8954)
  not u9351 (Nn0ju6, n2458);  // ../RTL/cortexm0ds_logic.v(8954)
  and u9352 (Bo0ju6, Io0ju6, Po0ju6);  // ../RTL/cortexm0ds_logic.v(8955)
  and u9353 (Po0ju6, Wo0ju6, Dp0ju6);  // ../RTL/cortexm0ds_logic.v(8956)
  and u9354 (Dp0ju6, Kp0ju6, Rp0ju6);  // ../RTL/cortexm0ds_logic.v(8957)
  and u9355 (n2459, J9kiu6, Yp0ju6);  // ../RTL/cortexm0ds_logic.v(8958)
  not u9356 (Rp0ju6, n2459);  // ../RTL/cortexm0ds_logic.v(8958)
  and u9357 (n2460, Fq0ju6, Mq0ju6);  // ../RTL/cortexm0ds_logic.v(8959)
  not u9358 (Yp0ju6, n2460);  // ../RTL/cortexm0ds_logic.v(8959)
  and u9359 (Mq0ju6, Tq0ju6, Ar0ju6);  // ../RTL/cortexm0ds_logic.v(8960)
  buf u936 (Trgpw6[28], Elgax6);  // ../RTL/cortexm0ds_logic.v(2376)
  or u9360 (n2461, D7fpw6[14], D7fpw6[7]);  // ../RTL/cortexm0ds_logic.v(8961)
  not u9361 (Tq0ju6, n2461);  // ../RTL/cortexm0ds_logic.v(8961)
  and u9362 (Fq0ju6, Hr0ju6, D7fpw6[13]);  // ../RTL/cortexm0ds_logic.v(8962)
  and u9363 (Hr0ju6, D7fpw6[5], Or0ju6);  // ../RTL/cortexm0ds_logic.v(8963)
  and u9364 (n2462, Vr0ju6, Cs0ju6);  // ../RTL/cortexm0ds_logic.v(8964)
  not u9365 (Or0ju6, n2462);  // ../RTL/cortexm0ds_logic.v(8964)
  and u9366 (n2463, Js0ju6, Qs0ju6);  // ../RTL/cortexm0ds_logic.v(8965)
  not u9367 (Cs0ju6, n2463);  // ../RTL/cortexm0ds_logic.v(8965)
  or u9368 (Un9ow6, D7fpw6[4], D7fpw6[6]);  // ../RTL/cortexm0ds_logic.v(8966)
  not u9369 (Qs0ju6, Un9ow6);  // ../RTL/cortexm0ds_logic.v(8966)
  not u937 (Tugpw6[5], n1272[5]);  // ../RTL/cortexm0ds_logic.v(16030)
  and u9370 (Js0ju6, Wh0ju6, F6ziu6);  // ../RTL/cortexm0ds_logic.v(8967)
  and u9371 (n2464, Ak0ju6, Oviiu6);  // ../RTL/cortexm0ds_logic.v(8968)
  not u9372 (Vr0ju6, n2464);  // ../RTL/cortexm0ds_logic.v(8968)
  and u9373 (Kp0ju6, Xs0ju6, Et0ju6);  // ../RTL/cortexm0ds_logic.v(8969)
  and u9374 (Wo0ju6, Lt0ju6, St0ju6);  // ../RTL/cortexm0ds_logic.v(8970)
  and u9375 (n2465, Zt0ju6, S6aiu6);  // ../RTL/cortexm0ds_logic.v(8971)
  not u9376 (St0ju6, n2465);  // ../RTL/cortexm0ds_logic.v(8971)
  or u9377 (n2466, Ii0iu6, Cyfpw6[4]);  // ../RTL/cortexm0ds_logic.v(8972)
  not u9378 (Zt0ju6, n2466);  // ../RTL/cortexm0ds_logic.v(8972)
  and u9379 (n2467, Gu0ju6, Xe8iu6);  // ../RTL/cortexm0ds_logic.v(8973)
  buf u938 (Uthpw6[16], Cjwpw6);  // ../RTL/cortexm0ds_logic.v(1882)
  not u9380 (Lt0ju6, n2467);  // ../RTL/cortexm0ds_logic.v(8973)
  or u9381 (Gu0ju6, W8aiu6, M2piu6);  // ../RTL/cortexm0ds_logic.v(8974)
  and u9382 (Io0ju6, Nu0ju6, Uu0ju6);  // ../RTL/cortexm0ds_logic.v(8975)
  and u9383 (Uu0ju6, Bv0ju6, Iv0ju6);  // ../RTL/cortexm0ds_logic.v(8976)
  and u9384 (n2468, Pv0ju6, Mr0iu6);  // ../RTL/cortexm0ds_logic.v(8977)
  not u9385 (Iv0ju6, n2468);  // ../RTL/cortexm0ds_logic.v(8977)
  or u9386 (Pv0ju6, Hzziu6, N3ziu6);  // ../RTL/cortexm0ds_logic.v(8978)
  and u9387 (n2469, Bziiu6, D7fpw6[11]);  // ../RTL/cortexm0ds_logic.v(8979)
  not u9388 (Bv0ju6, n2469);  // ../RTL/cortexm0ds_logic.v(8979)
  and u9389 (Nu0ju6, Wv0ju6, Dw0ju6);  // ../RTL/cortexm0ds_logic.v(8980)
  buf u939 (E1hpw6[4], Jraax6);  // ../RTL/cortexm0ds_logic.v(2367)
  or u9390 (Dw0ju6, Kw0ju6, Wxyiu6);  // ../RTL/cortexm0ds_logic.v(8981)
  and u9391 (n2470, D7fpw6[14], Rw0ju6);  // ../RTL/cortexm0ds_logic.v(8982)
  not u9392 (Wv0ju6, n2470);  // ../RTL/cortexm0ds_logic.v(8982)
  and u9393 (n2471, Yw0ju6, Fx0ju6);  // ../RTL/cortexm0ds_logic.v(8983)
  not u9394 (Rw0ju6, n2471);  // ../RTL/cortexm0ds_logic.v(8983)
  and u9395 (Fx0ju6, Mx0ju6, Tx0ju6);  // ../RTL/cortexm0ds_logic.v(8984)
  and u9396 (n2472, Mtjiu6, Ay0ju6);  // ../RTL/cortexm0ds_logic.v(8985)
  not u9397 (Tx0ju6, n2472);  // ../RTL/cortexm0ds_logic.v(8985)
  and u9398 (n2473, Hy0ju6, Oy0ju6);  // ../RTL/cortexm0ds_logic.v(8986)
  not u9399 (Ay0ju6, n2473);  // ../RTL/cortexm0ds_logic.v(8986)
  buf u94 (vis_r2_o[31], A3qax6);  // ../RTL/cortexm0ds_logic.v(2551)
  buf u940 (Gfghu6, Kqhbx6);  // ../RTL/cortexm0ds_logic.v(3050)
  and u9400 (Oy0ju6, Vy0ju6, Oviiu6);  // ../RTL/cortexm0ds_logic.v(8987)
  and u9401 (n2474, Cz0ju6, Jz0ju6);  // ../RTL/cortexm0ds_logic.v(8988)
  not u9402 (Vy0ju6, n2474);  // ../RTL/cortexm0ds_logic.v(8988)
  or u9403 (n2475, Hk0ju6, D7fpw6[7]);  // ../RTL/cortexm0ds_logic.v(8989)
  not u9404 (Cz0ju6, n2475);  // ../RTL/cortexm0ds_logic.v(8989)
  and u9405 (Hy0ju6, Qz0ju6, Xz0ju6);  // ../RTL/cortexm0ds_logic.v(8990)
  and u9406 (n2476, E01ju6, D7fpw6[8]);  // ../RTL/cortexm0ds_logic.v(8991)
  not u9407 (Xz0ju6, n2476);  // ../RTL/cortexm0ds_logic.v(8991)
  AL_MUX u9408 (
    .i0(Dcziu6),
    .i1(L01ju6),
    .sel(Tniiu6),
    .o(E01ju6));  // ../RTL/cortexm0ds_logic.v(8992)
  or u9409 (Mx0ju6, S01ju6, Jjhiu6);  // ../RTL/cortexm0ds_logic.v(8993)
  not u941 (Jndpw6, Kshbx6);  // ../RTL/cortexm0ds_logic.v(3051)
  and u9410 (Yw0ju6, Z01ju6, G11ju6);  // ../RTL/cortexm0ds_logic.v(8994)
  or u9411 (G11ju6, Hk0ju6, H95iu6);  // ../RTL/cortexm0ds_logic.v(8995)
  and u9412 (Un0ju6, N11ju6, U11ju6);  // ../RTL/cortexm0ds_logic.v(8996)
  and u9413 (U11ju6, B21ju6, I21ju6);  // ../RTL/cortexm0ds_logic.v(8997)
  and u9414 (I21ju6, P21ju6, W21ju6);  // ../RTL/cortexm0ds_logic.v(8998)
  and u9415 (n2477, N3ziu6, Taaiu6);  // ../RTL/cortexm0ds_logic.v(8999)
  not u9416 (W21ju6, n2477);  // ../RTL/cortexm0ds_logic.v(8999)
  and u9417 (n2478, Y0jiu6, D31ju6);  // ../RTL/cortexm0ds_logic.v(9000)
  not u9418 (P21ju6, n2478);  // ../RTL/cortexm0ds_logic.v(9000)
  and u9419 (B21ju6, K31ju6, R31ju6);  // ../RTL/cortexm0ds_logic.v(9001)
  buf u942 (Gtgpw6[3], Phcax6);  // ../RTL/cortexm0ds_logic.v(2375)
  or u9420 (R31ju6, Nloiu6, Lkaiu6);  // ../RTL/cortexm0ds_logic.v(9002)
  or u9421 (K31ju6, Jjhiu6, Y31ju6);  // ../RTL/cortexm0ds_logic.v(9003)
  and u9422 (N11ju6, F41ju6, M41ju6);  // ../RTL/cortexm0ds_logic.v(9004)
  and u9423 (M41ju6, T41ju6, A51ju6);  // ../RTL/cortexm0ds_logic.v(9005)
  or u9424 (A51ju6, Wiliu6, Ftjiu6);  // ../RTL/cortexm0ds_logic.v(9006)
  or u9425 (n2479, H51ju6, O51ju6);  // ../RTL/cortexm0ds_logic.v(9007)
  not u9426 (F41ju6, n2479);  // ../RTL/cortexm0ds_logic.v(9007)
  AL_MUX u9427 (
    .i0(Yljiu6),
    .i1(V51ju6),
    .sel(Cyfpw6[6]),
    .o(O51ju6));  // ../RTL/cortexm0ds_logic.v(9008)
  or u9428 (n2480, Ccoiu6, R75iu6);  // ../RTL/cortexm0ds_logic.v(9009)
  not u9429 (V51ju6, n2480);  // ../RTL/cortexm0ds_logic.v(9009)
  not u943 (Tugpw6[6], n1272[6]);  // ../RTL/cortexm0ds_logic.v(16030)
  AL_MUX u9430 (
    .i0(M2piu6),
    .i1(C61ju6),
    .sel(Cyfpw6[7]),
    .o(H51ju6));  // ../RTL/cortexm0ds_logic.v(9010)
  and u9431 (n2481, J61ju6, Q61ju6);  // ../RTL/cortexm0ds_logic.v(9011)
  not u9432 (C61ju6, n2481);  // ../RTL/cortexm0ds_logic.v(9011)
  and u9433 (Q61ju6, X61ju6, E71ju6);  // ../RTL/cortexm0ds_logic.v(9012)
  and u9434 (n2482, I30ju6, Pxyiu6);  // ../RTL/cortexm0ds_logic.v(9013)
  not u9435 (E71ju6, n2482);  // ../RTL/cortexm0ds_logic.v(9013)
  and u9436 (n2483, Moaiu6, N2ghu6);  // ../RTL/cortexm0ds_logic.v(9014)
  not u9437 (X61ju6, n2483);  // ../RTL/cortexm0ds_logic.v(9014)
  and u9438 (J61ju6, L71ju6, S71ju6);  // ../RTL/cortexm0ds_logic.v(9015)
  or u9439 (S71ju6, X5oiu6, C0ehu6);  // ../RTL/cortexm0ds_logic.v(9016)
  buf u944 (Uthpw6[17], Pdbbx6);  // ../RTL/cortexm0ds_logic.v(1882)
  and u9440 (n2484, D1piu6, Pugiu6);  // ../RTL/cortexm0ds_logic.v(9017)
  not u9441 (L71ju6, n2484);  // ../RTL/cortexm0ds_logic.v(9017)
  or u9442 (Gn0ju6, Cyfpw6[7], HREADY);  // ../RTL/cortexm0ds_logic.v(9018)
  AL_MUX u9443 (
    .i0(Z71ju6),
    .i1(H2fpw6[1]),
    .sel(G81ju6),
    .o(Mwohu6));  // ../RTL/cortexm0ds_logic.v(9019)
  and u9444 (n2485, N81ju6, U81ju6);  // ../RTL/cortexm0ds_logic.v(9020)
  not u9445 (Z71ju6, n2485);  // ../RTL/cortexm0ds_logic.v(9020)
  and u9446 (U81ju6, B91ju6, I91ju6);  // ../RTL/cortexm0ds_logic.v(9021)
  and u9447 (n2486, P91ju6, D7fpw6[4]);  // ../RTL/cortexm0ds_logic.v(9022)
  not u9448 (I91ju6, n2486);  // ../RTL/cortexm0ds_logic.v(9022)
  and u9449 (B91ju6, W91ju6, Da1ju6);  // ../RTL/cortexm0ds_logic.v(9023)
  buf u945 (E1hpw6[5], Npaax6);  // ../RTL/cortexm0ds_logic.v(2367)
  and u9450 (n2487, Ka1ju6, Ra1ju6);  // ../RTL/cortexm0ds_logic.v(9024)
  not u9451 (Da1ju6, n2487);  // ../RTL/cortexm0ds_logic.v(9024)
  or u9452 (n2488, Jcaiu6, D7fpw6[11]);  // ../RTL/cortexm0ds_logic.v(9025)
  not u9453 (Ra1ju6, n2488);  // ../RTL/cortexm0ds_logic.v(9025)
  and u9454 (Ka1ju6, D7fpw6[13], Ya1ju6);  // ../RTL/cortexm0ds_logic.v(9026)
  and u9455 (n2489, Fb1ju6, D7fpw6[9]);  // ../RTL/cortexm0ds_logic.v(9027)
  not u9456 (W91ju6, n2489);  // ../RTL/cortexm0ds_logic.v(9027)
  and u9457 (N81ju6, Mb1ju6, Tb1ju6);  // ../RTL/cortexm0ds_logic.v(9028)
  and u9458 (n2490, D7fpw6[1], Ac1ju6);  // ../RTL/cortexm0ds_logic.v(9029)
  not u9459 (Tb1ju6, n2490);  // ../RTL/cortexm0ds_logic.v(9029)
  buf u946 (vis_r4_o[29], Wpuax6);  // ../RTL/cortexm0ds_logic.v(2626)
  and u9460 (Fwohu6, Rgnhu6, Hc1ju6);  // ../RTL/cortexm0ds_logic.v(9030)
  and u9461 (n2491, Aw3iu6, Oc1ju6);  // ../RTL/cortexm0ds_logic.v(9031)
  not u9462 (Hc1ju6, n2491);  // ../RTL/cortexm0ds_logic.v(9031)
  and u9463 (n2492, Tonhu6, Di1iu6);  // ../RTL/cortexm0ds_logic.v(9032)
  not u9464 (Oc1ju6, n2492);  // ../RTL/cortexm0ds_logic.v(9032)
  and u9465 (Di1iu6, Tezhu6, O8zhu6);  // ../RTL/cortexm0ds_logic.v(9033)
  and u9466 (Tezhu6, Vc1ju6, Cq3iu6);  // ../RTL/cortexm0ds_logic.v(9034)
  and u9467 (Cq3iu6, Cd1ju6, Fj1iu6);  // ../RTL/cortexm0ds_logic.v(9035)
  and u9468 (Fj1iu6, Jd1ju6, Qd1ju6);  // ../RTL/cortexm0ds_logic.v(9036)
  and u9469 (Qd1ju6, Omzhu6, Xj3iu6);  // ../RTL/cortexm0ds_logic.v(9037)
  buf u947 (Vxmhu6, F4ibx6);  // ../RTL/cortexm0ds_logic.v(3057)
  and u9470 (K7yhu6, Xd1ju6, Ow3iu6);  // ../RTL/cortexm0ds_logic.v(9038)
  not u9471 (Xj3iu6, K7yhu6);  // ../RTL/cortexm0ds_logic.v(9038)
  and u9472 (n2493, Ee1ju6, Yn3iu6);  // ../RTL/cortexm0ds_logic.v(9039)
  not u9473 (Ow3iu6, n2493);  // ../RTL/cortexm0ds_logic.v(9039)
  or u9474 (n2494, Ulnhu6, Mdhpw6[2]);  // ../RTL/cortexm0ds_logic.v(9040)
  not u9475 (Yn3iu6, n2494);  // ../RTL/cortexm0ds_logic.v(9040)
  and u9476 (Ee1ju6, Le1ju6, Qnzhu6);  // ../RTL/cortexm0ds_logic.v(9041)
  or u9477 (Qnzhu6, O8zhu6, Mdhpw6[0]);  // ../RTL/cortexm0ds_logic.v(9042)
  not u9478 (O8zhu6, Mdhpw6[1]);  // ../RTL/cortexm0ds_logic.v(9043)
  and u9479 (n2495, Pinhu6, Mdhpw6[1]);  // ../RTL/cortexm0ds_logic.v(9044)
  buf u948 (vis_r1_o[13], I5qpw6);  // ../RTL/cortexm0ds_logic.v(1876)
  not u9480 (Le1ju6, n2495);  // ../RTL/cortexm0ds_logic.v(9044)
  and u9481 (n2496, Se1ju6, Ze1ju6);  // ../RTL/cortexm0ds_logic.v(9045)
  not u9482 (Xd1ju6, n2496);  // ../RTL/cortexm0ds_logic.v(9045)
  or u9483 (n2497, Fanhu6, Jdnhu6);  // ../RTL/cortexm0ds_logic.v(9046)
  not u9484 (Ze1ju6, n2497);  // ../RTL/cortexm0ds_logic.v(9046)
  or u9485 (n2498, Ph1iu6, Q8nhu6);  // ../RTL/cortexm0ds_logic.v(9047)
  not u9486 (Se1ju6, n2498);  // ../RTL/cortexm0ds_logic.v(9047)
  and u9487 (Ph1iu6, Gf1ju6, X0ohu6);  // ../RTL/cortexm0ds_logic.v(9048)
  and u9488 (Gf1ju6, Mo3iu6, Aw3iu6);  // ../RTL/cortexm0ds_logic.v(9049)
  and u9489 (Mo3iu6, Nf1ju6, Uf1ju6);  // ../RTL/cortexm0ds_logic.v(9050)
  buf u949 (D7fpw6[10], Ssjax6);  // ../RTL/cortexm0ds_logic.v(2074)
  or u9490 (n2499, Z63iu6, Vmdpw6);  // ../RTL/cortexm0ds_logic.v(9051)
  not u9491 (Uf1ju6, n2499);  // ../RTL/cortexm0ds_logic.v(9051)
  xor u9492 (Z63iu6, G2ohu6, Rrnhu6);  // ../RTL/cortexm0ds_logic.v(9052)
  and u9493 (Nf1ju6, Rgnhu6, Fmyhu6);  // ../RTL/cortexm0ds_logic.v(9053)
  and u9494 (Fmyhu6, Bg1ju6, Mdhpw6[3]);  // ../RTL/cortexm0ds_logic.v(9055)
  not u9495 (N5yhu6, Fmyhu6);  // ../RTL/cortexm0ds_logic.v(9055)
  and u9496 (Bg1ju6, U5yhu6, Agyhu6);  // ../RTL/cortexm0ds_logic.v(9056)
  and u9497 (Agyhu6, Ig1ju6, Ighpw6[3]);  // ../RTL/cortexm0ds_logic.v(9057)
  or u9498 (n2500, Vmzhu6, Deyhu6);  // ../RTL/cortexm0ds_logic.v(9058)
  not u9499 (Ig1ju6, n2500);  // ../RTL/cortexm0ds_logic.v(9058)
  buf u95 (Shhpw6[0], I4rpw6);  // ../RTL/cortexm0ds_logic.v(1941)
  buf u950 (Tzfpw6[2], Kzabx6);  // ../RTL/cortexm0ds_logic.v(2007)
  or u9500 (Deyhu6, Zwyhu6, Ighpw6[0]);  // ../RTL/cortexm0ds_logic.v(9059)
  not u9501 (Zwyhu6, Ighpw6[1]);  // ../RTL/cortexm0ds_logic.v(9060)
  or u9502 (n2501, Ighpw6[0], Ighpw6[1]);  // ../RTL/cortexm0ds_logic.v(9061)
  not u9503 (Omzhu6, n2501);  // ../RTL/cortexm0ds_logic.v(9061)
  and u9504 (Jd1ju6, Iyyhu6, U5yhu6);  // ../RTL/cortexm0ds_logic.v(9062)
  and u9505 (Iyyhu6, Ez2iu6, Wdyhu6);  // ../RTL/cortexm0ds_logic.v(9063)
  or u9506 (n2502, Ulnhu6, Mdhpw6[0]);  // ../RTL/cortexm0ds_logic.v(9064)
  not u9507 (Cd1ju6, n2502);  // ../RTL/cortexm0ds_logic.v(9064)
  or u9508 (n2503, Vp3iu6, Mdhpw6[2]);  // ../RTL/cortexm0ds_logic.v(9065)
  not u9509 (Vc1ju6, n2503);  // ../RTL/cortexm0ds_logic.v(9065)
  buf u951 (vis_r12_o[15], Zf8bx6);  // ../RTL/cortexm0ds_logic.v(2599)
  xor u9510 (Ofzhu6, Rzyhu6, Mdhpw6[3]);  // ../RTL/cortexm0ds_logic.v(9066)
  not u9511 (Vp3iu6, Ofzhu6);  // ../RTL/cortexm0ds_logic.v(9066)
  not u9512 (Rzyhu6, Hknhu6);  // ../RTL/cortexm0ds_logic.v(9067)
  not u9513 (Aw3iu6, Yenhu6);  // ../RTL/cortexm0ds_logic.v(9068)
  AL_MUX u9514 (
    .i0(Mdhpw6[2]),
    .i1(Mdhpw6[3]),
    .sel(Y14iu6),
    .o(Yvohu6));  // ../RTL/cortexm0ds_logic.v(9069)
  AL_MUX u9515 (
    .i0(Mdhpw6[1]),
    .i1(Mdhpw6[2]),
    .sel(Y14iu6),
    .o(Rvohu6));  // ../RTL/cortexm0ds_logic.v(9070)
  not u9516 (Y14iu6, U03iu6);  // ../RTL/cortexm0ds_logic.v(9071)
  AL_MUX u9517 (
    .i0(Mdhpw6[1]),
    .i1(Mdhpw6[0]),
    .sel(U03iu6),
    .o(Kvohu6));  // ../RTL/cortexm0ds_logic.v(9072)
  AL_MUX u9518 (
    .i0(Mdhpw6[0]),
    .i1(Ulnhu6),
    .sel(U03iu6),
    .o(Dvohu6));  // ../RTL/cortexm0ds_logic.v(9073)
  and u9519 (U03iu6, Pg1ju6, Wg1ju6);  // ../RTL/cortexm0ds_logic.v(9074)
  buf u952 (vis_r0_o[14], Sx7ax6);  // ../RTL/cortexm0ds_logic.v(1875)
  and u9520 (n2504, Dh1ju6, Ijzhu6);  // ../RTL/cortexm0ds_logic.v(9075)
  not u9521 (Wg1ju6, n2504);  // ../RTL/cortexm0ds_logic.v(9075)
  or u9522 (n2505, Ighpw6[3], Ighpw6[4]);  // ../RTL/cortexm0ds_logic.v(9076)
  not u9523 (Ijzhu6, n2505);  // ../RTL/cortexm0ds_logic.v(9076)
  and u9524 (Dh1ju6, U5yhu6, Vmzhu6);  // ../RTL/cortexm0ds_logic.v(9077)
  not u9525 (Vmzhu6, Ez2iu6);  // ../RTL/cortexm0ds_logic.v(9078)
  and u9526 (Ez2iu6, Vuyhu6, Eiyhu6);  // ../RTL/cortexm0ds_logic.v(9079)
  not u9527 (Eiyhu6, Ighpw6[4]);  // ../RTL/cortexm0ds_logic.v(9080)
  not u9528 (Vuyhu6, Ighpw6[2]);  // ../RTL/cortexm0ds_logic.v(9081)
  and u9529 (n2506, Kh1ju6, Rh1ju6);  // ../RTL/cortexm0ds_logic.v(9082)
  buf u953 (Tzfpw6[21], Tjkpw6);  // ../RTL/cortexm0ds_logic.v(2007)
  not u9530 (Pg1ju6, n2506);  // ../RTL/cortexm0ds_logic.v(9082)
  and u9531 (Rh1ju6, Yh1ju6, Pdyhu6);  // ../RTL/cortexm0ds_logic.v(9083)
  not u9532 (Pdyhu6, Pkyhu6);  // ../RTL/cortexm0ds_logic.v(9084)
  and u9533 (Pkyhu6, Ighpw6[2], Cvyhu6);  // ../RTL/cortexm0ds_logic.v(9085)
  or u9534 (Yh1ju6, Cvyhu6, Ighpw6[2]);  // ../RTL/cortexm0ds_logic.v(9086)
  and u9535 (Cvyhu6, Ighpw6[0], Ighpw6[1]);  // ../RTL/cortexm0ds_logic.v(9087)
  and u9536 (Kh1ju6, Epyhu6, U5yhu6);  // ../RTL/cortexm0ds_logic.v(9088)
  and u9537 (U5yhu6, Vx2iu6, Ujyhu6);  // ../RTL/cortexm0ds_logic.v(9089)
  not u9538 (Vx2iu6, Fnnhu6);  // ../RTL/cortexm0ds_logic.v(9090)
  and u9539 (Epyhu6, Ighpw6[4], Wdyhu6);  // ../RTL/cortexm0ds_logic.v(9091)
  not u954 (Zehpw6[1], n7[1]);  // ../RTL/cortexm0ds_logic.v(3185)
  not u9540 (Wdyhu6, Ighpw6[3]);  // ../RTL/cortexm0ds_logic.v(9092)
  AL_MUX u9541 (
    .i0(Fi1ju6),
    .i1(X3fpw6[2]),
    .sel(O25iu6),
    .o(Wuohu6));  // ../RTL/cortexm0ds_logic.v(9093)
  and u9542 (n2507, Mi1ju6, Ti1ju6);  // ../RTL/cortexm0ds_logic.v(9094)
  not u9543 (Fi1ju6, n2507);  // ../RTL/cortexm0ds_logic.v(9094)
  and u9544 (Ti1ju6, Aj1ju6, Hj1ju6);  // ../RTL/cortexm0ds_logic.v(9095)
  and u9545 (n2508, Omyiu6, S8fpw6[10]);  // ../RTL/cortexm0ds_logic.v(9096)
  not u9546 (Hj1ju6, n2508);  // ../RTL/cortexm0ds_logic.v(9096)
  and u9547 (Aj1ju6, Oj1ju6, Vj1ju6);  // ../RTL/cortexm0ds_logic.v(9097)
  and u9548 (n2509, D7fpw6[5], K75iu6);  // ../RTL/cortexm0ds_logic.v(9098)
  not u9549 (Vj1ju6, n2509);  // ../RTL/cortexm0ds_logic.v(9098)
  buf u955 (Shhpw6[3], L03qw6);  // ../RTL/cortexm0ds_logic.v(1941)
  and u9550 (n2510, L45iu6, N55iu6);  // ../RTL/cortexm0ds_logic.v(9099)
  not u9551 (Oj1ju6, n2510);  // ../RTL/cortexm0ds_logic.v(9099)
  and u9552 (Mi1ju6, Ck1ju6, Gpyiu6);  // ../RTL/cortexm0ds_logic.v(9100)
  and u9553 (Ck1ju6, Jk1ju6, Qk1ju6);  // ../RTL/cortexm0ds_logic.v(9101)
  and u9554 (n2511, A95iu6, D7fpw6[2]);  // ../RTL/cortexm0ds_logic.v(9102)
  not u9555 (Qk1ju6, n2511);  // ../RTL/cortexm0ds_logic.v(9102)
  or u9556 (Jk1ju6, Ndiiu6, H95iu6);  // ../RTL/cortexm0ds_logic.v(9103)
  not u9557 (Puohu6, Xk1ju6);  // ../RTL/cortexm0ds_logic.v(9104)
  AL_MUX u9558 (
    .i0(El1ju6),
    .i1(Ll1ju6),
    .sel(HREADY),
    .o(Xk1ju6));  // ../RTL/cortexm0ds_logic.v(9105)
  and u9559 (Ll1ju6, Sl1ju6, Zl1ju6);  // ../RTL/cortexm0ds_logic.v(9106)
  buf u956 (vis_r9_o[16], C9wpw6);  // ../RTL/cortexm0ds_logic.v(1898)
  not u9560 (Iuohu6, Gm1ju6);  // ../RTL/cortexm0ds_logic.v(9107)
  AL_MUX u9561 (
    .i0(Nm1ju6),
    .i1(Um1ju6),
    .sel(HREADY),
    .o(Gm1ju6));  // ../RTL/cortexm0ds_logic.v(9108)
  and u9562 (Um1ju6, Bn1ju6, In1ju6);  // ../RTL/cortexm0ds_logic.v(9109)
  and u9563 (In1ju6, Pn1ju6, Wn1ju6);  // ../RTL/cortexm0ds_logic.v(9110)
  and u9564 (Wn1ju6, Do1ju6, Ko1ju6);  // ../RTL/cortexm0ds_logic.v(9111)
  and u9565 (n2512, Ro1ju6, Yo1ju6);  // ../RTL/cortexm0ds_logic.v(9112)
  not u9566 (Ko1ju6, n2512);  // ../RTL/cortexm0ds_logic.v(9112)
  and u9567 (Ro1ju6, Fp1ju6, Mp1ju6);  // ../RTL/cortexm0ds_logic.v(9113)
  and u9568 (n2513, Ph0ju6, Tp1ju6);  // ../RTL/cortexm0ds_logic.v(9114)
  not u9569 (Mp1ju6, n2513);  // ../RTL/cortexm0ds_logic.v(9114)
  buf u957 (vis_r3_o[21], D46bx6);  // ../RTL/cortexm0ds_logic.v(2694)
  and u9570 (n2514, D7fpw6[7], Aq1ju6);  // ../RTL/cortexm0ds_logic.v(9115)
  not u9571 (Tp1ju6, n2514);  // ../RTL/cortexm0ds_logic.v(9115)
  and u9572 (Do1ju6, Hq1ju6, Oq1ju6);  // ../RTL/cortexm0ds_logic.v(9116)
  and u9573 (Pn1ju6, Vq1ju6, Cr1ju6);  // ../RTL/cortexm0ds_logic.v(9117)
  and u9574 (n2515, Oiaiu6, Jr1ju6);  // ../RTL/cortexm0ds_logic.v(9118)
  not u9575 (Cr1ju6, n2515);  // ../RTL/cortexm0ds_logic.v(9118)
  and u9576 (n2516, Qr1ju6, Xr1ju6);  // ../RTL/cortexm0ds_logic.v(9119)
  not u9577 (Jr1ju6, n2516);  // ../RTL/cortexm0ds_logic.v(9119)
  and u9578 (n2517, Es1ju6, Qe8iu6);  // ../RTL/cortexm0ds_logic.v(9120)
  not u9579 (Xr1ju6, n2517);  // ../RTL/cortexm0ds_logic.v(9120)
  buf u958 (vis_msp_o[16], Tc0qw6);  // ../RTL/cortexm0ds_logic.v(2097)
  and u9580 (n2518, Toaiu6, Ls1ju6);  // ../RTL/cortexm0ds_logic.v(9121)
  not u9581 (Qr1ju6, n2518);  // ../RTL/cortexm0ds_logic.v(9121)
  and u9582 (Vq1ju6, Ss1ju6, Zs1ju6);  // ../RTL/cortexm0ds_logic.v(9122)
  and u9583 (n2519, Gt1ju6, M2piu6);  // ../RTL/cortexm0ds_logic.v(9123)
  not u9584 (Zs1ju6, n2519);  // ../RTL/cortexm0ds_logic.v(9123)
  or u9585 (n2520, Ccoiu6, Cyfpw6[0]);  // ../RTL/cortexm0ds_logic.v(9124)
  not u9586 (Gt1ju6, n2520);  // ../RTL/cortexm0ds_logic.v(9124)
  and u9587 (n2521, K2aiu6, Nt1ju6);  // ../RTL/cortexm0ds_logic.v(9125)
  not u9588 (Ss1ju6, n2521);  // ../RTL/cortexm0ds_logic.v(9125)
  and u9589 (n2522, Ut1ju6, Bu1ju6);  // ../RTL/cortexm0ds_logic.v(9126)
  buf u959 (vis_r11_o[13], Vlkpw6);  // ../RTL/cortexm0ds_logic.v(1874)
  not u9590 (Nt1ju6, n2522);  // ../RTL/cortexm0ds_logic.v(9126)
  and u9591 (n2523, Iu1ju6, Pu1ju6);  // ../RTL/cortexm0ds_logic.v(9127)
  not u9592 (Bu1ju6, n2523);  // ../RTL/cortexm0ds_logic.v(9127)
  and u9593 (Iu1ju6, Md0iu6, Sijiu6);  // ../RTL/cortexm0ds_logic.v(9128)
  and u9594 (Qdaow6, Qe8iu6, Mr0iu6);  // ../RTL/cortexm0ds_logic.v(9129)
  not u9595 (Ut1ju6, Qdaow6);  // ../RTL/cortexm0ds_logic.v(9129)
  and u9596 (Bn1ju6, Wu1ju6, Dv1ju6);  // ../RTL/cortexm0ds_logic.v(9130)
  and u9597 (Dv1ju6, Kv1ju6, Rv1ju6);  // ../RTL/cortexm0ds_logic.v(9131)
  and u9598 (n2524, Yv1ju6, Wliiu6);  // ../RTL/cortexm0ds_logic.v(9132)
  not u9599 (Rv1ju6, n2524);  // ../RTL/cortexm0ds_logic.v(9132)
  buf u96 (vis_r12_o[0], Kssax6);  // ../RTL/cortexm0ds_logic.v(2599)
  buf u960 (Hrfpw6[8], Qyjax6);  // ../RTL/cortexm0ds_logic.v(2428)
  and u9600 (Kv1ju6, Fw1ju6, Mw1ju6);  // ../RTL/cortexm0ds_logic.v(9133)
  and u9601 (n2525, Tw1ju6, Oviiu6);  // ../RTL/cortexm0ds_logic.v(9134)
  not u9602 (Mw1ju6, n2525);  // ../RTL/cortexm0ds_logic.v(9134)
  and u9603 (n2526, Ax1ju6, Hx1ju6);  // ../RTL/cortexm0ds_logic.v(9135)
  not u9604 (Tw1ju6, n2526);  // ../RTL/cortexm0ds_logic.v(9135)
  and u9605 (Pv9ow6, Yv1ju6, Nbkiu6);  // ../RTL/cortexm0ds_logic.v(9136)
  not u9606 (Hx1ju6, Pv9ow6);  // ../RTL/cortexm0ds_logic.v(9136)
  and u9607 (n2527, Pugiu6, Ox1ju6);  // ../RTL/cortexm0ds_logic.v(9137)
  not u9608 (Fw1ju6, n2527);  // ../RTL/cortexm0ds_logic.v(9137)
  and u9609 (n2528, Vx1ju6, Cy1ju6);  // ../RTL/cortexm0ds_logic.v(9138)
  buf u961 (Gqgpw6[8], R1eax6);  // ../RTL/cortexm0ds_logic.v(2377)
  not u9610 (Ox1ju6, n2528);  // ../RTL/cortexm0ds_logic.v(9138)
  and u9611 (n2529, M2piu6, Jy1ju6);  // ../RTL/cortexm0ds_logic.v(9139)
  not u9612 (Cy1ju6, n2529);  // ../RTL/cortexm0ds_logic.v(9139)
  and u9613 (n2530, Xojiu6, Qy1ju6);  // ../RTL/cortexm0ds_logic.v(9140)
  not u9614 (Jy1ju6, n2530);  // ../RTL/cortexm0ds_logic.v(9140)
  or u9615 (Qy1ju6, Mmjiu6, Ae0iu6);  // ../RTL/cortexm0ds_logic.v(9141)
  and u9616 (Wu1ju6, Xy1ju6, Ez1ju6);  // ../RTL/cortexm0ds_logic.v(9142)
  and u9617 (Xy1ju6, Lz1ju6, Sz1ju6);  // ../RTL/cortexm0ds_logic.v(9143)
  and u9618 (n2531, U98iu6, Vxniu6);  // ../RTL/cortexm0ds_logic.v(9144)
  not u9619 (Sz1ju6, n2531);  // ../RTL/cortexm0ds_logic.v(9144)
  buf u962 (Shhpw6[13], Fj8ax6);  // ../RTL/cortexm0ds_logic.v(1941)
  or u9620 (Lz1ju6, Ax1ju6, L01ju6);  // ../RTL/cortexm0ds_logic.v(9145)
  and u9621 (n2532, Zz1ju6, G02ju6);  // ../RTL/cortexm0ds_logic.v(9146)
  not u9622 (Buohu6, n2532);  // ../RTL/cortexm0ds_logic.v(9146)
  and u9623 (n2533, C0ehu6, N02ju6);  // ../RTL/cortexm0ds_logic.v(9147)
  not u9624 (G02ju6, n2533);  // ../RTL/cortexm0ds_logic.v(9147)
  or u9625 (N02ju6, Eh6iu6, Yv1ju6);  // ../RTL/cortexm0ds_logic.v(9148)
  and u9626 (n2534, HREADY, U02ju6);  // ../RTL/cortexm0ds_logic.v(9149)
  not u9627 (Zz1ju6, n2534);  // ../RTL/cortexm0ds_logic.v(9149)
  and u9628 (n2535, B12ju6, I12ju6);  // ../RTL/cortexm0ds_logic.v(9150)
  not u9629 (U02ju6, n2535);  // ../RTL/cortexm0ds_logic.v(9150)
  not u963 (Cndpw6, Pgjbx6);  // ../RTL/cortexm0ds_logic.v(3082)
  and u9630 (I12ju6, P12ju6, W12ju6);  // ../RTL/cortexm0ds_logic.v(9151)
  and u9631 (W12ju6, D22ju6, K22ju6);  // ../RTL/cortexm0ds_logic.v(9152)
  and u9632 (n2536, U98iu6, R22ju6);  // ../RTL/cortexm0ds_logic.v(9153)
  not u9633 (K22ju6, n2536);  // ../RTL/cortexm0ds_logic.v(9153)
  and u9634 (n2537, Y22ju6, F32ju6);  // ../RTL/cortexm0ds_logic.v(9154)
  not u9635 (R22ju6, n2537);  // ../RTL/cortexm0ds_logic.v(9154)
  or u9636 (F32ju6, M32ju6, Xmliu6);  // ../RTL/cortexm0ds_logic.v(9155)
  and u9637 (n2538, Pthiu6, Cyfpw6[1]);  // ../RTL/cortexm0ds_logic.v(9156)
  not u9638 (Y22ju6, n2538);  // ../RTL/cortexm0ds_logic.v(9156)
  and u9639 (D22ju6, T32ju6, A42ju6);  // ../RTL/cortexm0ds_logic.v(9157)
  buf u964 (Trgpw6[23], Q1hbx6);  // ../RTL/cortexm0ds_logic.v(2376)
  and u9640 (n2539, H42ju6, Neoiu6);  // ../RTL/cortexm0ds_logic.v(9158)
  not u9641 (T32ju6, n2539);  // ../RTL/cortexm0ds_logic.v(9158)
  and u9642 (H42ju6, Omyiu6, O42ju6);  // ../RTL/cortexm0ds_logic.v(9159)
  and u9643 (n2540, V42ju6, C52ju6);  // ../RTL/cortexm0ds_logic.v(9160)
  not u9644 (O42ju6, n2540);  // ../RTL/cortexm0ds_logic.v(9160)
  and u9645 (C52ju6, J52ju6, Q52ju6);  // ../RTL/cortexm0ds_logic.v(9161)
  or u9646 (Q52ju6, As0iu6, Xe8iu6);  // ../RTL/cortexm0ds_logic.v(9162)
  and u9647 (J52ju6, X52ju6, E62ju6);  // ../RTL/cortexm0ds_logic.v(9163)
  or u9648 (X52ju6, L62ju6, Cyfpw6[6]);  // ../RTL/cortexm0ds_logic.v(9164)
  and u9649 (V42ju6, Cyfpw6[0], S62ju6);  // ../RTL/cortexm0ds_logic.v(9165)
  buf u965 (Gtgpw6[28], Hjgax6);  // ../RTL/cortexm0ds_logic.v(2375)
  and u9650 (P12ju6, Z62ju6, G72ju6);  // ../RTL/cortexm0ds_logic.v(9166)
  and u9651 (n2541, Dxziu6, N72ju6);  // ../RTL/cortexm0ds_logic.v(9167)
  not u9652 (G72ju6, n2541);  // ../RTL/cortexm0ds_logic.v(9167)
  and u9653 (n2542, U72ju6, B82ju6);  // ../RTL/cortexm0ds_logic.v(9168)
  not u9654 (N72ju6, n2542);  // ../RTL/cortexm0ds_logic.v(9168)
  and u9655 (n2543, Ls1ju6, Xzmiu6);  // ../RTL/cortexm0ds_logic.v(9169)
  not u9656 (B82ju6, n2543);  // ../RTL/cortexm0ds_logic.v(9169)
  and u9657 (n2544, I82ju6, Nlaiu6);  // ../RTL/cortexm0ds_logic.v(9170)
  not u9658 (U72ju6, n2544);  // ../RTL/cortexm0ds_logic.v(9170)
  or u9659 (Z62ju6, P82ju6, W82ju6);  // ../RTL/cortexm0ds_logic.v(9171)
  buf u966 (Uthpw6[11], Bu6bx6);  // ../RTL/cortexm0ds_logic.v(1882)
  and u9660 (B12ju6, D92ju6, K92ju6);  // ../RTL/cortexm0ds_logic.v(9172)
  and u9661 (K92ju6, R92ju6, Y92ju6);  // ../RTL/cortexm0ds_logic.v(9173)
  and u9662 (n2545, Qe8iu6, Fa2ju6);  // ../RTL/cortexm0ds_logic.v(9174)
  not u9663 (Y92ju6, n2545);  // ../RTL/cortexm0ds_logic.v(9174)
  and u9664 (n2546, Ma2ju6, Ta2ju6);  // ../RTL/cortexm0ds_logic.v(9175)
  not u9665 (Fa2ju6, n2546);  // ../RTL/cortexm0ds_logic.v(9175)
  AL_MUX u9666 (
    .i0(Ab2ju6),
    .i1(Hb2ju6),
    .sel(H4ghu6),
    .o(Ta2ju6));  // ../RTL/cortexm0ds_logic.v(9176)
  and u9667 (n2547, Dxziu6, Ob2ju6);  // ../RTL/cortexm0ds_logic.v(9177)
  not u9668 (Hb2ju6, n2547);  // ../RTL/cortexm0ds_logic.v(9177)
  and u9669 (n2548, Cyfpw6[5], Vb2ju6);  // ../RTL/cortexm0ds_logic.v(9178)
  buf u967 (G4hpw6[1], X5bax6);  // ../RTL/cortexm0ds_logic.v(2274)
  not u9670 (Ob2ju6, n2548);  // ../RTL/cortexm0ds_logic.v(9178)
  and u9671 (n2549, Cc2ju6, Eoyiu6);  // ../RTL/cortexm0ds_logic.v(9179)
  not u9672 (Vb2ju6, n2549);  // ../RTL/cortexm0ds_logic.v(9179)
  or u9673 (n2550, Nlaiu6, Cyfpw6[3]);  // ../RTL/cortexm0ds_logic.v(9180)
  not u9674 (Cc2ju6, n2550);  // ../RTL/cortexm0ds_logic.v(9180)
  and u9675 (Ab2ju6, Jc2ju6, Qc2ju6);  // ../RTL/cortexm0ds_logic.v(9181)
  and u9676 (n2551, Xc2ju6, Ed2ju6);  // ../RTL/cortexm0ds_logic.v(9182)
  not u9677 (Qc2ju6, n2551);  // ../RTL/cortexm0ds_logic.v(9182)
  or u9678 (n2552, Xojiu6, Sbghu6);  // ../RTL/cortexm0ds_logic.v(9183)
  not u9679 (Ed2ju6, n2552);  // ../RTL/cortexm0ds_logic.v(9183)
  buf u968 (E1hpw6[29], Tchbx6);  // ../RTL/cortexm0ds_logic.v(2367)
  or u9680 (Er2ju6, Nlaiu6, Lkaiu6);  // ../RTL/cortexm0ds_logic.v(9184)
  not u9681 (Xc2ju6, Er2ju6);  // ../RTL/cortexm0ds_logic.v(9184)
  and u9682 (Ma2ju6, Ld2ju6, M32ju6);  // ../RTL/cortexm0ds_logic.v(9185)
  and u9683 (n2553, Sd2ju6, Hs0iu6);  // ../RTL/cortexm0ds_logic.v(9186)
  not u9684 (Ld2ju6, n2553);  // ../RTL/cortexm0ds_logic.v(9186)
  and u9685 (n2554, Q5aiu6, Zd2ju6);  // ../RTL/cortexm0ds_logic.v(9187)
  not u9686 (Sd2ju6, n2554);  // ../RTL/cortexm0ds_logic.v(9187)
  and u9687 (n2555, Fsdhu6, Xbopw6);  // ../RTL/cortexm0ds_logic.v(9188)
  not u9688 (Zd2ju6, n2555);  // ../RTL/cortexm0ds_logic.v(9188)
  and u9689 (n2556, Yo1ju6, I6jiu6);  // ../RTL/cortexm0ds_logic.v(9189)
  buf u969 (E1hpw6[30], Z2aax6);  // ../RTL/cortexm0ds_logic.v(2367)
  not u9690 (R92ju6, n2556);  // ../RTL/cortexm0ds_logic.v(9189)
  and u9691 (D92ju6, Ge2ju6, Ne2ju6);  // ../RTL/cortexm0ds_logic.v(9190)
  and u9692 (n2557, W8aiu6, Whfiu6);  // ../RTL/cortexm0ds_logic.v(9191)
  not u9693 (Ne2ju6, n2557);  // ../RTL/cortexm0ds_logic.v(9191)
  AL_MUX u9694 (
    .i0(Ue2ju6),
    .i1(Bf2ju6),
    .sel(D7fpw6[8]),
    .o(Ge2ju6));  // ../RTL/cortexm0ds_logic.v(9192)
  and u9695 (Bf2ju6, If2ju6, Pf2ju6);  // ../RTL/cortexm0ds_logic.v(9193)
  and u9696 (n2558, Wf2ju6, Y5ziu6);  // ../RTL/cortexm0ds_logic.v(9194)
  not u9697 (Pf2ju6, n2558);  // ../RTL/cortexm0ds_logic.v(9194)
  and u9698 (n2559, Yo1ju6, Tniiu6);  // ../RTL/cortexm0ds_logic.v(9195)
  not u9699 (If2ju6, n2559);  // ../RTL/cortexm0ds_logic.v(9195)
  buf u97 (vis_r1_o[0], M2lax6);  // ../RTL/cortexm0ds_logic.v(1876)
  buf u970 (E1hpw6[31], N4gax6);  // ../RTL/cortexm0ds_logic.v(2367)
  and u9700 (Ue2ju6, Dg2ju6, Kg2ju6);  // ../RTL/cortexm0ds_logic.v(9196)
  and u9701 (n2560, Yo1ju6, Rg2ju6);  // ../RTL/cortexm0ds_logic.v(9197)
  not u9702 (Kg2ju6, n2560);  // ../RTL/cortexm0ds_logic.v(9197)
  and u9703 (Dg2ju6, Yg2ju6, Fh2ju6);  // ../RTL/cortexm0ds_logic.v(9198)
  and u9704 (n2561, Mh2ju6, Htyiu6);  // ../RTL/cortexm0ds_logic.v(9199)
  not u9705 (Fh2ju6, n2561);  // ../RTL/cortexm0ds_logic.v(9199)
  and u9706 (Mh2ju6, Th2ju6, Ai2ju6);  // ../RTL/cortexm0ds_logic.v(9200)
  and u9707 (n2562, Xe0ju6, Hi2ju6);  // ../RTL/cortexm0ds_logic.v(9201)
  not u9708 (Ai2ju6, n2562);  // ../RTL/cortexm0ds_logic.v(9201)
  and u9709 (n2563, Zroiu6, Cwiiu6);  // ../RTL/cortexm0ds_logic.v(9202)
  buf u971 (E1hpw6[18], Naaax6);  // ../RTL/cortexm0ds_logic.v(2367)
  not u9710 (Hi2ju6, n2563);  // ../RTL/cortexm0ds_logic.v(9202)
  or u9711 (Yg2ju6, Oi2ju6, Y5ziu6);  // ../RTL/cortexm0ds_logic.v(9203)
  and u9712 (Y5ziu6, Vi2ju6, Cj2ju6);  // ../RTL/cortexm0ds_logic.v(9204)
  xor u9713 (Cj2ju6, Jj2ju6, Qj2ju6);  // ../RTL/cortexm0ds_logic.v(9205)
  and u9714 (Qj2ju6, Xj2ju6, Ek2ju6);  // ../RTL/cortexm0ds_logic.v(9206)
  or u9715 (n2564, G8niu6, Fp1ju6);  // ../RTL/cortexm0ds_logic.v(9207)
  not u9716 (Ek2ju6, n2564);  // ../RTL/cortexm0ds_logic.v(9207)
  and u9717 (G8niu6, P9niu6, vis_apsr_o[0]);  // ../RTL/cortexm0ds_logic.v(9208)
  and u9718 (Xj2ju6, Lk2ju6, Sk2ju6);  // ../RTL/cortexm0ds_logic.v(9209)
  or u9719 (Sk2ju6, D7fpw6[11], Qxoiu6);  // ../RTL/cortexm0ds_logic.v(9210)
  buf u972 (Mdhpw6[2], Golpw6);  // ../RTL/cortexm0ds_logic.v(1838)
  or u9720 (Lk2ju6, Zk2ju6, Gl2ju6);  // ../RTL/cortexm0ds_logic.v(9211)
  AL_MUX u9721 (
    .i0(Eafpw6[31]),
    .i1(Idfpw6[31]),
    .sel(Nl2ju6),
    .o(Gl2ju6));  // ../RTL/cortexm0ds_logic.v(9212)
  or u9722 (Zk2ju6, Ul2ju6, P9niu6);  // ../RTL/cortexm0ds_logic.v(9213)
  and u9723 (P9niu6, Bm2ju6, Im2ju6);  // ../RTL/cortexm0ds_logic.v(9214)
  and u9724 (Bm2ju6, Pm2ju6, Wm2ju6);  // ../RTL/cortexm0ds_logic.v(9215)
  and u9725 (n2565, Dn2ju6, Kn2ju6);  // ../RTL/cortexm0ds_logic.v(9216)
  not u9726 (Wm2ju6, n2565);  // ../RTL/cortexm0ds_logic.v(9216)
  or u9727 (n2566, Y2oiu6, Tfjiu6);  // ../RTL/cortexm0ds_logic.v(9217)
  not u9728 (Kn2ju6, n2566);  // ../RTL/cortexm0ds_logic.v(9217)
  or u9729 (n2567, Rn2ju6, Yn2ju6);  // ../RTL/cortexm0ds_logic.v(9218)
  buf u973 (Cyfpw6[0], Vzupw6);  // ../RTL/cortexm0ds_logic.v(1807)
  not u9730 (Dn2ju6, n2567);  // ../RTL/cortexm0ds_logic.v(9218)
  and u9731 (n2568, Fo2ju6, Mo2ju6);  // ../RTL/cortexm0ds_logic.v(9219)
  not u9732 (Pm2ju6, n2568);  // ../RTL/cortexm0ds_logic.v(9219)
  or u9733 (n2569, Jjhiu6, As0iu6);  // ../RTL/cortexm0ds_logic.v(9220)
  not u9734 (Fo2ju6, n2569);  // ../RTL/cortexm0ds_logic.v(9220)
  or u9735 (n2570, Idfpw6[31], Eafpw6[31]);  // ../RTL/cortexm0ds_logic.v(9221)
  not u9736 (Ul2ju6, n2570);  // ../RTL/cortexm0ds_logic.v(9221)
  or u9737 (n114[0], Hl0iu6, Cf0iu6);  // ../RTL/cortexm0ds_logic.v(3453)
  and u9738 (Cf0iu6, Ap2ju6, Hp2ju6);  // ../RTL/cortexm0ds_logic.v(9223)
  not u9739 (Oe0iu6, Cf0iu6);  // ../RTL/cortexm0ds_logic.v(9223)
  buf u974 (Krghu6, T2kbx6);  // ../RTL/cortexm0ds_logic.v(3093)
  and u9740 (Hp2ju6, Op2ju6, Vp2ju6);  // ../RTL/cortexm0ds_logic.v(9224)
  and u9741 (Vp2ju6, Cq2ju6, Owaiu6);  // ../RTL/cortexm0ds_logic.v(9225)
  and u9742 (n2571, Jq2ju6, K9aiu6);  // ../RTL/cortexm0ds_logic.v(9226)
  not u9743 (Cq2ju6, n2571);  // ../RTL/cortexm0ds_logic.v(9226)
  and u9744 (n2572, Knaiu6, Qq2ju6);  // ../RTL/cortexm0ds_logic.v(9227)
  not u9745 (Jq2ju6, n2572);  // ../RTL/cortexm0ds_logic.v(9227)
  or u9746 (Qq2ju6, Xe8iu6, Cyfpw6[4]);  // ../RTL/cortexm0ds_logic.v(9228)
  and u9747 (Op2ju6, Xq2ju6, Er2ju6);  // ../RTL/cortexm0ds_logic.v(9229)
  buf u9748 (Qvehu6, Ozkbx6[20]);  // ../RTL/cortexm0ds_logic.v(3176)
  and u9749 (n2573, F3aiu6, Ldoiu6);  // ../RTL/cortexm0ds_logic.v(9231)
  buf u975 (E1hpw6[15], Heaax6);  // ../RTL/cortexm0ds_logic.v(2367)
  not u9750 (Xq2ju6, n2573);  // ../RTL/cortexm0ds_logic.v(9231)
  and u9751 (Ap2ju6, Lr2ju6, Sr2ju6);  // ../RTL/cortexm0ds_logic.v(9232)
  and u9752 (Sr2ju6, H6ghu6, Zr2ju6);  // ../RTL/cortexm0ds_logic.v(9233)
  and u9753 (n2574, Pthiu6, H4ghu6);  // ../RTL/cortexm0ds_logic.v(9234)
  not u9754 (Zr2ju6, n2574);  // ../RTL/cortexm0ds_logic.v(9234)
  or u9755 (n2575, Gs2ju6, Ns2ju6);  // ../RTL/cortexm0ds_logic.v(9235)
  not u9756 (Lr2ju6, n2575);  // ../RTL/cortexm0ds_logic.v(9235)
  AL_MUX u9757 (
    .i0(Us2ju6),
    .i1(Bt2ju6),
    .sel(Cyfpw6[4]),
    .o(Ns2ju6));  // ../RTL/cortexm0ds_logic.v(9236)
  or u9758 (n2576, Wfoiu6, R75iu6);  // ../RTL/cortexm0ds_logic.v(9237)
  not u9759 (Bt2ju6, n2576);  // ../RTL/cortexm0ds_logic.v(9237)
  buf u976 (Mdhpw6[1], Vplpw6);  // ../RTL/cortexm0ds_logic.v(1838)
  AL_MUX u9760 (
    .i0(It2ju6),
    .i1(Pt2ju6),
    .sel(Cyfpw6[6]),
    .o(Gs2ju6));  // ../RTL/cortexm0ds_logic.v(9238)
  and u9761 (n2577, Wt2ju6, Du2ju6);  // ../RTL/cortexm0ds_logic.v(9239)
  not u9762 (Jj2ju6, n2577);  // ../RTL/cortexm0ds_logic.v(9239)
  AL_MUX u9763 (
    .i0(Vioiu6),
    .i1(Ku2ju6),
    .sel(Fhoiu6),
    .o(Du2ju6));  // ../RTL/cortexm0ds_logic.v(9240)
  not u9764 (Ku2ju6, vis_apsr_o[3]);  // ../RTL/cortexm0ds_logic.v(9241)
  AL_MUX u9765 (
    .i0(Bbliu6),
    .i1(Ru2ju6),
    .sel(E5ehu6),
    .o(Vioiu6));  // ../RTL/cortexm0ds_logic.v(9242)
  or u9766 (n2578, Fp1ju6, Zroiu6);  // ../RTL/cortexm0ds_logic.v(9243)
  not u9767 (Wt2ju6, n2578);  // ../RTL/cortexm0ds_logic.v(9243)
  and u9768 (Vi2ju6, Yu2ju6, Fv2ju6);  // ../RTL/cortexm0ds_logic.v(9244)
  or u9769 (Fv2ju6, Mv2ju6, Tv2ju6);  // ../RTL/cortexm0ds_logic.v(9245)
  buf u977 (Righu6, T8kbx6);  // ../RTL/cortexm0ds_logic.v(3096)
  AL_MUX u9770 (
    .i0(Ri8iu6),
    .i1(vis_apsr_o[1]),
    .sel(Ng8iu6),
    .o(Tv2ju6));  // ../RTL/cortexm0ds_logic.v(9246)
  and u9771 (Ng8iu6, Aw2ju6, Im2ju6);  // ../RTL/cortexm0ds_logic.v(9247)
  and u9772 (Im2ju6, Hw2ju6, Ow2ju6);  // ../RTL/cortexm0ds_logic.v(9248)
  and u9773 (n2579, Vw2ju6, Cx2ju6);  // ../RTL/cortexm0ds_logic.v(9249)
  not u9774 (Ow2ju6, n2579);  // ../RTL/cortexm0ds_logic.v(9249)
  and u9775 (Cx2ju6, Jx2ju6, Qx2ju6);  // ../RTL/cortexm0ds_logic.v(9250)
  and u9776 (n2580, Xx2ju6, Ey2ju6);  // ../RTL/cortexm0ds_logic.v(9251)
  not u9777 (Qx2ju6, n2580);  // ../RTL/cortexm0ds_logic.v(9251)
  or u9778 (Xx2ju6, Mr0iu6, Ly2ju6);  // ../RTL/cortexm0ds_logic.v(9252)
  or u9779 (n2581, Sy2ju6, Oiaiu6);  // ../RTL/cortexm0ds_logic.v(9253)
  buf u978 (Jydhu6, Qakbx6);  // ../RTL/cortexm0ds_logic.v(3097)
  not u9780 (Jx2ju6, n2581);  // ../RTL/cortexm0ds_logic.v(9253)
  and u9781 (Vw2ju6, C0ehu6, Zy2ju6);  // ../RTL/cortexm0ds_logic.v(9254)
  or u9782 (Zy2ju6, Y2oiu6, Qxaiu6);  // ../RTL/cortexm0ds_logic.v(9255)
  or u9783 (n2582, Gz2ju6, Nz2ju6);  // ../RTL/cortexm0ds_logic.v(9256)
  not u9784 (Hw2ju6, n2582);  // ../RTL/cortexm0ds_logic.v(9256)
  and u9785 (Aw2ju6, Uz2ju6, B03ju6);  // ../RTL/cortexm0ds_logic.v(9257)
  and u9786 (n2583, C0ehu6, I03ju6);  // ../RTL/cortexm0ds_logic.v(9258)
  not u9787 (B03ju6, n2583);  // ../RTL/cortexm0ds_logic.v(9258)
  and u9788 (n2584, P03ju6, O60ju6);  // ../RTL/cortexm0ds_logic.v(9259)
  not u9789 (I03ju6, n2584);  // ../RTL/cortexm0ds_logic.v(9259)
  buf u979 (vis_r4_o[16], V5vax6);  // ../RTL/cortexm0ds_logic.v(2626)
  and u9790 (n2585, Cyfpw6[4], W03ju6);  // ../RTL/cortexm0ds_logic.v(9260)
  not u9791 (Uz2ju6, n2585);  // ../RTL/cortexm0ds_logic.v(9260)
  and u9792 (n2586, D13ju6, K13ju6);  // ../RTL/cortexm0ds_logic.v(9261)
  not u9793 (W03ju6, n2586);  // ../RTL/cortexm0ds_logic.v(9261)
  or u9794 (K13ju6, Mr0iu6, Cyfpw6[7]);  // ../RTL/cortexm0ds_logic.v(9262)
  and u9795 (D13ju6, R13ju6, Y13ju6);  // ../RTL/cortexm0ds_logic.v(9263)
  and u9796 (n2587, F23ju6, M23ju6);  // ../RTL/cortexm0ds_logic.v(9264)
  not u9797 (Y13ju6, n2587);  // ../RTL/cortexm0ds_logic.v(9264)
  or u9798 (M23ju6, Ii0iu6, Pugiu6);  // ../RTL/cortexm0ds_logic.v(9265)
  and u9799 (n2588, T23ju6, Pfoiu6);  // ../RTL/cortexm0ds_logic.v(9266)
  buf u98 (vis_r2_o[0], A5qax6);  // ../RTL/cortexm0ds_logic.v(2551)
  buf u980 (SYSRESETREQ, Rekbx6);  // ../RTL/cortexm0ds_logic.v(3099)
  not u9800 (R13ju6, n2588);  // ../RTL/cortexm0ds_logic.v(9266)
  AL_MUX u9801 (
    .i0(Caehu6),
    .i1(A33ju6),
    .sel(E5ehu6),
    .o(Ri8iu6));  // ../RTL/cortexm0ds_logic.v(9267)
  and u9802 (n2589, H33ju6, O33ju6);  // ../RTL/cortexm0ds_logic.v(9268)
  not u9803 (A33ju6, n2589);  // ../RTL/cortexm0ds_logic.v(9268)
  and u9804 (n2590, V33ju6, C43ju6);  // ../RTL/cortexm0ds_logic.v(9269)
  not u9805 (O33ju6, n2590);  // ../RTL/cortexm0ds_logic.v(9269)
  and u9806 (C43ju6, J43ju6, vis_apsr_o[1]);  // ../RTL/cortexm0ds_logic.v(9270)
  or u9807 (n2591, Q43ju6, X43ju6);  // ../RTL/cortexm0ds_logic.v(9271)
  not u9808 (V33ju6, n2591);  // ../RTL/cortexm0ds_logic.v(9271)
  and u9809 (n2592, E53ju6, L53ju6);  // ../RTL/cortexm0ds_logic.v(9272)
  not u981 (Kaohu6, Rekbx6);  // ../RTL/cortexm0ds_logic.v(3100)
  not u9810 (H33ju6, n2592);  // ../RTL/cortexm0ds_logic.v(9272)
  and u9811 (n2593, S53ju6, Z53ju6);  // ../RTL/cortexm0ds_logic.v(9273)
  not u9812 (L53ju6, n2593);  // ../RTL/cortexm0ds_logic.v(9273)
  or u9813 (n2594, X43ju6, G63ju6);  // ../RTL/cortexm0ds_logic.v(9274)
  not u9814 (S53ju6, n2594);  // ../RTL/cortexm0ds_logic.v(9274)
  and u9815 (n2595, N63ju6, U63ju6);  // ../RTL/cortexm0ds_logic.v(9275)
  not u9816 (E53ju6, n2595);  // ../RTL/cortexm0ds_logic.v(9275)
  and u9817 (n2596, B73ju6, I73ju6);  // ../RTL/cortexm0ds_logic.v(9276)
  not u9818 (U63ju6, n2596);  // ../RTL/cortexm0ds_logic.v(9276)
  and u9819 (n2597, P73ju6, Cyfpw6[3]);  // ../RTL/cortexm0ds_logic.v(9277)
  buf u982 (Aygpw6[2], Dfbax6);  // ../RTL/cortexm0ds_logic.v(2278)
  not u9820 (I73ju6, n2597);  // ../RTL/cortexm0ds_logic.v(9277)
  and u9821 (B73ju6, W73ju6, Mr0iu6);  // ../RTL/cortexm0ds_logic.v(9278)
  and u9822 (n2598, D83ju6, K83ju6);  // ../RTL/cortexm0ds_logic.v(9279)
  not u9823 (W73ju6, n2598);  // ../RTL/cortexm0ds_logic.v(9279)
  and u9824 (n2599, R83ju6, Y83ju6);  // ../RTL/cortexm0ds_logic.v(9280)
  not u9825 (K83ju6, n2599);  // ../RTL/cortexm0ds_logic.v(9280)
  or u9826 (n2600, F93ju6, M93ju6);  // ../RTL/cortexm0ds_logic.v(9281)
  not u9827 (R83ju6, n2600);  // ../RTL/cortexm0ds_logic.v(9281)
  and u9828 (n2601, T93ju6, Aa3ju6);  // ../RTL/cortexm0ds_logic.v(9282)
  not u9829 (D83ju6, n2601);  // ../RTL/cortexm0ds_logic.v(9282)
  buf u983 (vis_r7_o[2], Tjvax6);  // ../RTL/cortexm0ds_logic.v(2654)
  and u9830 (n2602, Ha3ju6, Oa3ju6);  // ../RTL/cortexm0ds_logic.v(9283)
  not u9831 (Aa3ju6, n2602);  // ../RTL/cortexm0ds_logic.v(9283)
  AL_MUX u9832 (
    .i0(Va3ju6),
    .i1(Cb3ju6),
    .sel(F93ju6),
    .o(T93ju6));  // ../RTL/cortexm0ds_logic.v(9284)
  or u9833 (Cb3ju6, Jb3ju6, Oa3ju6);  // ../RTL/cortexm0ds_logic.v(9285)
  and u9834 (Va3ju6, Qb3ju6, M93ju6);  // ../RTL/cortexm0ds_logic.v(9286)
  AL_MUX u9835 (
    .i0(Xb3ju6),
    .i1(Ru2ju6),
    .sel(P73ju6),
    .o(N63ju6));  // ../RTL/cortexm0ds_logic.v(9287)
  and u9836 (P73ju6, Ec3ju6, Q43ju6);  // ../RTL/cortexm0ds_logic.v(9288)
  and u9837 (n2603, Lc3ju6, Sc3ju6);  // ../RTL/cortexm0ds_logic.v(9289)
  not u9838 (Ec3ju6, n2603);  // ../RTL/cortexm0ds_logic.v(9289)
  and u9839 (Lc3ju6, J43ju6, Zc3ju6);  // ../RTL/cortexm0ds_logic.v(9290)
  buf u984 (vis_r9_o[28], Rdibx6);  // ../RTL/cortexm0ds_logic.v(1898)
  not u9840 (J43ju6, G63ju6);  // ../RTL/cortexm0ds_logic.v(9291)
  and u9841 (Ru2ju6, Gd3ju6, Nd3ju6);  // ../RTL/cortexm0ds_logic.v(9292)
  and u9842 (Nd3ju6, Ud3ju6, Be3ju6);  // ../RTL/cortexm0ds_logic.v(9293)
  and u9843 (n2604, Ie3ju6, Pe3ju6);  // ../RTL/cortexm0ds_logic.v(9294)
  not u9844 (Be3ju6, n2604);  // ../RTL/cortexm0ds_logic.v(9294)
  or u9845 (n2605, We3ju6, Df3ju6);  // ../RTL/cortexm0ds_logic.v(9295)
  not u9846 (Ie3ju6, n2605);  // ../RTL/cortexm0ds_logic.v(9295)
  or u9847 (Ud3ju6, Kf3ju6, Ha3ju6);  // ../RTL/cortexm0ds_logic.v(9296)
  or u9848 (n2606, Rf3ju6, Yf3ju6);  // ../RTL/cortexm0ds_logic.v(9297)
  not u9849 (Gd3ju6, n2606);  // ../RTL/cortexm0ds_logic.v(9297)
  buf u985 (Gqgpw6[23], N3hbx6);  // ../RTL/cortexm0ds_logic.v(2377)
  or u9850 (n2607, Fg3ju6, Mg3ju6);  // ../RTL/cortexm0ds_logic.v(9298)
  not u9851 (Yf3ju6, n2607);  // ../RTL/cortexm0ds_logic.v(9298)
  AL_MUX u9852 (
    .i0(Jb3ju6),
    .i1(Tg3ju6),
    .sel(Ah3ju6),
    .o(Rf3ju6));  // ../RTL/cortexm0ds_logic.v(9299)
  and u9853 (Tg3ju6, Hh3ju6, Oh3ju6);  // ../RTL/cortexm0ds_logic.v(9300)
  and u9854 (Hh3ju6, Vh3ju6, Fg3ju6);  // ../RTL/cortexm0ds_logic.v(9301)
  and u9855 (n2608, H4ghu6, Ci3ju6);  // ../RTL/cortexm0ds_logic.v(9302)
  not u9856 (Xb3ju6, n2608);  // ../RTL/cortexm0ds_logic.v(9302)
  and u9857 (n2609, Ji3ju6, Qi3ju6);  // ../RTL/cortexm0ds_logic.v(9303)
  not u9858 (Ci3ju6, n2609);  // ../RTL/cortexm0ds_logic.v(9303)
  and u9859 (n2610, Xi3ju6, Ej3ju6);  // ../RTL/cortexm0ds_logic.v(9304)
  buf u986 (Qnghu6, Cokbx6);  // ../RTL/cortexm0ds_logic.v(3105)
  not u9860 (Qi3ju6, n2610);  // ../RTL/cortexm0ds_logic.v(9304)
  and u9861 (Xi3ju6, Lj3ju6, M93ju6);  // ../RTL/cortexm0ds_logic.v(9305)
  AL_MUX u9862 (
    .i0(Sj3ju6),
    .i1(Zj3ju6),
    .sel(M93ju6),
    .o(Ji3ju6));  // ../RTL/cortexm0ds_logic.v(9306)
  and u9863 (n2611, F93ju6, Gk3ju6);  // ../RTL/cortexm0ds_logic.v(9307)
  not u9864 (Zj3ju6, n2611);  // ../RTL/cortexm0ds_logic.v(9307)
  AL_MUX u9865 (
    .i0(Nk3ju6),
    .i1(Uk3ju6),
    .sel(Ej3ju6),
    .o(Sj3ju6));  // ../RTL/cortexm0ds_logic.v(9308)
  and u9866 (n2612, Bl3ju6, I6jiu6);  // ../RTL/cortexm0ds_logic.v(9309)
  not u9867 (Mv2ju6, n2612);  // ../RTL/cortexm0ds_logic.v(9309)
  or u9868 (Bl3ju6, Zroiu6, Il3ju6);  // ../RTL/cortexm0ds_logic.v(9310)
  and u9869 (n2613, Pl3ju6, Wl3ju6);  // ../RTL/cortexm0ds_logic.v(9311)
  buf u987 (SWDOEN, Dqkbx6);  // ../RTL/cortexm0ds_logic.v(3106)
  not u9870 (Yu2ju6, n2613);  // ../RTL/cortexm0ds_logic.v(9311)
  or u9871 (Wl3ju6, Fp1ju6, Il3ju6);  // ../RTL/cortexm0ds_logic.v(9312)
  xor u9872 (Pl3ju6, Xe0ju6, Dm3ju6);  // ../RTL/cortexm0ds_logic.v(9313)
  AL_MUX u9873 (
    .i0(V7liu6),
    .i1(Km3ju6),
    .sel(Fhoiu6),
    .o(Dm3ju6));  // ../RTL/cortexm0ds_logic.v(9314)
  and u9874 (Fhoiu6, Rm3ju6, Mwniu6);  // ../RTL/cortexm0ds_logic.v(9315)
  or u9875 (Mwniu6, Szniu6, Yn2ju6);  // ../RTL/cortexm0ds_logic.v(9316)
  and u9876 (n2614, C0ehu6, Ym3ju6);  // ../RTL/cortexm0ds_logic.v(9317)
  not u9877 (Rm3ju6, n2614);  // ../RTL/cortexm0ds_logic.v(9317)
  and u9878 (n2615, Fn3ju6, Mn3ju6);  // ../RTL/cortexm0ds_logic.v(9318)
  not u9879 (Ym3ju6, n2615);  // ../RTL/cortexm0ds_logic.v(9318)
  buf u988 (R4gpw6[37], Nazax6);  // ../RTL/cortexm0ds_logic.v(2815)
  and u9880 (Mn3ju6, Tn3ju6, Ao3ju6);  // ../RTL/cortexm0ds_logic.v(9319)
  and u9881 (n2616, H4ghu6, Ho3ju6);  // ../RTL/cortexm0ds_logic.v(9320)
  not u9882 (Ao3ju6, n2616);  // ../RTL/cortexm0ds_logic.v(9320)
  and u9883 (n2617, Oo3ju6, Vo3ju6);  // ../RTL/cortexm0ds_logic.v(9321)
  not u9884 (Ho3ju6, n2617);  // ../RTL/cortexm0ds_logic.v(9321)
  or u9885 (n2618, Hs0iu6, Cp3ju6);  // ../RTL/cortexm0ds_logic.v(9322)
  not u9886 (Oo3ju6, n2618);  // ../RTL/cortexm0ds_logic.v(9322)
  and u9887 (Tn3ju6, Jp3ju6, Qp3ju6);  // ../RTL/cortexm0ds_logic.v(9323)
  and u9888 (n2619, Ly2ju6, Cyfpw6[4]);  // ../RTL/cortexm0ds_logic.v(9324)
  not u9889 (Jp3ju6, n2619);  // ../RTL/cortexm0ds_logic.v(9324)
  buf u989 (R4gpw6[38], Pczax6);  // ../RTL/cortexm0ds_logic.v(2815)
  and u9890 (Fn3ju6, Xp3ju6, Eq3ju6);  // ../RTL/cortexm0ds_logic.v(9325)
  or u9891 (Eq3ju6, Ezniu6, Cyfpw6[6]);  // ../RTL/cortexm0ds_logic.v(9326)
  and u9892 (Xp3ju6, Lq3ju6, P03ju6);  // ../RTL/cortexm0ds_logic.v(9327)
  and u9893 (n2620, Sq3ju6, Hs0iu6);  // ../RTL/cortexm0ds_logic.v(9328)
  not u9894 (P03ju6, n2620);  // ../RTL/cortexm0ds_logic.v(9328)
  or u9895 (Lq3ju6, Ey2ju6, As0iu6);  // ../RTL/cortexm0ds_logic.v(9329)
  not u9896 (Km3ju6, vis_apsr_o[2]);  // ../RTL/cortexm0ds_logic.v(9330)
  AL_MUX u9897 (
    .i0(Zq3ju6),
    .i1(Gr3ju6),
    .sel(E5ehu6),
    .o(V7liu6));  // ../RTL/cortexm0ds_logic.v(9331)
  and u9898 (n2621, Nr3ju6, Ur3ju6);  // ../RTL/cortexm0ds_logic.v(9332)
  not u9899 (Gr3ju6, n2621);  // ../RTL/cortexm0ds_logic.v(9332)
  buf u99 (Stdhu6, Fnnpw6);  // ../RTL/cortexm0ds_logic.v(1878)
  buf u990 (R4gpw6[39], Rezax6);  // ../RTL/cortexm0ds_logic.v(2815)
  and u9900 (Ur3ju6, Bs3ju6, Is3ju6);  // ../RTL/cortexm0ds_logic.v(9333)
  and u9901 (n2622, Ps3ju6, Ws3ju6);  // ../RTL/cortexm0ds_logic.v(9334)
  not u9902 (Is3ju6, n2622);  // ../RTL/cortexm0ds_logic.v(9334)
  and u9903 (n2623, Dt3ju6, Kt3ju6);  // ../RTL/cortexm0ds_logic.v(9335)
  not u9904 (Ws3ju6, n2623);  // ../RTL/cortexm0ds_logic.v(9335)
  and u9905 (Kt3ju6, Rt3ju6, Yt3ju6);  // ../RTL/cortexm0ds_logic.v(9336)
  or u9906 (n2624, Lj3ju6, Jb3ju6);  // ../RTL/cortexm0ds_logic.v(9337)
  not u9907 (Rt3ju6, n2624);  // ../RTL/cortexm0ds_logic.v(9337)
  and u9908 (Dt3ju6, Fu3ju6, Mu3ju6);  // ../RTL/cortexm0ds_logic.v(9338)
  AL_MUX u9909 (
    .i0(Tu3ju6),
    .i1(Av3ju6),
    .sel(Hv3ju6),
    .o(Fu3ju6));  // ../RTL/cortexm0ds_logic.v(9339)
  buf u991 (R4gpw6[40], T3abx6);  // ../RTL/cortexm0ds_logic.v(2815)
  and u9910 (Av3ju6, Ov3ju6, Vv3ju6);  // ../RTL/cortexm0ds_logic.v(9340)
  or u9911 (n2625, Cw3ju6, Jw3ju6);  // ../RTL/cortexm0ds_logic.v(9341)
  not u9912 (Vv3ju6, n2625);  // ../RTL/cortexm0ds_logic.v(9341)
  and u9913 (Tu3ju6, Qw3ju6, Xw3ju6);  // ../RTL/cortexm0ds_logic.v(9342)
  or u9914 (n2626, Ex3ju6, Lx3ju6);  // ../RTL/cortexm0ds_logic.v(9343)
  not u9915 (Xw3ju6, n2626);  // ../RTL/cortexm0ds_logic.v(9343)
  or u9916 (n2627, Sx3ju6, Zx3ju6);  // ../RTL/cortexm0ds_logic.v(9344)
  not u9917 (Qw3ju6, n2627);  // ../RTL/cortexm0ds_logic.v(9344)
  and u9918 (n2628, Gy3ju6, Oh3ju6);  // ../RTL/cortexm0ds_logic.v(9345)
  not u9919 (Ps3ju6, n2628);  // ../RTL/cortexm0ds_logic.v(9345)
  buf u992 (R4gpw6[41], Mfyax6);  // ../RTL/cortexm0ds_logic.v(2815)
  and u9920 (Gy3ju6, Ah3ju6, Ny3ju6);  // ../RTL/cortexm0ds_logic.v(9346)
  and u9921 (Bs3ju6, Uy3ju6, Bz3ju6);  // ../RTL/cortexm0ds_logic.v(9347)
  and u9922 (n2629, Iz3ju6, Pz3ju6);  // ../RTL/cortexm0ds_logic.v(9348)
  not u9923 (Uy3ju6, n2629);  // ../RTL/cortexm0ds_logic.v(9348)
  and u9924 (n2630, Wz3ju6, D04ju6);  // ../RTL/cortexm0ds_logic.v(9349)
  not u9925 (Pz3ju6, n2630);  // ../RTL/cortexm0ds_logic.v(9349)
  and u9926 (D04ju6, K04ju6, R04ju6);  // ../RTL/cortexm0ds_logic.v(9350)
  and u9927 (K04ju6, Ha3ju6, Uk3ju6);  // ../RTL/cortexm0ds_logic.v(9351)
  and u9928 (Wz3ju6, Y04ju6, F14ju6);  // ../RTL/cortexm0ds_logic.v(9352)
  AL_MUX u9929 (
    .i0(M14ju6),
    .i1(T14ju6),
    .sel(Hv3ju6),
    .o(Y04ju6));  // ../RTL/cortexm0ds_logic.v(9353)
  buf u993 (R4gpw6[42], Ohyax6);  // ../RTL/cortexm0ds_logic.v(2815)
  and u9930 (T14ju6, A24ju6, H24ju6);  // ../RTL/cortexm0ds_logic.v(9354)
  or u9931 (n2631, O24ju6, V24ju6);  // ../RTL/cortexm0ds_logic.v(9355)
  not u9932 (H24ju6, n2631);  // ../RTL/cortexm0ds_logic.v(9355)
  and u9933 (A24ju6, C34ju6, J34ju6);  // ../RTL/cortexm0ds_logic.v(9356)
  and u9934 (M14ju6, Q34ju6, X34ju6);  // ../RTL/cortexm0ds_logic.v(9357)
  or u9935 (n2632, E44ju6, L44ju6);  // ../RTL/cortexm0ds_logic.v(9358)
  not u9936 (X34ju6, n2632);  // ../RTL/cortexm0ds_logic.v(9358)
  and u9937 (n2633, S44ju6, Kf3ju6);  // ../RTL/cortexm0ds_logic.v(9359)
  not u9938 (Iz3ju6, n2633);  // ../RTL/cortexm0ds_logic.v(9359)
  and u9939 (S44ju6, Z44ju6, Ny3ju6);  // ../RTL/cortexm0ds_logic.v(9360)
  buf u994 (R4gpw6[43], Qjyax6);  // ../RTL/cortexm0ds_logic.v(2815)
  and u9940 (Nr3ju6, G54ju6, N54ju6);  // ../RTL/cortexm0ds_logic.v(9361)
  and u9941 (n2634, U54ju6, B64ju6);  // ../RTL/cortexm0ds_logic.v(9362)
  not u9942 (N54ju6, n2634);  // ../RTL/cortexm0ds_logic.v(9362)
  and u9943 (n2635, I64ju6, P64ju6);  // ../RTL/cortexm0ds_logic.v(9363)
  not u9944 (B64ju6, n2635);  // ../RTL/cortexm0ds_logic.v(9363)
  and u9945 (P64ju6, W64ju6, D74ju6);  // ../RTL/cortexm0ds_logic.v(9364)
  and u9946 (D74ju6, K74ju6, R74ju6);  // ../RTL/cortexm0ds_logic.v(9365)
  and u9947 (n2636, Hv3ju6, Y74ju6);  // ../RTL/cortexm0ds_logic.v(9366)
  not u9948 (R74ju6, n2636);  // ../RTL/cortexm0ds_logic.v(9366)
  or u9949 (Y74ju6, F84ju6, M84ju6);  // ../RTL/cortexm0ds_logic.v(9367)
  buf u995 (R4gpw6[44], Lfgbx6);  // ../RTL/cortexm0ds_logic.v(2815)
  and u9950 (K74ju6, T84ju6, A94ju6);  // ../RTL/cortexm0ds_logic.v(9368)
  and u9951 (W64ju6, H94ju6, O94ju6);  // ../RTL/cortexm0ds_logic.v(9369)
  and u9952 (n2637, M84ju6, V94ju6);  // ../RTL/cortexm0ds_logic.v(9370)
  not u9953 (H94ju6, n2637);  // ../RTL/cortexm0ds_logic.v(9370)
  and u9954 (I64ju6, Ca4ju6, Ja4ju6);  // ../RTL/cortexm0ds_logic.v(9371)
  and u9955 (Ja4ju6, Mg3ju6, Qa4ju6);  // ../RTL/cortexm0ds_logic.v(9372)
  and u9956 (n2638, F84ju6, O24ju6);  // ../RTL/cortexm0ds_logic.v(9373)
  not u9957 (Qa4ju6, n2638);  // ../RTL/cortexm0ds_logic.v(9373)
  or u9958 (n2639, Xa4ju6, Eb4ju6);  // ../RTL/cortexm0ds_logic.v(9374)
  not u9959 (Ca4ju6, n2639);  // ../RTL/cortexm0ds_logic.v(9374)
  buf u996 (R4gpw6[45], Slyax6);  // ../RTL/cortexm0ds_logic.v(2815)
  and u9960 (n2640, Lb4ju6, Sb4ju6);  // ../RTL/cortexm0ds_logic.v(9375)
  not u9961 (G54ju6, n2640);  // ../RTL/cortexm0ds_logic.v(9375)
  and u9962 (n2641, Zb4ju6, Gc4ju6);  // ../RTL/cortexm0ds_logic.v(9376)
  not u9963 (Sb4ju6, n2641);  // ../RTL/cortexm0ds_logic.v(9376)
  and u9964 (Gc4ju6, Nc4ju6, Uc4ju6);  // ../RTL/cortexm0ds_logic.v(9377)
  or u9965 (n2642, Gk3ju6, Y83ju6);  // ../RTL/cortexm0ds_logic.v(9378)
  not u9966 (Nc4ju6, n2642);  // ../RTL/cortexm0ds_logic.v(9378)
  and u9967 (Zb4ju6, Bd4ju6, Id4ju6);  // ../RTL/cortexm0ds_logic.v(9379)
  AL_MUX u9968 (
    .i0(Pd4ju6),
    .i1(Wd4ju6),
    .sel(Hv3ju6),
    .o(Bd4ju6));  // ../RTL/cortexm0ds_logic.v(9380)
  and u9969 (Wd4ju6, Q34ju6, De4ju6);  // ../RTL/cortexm0ds_logic.v(9381)
  buf u997 (R4gpw6[46], Unyax6);  // ../RTL/cortexm0ds_logic.v(2815)
  or u9970 (n2643, Ke4ju6, Re4ju6);  // ../RTL/cortexm0ds_logic.v(9382)
  not u9971 (De4ju6, n2643);  // ../RTL/cortexm0ds_logic.v(9382)
  or u9972 (n2644, Ye4ju6, Ff4ju6);  // ../RTL/cortexm0ds_logic.v(9383)
  not u9973 (Q34ju6, n2644);  // ../RTL/cortexm0ds_logic.v(9383)
  and u9974 (Pd4ju6, Ov3ju6, Mf4ju6);  // ../RTL/cortexm0ds_logic.v(9384)
  or u9975 (n2645, Tf4ju6, Ag4ju6);  // ../RTL/cortexm0ds_logic.v(9385)
  not u9976 (Mf4ju6, n2645);  // ../RTL/cortexm0ds_logic.v(9385)
  or u9977 (n2646, Hg4ju6, Og4ju6);  // ../RTL/cortexm0ds_logic.v(9386)
  not u9978 (Ov3ju6, n2646);  // ../RTL/cortexm0ds_logic.v(9386)
  and u9979 (n2647, Vg4ju6, Oh3ju6);  // ../RTL/cortexm0ds_logic.v(9387)
  buf u998 (R4gpw6[47], Wpyax6);  // ../RTL/cortexm0ds_logic.v(2815)
  not u9980 (Lb4ju6, n2647);  // ../RTL/cortexm0ds_logic.v(9387)
  and u9981 (Vg4ju6, Ch4ju6, Ny3ju6);  // ../RTL/cortexm0ds_logic.v(9388)
  and u9982 (n2648, Jh4ju6, Qh4ju6);  // ../RTL/cortexm0ds_logic.v(9389)
  not u9983 (Zq3ju6, n2648);  // ../RTL/cortexm0ds_logic.v(9389)
  and u9984 (Qh4ju6, Xh4ju6, Ei4ju6);  // ../RTL/cortexm0ds_logic.v(9390)
  and u9985 (Ei4ju6, Li4ju6, Si4ju6);  // ../RTL/cortexm0ds_logic.v(9391)
  and u9986 (Si4ju6, Zi4ju6, Gj4ju6);  // ../RTL/cortexm0ds_logic.v(9392)
  and u9987 (Gj4ju6, Ibliu6, Kkkiu6);  // ../RTL/cortexm0ds_logic.v(9393)
  and u9988 (Kkkiu6, Nj4ju6, Uj4ju6);  // ../RTL/cortexm0ds_logic.v(9394)
  and u9989 (Uj4ju6, Bk4ju6, Ik4ju6);  // ../RTL/cortexm0ds_logic.v(9395)
  buf u999 (R4gpw6[48], R1abx6);  // ../RTL/cortexm0ds_logic.v(2815)
  and u9990 (n2649, Pk4ju6, vis_ipsr_o[4]);  // ../RTL/cortexm0ds_logic.v(9396)
  not u9991 (Ik4ju6, n2649);  // ../RTL/cortexm0ds_logic.v(9396)
  or u9992 (n2650, Affpw6[4], Wk4ju6);  // ../RTL/cortexm0ds_logic.v(9397)
  not u9993 (Bk4ju6, n2650);  // ../RTL/cortexm0ds_logic.v(9397)
  and u9994 (Nj4ju6, Dl4ju6, Kl4ju6);  // ../RTL/cortexm0ds_logic.v(9398)
  AL_MUX u9995 (
    .i0(Rl4ju6),
    .i1(Yl4ju6),
    .sel(Eg0iu6),
    .o(Kl4ju6));  // ../RTL/cortexm0ds_logic.v(9399)
  AL_MUX u9996 (
    .i0(V3iiu6),
    .i1(Fm4ju6),
    .sel(Mm4ju6),
    .o(Eg0iu6));  // ../RTL/cortexm0ds_logic.v(9400)
  and u9997 (Fm4ju6, Tm4ju6, An4ju6);  // ../RTL/cortexm0ds_logic.v(9401)
  and u9998 (An4ju6, Hn4ju6, On4ju6);  // ../RTL/cortexm0ds_logic.v(9402)
  and u9999 (On4ju6, Vn4ju6, Co4ju6);  // ../RTL/cortexm0ds_logic.v(9403)

endmodule 

module eq_w12
  (
  i0,
  i1,
  o
  );

  input [11:0] i0;
  input [11:0] i1;
  output o;



endmodule 

module reg_ar_as_w12
  (
  clk,
  d,
  en,
  reset,
  set,
  q
  );

  input clk;
  input [11:0] d;
  input en;
  input [11:0] reset;
  input [11:0] set;
  output [11:0] q;



endmodule 

module eq_w4
  (
  i0,
  i1,
  o
  );

  input [3:0] i0;
  input [3:0] i1;
  output o;



endmodule 

module binary_mux_s1_w8
  (
  i0,
  i1,
  sel,
  o
  );

  input [7:0] i0;
  input [7:0] i1;
  input sel;
  output [7:0] o;



endmodule 

module binary_mux_s1_w16
  (
  i0,
  i1,
  sel,
  o
  );

  input [15:0] i0;
  input [15:0] i1;
  input sel;
  output [15:0] o;



endmodule 

module reg_ar_as_w16
  (
  clk,
  d,
  en,
  reset,
  set,
  q
  );

  input clk;
  input [15:0] d;
  input en;
  input [15:0] reset;
  input [15:0] set;
  output [15:0] q;



endmodule 

module gpio_apbif  // ../RTL/gpio_apbif.v(39)
  (
  gpio_ext_porta_rb,
  gpio_intstatus,
  gpio_raw_intstatus,
  paddr,
  pclk,
  penable,
  presetn,
  psel,
  pwdata,
  pwrite,
  gpio_int_polarity,
  gpio_inten,
  gpio_intmask,
  gpio_inttype_level,
  gpio_ls_sync,
  gpio_porta_eoi,
  gpio_swporta_ctl,
  gpio_swporta_ddr,
  gpio_swporta_dr,
  prdata
  );

  input [7:0] gpio_ext_porta_rb;  // ../RTL/gpio_apbif.v(63)
  input [7:0] gpio_intstatus;  // ../RTL/gpio_apbif.v(64)
  input [7:0] gpio_raw_intstatus;  // ../RTL/gpio_apbif.v(65)
  input [6:2] paddr;  // ../RTL/gpio_apbif.v(66)
  input pclk;  // ../RTL/gpio_apbif.v(67)
  input penable;  // ../RTL/gpio_apbif.v(68)
  input presetn;  // ../RTL/gpio_apbif.v(69)
  input psel;  // ../RTL/gpio_apbif.v(70)
  input [31:0] pwdata;  // ../RTL/gpio_apbif.v(71)
  input pwrite;  // ../RTL/gpio_apbif.v(72)
  output [7:0] gpio_int_polarity;  // ../RTL/gpio_apbif.v(73)
  output [7:0] gpio_inten;  // ../RTL/gpio_apbif.v(74)
  output [7:0] gpio_intmask;  // ../RTL/gpio_apbif.v(75)
  output [7:0] gpio_inttype_level;  // ../RTL/gpio_apbif.v(76)
  output gpio_ls_sync;  // ../RTL/gpio_apbif.v(77)
  output [7:0] gpio_porta_eoi;  // ../RTL/gpio_apbif.v(78)
  output [7:0] gpio_swporta_ctl;  // ../RTL/gpio_apbif.v(79)
  output [7:0] gpio_swporta_ddr;  // ../RTL/gpio_apbif.v(80)
  output [7:0] gpio_swporta_dr;  // ../RTL/gpio_apbif.v(81)
  output [31:0] prdata;  // ../RTL/gpio_apbif.v(82)

  wire [3:0] gpio_int_polarity_wen;  // ../RTL/gpio_apbif.v(85)
  wire [3:0] gpio_inten_wen;  // ../RTL/gpio_apbif.v(86)
  wire [3:0] gpio_intmask_wen;  // ../RTL/gpio_apbif.v(87)
  wire [3:0] gpio_inttype_level_wen;  // ../RTL/gpio_apbif.v(88)
  wire [3:0] gpio_ls_sync_wen;  // ../RTL/gpio_apbif.v(89)
  wire [3:0] gpio_porta_eoi_wen;  // ../RTL/gpio_apbif.v(90)
  wire [3:0] gpio_swporta_ctl_wen;  // ../RTL/gpio_apbif.v(91)
  wire [3:0] gpio_swporta_ddr_wen;  // ../RTL/gpio_apbif.v(92)
  wire [3:0] gpio_swporta_dr_wen;  // ../RTL/gpio_apbif.v(93)
  wire [31:0] int_gpio_int_polarity;  // ../RTL/gpio_apbif.v(94)
  wire [31:0] int_gpio_inten;  // ../RTL/gpio_apbif.v(95)
  wire [31:0] int_gpio_intmask;  // ../RTL/gpio_apbif.v(96)
  wire [31:0] int_gpio_inttype_level;  // ../RTL/gpio_apbif.v(97)
  wire [31:0] int_gpio_ls_sync;  // ../RTL/gpio_apbif.v(98)
  wire [31:0] int_gpio_porta_eoi;  // ../RTL/gpio_apbif.v(99)
  wire [31:0] int_gpio_swporta_ctl;  // ../RTL/gpio_apbif.v(100)
  wire [31:0] int_gpio_swporta_ddr;  // ../RTL/gpio_apbif.v(101)
  wire [31:0] int_gpio_swporta_dr;  // ../RTL/gpio_apbif.v(102)
  wire [31:0] iprdata;  // ../RTL/gpio_apbif.v(103)
  wire [3:0] n13;
  wire [3:0] n14;
  wire [3:0] n15;
  wire [3:0] n19;
  wire [3:0] n20;
  wire [3:0] n21;
  wire [3:0] n26;
  wire [3:0] n27;
  wire [3:0] n28;
  wire [3:0] n29;
  wire [3:0] n34;
  wire [3:0] n35;
  wire [3:0] n36;
  wire [3:0] n37;
  wire [3:0] n38;
  wire [3:0] n4;
  wire [31:0] n41;
  wire [31:0] n44;
  wire [31:0] n47;
  wire [31:0] n50;
  wire [31:0] n53;
  wire [31:0] n56;
  wire [31:0] n59;
  wire [31:0] n62;
  wire [31:0] n81;
  wire [31:0] n82;
  wire [31:0] pwdata_int;  // ../RTL/gpio_apbif.v(105)
  wire [31:0] ri_gpio_ext_porta_rb;  // ../RTL/gpio_apbif.v(106)
  wire [31:0] ri_gpio_int_polarity;  // ../RTL/gpio_apbif.v(107)
  wire [31:0] ri_gpio_inten;  // ../RTL/gpio_apbif.v(108)
  wire [31:0] ri_gpio_intmask;  // ../RTL/gpio_apbif.v(109)
  wire [31:0] ri_gpio_intstatus;  // ../RTL/gpio_apbif.v(110)
  wire [31:0] ri_gpio_inttype_level;  // ../RTL/gpio_apbif.v(111)
  wire [31:0] ri_gpio_ls_sync;  // ../RTL/gpio_apbif.v(112)
  wire [31:0] ri_gpio_raw_intstatus;  // ../RTL/gpio_apbif.v(113)
  wire [31:0] ri_gpio_swporta_ctl;  // ../RTL/gpio_apbif.v(114)
  wire [31:0] ri_gpio_swporta_ddr;  // ../RTL/gpio_apbif.v(115)
  wire [31:0] ri_gpio_swporta_dr;  // ../RTL/gpio_apbif.v(116)
  wire n0;
  wire n1;
  wire n10;
  wire n11;
  wire n12;
  wire n16;
  wire n17;
  wire n18;
  wire n2;
  wire n22;
  wire n23;
  wire n24;
  wire n25;
  wire n3;
  wire n30;
  wire n31;
  wire n32;
  wire n33;
  wire n39;
  wire n40;
  wire n42;
  wire n43;
  wire n45;
  wire n46;
  wire n48;
  wire n49;
  wire n5;
  wire n51;
  wire n52;
  wire n54;
  wire n55;
  wire n57;
  wire n58;
  wire n6;
  wire n60;
  wire n61;
  wire n63;
  wire n64;
  wire n65;
  wire n66;
  wire n67;
  wire n68;
  wire n69;
  wire n7;
  wire n70;
  wire n71;
  wire n72;
  wire n73;
  wire n74;
  wire n75;
  wire n76;
  wire n77;
  wire n78;
  wire n79;
  wire n8;
  wire n80;
  wire n9;

  eq_w5 eq0 (
    .i0(paddr),
    .i1(5'b00000),
    .o(n2));  // ../RTL/gpio_apbif.v(164)
  eq_w5 eq1 (
    .i0(paddr),
    .i1(5'b00001),
    .o(n3));  // ../RTL/gpio_apbif.v(169)
  eq_w5 eq10 (
    .i0(paddr),
    .i1(5'b10001),
    .o(n77));  // ../RTL/gpio_apbif.v(449)
  eq_w5 eq11 (
    .i0(paddr),
    .i1(5'b10100),
    .o(n79));  // ../RTL/gpio_apbif.v(451)
  eq_w5 eq2 (
    .i0(paddr),
    .i1(5'b01100),
    .o(n7));  // ../RTL/gpio_apbif.v(202)
  eq_w5 eq3 (
    .i0(paddr),
    .i1(5'b01101),
    .o(n8));  // ../RTL/gpio_apbif.v(207)
  eq_w5 eq4 (
    .i0(paddr),
    .i1(5'b01110),
    .o(n9));  // ../RTL/gpio_apbif.v(212)
  eq_w5 eq5 (
    .i0(paddr),
    .i1(5'b01111),
    .o(n10));  // ../RTL/gpio_apbif.v(217)
  eq_w5 eq6 (
    .i0(paddr),
    .i1(5'b11000),
    .o(n11));  // ../RTL/gpio_apbif.v(222)
  eq_w5 eq7 (
    .i0(paddr),
    .i1(5'b10011),
    .o(n12));  // ../RTL/gpio_apbif.v(227)
  eq_w5 eq8 (
    .i0(paddr),
    .i1(5'b00010),
    .o(n71));  // ../RTL/gpio_apbif.v(443)
  eq_w5 eq9 (
    .i0(paddr),
    .i1(5'b10000),
    .o(n76));  // ../RTL/gpio_apbif.v(448)
  binary_mux_s1_w4 mux0 (
    .i0({n3,n3,n3,n3}),
    .i1(4'b0000),
    .sel(n2),
    .o(n4));  // ../RTL/gpio_apbif.v(177)
  binary_mux_s1_w4 mux1 (
    .i0(4'b0000),
    .i1({n2,n2,n2,n2}),
    .sel(n6),
    .o(gpio_swporta_dr_wen));  // ../RTL/gpio_apbif.v(178)
  binary_mux_s1_w4 mux10 (
    .i0(n19),
    .i1(4'b0000),
    .sel(n8),
    .o(n27));  // ../RTL/gpio_apbif.v(230)
  binary_mux_s1_w4 mux11 (
    .i0(n20),
    .i1(4'b0000),
    .sel(n8),
    .o(n28));  // ../RTL/gpio_apbif.v(230)
  binary_mux_s1_w4 mux12 (
    .i0(n21),
    .i1(4'b0000),
    .sel(n8),
    .o(n29));  // ../RTL/gpio_apbif.v(230)
  binary_mux_s1_w4 mux13 (
    .i0({n8,n8,n8,n8}),
    .i1(4'b0000),
    .sel(n7),
    .o(n34));  // ../RTL/gpio_apbif.v(230)
  binary_mux_s1_w4 mux14 (
    .i0(n26),
    .i1(4'b0000),
    .sel(n7),
    .o(n35));  // ../RTL/gpio_apbif.v(230)
  binary_mux_s1_w4 mux15 (
    .i0(n27),
    .i1(4'b0000),
    .sel(n7),
    .o(n36));  // ../RTL/gpio_apbif.v(230)
  binary_mux_s1_w4 mux16 (
    .i0(n28),
    .i1(4'b0000),
    .sel(n7),
    .o(n37));  // ../RTL/gpio_apbif.v(230)
  binary_mux_s1_w4 mux17 (
    .i0(n29),
    .i1(4'b0000),
    .sel(n7),
    .o(n38));  // ../RTL/gpio_apbif.v(230)
  binary_mux_s1_w4 mux18 (
    .i0(4'b0000),
    .i1({n7,n7,n7,n7}),
    .sel(n6),
    .o(gpio_inten_wen));  // ../RTL/gpio_apbif.v(231)
  binary_mux_s1_w4 mux19 (
    .i0(4'b0000),
    .i1(n34),
    .sel(n6),
    .o(gpio_intmask_wen));  // ../RTL/gpio_apbif.v(231)
  binary_mux_s1_w4 mux2 (
    .i0(4'b0000),
    .i1(n4),
    .sel(n6),
    .o(gpio_swporta_ddr_wen));  // ../RTL/gpio_apbif.v(178)
  binary_mux_s1_w4 mux20 (
    .i0(4'b0000),
    .i1(n35),
    .sel(n6),
    .o(gpio_inttype_level_wen));  // ../RTL/gpio_apbif.v(231)
  binary_mux_s1_w4 mux21 (
    .i0(4'b0000),
    .i1(n36),
    .sel(n6),
    .o(gpio_int_polarity_wen));  // ../RTL/gpio_apbif.v(231)
  binary_mux_s1_w4 mux22 (
    .i0(4'b0000),
    .i1(n37),
    .sel(n6),
    .o(gpio_ls_sync_wen));  // ../RTL/gpio_apbif.v(231)
  binary_mux_s1_w4 mux23 (
    .i0(4'b0000),
    .i1(n38),
    .sel(n6),
    .o(gpio_porta_eoi_wen));  // ../RTL/gpio_apbif.v(231)
  binary_mux_s1_w32 mux24 (
    .i0(int_gpio_swporta_dr),
    .i1(pwdata_int),
    .sel(n40),
    .o(n41));  // ../RTL/gpio_apbif.v(242)
  binary_mux_s1_w32 mux25 (
    .i0(int_gpio_swporta_ddr),
    .i1(pwdata_int),
    .sel(n43),
    .o(n44));  // ../RTL/gpio_apbif.v(262)
  binary_mux_s1_w32 mux26 (
    .i0(int_gpio_swporta_ctl),
    .i1(pwdata_int),
    .sel(n46),
    .o(n47));  // ../RTL/gpio_apbif.v(282)
  binary_mux_s1_w32 mux27 (
    .i0(int_gpio_inten),
    .i1(pwdata_int),
    .sel(n49),
    .o(n50));  // ../RTL/gpio_apbif.v(303)
  binary_mux_s1_w32 mux28 (
    .i0(int_gpio_intmask),
    .i1(pwdata_int),
    .sel(n52),
    .o(n53));  // ../RTL/gpio_apbif.v(323)
  binary_mux_s1_w32 mux29 (
    .i0(int_gpio_inttype_level),
    .i1(pwdata_int),
    .sel(n55),
    .o(n56));  // ../RTL/gpio_apbif.v(343)
  binary_mux_s1_w4 mux3 (
    .i0({n12,n12,n12,n12}),
    .i1(4'b0000),
    .sel(n11),
    .o(n13));  // ../RTL/gpio_apbif.v(230)
  binary_mux_s1_w32 mux30 (
    .i0(int_gpio_int_polarity),
    .i1(pwdata_int),
    .sel(n58),
    .o(n59));  // ../RTL/gpio_apbif.v(363)
  binary_mux_s1_w32 mux31 (
    .i0(int_gpio_ls_sync),
    .i1(pwdata_int),
    .sel(n61),
    .o(n62));  // ../RTL/gpio_apbif.v(383)
  binary_mux_s1_w32 mux32 (
    .i0(32'b00000000000000000000000000000000),
    .i1(pwdata_int),
    .sel(n63),
    .o({open_n0,open_n1,open_n2,open_n3,open_n4,open_n5,open_n6,open_n7,open_n8,open_n9,open_n10,open_n11,open_n12,open_n13,open_n14,open_n15,open_n16,open_n17,open_n18,open_n19,open_n20,open_n21,open_n22,open_n23,int_gpio_porta_eoi[7:0]}));  // ../RTL/gpio_apbif.v(404)
  binary_mux_s1_w32 mux33 (
    .i0(iprdata),
    .i1(n81),
    .sel(n68),
    .o(n82));  // ../RTL/gpio_apbif.v(453)
  binary_mux_s1_w4 mux4 (
    .i0({n11,n11,n11,n11}),
    .i1(4'b0000),
    .sel(n10),
    .o(n14));  // ../RTL/gpio_apbif.v(230)
  binary_mux_s1_w4 mux5 (
    .i0(n13),
    .i1(4'b0000),
    .sel(n10),
    .o(n15));  // ../RTL/gpio_apbif.v(230)
  binary_mux_s1_w4 mux6 (
    .i0({n10,n10,n10,n10}),
    .i1(4'b0000),
    .sel(n9),
    .o(n19));  // ../RTL/gpio_apbif.v(230)
  binary_mux_s1_w4 mux7 (
    .i0(n14),
    .i1(4'b0000),
    .sel(n9),
    .o(n20));  // ../RTL/gpio_apbif.v(230)
  binary_mux_s1_w4 mux8 (
    .i0(n15),
    .i1(4'b0000),
    .sel(n9),
    .o(n21));  // ../RTL/gpio_apbif.v(230)
  binary_mux_s1_w4 mux9 (
    .i0({n9,n9,n9,n9}),
    .i1(4'b0000),
    .sel(n8),
    .o(n26));  // ../RTL/gpio_apbif.v(230)
  reg_ar_as_w32 reg0 (
    .clk(pclk),
    .d(n44),
    .reset({n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39}),
    .set(32'b00000000000000000000000000000000),
    .q(int_gpio_swporta_ddr));  // ../RTL/gpio_apbif.v(262)
  reg_ar_as_w32 reg1 (
    .clk(pclk),
    .d(n47),
    .reset({n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39}),
    .set(32'b00000000000000000000000000000000),
    .q(int_gpio_swporta_ctl));  // ../RTL/gpio_apbif.v(282)
  reg_ar_as_w32 reg2 (
    .clk(pclk),
    .d(n50),
    .reset({n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39}),
    .set(32'b00000000000000000000000000000000),
    .q(int_gpio_inten));  // ../RTL/gpio_apbif.v(303)
  reg_ar_as_w32 reg3 (
    .clk(pclk),
    .d(n53),
    .reset({n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39}),
    .set(32'b00000000000000000000000000000000),
    .q(int_gpio_intmask));  // ../RTL/gpio_apbif.v(323)
  reg_ar_as_w32 reg4 (
    .clk(pclk),
    .d(n56),
    .reset({n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39}),
    .set(32'b00000000000000000000000000000000),
    .q(int_gpio_inttype_level));  // ../RTL/gpio_apbif.v(343)
  reg_ar_as_w32 reg5 (
    .clk(pclk),
    .d(n59),
    .reset({n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39}),
    .set(32'b00000000000000000000000000000000),
    .q(int_gpio_int_polarity));  // ../RTL/gpio_apbif.v(363)
  reg_ar_as_w32 reg6 (
    .clk(pclk),
    .d(n62),
    .reset({n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39}),
    .set(32'b00000000000000000000000000000000),
    .q(int_gpio_ls_sync));  // ../RTL/gpio_apbif.v(383)
  reg_ar_as_w32 reg7 (
    .clk(pclk),
    .d(n82),
    .reset({n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39}),
    .set(32'b00000000000000000000000000000000),
    .q(iprdata));  // ../RTL/gpio_apbif.v(453)
  reg_ar_as_w32 reg8 (
    .clk(pclk),
    .d(n41),
    .reset({n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39,n39}),
    .set(32'b00000000000000000000000000000000),
    .q(int_gpio_swporta_dr));  // ../RTL/gpio_apbif.v(242)
  onehot_mux_s12_w32 sel0 (
    .i0(32'b00000000000000000000000000000000),
    .i1(ri_gpio_ext_porta_rb),
    .i10(ri_gpio_swporta_ddr),
    .i11(ri_gpio_swporta_dr),
    .i2(ri_gpio_ls_sync),
    .i3(ri_gpio_raw_intstatus),
    .i4(ri_gpio_intstatus),
    .i5(ri_gpio_int_polarity),
    .i6(ri_gpio_inttype_level),
    .i7(ri_gpio_intmask),
    .i8(ri_gpio_inten),
    .i9(ri_gpio_swporta_ctl),
    .sel({n2,n3,n71,n7,n8,n9,n10,n76,n77,n11,n79,n80}),
    .o(n81));  // ../RTL/gpio_apbif.v(453)
  buf u10 (prdata[24], 1'b0);  // ../RTL/gpio_apbif.v(462)
  buf u100 (ri_gpio_ext_porta_rb[18], 1'b0);  // ../RTL/gpio_apbif.v(430)
  buf u101 (ri_gpio_ext_porta_rb[19], 1'b0);  // ../RTL/gpio_apbif.v(430)
  buf u102 (ri_gpio_ext_porta_rb[20], 1'b0);  // ../RTL/gpio_apbif.v(430)
  buf u103 (ri_gpio_ext_porta_rb[21], 1'b0);  // ../RTL/gpio_apbif.v(430)
  buf u104 (ri_gpio_ext_porta_rb[22], 1'b0);  // ../RTL/gpio_apbif.v(430)
  buf u105 (ri_gpio_ext_porta_rb[23], 1'b0);  // ../RTL/gpio_apbif.v(430)
  buf u106 (ri_gpio_ext_porta_rb[24], 1'b0);  // ../RTL/gpio_apbif.v(430)
  buf u107 (ri_gpio_ext_porta_rb[25], 1'b0);  // ../RTL/gpio_apbif.v(430)
  buf u108 (ri_gpio_ext_porta_rb[26], 1'b0);  // ../RTL/gpio_apbif.v(430)
  buf u109 (ri_gpio_ext_porta_rb[27], 1'b0);  // ../RTL/gpio_apbif.v(430)
  buf u11 (prdata[23], 1'b0);  // ../RTL/gpio_apbif.v(462)
  buf u110 (ri_gpio_ext_porta_rb[28], 1'b0);  // ../RTL/gpio_apbif.v(430)
  buf u111 (ri_gpio_ext_porta_rb[29], 1'b0);  // ../RTL/gpio_apbif.v(430)
  buf u112 (ri_gpio_ext_porta_rb[30], 1'b0);  // ../RTL/gpio_apbif.v(430)
  buf u113 (ri_gpio_ext_porta_rb[31], 1'b0);  // ../RTL/gpio_apbif.v(430)
  buf u114 (ri_gpio_intstatus[1], gpio_intstatus[1]);  // ../RTL/gpio_apbif.v(421)
  buf u115 (ri_gpio_intstatus[2], gpio_intstatus[2]);  // ../RTL/gpio_apbif.v(421)
  buf u116 (ri_gpio_intstatus[3], gpio_intstatus[3]);  // ../RTL/gpio_apbif.v(421)
  buf u117 (ri_gpio_intstatus[4], gpio_intstatus[4]);  // ../RTL/gpio_apbif.v(421)
  buf u118 (ri_gpio_intstatus[5], gpio_intstatus[5]);  // ../RTL/gpio_apbif.v(421)
  buf u119 (ri_gpio_intstatus[6], gpio_intstatus[6]);  // ../RTL/gpio_apbif.v(421)
  buf u12 (pwdata_int[0], pwdata[0]);  // ../RTL/gpio_apbif.v(147)
  buf u120 (ri_gpio_intstatus[7], gpio_intstatus[7]);  // ../RTL/gpio_apbif.v(421)
  buf u121 (ri_gpio_intstatus[8], 1'b0);  // ../RTL/gpio_apbif.v(421)
  buf u122 (ri_gpio_intstatus[9], 1'b0);  // ../RTL/gpio_apbif.v(421)
  buf u123 (ri_gpio_intstatus[10], 1'b0);  // ../RTL/gpio_apbif.v(421)
  buf u124 (ri_gpio_intstatus[11], 1'b0);  // ../RTL/gpio_apbif.v(421)
  buf u125 (ri_gpio_intstatus[12], 1'b0);  // ../RTL/gpio_apbif.v(421)
  buf u126 (ri_gpio_intstatus[13], 1'b0);  // ../RTL/gpio_apbif.v(421)
  buf u127 (ri_gpio_intstatus[14], 1'b0);  // ../RTL/gpio_apbif.v(421)
  buf u128 (ri_gpio_intstatus[15], 1'b0);  // ../RTL/gpio_apbif.v(421)
  buf u129 (ri_gpio_intstatus[16], 1'b0);  // ../RTL/gpio_apbif.v(421)
  or u13 (n69, n3, n2);  // ../RTL/gpio_apbif.v(453)
  buf u130 (ri_gpio_intstatus[17], 1'b0);  // ../RTL/gpio_apbif.v(421)
  buf u131 (ri_gpio_intstatus[18], 1'b0);  // ../RTL/gpio_apbif.v(421)
  buf u132 (ri_gpio_intstatus[19], 1'b0);  // ../RTL/gpio_apbif.v(421)
  buf u133 (ri_gpio_intstatus[20], 1'b0);  // ../RTL/gpio_apbif.v(421)
  buf u134 (ri_gpio_intstatus[21], 1'b0);  // ../RTL/gpio_apbif.v(421)
  buf u135 (ri_gpio_intstatus[22], 1'b0);  // ../RTL/gpio_apbif.v(421)
  buf u136 (ri_gpio_intstatus[23], 1'b0);  // ../RTL/gpio_apbif.v(421)
  buf u137 (ri_gpio_intstatus[24], 1'b0);  // ../RTL/gpio_apbif.v(421)
  buf u138 (ri_gpio_intstatus[25], 1'b0);  // ../RTL/gpio_apbif.v(421)
  buf u139 (ri_gpio_intstatus[26], 1'b0);  // ../RTL/gpio_apbif.v(421)
  or u14 (n70, n9, n72);  // ../RTL/gpio_apbif.v(453)
  buf u140 (ri_gpio_intstatus[27], 1'b0);  // ../RTL/gpio_apbif.v(421)
  buf u141 (ri_gpio_intstatus[28], 1'b0);  // ../RTL/gpio_apbif.v(421)
  buf u142 (ri_gpio_intstatus[29], 1'b0);  // ../RTL/gpio_apbif.v(421)
  buf u143 (ri_gpio_intstatus[30], 1'b0);  // ../RTL/gpio_apbif.v(421)
  buf u144 (ri_gpio_intstatus[31], 1'b0);  // ../RTL/gpio_apbif.v(421)
  buf u145 (ri_gpio_raw_intstatus[1], gpio_raw_intstatus[1]);  // ../RTL/gpio_apbif.v(421)
  buf u146 (ri_gpio_raw_intstatus[2], gpio_raw_intstatus[2]);  // ../RTL/gpio_apbif.v(421)
  buf u147 (ri_gpio_raw_intstatus[3], gpio_raw_intstatus[3]);  // ../RTL/gpio_apbif.v(421)
  buf u148 (ri_gpio_raw_intstatus[4], gpio_raw_intstatus[4]);  // ../RTL/gpio_apbif.v(421)
  buf u149 (ri_gpio_raw_intstatus[5], gpio_raw_intstatus[5]);  // ../RTL/gpio_apbif.v(421)
  buf u15 (prdata[16], 1'b0);  // ../RTL/gpio_apbif.v(462)
  buf u150 (ri_gpio_raw_intstatus[6], gpio_raw_intstatus[6]);  // ../RTL/gpio_apbif.v(421)
  buf u151 (ri_gpio_raw_intstatus[7], gpio_raw_intstatus[7]);  // ../RTL/gpio_apbif.v(421)
  buf u152 (ri_gpio_raw_intstatus[8], 1'b0);  // ../RTL/gpio_apbif.v(421)
  buf u153 (ri_gpio_raw_intstatus[9], 1'b0);  // ../RTL/gpio_apbif.v(421)
  buf u154 (ri_gpio_raw_intstatus[10], 1'b0);  // ../RTL/gpio_apbif.v(421)
  buf u155 (ri_gpio_raw_intstatus[11], 1'b0);  // ../RTL/gpio_apbif.v(421)
  buf u156 (ri_gpio_raw_intstatus[12], 1'b0);  // ../RTL/gpio_apbif.v(421)
  buf u157 (ri_gpio_raw_intstatus[13], 1'b0);  // ../RTL/gpio_apbif.v(421)
  buf u158 (ri_gpio_raw_intstatus[14], 1'b0);  // ../RTL/gpio_apbif.v(421)
  buf u159 (ri_gpio_raw_intstatus[15], 1'b0);  // ../RTL/gpio_apbif.v(421)
  or u16 (n72, n8, n7);  // ../RTL/gpio_apbif.v(453)
  buf u160 (ri_gpio_raw_intstatus[16], 1'b0);  // ../RTL/gpio_apbif.v(421)
  buf u161 (ri_gpio_raw_intstatus[17], 1'b0);  // ../RTL/gpio_apbif.v(421)
  buf u162 (ri_gpio_raw_intstatus[18], 1'b0);  // ../RTL/gpio_apbif.v(421)
  buf u163 (ri_gpio_raw_intstatus[19], 1'b0);  // ../RTL/gpio_apbif.v(421)
  buf u164 (ri_gpio_raw_intstatus[20], 1'b0);  // ../RTL/gpio_apbif.v(421)
  buf u165 (ri_gpio_raw_intstatus[21], 1'b0);  // ../RTL/gpio_apbif.v(421)
  buf u166 (ri_gpio_raw_intstatus[22], 1'b0);  // ../RTL/gpio_apbif.v(421)
  buf u167 (ri_gpio_raw_intstatus[23], 1'b0);  // ../RTL/gpio_apbif.v(421)
  buf u168 (ri_gpio_raw_intstatus[24], 1'b0);  // ../RTL/gpio_apbif.v(421)
  buf u169 (ri_gpio_raw_intstatus[25], 1'b0);  // ../RTL/gpio_apbif.v(421)
  buf u17 (prdata[15], 1'b0);  // ../RTL/gpio_apbif.v(462)
  buf u170 (ri_gpio_raw_intstatus[26], 1'b0);  // ../RTL/gpio_apbif.v(421)
  buf u171 (ri_gpio_raw_intstatus[27], 1'b0);  // ../RTL/gpio_apbif.v(421)
  buf u172 (ri_gpio_raw_intstatus[28], 1'b0);  // ../RTL/gpio_apbif.v(421)
  buf u173 (ri_gpio_raw_intstatus[29], 1'b0);  // ../RTL/gpio_apbif.v(421)
  buf u174 (ri_gpio_raw_intstatus[30], 1'b0);  // ../RTL/gpio_apbif.v(421)
  buf u175 (ri_gpio_raw_intstatus[31], 1'b0);  // ../RTL/gpio_apbif.v(421)
  buf u176 (gpio_porta_eoi[1], int_gpio_porta_eoi[1]);  // ../RTL/gpio_apbif.v(408)
  buf u177 (gpio_porta_eoi[2], int_gpio_porta_eoi[2]);  // ../RTL/gpio_apbif.v(408)
  buf u178 (gpio_porta_eoi[3], int_gpio_porta_eoi[3]);  // ../RTL/gpio_apbif.v(408)
  buf u179 (gpio_porta_eoi[4], int_gpio_porta_eoi[4]);  // ../RTL/gpio_apbif.v(408)
  buf u18 (prdata[22], 1'b0);  // ../RTL/gpio_apbif.v(462)
  buf u180 (gpio_porta_eoi[5], int_gpio_porta_eoi[5]);  // ../RTL/gpio_apbif.v(408)
  buf u181 (gpio_porta_eoi[6], int_gpio_porta_eoi[6]);  // ../RTL/gpio_apbif.v(408)
  buf u182 (gpio_porta_eoi[7], int_gpio_porta_eoi[7]);  // ../RTL/gpio_apbif.v(408)
  and u183 (n51, gpio_porta_eoi_wen[2], gpio_porta_eoi_wen[3]);  // ../RTL/gpio_apbif.v(403)
  and u184 (n63, n54, n51);  // ../RTL/gpio_apbif.v(403)
  buf u185 (ri_gpio_ls_sync[1], int_gpio_ls_sync[1]);  // ../RTL/gpio_apbif.v(394)
  buf u186 (ri_gpio_ls_sync[2], int_gpio_ls_sync[2]);  // ../RTL/gpio_apbif.v(394)
  buf u187 (ri_gpio_ls_sync[3], int_gpio_ls_sync[3]);  // ../RTL/gpio_apbif.v(394)
  buf u188 (ri_gpio_ls_sync[4], int_gpio_ls_sync[4]);  // ../RTL/gpio_apbif.v(394)
  buf u189 (ri_gpio_ls_sync[5], int_gpio_ls_sync[5]);  // ../RTL/gpio_apbif.v(394)
  buf u19 (prdata[21], 1'b0);  // ../RTL/gpio_apbif.v(462)
  buf u190 (ri_gpio_ls_sync[6], int_gpio_ls_sync[6]);  // ../RTL/gpio_apbif.v(394)
  buf u191 (ri_gpio_ls_sync[7], int_gpio_ls_sync[7]);  // ../RTL/gpio_apbif.v(394)
  buf u192 (ri_gpio_ls_sync[8], 1'b0);  // ../RTL/gpio_apbif.v(394)
  buf u193 (ri_gpio_ls_sync[9], 1'b0);  // ../RTL/gpio_apbif.v(394)
  buf u194 (ri_gpio_ls_sync[10], 1'b0);  // ../RTL/gpio_apbif.v(394)
  buf u195 (ri_gpio_ls_sync[11], 1'b0);  // ../RTL/gpio_apbif.v(394)
  buf u196 (ri_gpio_ls_sync[12], 1'b0);  // ../RTL/gpio_apbif.v(394)
  buf u197 (ri_gpio_ls_sync[13], 1'b0);  // ../RTL/gpio_apbif.v(394)
  buf u198 (ri_gpio_ls_sync[14], 1'b0);  // ../RTL/gpio_apbif.v(394)
  buf u199 (ri_gpio_ls_sync[15], 1'b0);  // ../RTL/gpio_apbif.v(394)
  buf u2 (ri_gpio_ext_porta_rb[2], gpio_ext_porta_rb[2]);  // ../RTL/gpio_apbif.v(430)
  buf u20 (prdata[20], 1'b0);  // ../RTL/gpio_apbif.v(462)
  buf u200 (ri_gpio_ls_sync[16], 1'b0);  // ../RTL/gpio_apbif.v(394)
  buf u201 (ri_gpio_ls_sync[17], 1'b0);  // ../RTL/gpio_apbif.v(394)
  buf u202 (ri_gpio_ls_sync[18], 1'b0);  // ../RTL/gpio_apbif.v(394)
  buf u203 (ri_gpio_ls_sync[19], 1'b0);  // ../RTL/gpio_apbif.v(394)
  buf u204 (ri_gpio_ls_sync[20], 1'b0);  // ../RTL/gpio_apbif.v(394)
  buf u205 (ri_gpio_ls_sync[21], 1'b0);  // ../RTL/gpio_apbif.v(394)
  buf u206 (ri_gpio_ls_sync[22], 1'b0);  // ../RTL/gpio_apbif.v(394)
  buf u207 (ri_gpio_ls_sync[23], 1'b0);  // ../RTL/gpio_apbif.v(394)
  buf u208 (ri_gpio_ls_sync[24], 1'b0);  // ../RTL/gpio_apbif.v(394)
  buf u209 (ri_gpio_ls_sync[25], 1'b0);  // ../RTL/gpio_apbif.v(394)
  buf u21 (prdata[19], 1'b0);  // ../RTL/gpio_apbif.v(462)
  buf u210 (ri_gpio_ls_sync[26], 1'b0);  // ../RTL/gpio_apbif.v(394)
  buf u211 (ri_gpio_ls_sync[27], 1'b0);  // ../RTL/gpio_apbif.v(394)
  buf u212 (ri_gpio_ls_sync[28], 1'b0);  // ../RTL/gpio_apbif.v(394)
  buf u213 (ri_gpio_ls_sync[29], 1'b0);  // ../RTL/gpio_apbif.v(394)
  buf u214 (ri_gpio_ls_sync[30], 1'b0);  // ../RTL/gpio_apbif.v(394)
  buf u215 (ri_gpio_ls_sync[31], 1'b0);  // ../RTL/gpio_apbif.v(394)
  and u216 (n45, gpio_ls_sync_wen[2], gpio_ls_sync_wen[3]);  // ../RTL/gpio_apbif.v(382)
  and u217 (n61, n48, n45);  // ../RTL/gpio_apbif.v(382)
  buf u218 (ri_gpio_int_polarity[1], int_gpio_int_polarity[1]);  // ../RTL/gpio_apbif.v(374)
  buf u219 (ri_gpio_int_polarity[2], int_gpio_int_polarity[2]);  // ../RTL/gpio_apbif.v(374)
  buf u22 (prdata[18], 1'b0);  // ../RTL/gpio_apbif.v(462)
  buf u220 (ri_gpio_int_polarity[3], int_gpio_int_polarity[3]);  // ../RTL/gpio_apbif.v(374)
  buf u221 (ri_gpio_int_polarity[4], int_gpio_int_polarity[4]);  // ../RTL/gpio_apbif.v(374)
  buf u222 (ri_gpio_int_polarity[5], int_gpio_int_polarity[5]);  // ../RTL/gpio_apbif.v(374)
  buf u223 (ri_gpio_int_polarity[6], int_gpio_int_polarity[6]);  // ../RTL/gpio_apbif.v(374)
  buf u224 (ri_gpio_int_polarity[7], int_gpio_int_polarity[7]);  // ../RTL/gpio_apbif.v(374)
  buf u225 (ri_gpio_int_polarity[8], 1'b0);  // ../RTL/gpio_apbif.v(374)
  buf u226 (ri_gpio_int_polarity[9], 1'b0);  // ../RTL/gpio_apbif.v(374)
  buf u227 (ri_gpio_int_polarity[10], 1'b0);  // ../RTL/gpio_apbif.v(374)
  buf u228 (ri_gpio_int_polarity[11], 1'b0);  // ../RTL/gpio_apbif.v(374)
  buf u229 (ri_gpio_int_polarity[12], 1'b0);  // ../RTL/gpio_apbif.v(374)
  buf u23 (prdata[17], 1'b0);  // ../RTL/gpio_apbif.v(462)
  buf u230 (ri_gpio_int_polarity[13], 1'b0);  // ../RTL/gpio_apbif.v(374)
  buf u231 (ri_gpio_int_polarity[14], 1'b0);  // ../RTL/gpio_apbif.v(374)
  buf u232 (ri_gpio_int_polarity[15], 1'b0);  // ../RTL/gpio_apbif.v(374)
  buf u233 (ri_gpio_int_polarity[16], 1'b0);  // ../RTL/gpio_apbif.v(374)
  buf u234 (ri_gpio_int_polarity[17], 1'b0);  // ../RTL/gpio_apbif.v(374)
  buf u235 (ri_gpio_int_polarity[18], 1'b0);  // ../RTL/gpio_apbif.v(374)
  buf u236 (ri_gpio_int_polarity[19], 1'b0);  // ../RTL/gpio_apbif.v(374)
  buf u237 (ri_gpio_int_polarity[20], 1'b0);  // ../RTL/gpio_apbif.v(374)
  buf u238 (ri_gpio_int_polarity[21], 1'b0);  // ../RTL/gpio_apbif.v(374)
  buf u239 (ri_gpio_int_polarity[22], 1'b0);  // ../RTL/gpio_apbif.v(374)
  or u24 (n73, n78, n74);  // ../RTL/gpio_apbif.v(453)
  buf u240 (ri_gpio_int_polarity[23], 1'b0);  // ../RTL/gpio_apbif.v(374)
  buf u241 (ri_gpio_int_polarity[24], 1'b0);  // ../RTL/gpio_apbif.v(374)
  buf u242 (ri_gpio_int_polarity[25], 1'b0);  // ../RTL/gpio_apbif.v(374)
  buf u243 (ri_gpio_int_polarity[26], 1'b0);  // ../RTL/gpio_apbif.v(374)
  buf u244 (ri_gpio_int_polarity[27], 1'b0);  // ../RTL/gpio_apbif.v(374)
  buf u245 (ri_gpio_int_polarity[28], 1'b0);  // ../RTL/gpio_apbif.v(374)
  buf u246 (ri_gpio_int_polarity[29], 1'b0);  // ../RTL/gpio_apbif.v(374)
  buf u247 (ri_gpio_int_polarity[30], 1'b0);  // ../RTL/gpio_apbif.v(374)
  buf u248 (ri_gpio_int_polarity[31], 1'b0);  // ../RTL/gpio_apbif.v(374)
  buf u249 (gpio_int_polarity[1], int_gpio_int_polarity[1]);  // ../RTL/gpio_apbif.v(366)
  not u25 (n39, presetn);  // ../RTL/gpio_apbif.v(238)
  buf u250 (gpio_int_polarity[2], int_gpio_int_polarity[2]);  // ../RTL/gpio_apbif.v(366)
  buf u251 (gpio_int_polarity[3], int_gpio_int_polarity[3]);  // ../RTL/gpio_apbif.v(366)
  buf u252 (gpio_int_polarity[4], int_gpio_int_polarity[4]);  // ../RTL/gpio_apbif.v(366)
  buf u253 (gpio_int_polarity[5], int_gpio_int_polarity[5]);  // ../RTL/gpio_apbif.v(366)
  buf u254 (gpio_int_polarity[6], int_gpio_int_polarity[6]);  // ../RTL/gpio_apbif.v(366)
  buf u255 (gpio_int_polarity[7], int_gpio_int_polarity[7]);  // ../RTL/gpio_apbif.v(366)
  and u256 (n1, gpio_int_polarity_wen[2], gpio_int_polarity_wen[3]);  // ../RTL/gpio_apbif.v(362)
  and u257 (n58, n42, n1);  // ../RTL/gpio_apbif.v(362)
  buf u258 (ri_gpio_inttype_level[1], int_gpio_inttype_level[1]);  // ../RTL/gpio_apbif.v(354)
  buf u259 (ri_gpio_inttype_level[2], int_gpio_inttype_level[2]);  // ../RTL/gpio_apbif.v(354)
  buf u26 (gpio_swporta_ctl_wen[0], 1'b0);  // ../RTL/gpio_apbif.v(180)
  buf u260 (ri_gpio_inttype_level[3], int_gpio_inttype_level[3]);  // ../RTL/gpio_apbif.v(354)
  buf u261 (ri_gpio_inttype_level[4], int_gpio_inttype_level[4]);  // ../RTL/gpio_apbif.v(354)
  buf u262 (ri_gpio_inttype_level[5], int_gpio_inttype_level[5]);  // ../RTL/gpio_apbif.v(354)
  buf u263 (ri_gpio_inttype_level[6], int_gpio_inttype_level[6]);  // ../RTL/gpio_apbif.v(354)
  buf u264 (ri_gpio_inttype_level[7], int_gpio_inttype_level[7]);  // ../RTL/gpio_apbif.v(354)
  buf u265 (ri_gpio_inttype_level[8], 1'b0);  // ../RTL/gpio_apbif.v(354)
  buf u266 (ri_gpio_inttype_level[9], 1'b0);  // ../RTL/gpio_apbif.v(354)
  buf u267 (ri_gpio_inttype_level[10], 1'b0);  // ../RTL/gpio_apbif.v(354)
  buf u268 (ri_gpio_inttype_level[11], 1'b0);  // ../RTL/gpio_apbif.v(354)
  buf u269 (ri_gpio_inttype_level[12], 1'b0);  // ../RTL/gpio_apbif.v(354)
  and u27 (n17, gpio_swporta_dr_wen[0], gpio_swporta_dr_wen[1]);  // ../RTL/gpio_apbif.v(241)
  buf u270 (ri_gpio_inttype_level[13], 1'b0);  // ../RTL/gpio_apbif.v(354)
  buf u271 (ri_gpio_inttype_level[14], 1'b0);  // ../RTL/gpio_apbif.v(354)
  buf u272 (ri_gpio_inttype_level[15], 1'b0);  // ../RTL/gpio_apbif.v(354)
  buf u273 (ri_gpio_inttype_level[16], 1'b0);  // ../RTL/gpio_apbif.v(354)
  buf u274 (ri_gpio_inttype_level[17], 1'b0);  // ../RTL/gpio_apbif.v(354)
  buf u275 (ri_gpio_inttype_level[18], 1'b0);  // ../RTL/gpio_apbif.v(354)
  buf u276 (ri_gpio_inttype_level[19], 1'b0);  // ../RTL/gpio_apbif.v(354)
  buf u277 (ri_gpio_inttype_level[20], 1'b0);  // ../RTL/gpio_apbif.v(354)
  buf u278 (ri_gpio_inttype_level[21], 1'b0);  // ../RTL/gpio_apbif.v(354)
  buf u279 (ri_gpio_inttype_level[22], 1'b0);  // ../RTL/gpio_apbif.v(354)
  buf u28 (gpio_swporta_dr[0], int_gpio_swporta_dr[0]);  // ../RTL/gpio_apbif.v(245)
  buf u280 (ri_gpio_inttype_level[23], 1'b0);  // ../RTL/gpio_apbif.v(354)
  buf u281 (ri_gpio_inttype_level[24], 1'b0);  // ../RTL/gpio_apbif.v(354)
  buf u282 (ri_gpio_inttype_level[25], 1'b0);  // ../RTL/gpio_apbif.v(354)
  buf u283 (ri_gpio_inttype_level[26], 1'b0);  // ../RTL/gpio_apbif.v(354)
  buf u284 (ri_gpio_inttype_level[27], 1'b0);  // ../RTL/gpio_apbif.v(354)
  buf u285 (ri_gpio_inttype_level[28], 1'b0);  // ../RTL/gpio_apbif.v(354)
  buf u286 (ri_gpio_inttype_level[29], 1'b0);  // ../RTL/gpio_apbif.v(354)
  buf u287 (ri_gpio_inttype_level[30], 1'b0);  // ../RTL/gpio_apbif.v(354)
  buf u288 (ri_gpio_inttype_level[31], 1'b0);  // ../RTL/gpio_apbif.v(354)
  buf u289 (gpio_inttype_level[1], int_gpio_inttype_level[1]);  // ../RTL/gpio_apbif.v(346)
  or u29 (n74, n77, n75);  // ../RTL/gpio_apbif.v(453)
  buf u290 (gpio_inttype_level[2], int_gpio_inttype_level[2]);  // ../RTL/gpio_apbif.v(346)
  buf u291 (gpio_inttype_level[3], int_gpio_inttype_level[3]);  // ../RTL/gpio_apbif.v(346)
  buf u292 (gpio_inttype_level[4], int_gpio_inttype_level[4]);  // ../RTL/gpio_apbif.v(346)
  buf u293 (gpio_inttype_level[5], int_gpio_inttype_level[5]);  // ../RTL/gpio_apbif.v(346)
  buf u294 (gpio_inttype_level[6], int_gpio_inttype_level[6]);  // ../RTL/gpio_apbif.v(346)
  buf u295 (gpio_inttype_level[7], int_gpio_inttype_level[7]);  // ../RTL/gpio_apbif.v(346)
  and u296 (n33, gpio_inttype_level_wen[2], gpio_inttype_level_wen[3]);  // ../RTL/gpio_apbif.v(342)
  and u297 (n55, n5, n33);  // ../RTL/gpio_apbif.v(342)
  buf u298 (ri_gpio_intmask[1], int_gpio_intmask[1]);  // ../RTL/gpio_apbif.v(334)
  buf u299 (ri_gpio_intmask[2], int_gpio_intmask[2]);  // ../RTL/gpio_apbif.v(334)
  buf u3 (ri_gpio_ext_porta_rb[1], gpio_ext_porta_rb[1]);  // ../RTL/gpio_apbif.v(430)
  buf u30 (prdata[14], 1'b0);  // ../RTL/gpio_apbif.v(462)
  buf u300 (ri_gpio_intmask[3], int_gpio_intmask[3]);  // ../RTL/gpio_apbif.v(334)
  buf u301 (ri_gpio_intmask[4], int_gpio_intmask[4]);  // ../RTL/gpio_apbif.v(334)
  buf u302 (ri_gpio_intmask[5], int_gpio_intmask[5]);  // ../RTL/gpio_apbif.v(334)
  buf u303 (ri_gpio_intmask[6], int_gpio_intmask[6]);  // ../RTL/gpio_apbif.v(334)
  buf u304 (ri_gpio_intmask[7], int_gpio_intmask[7]);  // ../RTL/gpio_apbif.v(334)
  buf u305 (ri_gpio_intmask[8], 1'b0);  // ../RTL/gpio_apbif.v(334)
  buf u306 (ri_gpio_intmask[9], 1'b0);  // ../RTL/gpio_apbif.v(334)
  buf u307 (ri_gpio_intmask[10], 1'b0);  // ../RTL/gpio_apbif.v(334)
  buf u308 (ri_gpio_intmask[11], 1'b0);  // ../RTL/gpio_apbif.v(334)
  buf u309 (ri_gpio_intmask[12], 1'b0);  // ../RTL/gpio_apbif.v(334)
  buf u31 (ri_gpio_swporta_dr[0], int_gpio_swporta_dr[0]);  // ../RTL/gpio_apbif.v(253)
  buf u310 (ri_gpio_intmask[13], 1'b0);  // ../RTL/gpio_apbif.v(334)
  buf u311 (ri_gpio_intmask[14], 1'b0);  // ../RTL/gpio_apbif.v(334)
  buf u312 (ri_gpio_intmask[15], 1'b0);  // ../RTL/gpio_apbif.v(334)
  buf u313 (ri_gpio_intmask[16], 1'b0);  // ../RTL/gpio_apbif.v(334)
  buf u314 (ri_gpio_intmask[17], 1'b0);  // ../RTL/gpio_apbif.v(334)
  buf u315 (ri_gpio_intmask[18], 1'b0);  // ../RTL/gpio_apbif.v(334)
  buf u316 (ri_gpio_intmask[19], 1'b0);  // ../RTL/gpio_apbif.v(334)
  buf u317 (ri_gpio_intmask[20], 1'b0);  // ../RTL/gpio_apbif.v(334)
  buf u318 (ri_gpio_intmask[21], 1'b0);  // ../RTL/gpio_apbif.v(334)
  buf u319 (ri_gpio_intmask[22], 1'b0);  // ../RTL/gpio_apbif.v(334)
  and u32 (n22, gpio_swporta_ddr_wen[0], gpio_swporta_ddr_wen[1]);  // ../RTL/gpio_apbif.v(261)
  buf u320 (ri_gpio_intmask[23], 1'b0);  // ../RTL/gpio_apbif.v(334)
  buf u321 (ri_gpio_intmask[24], 1'b0);  // ../RTL/gpio_apbif.v(334)
  buf u322 (ri_gpio_intmask[25], 1'b0);  // ../RTL/gpio_apbif.v(334)
  buf u323 (ri_gpio_intmask[26], 1'b0);  // ../RTL/gpio_apbif.v(334)
  buf u324 (ri_gpio_intmask[27], 1'b0);  // ../RTL/gpio_apbif.v(334)
  buf u325 (ri_gpio_intmask[28], 1'b0);  // ../RTL/gpio_apbif.v(334)
  buf u326 (ri_gpio_intmask[29], 1'b0);  // ../RTL/gpio_apbif.v(334)
  buf u327 (ri_gpio_intmask[30], 1'b0);  // ../RTL/gpio_apbif.v(334)
  buf u328 (ri_gpio_intmask[31], 1'b0);  // ../RTL/gpio_apbif.v(334)
  buf u329 (gpio_intmask[1], int_gpio_intmask[1]);  // ../RTL/gpio_apbif.v(326)
  buf u33 (gpio_swporta_ddr[0], int_gpio_swporta_ddr[0]);  // ../RTL/gpio_apbif.v(265)
  buf u330 (gpio_intmask[2], int_gpio_intmask[2]);  // ../RTL/gpio_apbif.v(326)
  buf u331 (gpio_intmask[3], int_gpio_intmask[3]);  // ../RTL/gpio_apbif.v(326)
  buf u332 (gpio_intmask[4], int_gpio_intmask[4]);  // ../RTL/gpio_apbif.v(326)
  buf u333 (gpio_intmask[5], int_gpio_intmask[5]);  // ../RTL/gpio_apbif.v(326)
  buf u334 (gpio_intmask[6], int_gpio_intmask[6]);  // ../RTL/gpio_apbif.v(326)
  buf u335 (gpio_intmask[7], int_gpio_intmask[7]);  // ../RTL/gpio_apbif.v(326)
  and u336 (n31, gpio_intmask_wen[2], gpio_intmask_wen[3]);  // ../RTL/gpio_apbif.v(322)
  and u337 (n52, n32, n31);  // ../RTL/gpio_apbif.v(322)
  buf u338 (ri_gpio_inten[1], int_gpio_inten[1]);  // ../RTL/gpio_apbif.v(314)
  buf u339 (ri_gpio_inten[2], int_gpio_inten[2]);  // ../RTL/gpio_apbif.v(314)
  or u34 (n75, n76, n10);  // ../RTL/gpio_apbif.v(453)
  buf u340 (ri_gpio_inten[3], int_gpio_inten[3]);  // ../RTL/gpio_apbif.v(314)
  buf u341 (ri_gpio_inten[4], int_gpio_inten[4]);  // ../RTL/gpio_apbif.v(314)
  buf u342 (ri_gpio_inten[5], int_gpio_inten[5]);  // ../RTL/gpio_apbif.v(314)
  buf u343 (ri_gpio_inten[6], int_gpio_inten[6]);  // ../RTL/gpio_apbif.v(314)
  buf u344 (ri_gpio_inten[7], int_gpio_inten[7]);  // ../RTL/gpio_apbif.v(314)
  buf u345 (ri_gpio_inten[8], 1'b0);  // ../RTL/gpio_apbif.v(314)
  buf u346 (ri_gpio_inten[9], 1'b0);  // ../RTL/gpio_apbif.v(314)
  buf u347 (ri_gpio_inten[10], 1'b0);  // ../RTL/gpio_apbif.v(314)
  buf u348 (ri_gpio_inten[11], 1'b0);  // ../RTL/gpio_apbif.v(314)
  buf u349 (ri_gpio_inten[12], 1'b0);  // ../RTL/gpio_apbif.v(314)
  buf u35 (prdata[13], 1'b0);  // ../RTL/gpio_apbif.v(462)
  buf u350 (ri_gpio_inten[13], 1'b0);  // ../RTL/gpio_apbif.v(314)
  buf u351 (ri_gpio_inten[14], 1'b0);  // ../RTL/gpio_apbif.v(314)
  buf u352 (ri_gpio_inten[15], 1'b0);  // ../RTL/gpio_apbif.v(314)
  buf u353 (ri_gpio_inten[16], 1'b0);  // ../RTL/gpio_apbif.v(314)
  buf u354 (ri_gpio_inten[17], 1'b0);  // ../RTL/gpio_apbif.v(314)
  buf u355 (ri_gpio_inten[18], 1'b0);  // ../RTL/gpio_apbif.v(314)
  buf u356 (ri_gpio_inten[19], 1'b0);  // ../RTL/gpio_apbif.v(314)
  buf u357 (ri_gpio_inten[20], 1'b0);  // ../RTL/gpio_apbif.v(314)
  buf u358 (ri_gpio_inten[21], 1'b0);  // ../RTL/gpio_apbif.v(314)
  buf u359 (ri_gpio_inten[22], 1'b0);  // ../RTL/gpio_apbif.v(314)
  buf u36 (ri_gpio_swporta_ddr[0], int_gpio_swporta_ddr[0]);  // ../RTL/gpio_apbif.v(273)
  buf u360 (ri_gpio_inten[23], 1'b0);  // ../RTL/gpio_apbif.v(314)
  buf u361 (ri_gpio_inten[24], 1'b0);  // ../RTL/gpio_apbif.v(314)
  buf u362 (ri_gpio_inten[25], 1'b0);  // ../RTL/gpio_apbif.v(314)
  buf u363 (ri_gpio_inten[26], 1'b0);  // ../RTL/gpio_apbif.v(314)
  buf u364 (ri_gpio_inten[27], 1'b0);  // ../RTL/gpio_apbif.v(314)
  buf u365 (ri_gpio_inten[28], 1'b0);  // ../RTL/gpio_apbif.v(314)
  buf u366 (ri_gpio_inten[29], 1'b0);  // ../RTL/gpio_apbif.v(314)
  buf u367 (ri_gpio_inten[30], 1'b0);  // ../RTL/gpio_apbif.v(314)
  buf u368 (ri_gpio_inten[31], 1'b0);  // ../RTL/gpio_apbif.v(314)
  buf u369 (gpio_inten[1], int_gpio_inten[1]);  // ../RTL/gpio_apbif.v(306)
  and u37 (n24, gpio_swporta_ctl_wen[0], gpio_swporta_ctl_wen[1]);  // ../RTL/gpio_apbif.v(281)
  buf u370 (gpio_inten[2], int_gpio_inten[2]);  // ../RTL/gpio_apbif.v(306)
  buf u371 (gpio_inten[3], int_gpio_inten[3]);  // ../RTL/gpio_apbif.v(306)
  buf u372 (gpio_inten[4], int_gpio_inten[4]);  // ../RTL/gpio_apbif.v(306)
  buf u373 (gpio_inten[5], int_gpio_inten[5]);  // ../RTL/gpio_apbif.v(306)
  buf u374 (gpio_inten[6], int_gpio_inten[6]);  // ../RTL/gpio_apbif.v(306)
  buf u375 (gpio_inten[7], int_gpio_inten[7]);  // ../RTL/gpio_apbif.v(306)
  and u376 (n25, gpio_inten_wen[2], gpio_inten_wen[3]);  // ../RTL/gpio_apbif.v(302)
  and u377 (n49, n30, n25);  // ../RTL/gpio_apbif.v(302)
  buf u378 (ri_gpio_swporta_ctl[1], int_gpio_swporta_ctl[1]);  // ../RTL/gpio_apbif.v(293)
  buf u379 (ri_gpio_swporta_ctl[2], int_gpio_swporta_ctl[2]);  // ../RTL/gpio_apbif.v(293)
  buf u38 (gpio_swporta_ctl[0], int_gpio_swporta_ctl[0]);  // ../RTL/gpio_apbif.v(285)
  buf u380 (ri_gpio_swporta_ctl[3], int_gpio_swporta_ctl[3]);  // ../RTL/gpio_apbif.v(293)
  buf u381 (ri_gpio_swporta_ctl[4], int_gpio_swporta_ctl[4]);  // ../RTL/gpio_apbif.v(293)
  buf u382 (ri_gpio_swporta_ctl[5], int_gpio_swporta_ctl[5]);  // ../RTL/gpio_apbif.v(293)
  buf u383 (ri_gpio_swporta_ctl[6], int_gpio_swporta_ctl[6]);  // ../RTL/gpio_apbif.v(293)
  buf u384 (ri_gpio_swporta_ctl[7], int_gpio_swporta_ctl[7]);  // ../RTL/gpio_apbif.v(293)
  buf u385 (ri_gpio_swporta_ctl[8], 1'b0);  // ../RTL/gpio_apbif.v(293)
  buf u386 (ri_gpio_swporta_ctl[9], 1'b0);  // ../RTL/gpio_apbif.v(293)
  buf u387 (ri_gpio_swporta_ctl[10], 1'b0);  // ../RTL/gpio_apbif.v(293)
  buf u388 (ri_gpio_swporta_ctl[11], 1'b0);  // ../RTL/gpio_apbif.v(293)
  buf u389 (ri_gpio_swporta_ctl[12], 1'b0);  // ../RTL/gpio_apbif.v(293)
  buf u39 (prdata[31], 1'b0);  // ../RTL/gpio_apbif.v(462)
  buf u390 (ri_gpio_swporta_ctl[13], 1'b0);  // ../RTL/gpio_apbif.v(293)
  buf u391 (ri_gpio_swporta_ctl[14], 1'b0);  // ../RTL/gpio_apbif.v(293)
  buf u392 (ri_gpio_swporta_ctl[15], 1'b0);  // ../RTL/gpio_apbif.v(293)
  buf u393 (ri_gpio_swporta_ctl[16], 1'b0);  // ../RTL/gpio_apbif.v(293)
  buf u394 (ri_gpio_swporta_ctl[17], 1'b0);  // ../RTL/gpio_apbif.v(293)
  buf u395 (ri_gpio_swporta_ctl[18], 1'b0);  // ../RTL/gpio_apbif.v(293)
  buf u396 (ri_gpio_swporta_ctl[19], 1'b0);  // ../RTL/gpio_apbif.v(293)
  buf u397 (ri_gpio_swporta_ctl[20], 1'b0);  // ../RTL/gpio_apbif.v(293)
  buf u398 (ri_gpio_swporta_ctl[21], 1'b0);  // ../RTL/gpio_apbif.v(293)
  buf u399 (ri_gpio_swporta_ctl[22], 1'b0);  // ../RTL/gpio_apbif.v(293)
  not u4 (n80, n57);  // ../RTL/gpio_apbif.v(453)
  buf u40 (prdata[12], 1'b0);  // ../RTL/gpio_apbif.v(462)
  buf u400 (ri_gpio_swporta_ctl[23], 1'b0);  // ../RTL/gpio_apbif.v(293)
  buf u401 (ri_gpio_swporta_ctl[24], 1'b0);  // ../RTL/gpio_apbif.v(293)
  buf u402 (ri_gpio_swporta_ctl[25], 1'b0);  // ../RTL/gpio_apbif.v(293)
  buf u403 (ri_gpio_swporta_ctl[26], 1'b0);  // ../RTL/gpio_apbif.v(293)
  buf u404 (ri_gpio_swporta_ctl[27], 1'b0);  // ../RTL/gpio_apbif.v(293)
  buf u405 (ri_gpio_swporta_ctl[28], 1'b0);  // ../RTL/gpio_apbif.v(293)
  buf u406 (ri_gpio_swporta_ctl[29], 1'b0);  // ../RTL/gpio_apbif.v(293)
  buf u407 (ri_gpio_swporta_ctl[30], 1'b0);  // ../RTL/gpio_apbif.v(293)
  buf u408 (ri_gpio_swporta_ctl[31], 1'b0);  // ../RTL/gpio_apbif.v(293)
  buf u409 (gpio_swporta_ctl[1], int_gpio_swporta_ctl[1]);  // ../RTL/gpio_apbif.v(285)
  buf u41 (ri_gpio_swporta_ctl[0], int_gpio_swporta_ctl[0]);  // ../RTL/gpio_apbif.v(293)
  buf u410 (gpio_swporta_ctl[2], int_gpio_swporta_ctl[2]);  // ../RTL/gpio_apbif.v(285)
  buf u411 (gpio_swporta_ctl[3], int_gpio_swporta_ctl[3]);  // ../RTL/gpio_apbif.v(285)
  buf u412 (gpio_swporta_ctl[4], int_gpio_swporta_ctl[4]);  // ../RTL/gpio_apbif.v(285)
  buf u413 (gpio_swporta_ctl[5], int_gpio_swporta_ctl[5]);  // ../RTL/gpio_apbif.v(285)
  buf u414 (gpio_swporta_ctl[6], int_gpio_swporta_ctl[6]);  // ../RTL/gpio_apbif.v(285)
  buf u415 (gpio_swporta_ctl[7], int_gpio_swporta_ctl[7]);  // ../RTL/gpio_apbif.v(285)
  and u416 (n23, gpio_swporta_ctl_wen[2], gpio_swporta_ctl_wen[3]);  // ../RTL/gpio_apbif.v(281)
  and u417 (n46, n24, n23);  // ../RTL/gpio_apbif.v(281)
  buf u418 (ri_gpio_swporta_ddr[1], int_gpio_swporta_ddr[1]);  // ../RTL/gpio_apbif.v(273)
  buf u419 (ri_gpio_swporta_ddr[2], int_gpio_swporta_ddr[2]);  // ../RTL/gpio_apbif.v(273)
  and u42 (n30, gpio_inten_wen[0], gpio_inten_wen[1]);  // ../RTL/gpio_apbif.v(302)
  buf u420 (ri_gpio_swporta_ddr[3], int_gpio_swporta_ddr[3]);  // ../RTL/gpio_apbif.v(273)
  buf u421 (ri_gpio_swporta_ddr[4], int_gpio_swporta_ddr[4]);  // ../RTL/gpio_apbif.v(273)
  buf u422 (ri_gpio_swporta_ddr[5], int_gpio_swporta_ddr[5]);  // ../RTL/gpio_apbif.v(273)
  buf u423 (ri_gpio_swporta_ddr[6], int_gpio_swporta_ddr[6]);  // ../RTL/gpio_apbif.v(273)
  buf u424 (ri_gpio_swporta_ddr[7], int_gpio_swporta_ddr[7]);  // ../RTL/gpio_apbif.v(273)
  buf u425 (ri_gpio_swporta_ddr[8], 1'b0);  // ../RTL/gpio_apbif.v(273)
  buf u426 (ri_gpio_swporta_ddr[9], 1'b0);  // ../RTL/gpio_apbif.v(273)
  buf u427 (ri_gpio_swporta_ddr[10], 1'b0);  // ../RTL/gpio_apbif.v(273)
  buf u428 (ri_gpio_swporta_ddr[11], 1'b0);  // ../RTL/gpio_apbif.v(273)
  buf u429 (ri_gpio_swporta_ddr[12], 1'b0);  // ../RTL/gpio_apbif.v(273)
  buf u43 (gpio_inten[0], int_gpio_inten[0]);  // ../RTL/gpio_apbif.v(306)
  buf u430 (ri_gpio_swporta_ddr[13], 1'b0);  // ../RTL/gpio_apbif.v(273)
  buf u431 (ri_gpio_swporta_ddr[14], 1'b0);  // ../RTL/gpio_apbif.v(273)
  buf u432 (ri_gpio_swporta_ddr[15], 1'b0);  // ../RTL/gpio_apbif.v(273)
  buf u433 (ri_gpio_swporta_ddr[16], 1'b0);  // ../RTL/gpio_apbif.v(273)
  buf u434 (ri_gpio_swporta_ddr[17], 1'b0);  // ../RTL/gpio_apbif.v(273)
  buf u435 (ri_gpio_swporta_ddr[18], 1'b0);  // ../RTL/gpio_apbif.v(273)
  buf u436 (ri_gpio_swporta_ddr[19], 1'b0);  // ../RTL/gpio_apbif.v(273)
  buf u437 (ri_gpio_swporta_ddr[20], 1'b0);  // ../RTL/gpio_apbif.v(273)
  buf u438 (ri_gpio_swporta_ddr[21], 1'b0);  // ../RTL/gpio_apbif.v(273)
  buf u439 (ri_gpio_swporta_ddr[22], 1'b0);  // ../RTL/gpio_apbif.v(273)
  buf u44 (prdata[30], 1'b0);  // ../RTL/gpio_apbif.v(462)
  buf u440 (ri_gpio_swporta_ddr[23], 1'b0);  // ../RTL/gpio_apbif.v(273)
  buf u441 (ri_gpio_swporta_ddr[24], 1'b0);  // ../RTL/gpio_apbif.v(273)
  buf u442 (ri_gpio_swporta_ddr[25], 1'b0);  // ../RTL/gpio_apbif.v(273)
  buf u443 (ri_gpio_swporta_ddr[26], 1'b0);  // ../RTL/gpio_apbif.v(273)
  buf u444 (ri_gpio_swporta_ddr[27], 1'b0);  // ../RTL/gpio_apbif.v(273)
  buf u445 (ri_gpio_swporta_ddr[28], 1'b0);  // ../RTL/gpio_apbif.v(273)
  buf u446 (ri_gpio_swporta_ddr[29], 1'b0);  // ../RTL/gpio_apbif.v(273)
  buf u447 (ri_gpio_swporta_ddr[30], 1'b0);  // ../RTL/gpio_apbif.v(273)
  buf u448 (ri_gpio_swporta_ddr[31], 1'b0);  // ../RTL/gpio_apbif.v(273)
  buf u449 (gpio_swporta_ddr[1], int_gpio_swporta_ddr[1]);  // ../RTL/gpio_apbif.v(265)
  buf u45 (prdata[11], 1'b0);  // ../RTL/gpio_apbif.v(462)
  buf u450 (gpio_swporta_ddr[2], int_gpio_swporta_ddr[2]);  // ../RTL/gpio_apbif.v(265)
  buf u451 (gpio_swporta_ddr[3], int_gpio_swporta_ddr[3]);  // ../RTL/gpio_apbif.v(265)
  buf u452 (gpio_swporta_ddr[4], int_gpio_swporta_ddr[4]);  // ../RTL/gpio_apbif.v(265)
  buf u453 (gpio_swporta_ddr[5], int_gpio_swporta_ddr[5]);  // ../RTL/gpio_apbif.v(265)
  buf u454 (gpio_swporta_ddr[6], int_gpio_swporta_ddr[6]);  // ../RTL/gpio_apbif.v(265)
  buf u455 (gpio_swporta_ddr[7], int_gpio_swporta_ddr[7]);  // ../RTL/gpio_apbif.v(265)
  and u456 (n18, gpio_swporta_ddr_wen[2], gpio_swporta_ddr_wen[3]);  // ../RTL/gpio_apbif.v(261)
  and u457 (n43, n22, n18);  // ../RTL/gpio_apbif.v(261)
  buf u458 (ri_gpio_swporta_dr[1], int_gpio_swporta_dr[1]);  // ../RTL/gpio_apbif.v(253)
  buf u459 (ri_gpio_swporta_dr[2], int_gpio_swporta_dr[2]);  // ../RTL/gpio_apbif.v(253)
  buf u46 (ri_gpio_inten[0], int_gpio_inten[0]);  // ../RTL/gpio_apbif.v(314)
  buf u460 (ri_gpio_swporta_dr[3], int_gpio_swporta_dr[3]);  // ../RTL/gpio_apbif.v(253)
  buf u461 (ri_gpio_swporta_dr[4], int_gpio_swporta_dr[4]);  // ../RTL/gpio_apbif.v(253)
  buf u462 (ri_gpio_swporta_dr[5], int_gpio_swporta_dr[5]);  // ../RTL/gpio_apbif.v(253)
  buf u463 (ri_gpio_swporta_dr[6], int_gpio_swporta_dr[6]);  // ../RTL/gpio_apbif.v(253)
  buf u464 (ri_gpio_swporta_dr[7], int_gpio_swporta_dr[7]);  // ../RTL/gpio_apbif.v(253)
  buf u465 (ri_gpio_swporta_dr[8], 1'b0);  // ../RTL/gpio_apbif.v(253)
  buf u466 (ri_gpio_swporta_dr[9], 1'b0);  // ../RTL/gpio_apbif.v(253)
  buf u467 (ri_gpio_swporta_dr[10], 1'b0);  // ../RTL/gpio_apbif.v(253)
  buf u468 (ri_gpio_swporta_dr[11], 1'b0);  // ../RTL/gpio_apbif.v(253)
  buf u469 (ri_gpio_swporta_dr[12], 1'b0);  // ../RTL/gpio_apbif.v(253)
  and u47 (n32, gpio_intmask_wen[0], gpio_intmask_wen[1]);  // ../RTL/gpio_apbif.v(322)
  buf u470 (ri_gpio_swporta_dr[13], 1'b0);  // ../RTL/gpio_apbif.v(253)
  buf u471 (ri_gpio_swporta_dr[14], 1'b0);  // ../RTL/gpio_apbif.v(253)
  buf u472 (ri_gpio_swporta_dr[15], 1'b0);  // ../RTL/gpio_apbif.v(253)
  buf u473 (ri_gpio_swporta_dr[16], 1'b0);  // ../RTL/gpio_apbif.v(253)
  buf u474 (ri_gpio_swporta_dr[17], 1'b0);  // ../RTL/gpio_apbif.v(253)
  buf u475 (ri_gpio_swporta_dr[18], 1'b0);  // ../RTL/gpio_apbif.v(253)
  buf u476 (ri_gpio_swporta_dr[19], 1'b0);  // ../RTL/gpio_apbif.v(253)
  buf u477 (ri_gpio_swporta_dr[20], 1'b0);  // ../RTL/gpio_apbif.v(253)
  buf u478 (ri_gpio_swporta_dr[21], 1'b0);  // ../RTL/gpio_apbif.v(253)
  buf u479 (ri_gpio_swporta_dr[22], 1'b0);  // ../RTL/gpio_apbif.v(253)
  buf u48 (gpio_intmask[0], int_gpio_intmask[0]);  // ../RTL/gpio_apbif.v(326)
  buf u480 (ri_gpio_swporta_dr[23], 1'b0);  // ../RTL/gpio_apbif.v(253)
  buf u481 (ri_gpio_swporta_dr[24], 1'b0);  // ../RTL/gpio_apbif.v(253)
  buf u482 (ri_gpio_swporta_dr[25], 1'b0);  // ../RTL/gpio_apbif.v(253)
  buf u483 (ri_gpio_swporta_dr[26], 1'b0);  // ../RTL/gpio_apbif.v(253)
  buf u484 (ri_gpio_swporta_dr[27], 1'b0);  // ../RTL/gpio_apbif.v(253)
  buf u485 (ri_gpio_swporta_dr[28], 1'b0);  // ../RTL/gpio_apbif.v(253)
  buf u486 (ri_gpio_swporta_dr[29], 1'b0);  // ../RTL/gpio_apbif.v(253)
  buf u487 (ri_gpio_swporta_dr[30], 1'b0);  // ../RTL/gpio_apbif.v(253)
  buf u488 (ri_gpio_swporta_dr[31], 1'b0);  // ../RTL/gpio_apbif.v(253)
  buf u489 (gpio_swporta_dr[1], int_gpio_swporta_dr[1]);  // ../RTL/gpio_apbif.v(245)
  buf u49 (prdata[29], 1'b0);  // ../RTL/gpio_apbif.v(462)
  buf u490 (gpio_swporta_dr[2], int_gpio_swporta_dr[2]);  // ../RTL/gpio_apbif.v(245)
  buf u491 (gpio_swporta_dr[3], int_gpio_swporta_dr[3]);  // ../RTL/gpio_apbif.v(245)
  buf u492 (gpio_swporta_dr[4], int_gpio_swporta_dr[4]);  // ../RTL/gpio_apbif.v(245)
  buf u493 (gpio_swporta_dr[5], int_gpio_swporta_dr[5]);  // ../RTL/gpio_apbif.v(245)
  buf u494 (gpio_swporta_dr[6], int_gpio_swporta_dr[6]);  // ../RTL/gpio_apbif.v(245)
  buf u495 (gpio_swporta_dr[7], int_gpio_swporta_dr[7]);  // ../RTL/gpio_apbif.v(245)
  and u496 (n16, gpio_swporta_dr_wen[2], gpio_swporta_dr_wen[3]);  // ../RTL/gpio_apbif.v(241)
  and u497 (n40, n17, n16);  // ../RTL/gpio_apbif.v(241)
  buf u498 (gpio_swporta_ctl_wen[1], 1'b0);  // ../RTL/gpio_apbif.v(180)
  buf u499 (gpio_swporta_ctl_wen[2], 1'b0);  // ../RTL/gpio_apbif.v(180)
  or u5 (n57, n73, n60);  // ../RTL/gpio_apbif.v(453)
  buf u50 (prdata[10], 1'b0);  // ../RTL/gpio_apbif.v(462)
  buf u500 (gpio_swporta_ctl_wen[3], 1'b0);  // ../RTL/gpio_apbif.v(180)
  buf u501 (pwdata_int[1], pwdata[1]);  // ../RTL/gpio_apbif.v(147)
  buf u502 (pwdata_int[2], pwdata[2]);  // ../RTL/gpio_apbif.v(147)
  buf u503 (pwdata_int[3], pwdata[3]);  // ../RTL/gpio_apbif.v(147)
  buf u504 (pwdata_int[4], pwdata[4]);  // ../RTL/gpio_apbif.v(147)
  buf u505 (pwdata_int[5], pwdata[5]);  // ../RTL/gpio_apbif.v(147)
  buf u506 (pwdata_int[6], pwdata[6]);  // ../RTL/gpio_apbif.v(147)
  buf u507 (pwdata_int[7], pwdata[7]);  // ../RTL/gpio_apbif.v(147)
  buf u508 (pwdata_int[8], pwdata[8]);  // ../RTL/gpio_apbif.v(147)
  buf u509 (pwdata_int[9], pwdata[9]);  // ../RTL/gpio_apbif.v(147)
  buf u51 (ri_gpio_intmask[0], int_gpio_intmask[0]);  // ../RTL/gpio_apbif.v(334)
  buf u510 (pwdata_int[10], pwdata[10]);  // ../RTL/gpio_apbif.v(147)
  buf u511 (pwdata_int[11], pwdata[11]);  // ../RTL/gpio_apbif.v(147)
  buf u512 (pwdata_int[12], pwdata[12]);  // ../RTL/gpio_apbif.v(147)
  buf u513 (pwdata_int[13], pwdata[13]);  // ../RTL/gpio_apbif.v(147)
  buf u514 (pwdata_int[14], pwdata[14]);  // ../RTL/gpio_apbif.v(147)
  buf u515 (pwdata_int[15], pwdata[15]);  // ../RTL/gpio_apbif.v(147)
  buf u516 (pwdata_int[16], pwdata[16]);  // ../RTL/gpio_apbif.v(147)
  buf u517 (pwdata_int[17], pwdata[17]);  // ../RTL/gpio_apbif.v(147)
  buf u518 (pwdata_int[18], pwdata[18]);  // ../RTL/gpio_apbif.v(147)
  buf u519 (pwdata_int[19], pwdata[19]);  // ../RTL/gpio_apbif.v(147)
  and u52 (n5, gpio_inttype_level_wen[0], gpio_inttype_level_wen[1]);  // ../RTL/gpio_apbif.v(342)
  buf u520 (pwdata_int[20], pwdata[20]);  // ../RTL/gpio_apbif.v(147)
  buf u521 (pwdata_int[21], pwdata[21]);  // ../RTL/gpio_apbif.v(147)
  buf u522 (pwdata_int[22], pwdata[22]);  // ../RTL/gpio_apbif.v(147)
  buf u523 (pwdata_int[23], pwdata[23]);  // ../RTL/gpio_apbif.v(147)
  buf u524 (pwdata_int[24], pwdata[24]);  // ../RTL/gpio_apbif.v(147)
  buf u525 (pwdata_int[25], pwdata[25]);  // ../RTL/gpio_apbif.v(147)
  buf u526 (pwdata_int[26], pwdata[26]);  // ../RTL/gpio_apbif.v(147)
  buf u527 (pwdata_int[27], pwdata[27]);  // ../RTL/gpio_apbif.v(147)
  buf u528 (pwdata_int[28], pwdata[28]);  // ../RTL/gpio_apbif.v(147)
  buf u529 (pwdata_int[29], pwdata[29]);  // ../RTL/gpio_apbif.v(147)
  buf u53 (gpio_inttype_level[0], int_gpio_inttype_level[0]);  // ../RTL/gpio_apbif.v(346)
  buf u530 (pwdata_int[30], pwdata[30]);  // ../RTL/gpio_apbif.v(147)
  buf u531 (pwdata_int[31], pwdata[31]);  // ../RTL/gpio_apbif.v(147)
  buf u54 (prdata[28], 1'b0);  // ../RTL/gpio_apbif.v(462)
  buf u55 (prdata[9], 1'b0);  // ../RTL/gpio_apbif.v(462)
  buf u56 (ri_gpio_inttype_level[0], int_gpio_inttype_level[0]);  // ../RTL/gpio_apbif.v(354)
  and u57 (n42, gpio_int_polarity_wen[0], gpio_int_polarity_wen[1]);  // ../RTL/gpio_apbif.v(362)
  buf u58 (gpio_int_polarity[0], int_gpio_int_polarity[0]);  // ../RTL/gpio_apbif.v(366)
  buf u59 (prdata[27], 1'b0);  // ../RTL/gpio_apbif.v(462)
  and u6 (n0, psel, penable);  // ../RTL/gpio_apbif.v(161)
  buf u60 (prdata[8], 1'b0);  // ../RTL/gpio_apbif.v(462)
  buf u61 (ri_gpio_int_polarity[0], int_gpio_int_polarity[0]);  // ../RTL/gpio_apbif.v(374)
  buf u62 (gpio_ls_sync, int_gpio_ls_sync[0]);  // ../RTL/gpio_apbif.v(386)
  and u63 (n48, gpio_ls_sync_wen[0], gpio_ls_sync_wen[1]);  // ../RTL/gpio_apbif.v(382)
  buf u64 (ri_gpio_ls_sync[0], int_gpio_ls_sync[0]);  // ../RTL/gpio_apbif.v(394)
  and u65 (n54, gpio_porta_eoi_wen[0], gpio_porta_eoi_wen[1]);  // ../RTL/gpio_apbif.v(403)
  buf u66 (gpio_porta_eoi[0], int_gpio_porta_eoi[0]);  // ../RTL/gpio_apbif.v(408)
  buf u67 (ri_gpio_raw_intstatus[0], gpio_raw_intstatus[0]);  // ../RTL/gpio_apbif.v(421)
  buf u68 (ri_gpio_intstatus[0], gpio_intstatus[0]);  // ../RTL/gpio_apbif.v(421)
  buf u69 (prdata[26], 1'b0);  // ../RTL/gpio_apbif.v(462)
  or u7 (n60, n70, n64);  // ../RTL/gpio_apbif.v(453)
  buf u70 (prdata[7], iprdata[7]);  // ../RTL/gpio_apbif.v(462)
  not u71 (n65, pwrite);  // ../RTL/gpio_apbif.v(439)
  buf u72 (prdata[25], 1'b0);  // ../RTL/gpio_apbif.v(462)
  and u73 (n66, n65, psel);  // ../RTL/gpio_apbif.v(439)
  not u74 (n67, penable);  // ../RTL/gpio_apbif.v(439)
  and u75 (n68, n66, n67);  // ../RTL/gpio_apbif.v(439)
  buf u76 (prdata[6], iprdata[6]);  // ../RTL/gpio_apbif.v(462)
  buf u77 (prdata[5], iprdata[5]);  // ../RTL/gpio_apbif.v(462)
  buf u78 (prdata[4], iprdata[4]);  // ../RTL/gpio_apbif.v(462)
  buf u79 (prdata[3], iprdata[3]);  // ../RTL/gpio_apbif.v(462)
  and u8 (n6, n0, pwrite);  // ../RTL/gpio_apbif.v(161)
  buf u80 (prdata[2], iprdata[2]);  // ../RTL/gpio_apbif.v(462)
  buf u81 (prdata[1], iprdata[1]);  // ../RTL/gpio_apbif.v(462)
  buf u82 (prdata[0], iprdata[0]);  // ../RTL/gpio_apbif.v(462)
  buf u83 (ri_gpio_ext_porta_rb[0], gpio_ext_porta_rb[0]);  // ../RTL/gpio_apbif.v(430)
  buf u84 (ri_gpio_ext_porta_rb[3], gpio_ext_porta_rb[3]);  // ../RTL/gpio_apbif.v(430)
  or u85 (n78, n79, n11);  // ../RTL/gpio_apbif.v(453)
  buf u86 (ri_gpio_ext_porta_rb[4], gpio_ext_porta_rb[4]);  // ../RTL/gpio_apbif.v(430)
  buf u87 (ri_gpio_ext_porta_rb[5], gpio_ext_porta_rb[5]);  // ../RTL/gpio_apbif.v(430)
  buf u88 (ri_gpio_ext_porta_rb[6], gpio_ext_porta_rb[6]);  // ../RTL/gpio_apbif.v(430)
  buf u89 (ri_gpio_ext_porta_rb[7], gpio_ext_porta_rb[7]);  // ../RTL/gpio_apbif.v(430)
  or u9 (n64, n71, n69);  // ../RTL/gpio_apbif.v(453)
  buf u90 (ri_gpio_ext_porta_rb[8], 1'b0);  // ../RTL/gpio_apbif.v(430)
  buf u91 (ri_gpio_ext_porta_rb[9], 1'b0);  // ../RTL/gpio_apbif.v(430)
  buf u92 (ri_gpio_ext_porta_rb[10], 1'b0);  // ../RTL/gpio_apbif.v(430)
  buf u93 (ri_gpio_ext_porta_rb[11], 1'b0);  // ../RTL/gpio_apbif.v(430)
  buf u94 (ri_gpio_ext_porta_rb[12], 1'b0);  // ../RTL/gpio_apbif.v(430)
  buf u95 (ri_gpio_ext_porta_rb[13], 1'b0);  // ../RTL/gpio_apbif.v(430)
  buf u96 (ri_gpio_ext_porta_rb[14], 1'b0);  // ../RTL/gpio_apbif.v(430)
  buf u97 (ri_gpio_ext_porta_rb[15], 1'b0);  // ../RTL/gpio_apbif.v(430)
  buf u98 (ri_gpio_ext_porta_rb[16], 1'b0);  // ../RTL/gpio_apbif.v(430)
  buf u99 (ri_gpio_ext_porta_rb[17], 1'b0);  // ../RTL/gpio_apbif.v(430)

endmodule 

module gpio_ctrl  // ../RTL/gpio_ctrl.v(22)
  (
  gpio_ext_porta,
  gpio_int_polarity,
  gpio_inten,
  gpio_intmask,
  gpio_inttype_level,
  gpio_ls_sync,
  gpio_porta_eoi,
  gpio_swporta_ctl,
  gpio_swporta_ddr,
  gpio_swporta_dr,
  pclk,
  pclk_intr,
  presetn,
  gpio_ext_porta_rb,
  gpio_intr,
  gpio_intr_flag_int,
  gpio_intr_int,
  gpio_intrclk_en,
  gpio_porta_ddr,
  gpio_porta_dr,
  gpio_raw_intstatus
  );

  input [7:0] gpio_ext_porta;  // ../RTL/gpio_ctrl.v(47)
  input [7:0] gpio_int_polarity;  // ../RTL/gpio_ctrl.v(48)
  input [7:0] gpio_inten;  // ../RTL/gpio_ctrl.v(49)
  input [7:0] gpio_intmask;  // ../RTL/gpio_ctrl.v(50)
  input [7:0] gpio_inttype_level;  // ../RTL/gpio_ctrl.v(51)
  input gpio_ls_sync;  // ../RTL/gpio_ctrl.v(52)
  input [7:0] gpio_porta_eoi;  // ../RTL/gpio_ctrl.v(53)
  input [7:0] gpio_swporta_ctl;  // ../RTL/gpio_ctrl.v(54)
  input [7:0] gpio_swporta_ddr;  // ../RTL/gpio_ctrl.v(55)
  input [7:0] gpio_swporta_dr;  // ../RTL/gpio_ctrl.v(56)
  input pclk;  // ../RTL/gpio_ctrl.v(57)
  input pclk_intr;  // ../RTL/gpio_ctrl.v(58)
  input presetn;  // ../RTL/gpio_ctrl.v(59)
  output [7:0] gpio_ext_porta_rb;  // ../RTL/gpio_ctrl.v(60)
  output [7:0] gpio_intr;  // ../RTL/gpio_ctrl.v(61)
  output gpio_intr_flag_int;  // ../RTL/gpio_ctrl.v(62)
  output [7:0] gpio_intr_int;  // ../RTL/gpio_ctrl.v(63)
  output gpio_intrclk_en;  // ../RTL/gpio_ctrl.v(64)
  output [7:0] gpio_porta_ddr;  // ../RTL/gpio_ctrl.v(65)
  output [7:0] gpio_porta_dr;  // ../RTL/gpio_ctrl.v(66)
  output [7:0] gpio_raw_intstatus;  // ../RTL/gpio_ctrl.v(67)

  wire [7:0] ed_int_d1;  // ../RTL/gpio_ctrl.v(70)
  wire [7:0] ed_out;  // ../RTL/gpio_ctrl.v(71)
  wire [7:0] ed_rf;  // ../RTL/gpio_ctrl.v(86)
  wire [7:0] gpio_ext_porta_int;  // ../RTL/gpio_ctrl.v(72)
  wire [7:0] gpio_intr_ed_pm;  // ../RTL/gpio_ctrl.v(74)
  wire [7:0] gpio_swporta_ctl_internal;  // ../RTL/gpio_ctrl.v(100)
  wire [7:0] int_gpio_raw_intstatus;  // ../RTL/gpio_ctrl.v(78)
  wire [7:0] int_in;  // ../RTL/gpio_ctrl.v(103)
  wire [7:0] int_pre_in;  // ../RTL/gpio_ctrl.v(79)
  wire [7:0] int_s1;  // ../RTL/gpio_ctrl.v(80)
  wire [7:0] int_sy_in;  // ../RTL/gpio_ctrl.v(81)
  wire [7:0] intrclk_en;  // ../RTL/gpio_ctrl.v(82)
  wire [7:0] ls_int_in;  // ../RTL/gpio_ctrl.v(83)
  wire [7:0] n117;
  wire gpio_intrclk_en_int;  // ../RTL/gpio_ctrl.v(94)
  wire n0;
  wire n1;
  wire n10;
  wire n100;
  wire n101;
  wire n102;
  wire n103;
  wire n104;
  wire n105;
  wire n106;
  wire n107;
  wire n108;
  wire n109;
  wire n11;
  wire n110;
  wire n111;
  wire n112;
  wire n113;
  wire n114;
  wire n115;
  wire n116;
  wire n12;
  wire n13;
  wire n14;
  wire n15;
  wire n16;
  wire n17;
  wire n18;
  wire n19;
  wire n2;
  wire n20;
  wire n21;
  wire n22;
  wire n23;
  wire n24;
  wire n25;
  wire n26;
  wire n27;
  wire n28;
  wire n29;
  wire n3;
  wire n30;
  wire n31;
  wire n32;
  wire n33;
  wire n34;
  wire n35;
  wire n36;
  wire n37;
  wire n38;
  wire n39;
  wire n4;
  wire n40;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n5;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n6;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n65;
  wire n66;
  wire n67;
  wire n68;
  wire n69;
  wire n7;
  wire n70;
  wire n71;
  wire n72;
  wire n73;
  wire n74;
  wire n75;
  wire n76;
  wire n77;
  wire n78;
  wire n79;
  wire n8;
  wire n80;
  wire n81;
  wire n82;
  wire n83;
  wire n84;
  wire n85;
  wire n86;
  wire n87;
  wire n88;
  wire n89;
  wire n9;
  wire n90;
  wire n91;
  wire n92;
  wire n93;
  wire n94;
  wire n95;
  wire n96;
  wire n97;
  wire n98;
  wire n99;

  AL_DFF gpio_intrclk_en_reg (
    .clk(pclk),
    .d(gpio_intrclk_en_int),
    .reset(n17),
    .set(1'b0),
    .q(gpio_intrclk_en));  // ../RTL/gpio_ctrl.v(147)
  reg_ar_as_w8 reg0 (
    .clk(pclk_intr),
    .d(int_sy_in),
    .reset({n17,n17,n17,n17,n17,n17,n17,n17}),
    .set(8'b00000000),
    .q(int_s1));  // ../RTL/gpio_ctrl.v(184)
  reg_ar_as_w8 reg1 (
    .clk(pclk_intr),
    .d(int_s1),
    .reset({n17,n17,n17,n17,n17,n17,n17,n17}),
    .set(8'b00000000),
    .q(int_pre_in));  // ../RTL/gpio_ctrl.v(192)
  reg_ar_as_w8 reg2 (
    .clk(pclk_intr),
    .d(int_in),
    .reset({n17,n17,n17,n17,n17,n17,n17,n17}),
    .set(8'b00000000),
    .q(ed_int_d1));  // ../RTL/gpio_ctrl.v(203)
  reg_ar_as_w8 reg3 (
    .clk(pclk_intr),
    .d({n84,n76,n68,n60,n52,n44,n36,n28}),
    .reset({n17,n17,n17,n17,n17,n17,n17,n17}),
    .set(8'b00000000),
    .q(gpio_intr_ed_pm));  // ../RTL/gpio_ctrl.v(248)
  AL_MUX u10 (
    .i0(gpio_ls_sync),
    .i1(1'b1),
    .sel(gpio_inttype_level[4]),
    .o(n4));  // ../RTL/gpio_ctrl.v(133)
  not u100 (n56, gpio_swporta_ctl_internal[4]);  // ../RTL/gpio_ctrl.v(243)
  and u101 (n57, n55, n56);  // ../RTL/gpio_ctrl.v(243)
  buf u102 (int_sy_in[4], gpio_ext_porta_int[4]);  // ../RTL/gpio_ctrl.v(176)
  AL_MUX u103 (
    .i0(gpio_intr_ed_pm[4]),
    .i1(1'b0),
    .sel(gpio_porta_eoi[4]),
    .o(n58));  // ../RTL/gpio_ctrl.v(247)
  AL_MUX u104 (
    .i0(n58),
    .i1(1'b1),
    .sel(n57),
    .o(n59));  // ../RTL/gpio_ctrl.v(247)
  AL_MUX u105 (
    .i0(1'b0),
    .i1(n59),
    .sel(gpio_inten[4]),
    .o(n60));  // ../RTL/gpio_ctrl.v(247)
  buf u106 (gpio_porta_dr[7], gpio_swporta_dr[7]);  // ../RTL/gpio_ctrl.v(316)
  buf u107 (int_sy_in[3], gpio_ext_porta_int[3]);  // ../RTL/gpio_ctrl.v(176)
  buf u108 (int_sy_in[2], gpio_ext_porta_int[2]);  // ../RTL/gpio_ctrl.v(176)
  and u109 (n61, ed_out[5], gpio_inten[5]);  // ../RTL/gpio_ctrl.v(241)
  AL_MUX u11 (
    .i0(1'b0),
    .i1(n4),
    .sel(gpio_inten[4]),
    .o(intrclk_en[4]));  // ../RTL/gpio_ctrl.v(135)
  not u110 (n62, gpio_swporta_ddr[5]);  // ../RTL/gpio_ctrl.v(242)
  and u111 (n63, n61, n62);  // ../RTL/gpio_ctrl.v(242)
  not u112 (n64, gpio_swporta_ctl_internal[5]);  // ../RTL/gpio_ctrl.v(243)
  and u113 (n65, n63, n64);  // ../RTL/gpio_ctrl.v(243)
  buf u114 (int_sy_in[1], gpio_ext_porta_int[1]);  // ../RTL/gpio_ctrl.v(176)
  AL_MUX u115 (
    .i0(gpio_intr_ed_pm[5]),
    .i1(1'b0),
    .sel(gpio_porta_eoi[5]),
    .o(n66));  // ../RTL/gpio_ctrl.v(247)
  AL_MUX u116 (
    .i0(n66),
    .i1(1'b1),
    .sel(n65),
    .o(n67));  // ../RTL/gpio_ctrl.v(247)
  AL_MUX u117 (
    .i0(1'b0),
    .i1(n67),
    .sel(gpio_inten[5]),
    .o(n68));  // ../RTL/gpio_ctrl.v(247)
  buf u118 (gpio_porta_dr[6], gpio_swporta_dr[6]);  // ../RTL/gpio_ctrl.v(316)
  buf u119 (int_in[7], int_pre_in[7]);  // ../RTL/gpio_ctrl.v(195)
  AL_MUX u12 (
    .i0(gpio_ls_sync),
    .i1(1'b1),
    .sel(gpio_inttype_level[5]),
    .o(n5));  // ../RTL/gpio_ctrl.v(133)
  buf u120 (int_in[6], int_pre_in[6]);  // ../RTL/gpio_ctrl.v(195)
  and u121 (n69, ed_out[6], gpio_inten[6]);  // ../RTL/gpio_ctrl.v(241)
  not u122 (n70, gpio_swporta_ddr[6]);  // ../RTL/gpio_ctrl.v(242)
  and u123 (n71, n69, n70);  // ../RTL/gpio_ctrl.v(242)
  not u124 (n72, gpio_swporta_ctl_internal[6]);  // ../RTL/gpio_ctrl.v(243)
  and u125 (n73, n71, n72);  // ../RTL/gpio_ctrl.v(243)
  buf u126 (int_in[5], int_pre_in[5]);  // ../RTL/gpio_ctrl.v(195)
  AL_MUX u127 (
    .i0(gpio_intr_ed_pm[6]),
    .i1(1'b0),
    .sel(gpio_porta_eoi[6]),
    .o(n74));  // ../RTL/gpio_ctrl.v(247)
  AL_MUX u128 (
    .i0(n74),
    .i1(1'b1),
    .sel(n73),
    .o(n75));  // ../RTL/gpio_ctrl.v(247)
  AL_MUX u129 (
    .i0(1'b0),
    .i1(n75),
    .sel(gpio_inten[6]),
    .o(n76));  // ../RTL/gpio_ctrl.v(247)
  AL_MUX u13 (
    .i0(1'b0),
    .i1(n5),
    .sel(gpio_inten[5]),
    .o(intrclk_en[5]));  // ../RTL/gpio_ctrl.v(135)
  buf u130 (gpio_porta_dr[5], gpio_swporta_dr[5]);  // ../RTL/gpio_ctrl.v(316)
  buf u131 (int_in[4], int_pre_in[4]);  // ../RTL/gpio_ctrl.v(195)
  buf u132 (int_in[3], int_pre_in[3]);  // ../RTL/gpio_ctrl.v(195)
  and u133 (n77, ed_out[7], gpio_inten[7]);  // ../RTL/gpio_ctrl.v(241)
  not u134 (n78, gpio_swporta_ddr[7]);  // ../RTL/gpio_ctrl.v(242)
  and u135 (n79, n77, n78);  // ../RTL/gpio_ctrl.v(242)
  not u136 (n80, gpio_swporta_ctl_internal[7]);  // ../RTL/gpio_ctrl.v(243)
  and u137 (n81, n79, n80);  // ../RTL/gpio_ctrl.v(243)
  buf u138 (int_in[2], int_pre_in[2]);  // ../RTL/gpio_ctrl.v(195)
  AL_MUX u139 (
    .i0(gpio_intr_ed_pm[7]),
    .i1(1'b0),
    .sel(gpio_porta_eoi[7]),
    .o(n82));  // ../RTL/gpio_ctrl.v(247)
  AL_MUX u14 (
    .i0(gpio_ls_sync),
    .i1(1'b1),
    .sel(gpio_inttype_level[6]),
    .o(n6));  // ../RTL/gpio_ctrl.v(133)
  AL_MUX u140 (
    .i0(n82),
    .i1(1'b1),
    .sel(n81),
    .o(n83));  // ../RTL/gpio_ctrl.v(247)
  AL_MUX u141 (
    .i0(1'b0),
    .i1(n83),
    .sel(gpio_inten[7]),
    .o(n84));  // ../RTL/gpio_ctrl.v(247)
  buf u142 (gpio_swporta_ctl_internal[0], gpio_swporta_ctl[0]);  // ../RTL/gpio_ctrl.v(228)
  buf u143 (int_in[1], int_pre_in[1]);  // ../RTL/gpio_ctrl.v(195)
  xor u144 (ed_rf[7], int_in[7], ed_int_d1[7]);  // ../RTL/gpio_ctrl.v(206)
  or u145 (n85, gpio_swporta_ddr[0], gpio_swporta_ctl_internal[0]);  // ../RTL/gpio_ctrl.v(269)
  xor u146 (ed_rf[6], int_in[6], ed_int_d1[6]);  // ../RTL/gpio_ctrl.v(206)
  AL_MUX u147 (
    .i0(int_sy_in[0]),
    .i1(int_in[0]),
    .sel(gpio_ls_sync),
    .o(n86));  // ../RTL/gpio_ctrl.v(275)
  AL_MUX u148 (
    .i0(n86),
    .i1(1'b0),
    .sel(n85),
    .o(ls_int_in[0]));  // ../RTL/gpio_ctrl.v(275)
  xor u149 (ed_rf[5], int_in[5], ed_int_d1[5]);  // ../RTL/gpio_ctrl.v(206)
  AL_MUX u15 (
    .i0(1'b0),
    .i1(n6),
    .sel(gpio_inten[6]),
    .o(intrclk_en[6]));  // ../RTL/gpio_ctrl.v(135)
  xor u150 (ed_rf[4], int_in[4], ed_int_d1[4]);  // ../RTL/gpio_ctrl.v(206)
  or u151 (n87, gpio_swporta_ddr[1], gpio_swporta_ctl_internal[1]);  // ../RTL/gpio_ctrl.v(269)
  xor u152 (ed_rf[3], int_in[3], ed_int_d1[3]);  // ../RTL/gpio_ctrl.v(206)
  AL_MUX u153 (
    .i0(int_sy_in[1]),
    .i1(int_in[1]),
    .sel(gpio_ls_sync),
    .o(n88));  // ../RTL/gpio_ctrl.v(275)
  AL_MUX u154 (
    .i0(n88),
    .i1(1'b0),
    .sel(n87),
    .o(ls_int_in[1]));  // ../RTL/gpio_ctrl.v(275)
  xor u155 (ed_rf[2], int_in[2], ed_int_d1[2]);  // ../RTL/gpio_ctrl.v(206)
  xor u156 (ed_rf[1], int_in[1], ed_int_d1[1]);  // ../RTL/gpio_ctrl.v(206)
  or u157 (n89, gpio_swporta_ddr[2], gpio_swporta_ctl_internal[2]);  // ../RTL/gpio_ctrl.v(269)
  buf u158 (gpio_swporta_ctl_internal[7], gpio_swporta_ctl[7]);  // ../RTL/gpio_ctrl.v(228)
  AL_MUX u159 (
    .i0(int_sy_in[2]),
    .i1(int_in[2]),
    .sel(gpio_ls_sync),
    .o(n90));  // ../RTL/gpio_ctrl.v(275)
  AL_MUX u16 (
    .i0(gpio_ls_sync),
    .i1(1'b1),
    .sel(gpio_inttype_level[7]),
    .o(n7));  // ../RTL/gpio_ctrl.v(133)
  AL_MUX u160 (
    .i0(n90),
    .i1(1'b0),
    .sel(n89),
    .o(ls_int_in[2]));  // ../RTL/gpio_ctrl.v(275)
  buf u161 (gpio_swporta_ctl_internal[6], gpio_swporta_ctl[6]);  // ../RTL/gpio_ctrl.v(228)
  buf u162 (gpio_swporta_ctl_internal[5], gpio_swporta_ctl[5]);  // ../RTL/gpio_ctrl.v(228)
  or u163 (n91, gpio_swporta_ddr[3], gpio_swporta_ctl_internal[3]);  // ../RTL/gpio_ctrl.v(269)
  buf u164 (gpio_swporta_ctl_internal[4], gpio_swporta_ctl[4]);  // ../RTL/gpio_ctrl.v(228)
  AL_MUX u165 (
    .i0(int_sy_in[3]),
    .i1(int_in[3]),
    .sel(gpio_ls_sync),
    .o(n92));  // ../RTL/gpio_ctrl.v(275)
  AL_MUX u166 (
    .i0(n92),
    .i1(1'b0),
    .sel(n91),
    .o(ls_int_in[3]));  // ../RTL/gpio_ctrl.v(275)
  buf u167 (gpio_swporta_ctl_internal[3], gpio_swporta_ctl[3]);  // ../RTL/gpio_ctrl.v(228)
  buf u168 (gpio_swporta_ctl_internal[2], gpio_swporta_ctl[2]);  // ../RTL/gpio_ctrl.v(228)
  or u169 (n93, gpio_swporta_ddr[4], gpio_swporta_ctl_internal[4]);  // ../RTL/gpio_ctrl.v(269)
  AL_MUX u17 (
    .i0(1'b0),
    .i1(n7),
    .sel(gpio_inten[7]),
    .o(intrclk_en[7]));  // ../RTL/gpio_ctrl.v(135)
  buf u170 (gpio_swporta_ctl_internal[1], gpio_swporta_ctl[1]);  // ../RTL/gpio_ctrl.v(228)
  AL_MUX u171 (
    .i0(int_sy_in[4]),
    .i1(int_in[4]),
    .sel(gpio_ls_sync),
    .o(n94));  // ../RTL/gpio_ctrl.v(275)
  AL_MUX u172 (
    .i0(n94),
    .i1(1'b0),
    .sel(n93),
    .o(ls_int_in[4]));  // ../RTL/gpio_ctrl.v(275)
  and u173 (ed_out[7], ed_rf[7], int_in[7]);  // ../RTL/gpio_ctrl.v(218)
  and u174 (ed_out[6], ed_rf[6], int_in[6]);  // ../RTL/gpio_ctrl.v(218)
  or u175 (n95, gpio_swporta_ddr[5], gpio_swporta_ctl_internal[5]);  // ../RTL/gpio_ctrl.v(269)
  and u176 (ed_out[5], ed_rf[5], int_in[5]);  // ../RTL/gpio_ctrl.v(218)
  AL_MUX u177 (
    .i0(int_sy_in[5]),
    .i1(int_in[5]),
    .sel(gpio_ls_sync),
    .o(n96));  // ../RTL/gpio_ctrl.v(275)
  AL_MUX u178 (
    .i0(n96),
    .i1(1'b0),
    .sel(n95),
    .o(ls_int_in[5]));  // ../RTL/gpio_ctrl.v(275)
  and u179 (ed_out[4], ed_rf[4], int_in[4]);  // ../RTL/gpio_ctrl.v(218)
  not u18 (n17, presetn);  // ../RTL/gpio_ctrl.v(144)
  and u180 (ed_out[3], ed_rf[3], int_in[3]);  // ../RTL/gpio_ctrl.v(218)
  or u181 (n97, gpio_swporta_ddr[6], gpio_swporta_ctl_internal[6]);  // ../RTL/gpio_ctrl.v(269)
  and u182 (ed_out[2], ed_rf[2], int_in[2]);  // ../RTL/gpio_ctrl.v(218)
  AL_MUX u183 (
    .i0(int_sy_in[6]),
    .i1(int_in[6]),
    .sel(gpio_ls_sync),
    .o(n98));  // ../RTL/gpio_ctrl.v(275)
  AL_MUX u184 (
    .i0(n98),
    .i1(1'b0),
    .sel(n97),
    .o(ls_int_in[6]));  // ../RTL/gpio_ctrl.v(275)
  and u185 (ed_out[1], ed_rf[1], int_in[1]);  // ../RTL/gpio_ctrl.v(218)
  buf u186 (gpio_raw_intstatus[7], int_gpio_raw_intstatus[7]);  // ../RTL/gpio_ctrl.v(305)
  or u187 (n99, gpio_swporta_ddr[7], gpio_swporta_ctl_internal[7]);  // ../RTL/gpio_ctrl.v(269)
  buf u188 (gpio_raw_intstatus[6], int_gpio_raw_intstatus[6]);  // ../RTL/gpio_ctrl.v(305)
  AL_MUX u189 (
    .i0(int_sy_in[7]),
    .i1(int_in[7]),
    .sel(gpio_ls_sync),
    .o(n100));  // ../RTL/gpio_ctrl.v(275)
  buf u19 (gpio_intr[7], gpio_intr_int[7]);  // ../RTL/gpio_ctrl.v(307)
  AL_MUX u190 (
    .i0(n100),
    .i1(1'b0),
    .sel(n99),
    .o(ls_int_in[7]));  // ../RTL/gpio_ctrl.v(275)
  buf u191 (gpio_raw_intstatus[5], int_gpio_raw_intstatus[5]);  // ../RTL/gpio_ctrl.v(305)
  buf u192 (gpio_porta_dr[4], gpio_swporta_dr[4]);  // ../RTL/gpio_ctrl.v(316)
  buf u193 (gpio_raw_intstatus[4], int_gpio_raw_intstatus[4]);  // ../RTL/gpio_ctrl.v(305)
  AL_MUX u194 (
    .i0(ls_int_in[0]),
    .i1(gpio_intr_ed_pm[0]),
    .sel(gpio_inttype_level[0]),
    .o(n102));  // ../RTL/gpio_ctrl.v(300)
  AL_MUX u195 (
    .i0(1'b0),
    .i1(n102),
    .sel(gpio_inten[0]),
    .o(int_gpio_raw_intstatus[0]));  // ../RTL/gpio_ctrl.v(300)
  buf u196 (gpio_porta_dr[3], gpio_swporta_dr[3]);  // ../RTL/gpio_ctrl.v(316)
  buf u197 (gpio_raw_intstatus[3], int_gpio_raw_intstatus[3]);  // ../RTL/gpio_ctrl.v(305)
  AL_MUX u198 (
    .i0(ls_int_in[1]),
    .i1(gpio_intr_ed_pm[1]),
    .sel(gpio_inttype_level[1]),
    .o(n104));  // ../RTL/gpio_ctrl.v(300)
  AL_MUX u199 (
    .i0(1'b0),
    .i1(n104),
    .sel(gpio_inten[1]),
    .o(int_gpio_raw_intstatus[1]));  // ../RTL/gpio_ctrl.v(300)
  AL_MUX u2 (
    .i0(gpio_ls_sync),
    .i1(1'b1),
    .sel(gpio_inttype_level[0]),
    .o(n0));  // ../RTL/gpio_ctrl.v(133)
  not u20 (n9, gpio_ext_porta[0]);  // ../RTL/gpio_ctrl.v(163)
  buf u200 (gpio_porta_dr[2], gpio_swporta_dr[2]);  // ../RTL/gpio_ctrl.v(316)
  buf u201 (gpio_raw_intstatus[2], int_gpio_raw_intstatus[2]);  // ../RTL/gpio_ctrl.v(305)
  AL_MUX u202 (
    .i0(ls_int_in[2]),
    .i1(gpio_intr_ed_pm[2]),
    .sel(gpio_inttype_level[2]),
    .o(n106));  // ../RTL/gpio_ctrl.v(300)
  AL_MUX u203 (
    .i0(1'b0),
    .i1(n106),
    .sel(gpio_inten[2]),
    .o(int_gpio_raw_intstatus[2]));  // ../RTL/gpio_ctrl.v(300)
  buf u204 (gpio_porta_dr[1], gpio_swporta_dr[1]);  // ../RTL/gpio_ctrl.v(316)
  buf u205 (gpio_raw_intstatus[1], int_gpio_raw_intstatus[1]);  // ../RTL/gpio_ctrl.v(305)
  AL_MUX u206 (
    .i0(ls_int_in[3]),
    .i1(gpio_intr_ed_pm[3]),
    .sel(gpio_inttype_level[3]),
    .o(n108));  // ../RTL/gpio_ctrl.v(300)
  AL_MUX u207 (
    .i0(1'b0),
    .i1(n108),
    .sel(gpio_inten[3]),
    .o(int_gpio_raw_intstatus[3]));  // ../RTL/gpio_ctrl.v(300)
  buf u208 (gpio_porta_ddr[7], gpio_swporta_ddr[7]);  // ../RTL/gpio_ctrl.v(324)
  not u209 (n117[7], gpio_intmask[7]);  // ../RTL/gpio_ctrl.v(306)
  AL_MUX u21 (
    .i0(n9),
    .i1(gpio_ext_porta[0]),
    .sel(gpio_int_polarity[0]),
    .o(gpio_ext_porta_int[0]));  // ../RTL/gpio_ctrl.v(165)
  AL_MUX u210 (
    .i0(ls_int_in[4]),
    .i1(gpio_intr_ed_pm[4]),
    .sel(gpio_inttype_level[4]),
    .o(n110));  // ../RTL/gpio_ctrl.v(300)
  AL_MUX u211 (
    .i0(1'b0),
    .i1(n110),
    .sel(gpio_inten[4]),
    .o(int_gpio_raw_intstatus[4]));  // ../RTL/gpio_ctrl.v(300)
  buf u212 (gpio_porta_ddr[6], gpio_swporta_ddr[6]);  // ../RTL/gpio_ctrl.v(324)
  not u213 (n117[6], gpio_intmask[6]);  // ../RTL/gpio_ctrl.v(306)
  AL_MUX u214 (
    .i0(ls_int_in[5]),
    .i1(gpio_intr_ed_pm[5]),
    .sel(gpio_inttype_level[5]),
    .o(n112));  // ../RTL/gpio_ctrl.v(300)
  AL_MUX u215 (
    .i0(1'b0),
    .i1(n112),
    .sel(gpio_inten[5]),
    .o(int_gpio_raw_intstatus[5]));  // ../RTL/gpio_ctrl.v(300)
  buf u216 (gpio_porta_ddr[5], gpio_swporta_ddr[5]);  // ../RTL/gpio_ctrl.v(324)
  not u217 (n117[5], gpio_intmask[5]);  // ../RTL/gpio_ctrl.v(306)
  AL_MUX u218 (
    .i0(ls_int_in[6]),
    .i1(gpio_intr_ed_pm[6]),
    .sel(gpio_inttype_level[6]),
    .o(n114));  // ../RTL/gpio_ctrl.v(300)
  AL_MUX u219 (
    .i0(1'b0),
    .i1(n114),
    .sel(gpio_inten[6]),
    .o(int_gpio_raw_intstatus[6]));  // ../RTL/gpio_ctrl.v(300)
  buf u22 (gpio_intr[6], gpio_intr_int[6]);  // ../RTL/gpio_ctrl.v(307)
  buf u220 (gpio_porta_ddr[4], gpio_swporta_ddr[4]);  // ../RTL/gpio_ctrl.v(324)
  not u221 (n117[4], gpio_intmask[4]);  // ../RTL/gpio_ctrl.v(306)
  AL_MUX u222 (
    .i0(ls_int_in[7]),
    .i1(gpio_intr_ed_pm[7]),
    .sel(gpio_inttype_level[7]),
    .o(n116));  // ../RTL/gpio_ctrl.v(300)
  AL_MUX u223 (
    .i0(1'b0),
    .i1(n116),
    .sel(gpio_inten[7]),
    .o(int_gpio_raw_intstatus[7]));  // ../RTL/gpio_ctrl.v(300)
  not u224 (n117[3], gpio_intmask[3]);  // ../RTL/gpio_ctrl.v(306)
  and u225 (ed_out[0], ed_rf[0], int_in[0]);  // ../RTL/gpio_ctrl.v(218)
  buf u226 (gpio_raw_intstatus[0], int_gpio_raw_intstatus[0]);  // ../RTL/gpio_ctrl.v(305)
  not u227 (n117[0], gpio_intmask[0]);  // ../RTL/gpio_ctrl.v(306)
  and u228 (gpio_intr_int[0], gpio_raw_intstatus[0], n117[0]);  // ../RTL/gpio_ctrl.v(306)
  buf u229 (gpio_intr[0], gpio_intr_int[0]);  // ../RTL/gpio_ctrl.v(307)
  not u23 (n10, gpio_ext_porta[1]);  // ../RTL/gpio_ctrl.v(163)
  or u230 (n20, gpio_intr_int[0], gpio_intr_int[1]);  // ../RTL/gpio_ctrl.v(309)
  buf u231 (gpio_porta_dr[0], gpio_swporta_dr[0]);  // ../RTL/gpio_ctrl.v(316)
  not u232 (n117[2], gpio_intmask[2]);  // ../RTL/gpio_ctrl.v(306)
  AL_MUX u233 (
    .i0(gpio_ext_porta[0]),
    .i1(gpio_swporta_dr[0]),
    .sel(gpio_porta_ddr[0]),
    .o(gpio_ext_porta_rb[0]));  // ../RTL/gpio_ctrl.v(340)
  not u234 (n117[1], gpio_intmask[1]);  // ../RTL/gpio_ctrl.v(306)
  AL_MUX u235 (
    .i0(gpio_ext_porta[1]),
    .i1(gpio_swporta_dr[1]),
    .sel(gpio_porta_ddr[1]),
    .o(gpio_ext_porta_rb[1]));  // ../RTL/gpio_ctrl.v(340)
  and u236 (gpio_intr_int[7], gpio_raw_intstatus[7], n117[7]);  // ../RTL/gpio_ctrl.v(306)
  AL_MUX u237 (
    .i0(gpio_ext_porta[2]),
    .i1(gpio_swporta_dr[2]),
    .sel(gpio_porta_ddr[2]),
    .o(gpio_ext_porta_rb[2]));  // ../RTL/gpio_ctrl.v(340)
  and u238 (gpio_intr_int[6], gpio_raw_intstatus[6], n117[6]);  // ../RTL/gpio_ctrl.v(306)
  AL_MUX u239 (
    .i0(gpio_ext_porta[3]),
    .i1(gpio_swporta_dr[3]),
    .sel(gpio_porta_ddr[3]),
    .o(gpio_ext_porta_rb[3]));  // ../RTL/gpio_ctrl.v(340)
  AL_MUX u24 (
    .i0(n10),
    .i1(gpio_ext_porta[1]),
    .sel(gpio_int_polarity[1]),
    .o(gpio_ext_porta_int[1]));  // ../RTL/gpio_ctrl.v(165)
  and u240 (gpio_intr_int[5], gpio_raw_intstatus[5], n117[5]);  // ../RTL/gpio_ctrl.v(306)
  AL_MUX u241 (
    .i0(gpio_ext_porta[4]),
    .i1(gpio_swporta_dr[4]),
    .sel(gpio_porta_ddr[4]),
    .o(gpio_ext_porta_rb[4]));  // ../RTL/gpio_ctrl.v(340)
  and u242 (gpio_intr_int[4], gpio_raw_intstatus[4], n117[4]);  // ../RTL/gpio_ctrl.v(306)
  AL_MUX u243 (
    .i0(gpio_ext_porta[5]),
    .i1(gpio_swporta_dr[5]),
    .sel(gpio_porta_ddr[5]),
    .o(gpio_ext_porta_rb[5]));  // ../RTL/gpio_ctrl.v(340)
  and u244 (gpio_intr_int[3], gpio_raw_intstatus[3], n117[3]);  // ../RTL/gpio_ctrl.v(306)
  AL_MUX u245 (
    .i0(gpio_ext_porta[6]),
    .i1(gpio_swporta_dr[6]),
    .sel(gpio_porta_ddr[6]),
    .o(gpio_ext_porta_rb[6]));  // ../RTL/gpio_ctrl.v(340)
  and u246 (gpio_intr_int[2], gpio_raw_intstatus[2], n117[2]);  // ../RTL/gpio_ctrl.v(306)
  AL_MUX u247 (
    .i0(gpio_ext_porta[7]),
    .i1(gpio_swporta_dr[7]),
    .sel(gpio_porta_ddr[7]),
    .o(gpio_ext_porta_rb[7]));  // ../RTL/gpio_ctrl.v(340)
  and u248 (gpio_intr_int[1], gpio_raw_intstatus[1], n117[1]);  // ../RTL/gpio_ctrl.v(306)
  buf u25 (gpio_intr[5], gpio_intr_int[5]);  // ../RTL/gpio_ctrl.v(307)
  not u26 (n11, gpio_ext_porta[2]);  // ../RTL/gpio_ctrl.v(163)
  AL_MUX u27 (
    .i0(n11),
    .i1(gpio_ext_porta[2]),
    .sel(gpio_int_polarity[2]),
    .o(gpio_ext_porta_int[2]));  // ../RTL/gpio_ctrl.v(165)
  buf u28 (gpio_intr[4], gpio_intr_int[4]);  // ../RTL/gpio_ctrl.v(307)
  not u29 (n12, gpio_ext_porta[3]);  // ../RTL/gpio_ctrl.v(163)
  AL_MUX u3 (
    .i0(1'b0),
    .i1(n0),
    .sel(gpio_inten[0]),
    .o(intrclk_en[0]));  // ../RTL/gpio_ctrl.v(135)
  AL_MUX u30 (
    .i0(n12),
    .i1(gpio_ext_porta[3]),
    .sel(gpio_int_polarity[3]),
    .o(gpio_ext_porta_int[3]));  // ../RTL/gpio_ctrl.v(165)
  buf u31 (gpio_intr[3], gpio_intr_int[3]);  // ../RTL/gpio_ctrl.v(307)
  not u32 (n13, gpio_ext_porta[4]);  // ../RTL/gpio_ctrl.v(163)
  AL_MUX u33 (
    .i0(n13),
    .i1(gpio_ext_porta[4]),
    .sel(gpio_int_polarity[4]),
    .o(gpio_ext_porta_int[4]));  // ../RTL/gpio_ctrl.v(165)
  buf u34 (gpio_intr[2], gpio_intr_int[2]);  // ../RTL/gpio_ctrl.v(307)
  not u35 (n14, gpio_ext_porta[5]);  // ../RTL/gpio_ctrl.v(163)
  AL_MUX u36 (
    .i0(n14),
    .i1(gpio_ext_porta[5]),
    .sel(gpio_int_polarity[5]),
    .o(gpio_ext_porta_int[5]));  // ../RTL/gpio_ctrl.v(165)
  buf u37 (gpio_intr[1], gpio_intr_int[1]);  // ../RTL/gpio_ctrl.v(307)
  not u38 (n15, gpio_ext_porta[6]);  // ../RTL/gpio_ctrl.v(163)
  AL_MUX u39 (
    .i0(n15),
    .i1(gpio_ext_porta[6]),
    .sel(gpio_int_polarity[6]),
    .o(gpio_ext_porta_int[6]));  // ../RTL/gpio_ctrl.v(165)
  AL_MUX u4 (
    .i0(gpio_ls_sync),
    .i1(1'b1),
    .sel(gpio_inttype_level[1]),
    .o(n1));  // ../RTL/gpio_ctrl.v(133)
  or u40 (gpio_intr_flag_int, n18, n113);  // ../RTL/gpio_ctrl.v(309)
  not u41 (n16, gpio_ext_porta[7]);  // ../RTL/gpio_ctrl.v(163)
  AL_MUX u42 (
    .i0(n16),
    .i1(gpio_ext_porta[7]),
    .sel(gpio_int_polarity[7]),
    .o(gpio_ext_porta_int[7]));  // ../RTL/gpio_ctrl.v(165)
  or u43 (n111, intrclk_en[0], intrclk_en[1]);  // ../RTL/gpio_ctrl.v(140)
  buf u44 (gpio_porta_ddr[3], gpio_swporta_ddr[3]);  // ../RTL/gpio_ctrl.v(324)
  buf u45 (gpio_porta_ddr[2], gpio_swporta_ddr[2]);  // ../RTL/gpio_ctrl.v(324)
  buf u46 (int_sy_in[0], gpio_ext_porta_int[0]);  // ../RTL/gpio_ctrl.v(176)
  buf u47 (gpio_porta_ddr[1], gpio_swporta_ddr[1]);  // ../RTL/gpio_ctrl.v(324)
  buf u48 (int_in[0], int_pre_in[0]);  // ../RTL/gpio_ctrl.v(195)
  xor u49 (ed_rf[0], int_in[0], ed_int_d1[0]);  // ../RTL/gpio_ctrl.v(206)
  AL_MUX u5 (
    .i0(1'b0),
    .i1(n1),
    .sel(gpio_inten[1]),
    .o(intrclk_en[1]));  // ../RTL/gpio_ctrl.v(135)
  buf u50 (gpio_porta_ddr[0], gpio_swporta_ddr[0]);  // ../RTL/gpio_ctrl.v(324)
  or u51 (n113, n8, n115);  // ../RTL/gpio_ctrl.v(309)
  and u52 (n21, ed_out[0], gpio_inten[0]);  // ../RTL/gpio_ctrl.v(241)
  not u53 (n22, gpio_swporta_ddr[0]);  // ../RTL/gpio_ctrl.v(242)
  and u54 (n23, n21, n22);  // ../RTL/gpio_ctrl.v(242)
  not u55 (n24, gpio_swporta_ctl_internal[0]);  // ../RTL/gpio_ctrl.v(243)
  and u56 (n25, n23, n24);  // ../RTL/gpio_ctrl.v(243)
  AL_MUX u57 (
    .i0(gpio_intr_ed_pm[0]),
    .i1(1'b0),
    .sel(gpio_porta_eoi[0]),
    .o(n26));  // ../RTL/gpio_ctrl.v(247)
  AL_MUX u58 (
    .i0(n26),
    .i1(1'b1),
    .sel(n25),
    .o(n27));  // ../RTL/gpio_ctrl.v(247)
  AL_MUX u59 (
    .i0(1'b0),
    .i1(n27),
    .sel(gpio_inten[0]),
    .o(n28));  // ../RTL/gpio_ctrl.v(247)
  AL_MUX u6 (
    .i0(gpio_ls_sync),
    .i1(1'b1),
    .sel(gpio_inttype_level[2]),
    .o(n2));  // ../RTL/gpio_ctrl.v(133)
  or u60 (n115, gpio_intr_int[6], gpio_intr_int[7]);  // ../RTL/gpio_ctrl.v(309)
  and u61 (n29, ed_out[1], gpio_inten[1]);  // ../RTL/gpio_ctrl.v(241)
  not u62 (n30, gpio_swporta_ddr[1]);  // ../RTL/gpio_ctrl.v(242)
  and u63 (n31, n29, n30);  // ../RTL/gpio_ctrl.v(242)
  not u64 (n32, gpio_swporta_ctl_internal[1]);  // ../RTL/gpio_ctrl.v(243)
  and u65 (n33, n31, n32);  // ../RTL/gpio_ctrl.v(243)
  or u66 (gpio_intrclk_en_int, n107, n101);  // ../RTL/gpio_ctrl.v(140)
  AL_MUX u67 (
    .i0(gpio_intr_ed_pm[1]),
    .i1(1'b0),
    .sel(gpio_porta_eoi[1]),
    .o(n34));  // ../RTL/gpio_ctrl.v(247)
  AL_MUX u68 (
    .i0(n34),
    .i1(1'b1),
    .sel(n33),
    .o(n35));  // ../RTL/gpio_ctrl.v(247)
  AL_MUX u69 (
    .i0(1'b0),
    .i1(n35),
    .sel(gpio_inten[1]),
    .o(n36));  // ../RTL/gpio_ctrl.v(247)
  AL_MUX u7 (
    .i0(1'b0),
    .i1(n2),
    .sel(gpio_inten[2]),
    .o(intrclk_en[2]));  // ../RTL/gpio_ctrl.v(135)
  or u70 (n8, gpio_intr_int[4], gpio_intr_int[5]);  // ../RTL/gpio_ctrl.v(309)
  or u71 (n101, n105, n103);  // ../RTL/gpio_ctrl.v(140)
  or u72 (n103, intrclk_en[6], intrclk_en[7]);  // ../RTL/gpio_ctrl.v(140)
  and u73 (n37, ed_out[2], gpio_inten[2]);  // ../RTL/gpio_ctrl.v(241)
  not u74 (n38, gpio_swporta_ddr[2]);  // ../RTL/gpio_ctrl.v(242)
  and u75 (n39, n37, n38);  // ../RTL/gpio_ctrl.v(242)
  not u76 (n40, gpio_swporta_ctl_internal[2]);  // ../RTL/gpio_ctrl.v(243)
  and u77 (n41, n39, n40);  // ../RTL/gpio_ctrl.v(243)
  or u78 (n105, intrclk_en[4], intrclk_en[5]);  // ../RTL/gpio_ctrl.v(140)
  AL_MUX u79 (
    .i0(gpio_intr_ed_pm[2]),
    .i1(1'b0),
    .sel(gpio_porta_eoi[2]),
    .o(n42));  // ../RTL/gpio_ctrl.v(247)
  AL_MUX u8 (
    .i0(gpio_ls_sync),
    .i1(1'b1),
    .sel(gpio_inttype_level[3]),
    .o(n3));  // ../RTL/gpio_ctrl.v(133)
  AL_MUX u80 (
    .i0(n42),
    .i1(1'b1),
    .sel(n41),
    .o(n43));  // ../RTL/gpio_ctrl.v(247)
  AL_MUX u81 (
    .i0(1'b0),
    .i1(n43),
    .sel(gpio_inten[2]),
    .o(n44));  // ../RTL/gpio_ctrl.v(247)
  or u82 (n18, n20, n19);  // ../RTL/gpio_ctrl.v(309)
  or u83 (n107, n111, n109);  // ../RTL/gpio_ctrl.v(140)
  or u84 (n109, intrclk_en[2], intrclk_en[3]);  // ../RTL/gpio_ctrl.v(140)
  and u85 (n45, ed_out[3], gpio_inten[3]);  // ../RTL/gpio_ctrl.v(241)
  not u86 (n46, gpio_swporta_ddr[3]);  // ../RTL/gpio_ctrl.v(242)
  and u87 (n47, n45, n46);  // ../RTL/gpio_ctrl.v(242)
  not u88 (n48, gpio_swporta_ctl_internal[3]);  // ../RTL/gpio_ctrl.v(243)
  and u89 (n49, n47, n48);  // ../RTL/gpio_ctrl.v(243)
  AL_MUX u9 (
    .i0(1'b0),
    .i1(n3),
    .sel(gpio_inten[3]),
    .o(intrclk_en[3]));  // ../RTL/gpio_ctrl.v(135)
  buf u90 (int_sy_in[7], gpio_ext_porta_int[7]);  // ../RTL/gpio_ctrl.v(176)
  AL_MUX u91 (
    .i0(gpio_intr_ed_pm[3]),
    .i1(1'b0),
    .sel(gpio_porta_eoi[3]),
    .o(n50));  // ../RTL/gpio_ctrl.v(247)
  AL_MUX u92 (
    .i0(n50),
    .i1(1'b1),
    .sel(n49),
    .o(n51));  // ../RTL/gpio_ctrl.v(247)
  AL_MUX u93 (
    .i0(1'b0),
    .i1(n51),
    .sel(gpio_inten[3]),
    .o(n52));  // ../RTL/gpio_ctrl.v(247)
  or u94 (n19, gpio_intr_int[2], gpio_intr_int[3]);  // ../RTL/gpio_ctrl.v(309)
  buf u95 (int_sy_in[6], gpio_ext_porta_int[6]);  // ../RTL/gpio_ctrl.v(176)
  buf u96 (int_sy_in[5], gpio_ext_porta_int[5]);  // ../RTL/gpio_ctrl.v(176)
  and u97 (n53, ed_out[4], gpio_inten[4]);  // ../RTL/gpio_ctrl.v(241)
  not u98 (n54, gpio_swporta_ddr[4]);  // ../RTL/gpio_ctrl.v(242)
  and u99 (n55, n53, n54);  // ../RTL/gpio_ctrl.v(242)

endmodule 

module add_pu4_pu4_o5
  (
  i0,
  i1,
  o
  );

  input [3:0] i0;
  input [3:0] i1;
  output [4:0] o;



endmodule 

module eq_w15
  (
  i0,
  i1,
  o
  );

  input [14:0] i0;
  input [14:0] i1;
  output o;



endmodule 

module lt_u4_u4
  (
  ci,
  i0,
  i1,
  o
  );

  input ci;
  input [3:0] i0;
  input [3:0] i1;
  output o;



endmodule 

module binary_mux_s1_w7
  (
  i0,
  i1,
  sel,
  o
  );

  input [6:0] i0;
  input [6:0] i1;
  input sel;
  output [6:0] o;



endmodule 

module binary_mux_s1_w5
  (
  i0,
  i1,
  sel,
  o
  );

  input [4:0] i0;
  input [4:0] i1;
  input sel;
  output [4:0] o;



endmodule 

module binary_mux_s4_w5
  (
  i0,
  i1,
  i10,
  i11,
  i12,
  i13,
  i14,
  i15,
  i2,
  i3,
  i4,
  i5,
  i6,
  i7,
  i8,
  i9,
  sel,
  o
  );

  input [4:0] i0;
  input [4:0] i1;
  input [4:0] i10;
  input [4:0] i11;
  input [4:0] i12;
  input [4:0] i13;
  input [4:0] i14;
  input [4:0] i15;
  input [4:0] i2;
  input [4:0] i3;
  input [4:0] i4;
  input [4:0] i5;
  input [4:0] i6;
  input [4:0] i7;
  input [4:0] i8;
  input [4:0] i9;
  input [3:0] sel;
  output [4:0] o;



endmodule 

module binary_mux_s1_w20
  (
  i0,
  i1,
  sel,
  o
  );

  input [19:0] i0;
  input [19:0] i1;
  input sel;
  output [19:0] o;



endmodule 

module binary_mux_s3_w8
  (
  i0,
  i1,
  i2,
  i3,
  i4,
  i5,
  i6,
  i7,
  sel,
  o
  );

  input [7:0] i0;
  input [7:0] i1;
  input [7:0] i2;
  input [7:0] i3;
  input [7:0] i4;
  input [7:0] i5;
  input [7:0] i6;
  input [7:0] i7;
  input [2:0] sel;
  output [7:0] o;



endmodule 

module binary_mux_s4_w8
  (
  i0,
  i1,
  i10,
  i11,
  i12,
  i13,
  i14,
  i15,
  i2,
  i3,
  i4,
  i5,
  i6,
  i7,
  i8,
  i9,
  sel,
  o
  );

  input [7:0] i0;
  input [7:0] i1;
  input [7:0] i10;
  input [7:0] i11;
  input [7:0] i12;
  input [7:0] i13;
  input [7:0] i14;
  input [7:0] i15;
  input [7:0] i2;
  input [7:0] i3;
  input [7:0] i4;
  input [7:0] i5;
  input [7:0] i6;
  input [7:0] i7;
  input [7:0] i8;
  input [7:0] i9;
  input [3:0] sel;
  output [7:0] o;



endmodule 

module binary_mux_s1_w12
  (
  i0,
  i1,
  sel,
  o
  );

  input [11:0] i0;
  input [11:0] i1;
  input sel;
  output [11:0] o;



endmodule 

module reg_ar_as_w7
  (
  clk,
  d,
  en,
  reset,
  set,
  q
  );

  input clk;
  input [6:0] d;
  input en;
  input [6:0] reset;
  input [6:0] set;
  output [6:0] q;



endmodule 

module reg_ar_as_w20
  (
  clk,
  d,
  en,
  reset,
  set,
  q
  );

  input clk;
  input [19:0] d;
  input en;
  input [19:0] reset;
  input [19:0] set;
  output [19:0] q;



endmodule 

module reg_ar_as_w8
  (
  clk,
  d,
  en,
  reset,
  set,
  q
  );

  input clk;
  input [7:0] d;
  input en;
  input [7:0] reset;
  input [7:0] set;
  output [7:0] q;



endmodule 

module add_pu16_mu16_o16
  (
  i0,
  i1,
  o
  );

  input [15:0] i0;
  input [15:0] i1;
  output [15:0] o;



endmodule 

module add_pu4_mu4_o4
  (
  i0,
  i1,
  o
  );

  input [3:0] i0;
  input [3:0] i1;
  output [3:0] o;



endmodule 

module eq_w3
  (
  i0,
  i1,
  o
  );

  input [2:0] i0;
  input [2:0] i1;
  output o;



endmodule 

module binary_mux_s1_w14
  (
  i0,
  i1,
  sel,
  o
  );

  input [13:0] i0;
  input [13:0] i1;
  input sel;
  output [13:0] o;



endmodule 

module binary_mux_s3_w1
  (
  i0,
  i1,
  i2,
  i3,
  i4,
  i5,
  i6,
  i7,
  sel,
  o
  );

  input i0;
  input i1;
  input i2;
  input i3;
  input i4;
  input i5;
  input i6;
  input i7;
  input [2:0] sel;
  output o;



endmodule 

module binary_mux_s3_w3
  (
  i0,
  i1,
  i2,
  i3,
  i4,
  i5,
  i6,
  i7,
  sel,
  o
  );

  input [2:0] i0;
  input [2:0] i1;
  input [2:0] i2;
  input [2:0] i3;
  input [2:0] i4;
  input [2:0] i5;
  input [2:0] i6;
  input [2:0] i7;
  input [2:0] sel;
  output [2:0] o;



endmodule 

module reg_ar_as_w14
  (
  clk,
  d,
  en,
  reset,
  set,
  q
  );

  input clk;
  input [13:0] d;
  input en;
  input [13:0] reset;
  input [13:0] set;
  output [13:0] q;



endmodule 

module add_pu10_pu10_o10
  (
  i0,
  i1,
  o
  );

  input [9:0] i0;
  input [9:0] i1;
  output [9:0] o;



endmodule 

module add_pu31_pu31_o31
  (
  i0,
  i1,
  o
  );

  input [30:0] i0;
  input [30:0] i1;
  output [30:0] o;



endmodule 

module add_pu30_pu30_o30
  (
  i0,
  i1,
  o
  );

  input [29:0] i0;
  input [29:0] i1;
  output [29:0] o;



endmodule 

module add_pu33_pu33_o33
  (
  i0,
  i1,
  o
  );

  input [32:0] i0;
  input [32:0] i1;
  output [32:0] o;



endmodule 

module add_pu32_pu32_o33
  (
  i0,
  i1,
  o
  );

  input [31:0] i0;
  input [31:0] i1;
  output [32:0] o;



endmodule 

module eq_w32
  (
  i0,
  i1,
  o
  );

  input [31:0] i0;
  input [31:0] i1;
  output o;



endmodule 

module eq_w27
  (
  i0,
  i1,
  o
  );

  input [26:0] i0;
  input [26:0] i1;
  output o;



endmodule 

module mult_u32_u32_o64
  (
  i0,
  i1,
  o
  );

  input [31:0] i0;
  input [31:0] i1;
  output [63:0] o;



endmodule 

module binary_mux_s1_w19
  (
  i0,
  i1,
  sel,
  o
  );

  input [18:0] i0;
  input [18:0] i1;
  input sel;
  output [18:0] o;



endmodule 

module binary_mux_s1_w11
  (
  i0,
  i1,
  sel,
  o
  );

  input [10:0] i0;
  input [10:0] i1;
  input sel;
  output [10:0] o;



endmodule 

module add_pu24_mu24_o24
  (
  i0,
  i1,
  o
  );

  input [23:0] i0;
  input [23:0] i1;
  output [23:0] o;



endmodule 

module add_pu9_mu9_o9
  (
  i0,
  i1,
  o
  );

  input [8:0] i0;
  input [8:0] i1;
  output [8:0] o;



endmodule 

module eq_w5
  (
  i0,
  i1,
  o
  );

  input [4:0] i0;
  input [4:0] i1;
  output o;



endmodule 

module onehot_mux_s12_w32
  (
  i0,
  i1,
  i10,
  i11,
  i2,
  i3,
  i4,
  i5,
  i6,
  i7,
  i8,
  i9,
  sel,
  o
  );

  input [31:0] i0;
  input [31:0] i1;
  input [31:0] i10;
  input [31:0] i11;
  input [31:0] i2;
  input [31:0] i3;
  input [31:0] i4;
  input [31:0] i5;
  input [31:0] i6;
  input [31:0] i7;
  input [31:0] i8;
  input [31:0] i9;
  input [11:0] sel;
  output [31:0] o;



endmodule 

module AL_MUX
  (
  input i0,
  input i1,
  input sel,
  output o
  );

  wire not_sel, sel_i0, sel_i1;
  not u0 (not_sel, sel);
  and u1 (sel_i1, sel, i1);
  and u2 (sel_i0, not_sel, i0);
  or u3 (o, sel_i1, sel_i0);

endmodule

module AL_DFF
  (
  input reset,
  input set,
  input clk,
  input d,
  output reg q
  );

  parameter INI = 1'b0;

  always @(posedge reset or posedge set or posedge clk)
  begin
    if (reset)
      q <= 1'b0;
    else if (set)
      q <= 1'b1;
    else
      q <= d;
  end

endmodule

