// Verilog netlist created by TD v4.6.12906
// Mon Jul 29 11:09:07 2019

`timescale 1ns / 1ps
module img_cache  // al_ip/ip_ram.v(14)
  (
  addra,
  addrb,
  cea,
  ceb,
  clka,
  clkb,
  dia,
  rstb,
  dob
  );

  input [15:0] addra;  // al_ip/ip_ram.v(23)
  input [15:0] addrb;  // al_ip/ip_ram.v(24)
  input cea;  // al_ip/ip_ram.v(25)
  input ceb;  // al_ip/ip_ram.v(26)
  input clka;  // al_ip/ip_ram.v(27)
  input clkb;  // al_ip/ip_ram.v(28)
  input [15:0] dia;  // al_ip/ip_ram.v(22)
  input rstb;  // al_ip/ip_ram.v(29)
  output [15:0] dob;  // al_ip/ip_ram.v(19)

  wire [0:6] addrb_piped;
  wire [0:6] addrb_piped_piped;
  wire  \inst_dob_mux_b0/B0_0 ;
  wire  \inst_dob_mux_b0/B0_1 ;
  wire  \inst_dob_mux_b0/B0_10 ;
  wire  \inst_dob_mux_b0/B0_11 ;
  wire  \inst_dob_mux_b0/B0_12 ;
  wire  \inst_dob_mux_b0/B0_13 ;
  wire  \inst_dob_mux_b0/B0_14 ;
  wire  \inst_dob_mux_b0/B0_15 ;
  wire  \inst_dob_mux_b0/B0_16 ;
  wire  \inst_dob_mux_b0/B0_17 ;
  wire  \inst_dob_mux_b0/B0_18 ;
  wire  \inst_dob_mux_b0/B0_19 ;
  wire  \inst_dob_mux_b0/B0_2 ;
  wire  \inst_dob_mux_b0/B0_20 ;
  wire  \inst_dob_mux_b0/B0_21 ;
  wire  \inst_dob_mux_b0/B0_22 ;
  wire  \inst_dob_mux_b0/B0_23 ;
  wire  \inst_dob_mux_b0/B0_24 ;
  wire  \inst_dob_mux_b0/B0_25 ;
  wire  \inst_dob_mux_b0/B0_26 ;
  wire  \inst_dob_mux_b0/B0_27 ;
  wire  \inst_dob_mux_b0/B0_28 ;
  wire  \inst_dob_mux_b0/B0_29 ;
  wire  \inst_dob_mux_b0/B0_3 ;
  wire  \inst_dob_mux_b0/B0_30 ;
  wire  \inst_dob_mux_b0/B0_31 ;
  wire  \inst_dob_mux_b0/B0_32 ;
  wire  \inst_dob_mux_b0/B0_33 ;
  wire  \inst_dob_mux_b0/B0_34 ;
  wire  \inst_dob_mux_b0/B0_35 ;
  wire  \inst_dob_mux_b0/B0_36 ;
  wire  \inst_dob_mux_b0/B0_37 ;
  wire  \inst_dob_mux_b0/B0_38 ;
  wire  \inst_dob_mux_b0/B0_39 ;
  wire  \inst_dob_mux_b0/B0_4 ;
  wire  \inst_dob_mux_b0/B0_40 ;
  wire  \inst_dob_mux_b0/B0_41 ;
  wire  \inst_dob_mux_b0/B0_42 ;
  wire  \inst_dob_mux_b0/B0_43 ;
  wire  \inst_dob_mux_b0/B0_44 ;
  wire  \inst_dob_mux_b0/B0_45 ;
  wire  \inst_dob_mux_b0/B0_46 ;
  wire  \inst_dob_mux_b0/B0_47 ;
  wire  \inst_dob_mux_b0/B0_48 ;
  wire  \inst_dob_mux_b0/B0_49 ;
  wire  \inst_dob_mux_b0/B0_5 ;
  wire  \inst_dob_mux_b0/B0_50 ;
  wire  \inst_dob_mux_b0/B0_51 ;
  wire  \inst_dob_mux_b0/B0_52 ;
  wire  \inst_dob_mux_b0/B0_53 ;
  wire  \inst_dob_mux_b0/B0_54 ;
  wire  \inst_dob_mux_b0/B0_55 ;
  wire  \inst_dob_mux_b0/B0_56 ;
  wire  \inst_dob_mux_b0/B0_57 ;
  wire  \inst_dob_mux_b0/B0_58 ;
  wire  \inst_dob_mux_b0/B0_59 ;
  wire  \inst_dob_mux_b0/B0_6 ;
  wire  \inst_dob_mux_b0/B0_60 ;
  wire  \inst_dob_mux_b0/B0_61 ;
  wire  \inst_dob_mux_b0/B0_62 ;
  wire  \inst_dob_mux_b0/B0_63 ;
  wire  \inst_dob_mux_b0/B0_7 ;
  wire  \inst_dob_mux_b0/B0_8 ;
  wire  \inst_dob_mux_b0/B0_9 ;
  wire  \inst_dob_mux_b0/B1_0 ;
  wire  \inst_dob_mux_b0/B1_1 ;
  wire  \inst_dob_mux_b0/B1_10 ;
  wire  \inst_dob_mux_b0/B1_11 ;
  wire  \inst_dob_mux_b0/B1_12 ;
  wire  \inst_dob_mux_b0/B1_13 ;
  wire  \inst_dob_mux_b0/B1_14 ;
  wire  \inst_dob_mux_b0/B1_15 ;
  wire  \inst_dob_mux_b0/B1_16 ;
  wire  \inst_dob_mux_b0/B1_17 ;
  wire  \inst_dob_mux_b0/B1_18 ;
  wire  \inst_dob_mux_b0/B1_19 ;
  wire  \inst_dob_mux_b0/B1_2 ;
  wire  \inst_dob_mux_b0/B1_20 ;
  wire  \inst_dob_mux_b0/B1_21 ;
  wire  \inst_dob_mux_b0/B1_22 ;
  wire  \inst_dob_mux_b0/B1_23 ;
  wire  \inst_dob_mux_b0/B1_24 ;
  wire  \inst_dob_mux_b0/B1_25 ;
  wire  \inst_dob_mux_b0/B1_26 ;
  wire  \inst_dob_mux_b0/B1_27 ;
  wire  \inst_dob_mux_b0/B1_28 ;
  wire  \inst_dob_mux_b0/B1_29 ;
  wire  \inst_dob_mux_b0/B1_3 ;
  wire  \inst_dob_mux_b0/B1_30 ;
  wire  \inst_dob_mux_b0/B1_31 ;
  wire  \inst_dob_mux_b0/B1_4 ;
  wire  \inst_dob_mux_b0/B1_5 ;
  wire  \inst_dob_mux_b0/B1_6 ;
  wire  \inst_dob_mux_b0/B1_7 ;
  wire  \inst_dob_mux_b0/B1_8 ;
  wire  \inst_dob_mux_b0/B1_9 ;
  wire  \inst_dob_mux_b0/B2_0 ;
  wire  \inst_dob_mux_b0/B2_1 ;
  wire  \inst_dob_mux_b0/B2_10 ;
  wire  \inst_dob_mux_b0/B2_11 ;
  wire  \inst_dob_mux_b0/B2_12 ;
  wire  \inst_dob_mux_b0/B2_13 ;
  wire  \inst_dob_mux_b0/B2_14 ;
  wire  \inst_dob_mux_b0/B2_15 ;
  wire  \inst_dob_mux_b0/B2_2 ;
  wire  \inst_dob_mux_b0/B2_3 ;
  wire  \inst_dob_mux_b0/B2_4 ;
  wire  \inst_dob_mux_b0/B2_5 ;
  wire  \inst_dob_mux_b0/B2_6 ;
  wire  \inst_dob_mux_b0/B2_7 ;
  wire  \inst_dob_mux_b0/B2_8 ;
  wire  \inst_dob_mux_b0/B2_9 ;
  wire  \inst_dob_mux_b0/B3_0 ;
  wire  \inst_dob_mux_b0/B3_1 ;
  wire  \inst_dob_mux_b0/B3_2 ;
  wire  \inst_dob_mux_b0/B3_3 ;
  wire  \inst_dob_mux_b0/B3_4 ;
  wire  \inst_dob_mux_b0/B3_5 ;
  wire  \inst_dob_mux_b0/B3_6 ;
  wire  \inst_dob_mux_b0/B3_7 ;
  wire  \inst_dob_mux_b0/B4_0 ;
  wire  \inst_dob_mux_b0/B4_1 ;
  wire  \inst_dob_mux_b0/B4_2 ;
  wire  \inst_dob_mux_b0/B4_3 ;
  wire  \inst_dob_mux_b0/B5_0 ;
  wire  \inst_dob_mux_b0/B5_1 ;
  wire  \inst_dob_mux_b1/B0_0 ;
  wire  \inst_dob_mux_b1/B0_1 ;
  wire  \inst_dob_mux_b1/B0_10 ;
  wire  \inst_dob_mux_b1/B0_11 ;
  wire  \inst_dob_mux_b1/B0_12 ;
  wire  \inst_dob_mux_b1/B0_13 ;
  wire  \inst_dob_mux_b1/B0_14 ;
  wire  \inst_dob_mux_b1/B0_15 ;
  wire  \inst_dob_mux_b1/B0_16 ;
  wire  \inst_dob_mux_b1/B0_17 ;
  wire  \inst_dob_mux_b1/B0_18 ;
  wire  \inst_dob_mux_b1/B0_19 ;
  wire  \inst_dob_mux_b1/B0_2 ;
  wire  \inst_dob_mux_b1/B0_20 ;
  wire  \inst_dob_mux_b1/B0_21 ;
  wire  \inst_dob_mux_b1/B0_22 ;
  wire  \inst_dob_mux_b1/B0_23 ;
  wire  \inst_dob_mux_b1/B0_24 ;
  wire  \inst_dob_mux_b1/B0_25 ;
  wire  \inst_dob_mux_b1/B0_26 ;
  wire  \inst_dob_mux_b1/B0_27 ;
  wire  \inst_dob_mux_b1/B0_28 ;
  wire  \inst_dob_mux_b1/B0_29 ;
  wire  \inst_dob_mux_b1/B0_3 ;
  wire  \inst_dob_mux_b1/B0_30 ;
  wire  \inst_dob_mux_b1/B0_31 ;
  wire  \inst_dob_mux_b1/B0_32 ;
  wire  \inst_dob_mux_b1/B0_33 ;
  wire  \inst_dob_mux_b1/B0_34 ;
  wire  \inst_dob_mux_b1/B0_35 ;
  wire  \inst_dob_mux_b1/B0_36 ;
  wire  \inst_dob_mux_b1/B0_37 ;
  wire  \inst_dob_mux_b1/B0_38 ;
  wire  \inst_dob_mux_b1/B0_39 ;
  wire  \inst_dob_mux_b1/B0_4 ;
  wire  \inst_dob_mux_b1/B0_40 ;
  wire  \inst_dob_mux_b1/B0_41 ;
  wire  \inst_dob_mux_b1/B0_42 ;
  wire  \inst_dob_mux_b1/B0_43 ;
  wire  \inst_dob_mux_b1/B0_44 ;
  wire  \inst_dob_mux_b1/B0_45 ;
  wire  \inst_dob_mux_b1/B0_46 ;
  wire  \inst_dob_mux_b1/B0_47 ;
  wire  \inst_dob_mux_b1/B0_48 ;
  wire  \inst_dob_mux_b1/B0_49 ;
  wire  \inst_dob_mux_b1/B0_5 ;
  wire  \inst_dob_mux_b1/B0_50 ;
  wire  \inst_dob_mux_b1/B0_51 ;
  wire  \inst_dob_mux_b1/B0_52 ;
  wire  \inst_dob_mux_b1/B0_53 ;
  wire  \inst_dob_mux_b1/B0_54 ;
  wire  \inst_dob_mux_b1/B0_55 ;
  wire  \inst_dob_mux_b1/B0_56 ;
  wire  \inst_dob_mux_b1/B0_57 ;
  wire  \inst_dob_mux_b1/B0_58 ;
  wire  \inst_dob_mux_b1/B0_59 ;
  wire  \inst_dob_mux_b1/B0_6 ;
  wire  \inst_dob_mux_b1/B0_60 ;
  wire  \inst_dob_mux_b1/B0_61 ;
  wire  \inst_dob_mux_b1/B0_62 ;
  wire  \inst_dob_mux_b1/B0_63 ;
  wire  \inst_dob_mux_b1/B0_7 ;
  wire  \inst_dob_mux_b1/B0_8 ;
  wire  \inst_dob_mux_b1/B0_9 ;
  wire  \inst_dob_mux_b1/B1_0 ;
  wire  \inst_dob_mux_b1/B1_1 ;
  wire  \inst_dob_mux_b1/B1_10 ;
  wire  \inst_dob_mux_b1/B1_11 ;
  wire  \inst_dob_mux_b1/B1_12 ;
  wire  \inst_dob_mux_b1/B1_13 ;
  wire  \inst_dob_mux_b1/B1_14 ;
  wire  \inst_dob_mux_b1/B1_15 ;
  wire  \inst_dob_mux_b1/B1_16 ;
  wire  \inst_dob_mux_b1/B1_17 ;
  wire  \inst_dob_mux_b1/B1_18 ;
  wire  \inst_dob_mux_b1/B1_19 ;
  wire  \inst_dob_mux_b1/B1_2 ;
  wire  \inst_dob_mux_b1/B1_20 ;
  wire  \inst_dob_mux_b1/B1_21 ;
  wire  \inst_dob_mux_b1/B1_22 ;
  wire  \inst_dob_mux_b1/B1_23 ;
  wire  \inst_dob_mux_b1/B1_24 ;
  wire  \inst_dob_mux_b1/B1_25 ;
  wire  \inst_dob_mux_b1/B1_26 ;
  wire  \inst_dob_mux_b1/B1_27 ;
  wire  \inst_dob_mux_b1/B1_28 ;
  wire  \inst_dob_mux_b1/B1_29 ;
  wire  \inst_dob_mux_b1/B1_3 ;
  wire  \inst_dob_mux_b1/B1_30 ;
  wire  \inst_dob_mux_b1/B1_31 ;
  wire  \inst_dob_mux_b1/B1_4 ;
  wire  \inst_dob_mux_b1/B1_5 ;
  wire  \inst_dob_mux_b1/B1_6 ;
  wire  \inst_dob_mux_b1/B1_7 ;
  wire  \inst_dob_mux_b1/B1_8 ;
  wire  \inst_dob_mux_b1/B1_9 ;
  wire  \inst_dob_mux_b1/B2_0 ;
  wire  \inst_dob_mux_b1/B2_1 ;
  wire  \inst_dob_mux_b1/B2_10 ;
  wire  \inst_dob_mux_b1/B2_11 ;
  wire  \inst_dob_mux_b1/B2_12 ;
  wire  \inst_dob_mux_b1/B2_13 ;
  wire  \inst_dob_mux_b1/B2_14 ;
  wire  \inst_dob_mux_b1/B2_15 ;
  wire  \inst_dob_mux_b1/B2_2 ;
  wire  \inst_dob_mux_b1/B2_3 ;
  wire  \inst_dob_mux_b1/B2_4 ;
  wire  \inst_dob_mux_b1/B2_5 ;
  wire  \inst_dob_mux_b1/B2_6 ;
  wire  \inst_dob_mux_b1/B2_7 ;
  wire  \inst_dob_mux_b1/B2_8 ;
  wire  \inst_dob_mux_b1/B2_9 ;
  wire  \inst_dob_mux_b1/B3_0 ;
  wire  \inst_dob_mux_b1/B3_1 ;
  wire  \inst_dob_mux_b1/B3_2 ;
  wire  \inst_dob_mux_b1/B3_3 ;
  wire  \inst_dob_mux_b1/B3_4 ;
  wire  \inst_dob_mux_b1/B3_5 ;
  wire  \inst_dob_mux_b1/B3_6 ;
  wire  \inst_dob_mux_b1/B3_7 ;
  wire  \inst_dob_mux_b1/B4_0 ;
  wire  \inst_dob_mux_b1/B4_1 ;
  wire  \inst_dob_mux_b1/B4_2 ;
  wire  \inst_dob_mux_b1/B4_3 ;
  wire  \inst_dob_mux_b1/B5_0 ;
  wire  \inst_dob_mux_b1/B5_1 ;
  wire  \inst_dob_mux_b10/B0_0 ;
  wire  \inst_dob_mux_b10/B0_1 ;
  wire  \inst_dob_mux_b10/B0_10 ;
  wire  \inst_dob_mux_b10/B0_11 ;
  wire  \inst_dob_mux_b10/B0_12 ;
  wire  \inst_dob_mux_b10/B0_13 ;
  wire  \inst_dob_mux_b10/B0_14 ;
  wire  \inst_dob_mux_b10/B0_15 ;
  wire  \inst_dob_mux_b10/B0_16 ;
  wire  \inst_dob_mux_b10/B0_17 ;
  wire  \inst_dob_mux_b10/B0_18 ;
  wire  \inst_dob_mux_b10/B0_19 ;
  wire  \inst_dob_mux_b10/B0_2 ;
  wire  \inst_dob_mux_b10/B0_20 ;
  wire  \inst_dob_mux_b10/B0_21 ;
  wire  \inst_dob_mux_b10/B0_22 ;
  wire  \inst_dob_mux_b10/B0_23 ;
  wire  \inst_dob_mux_b10/B0_24 ;
  wire  \inst_dob_mux_b10/B0_25 ;
  wire  \inst_dob_mux_b10/B0_26 ;
  wire  \inst_dob_mux_b10/B0_27 ;
  wire  \inst_dob_mux_b10/B0_28 ;
  wire  \inst_dob_mux_b10/B0_29 ;
  wire  \inst_dob_mux_b10/B0_3 ;
  wire  \inst_dob_mux_b10/B0_30 ;
  wire  \inst_dob_mux_b10/B0_31 ;
  wire  \inst_dob_mux_b10/B0_32 ;
  wire  \inst_dob_mux_b10/B0_33 ;
  wire  \inst_dob_mux_b10/B0_34 ;
  wire  \inst_dob_mux_b10/B0_35 ;
  wire  \inst_dob_mux_b10/B0_36 ;
  wire  \inst_dob_mux_b10/B0_37 ;
  wire  \inst_dob_mux_b10/B0_38 ;
  wire  \inst_dob_mux_b10/B0_39 ;
  wire  \inst_dob_mux_b10/B0_4 ;
  wire  \inst_dob_mux_b10/B0_40 ;
  wire  \inst_dob_mux_b10/B0_41 ;
  wire  \inst_dob_mux_b10/B0_42 ;
  wire  \inst_dob_mux_b10/B0_43 ;
  wire  \inst_dob_mux_b10/B0_44 ;
  wire  \inst_dob_mux_b10/B0_45 ;
  wire  \inst_dob_mux_b10/B0_46 ;
  wire  \inst_dob_mux_b10/B0_47 ;
  wire  \inst_dob_mux_b10/B0_48 ;
  wire  \inst_dob_mux_b10/B0_49 ;
  wire  \inst_dob_mux_b10/B0_5 ;
  wire  \inst_dob_mux_b10/B0_50 ;
  wire  \inst_dob_mux_b10/B0_51 ;
  wire  \inst_dob_mux_b10/B0_52 ;
  wire  \inst_dob_mux_b10/B0_53 ;
  wire  \inst_dob_mux_b10/B0_54 ;
  wire  \inst_dob_mux_b10/B0_55 ;
  wire  \inst_dob_mux_b10/B0_56 ;
  wire  \inst_dob_mux_b10/B0_57 ;
  wire  \inst_dob_mux_b10/B0_58 ;
  wire  \inst_dob_mux_b10/B0_59 ;
  wire  \inst_dob_mux_b10/B0_6 ;
  wire  \inst_dob_mux_b10/B0_60 ;
  wire  \inst_dob_mux_b10/B0_61 ;
  wire  \inst_dob_mux_b10/B0_62 ;
  wire  \inst_dob_mux_b10/B0_63 ;
  wire  \inst_dob_mux_b10/B0_7 ;
  wire  \inst_dob_mux_b10/B0_8 ;
  wire  \inst_dob_mux_b10/B0_9 ;
  wire  \inst_dob_mux_b10/B1_0 ;
  wire  \inst_dob_mux_b10/B1_1 ;
  wire  \inst_dob_mux_b10/B1_10 ;
  wire  \inst_dob_mux_b10/B1_11 ;
  wire  \inst_dob_mux_b10/B1_12 ;
  wire  \inst_dob_mux_b10/B1_13 ;
  wire  \inst_dob_mux_b10/B1_14 ;
  wire  \inst_dob_mux_b10/B1_15 ;
  wire  \inst_dob_mux_b10/B1_16 ;
  wire  \inst_dob_mux_b10/B1_17 ;
  wire  \inst_dob_mux_b10/B1_18 ;
  wire  \inst_dob_mux_b10/B1_19 ;
  wire  \inst_dob_mux_b10/B1_2 ;
  wire  \inst_dob_mux_b10/B1_20 ;
  wire  \inst_dob_mux_b10/B1_21 ;
  wire  \inst_dob_mux_b10/B1_22 ;
  wire  \inst_dob_mux_b10/B1_23 ;
  wire  \inst_dob_mux_b10/B1_24 ;
  wire  \inst_dob_mux_b10/B1_25 ;
  wire  \inst_dob_mux_b10/B1_26 ;
  wire  \inst_dob_mux_b10/B1_27 ;
  wire  \inst_dob_mux_b10/B1_28 ;
  wire  \inst_dob_mux_b10/B1_29 ;
  wire  \inst_dob_mux_b10/B1_3 ;
  wire  \inst_dob_mux_b10/B1_30 ;
  wire  \inst_dob_mux_b10/B1_31 ;
  wire  \inst_dob_mux_b10/B1_4 ;
  wire  \inst_dob_mux_b10/B1_5 ;
  wire  \inst_dob_mux_b10/B1_6 ;
  wire  \inst_dob_mux_b10/B1_7 ;
  wire  \inst_dob_mux_b10/B1_8 ;
  wire  \inst_dob_mux_b10/B1_9 ;
  wire  \inst_dob_mux_b10/B2_0 ;
  wire  \inst_dob_mux_b10/B2_1 ;
  wire  \inst_dob_mux_b10/B2_10 ;
  wire  \inst_dob_mux_b10/B2_11 ;
  wire  \inst_dob_mux_b10/B2_12 ;
  wire  \inst_dob_mux_b10/B2_13 ;
  wire  \inst_dob_mux_b10/B2_14 ;
  wire  \inst_dob_mux_b10/B2_15 ;
  wire  \inst_dob_mux_b10/B2_2 ;
  wire  \inst_dob_mux_b10/B2_3 ;
  wire  \inst_dob_mux_b10/B2_4 ;
  wire  \inst_dob_mux_b10/B2_5 ;
  wire  \inst_dob_mux_b10/B2_6 ;
  wire  \inst_dob_mux_b10/B2_7 ;
  wire  \inst_dob_mux_b10/B2_8 ;
  wire  \inst_dob_mux_b10/B2_9 ;
  wire  \inst_dob_mux_b10/B3_0 ;
  wire  \inst_dob_mux_b10/B3_1 ;
  wire  \inst_dob_mux_b10/B3_2 ;
  wire  \inst_dob_mux_b10/B3_3 ;
  wire  \inst_dob_mux_b10/B3_4 ;
  wire  \inst_dob_mux_b10/B3_5 ;
  wire  \inst_dob_mux_b10/B3_6 ;
  wire  \inst_dob_mux_b10/B3_7 ;
  wire  \inst_dob_mux_b10/B4_0 ;
  wire  \inst_dob_mux_b10/B4_1 ;
  wire  \inst_dob_mux_b10/B4_2 ;
  wire  \inst_dob_mux_b10/B4_3 ;
  wire  \inst_dob_mux_b10/B5_0 ;
  wire  \inst_dob_mux_b10/B5_1 ;
  wire  \inst_dob_mux_b11/B0_0 ;
  wire  \inst_dob_mux_b11/B0_1 ;
  wire  \inst_dob_mux_b11/B0_10 ;
  wire  \inst_dob_mux_b11/B0_11 ;
  wire  \inst_dob_mux_b11/B0_12 ;
  wire  \inst_dob_mux_b11/B0_13 ;
  wire  \inst_dob_mux_b11/B0_14 ;
  wire  \inst_dob_mux_b11/B0_15 ;
  wire  \inst_dob_mux_b11/B0_16 ;
  wire  \inst_dob_mux_b11/B0_17 ;
  wire  \inst_dob_mux_b11/B0_18 ;
  wire  \inst_dob_mux_b11/B0_19 ;
  wire  \inst_dob_mux_b11/B0_2 ;
  wire  \inst_dob_mux_b11/B0_20 ;
  wire  \inst_dob_mux_b11/B0_21 ;
  wire  \inst_dob_mux_b11/B0_22 ;
  wire  \inst_dob_mux_b11/B0_23 ;
  wire  \inst_dob_mux_b11/B0_24 ;
  wire  \inst_dob_mux_b11/B0_25 ;
  wire  \inst_dob_mux_b11/B0_26 ;
  wire  \inst_dob_mux_b11/B0_27 ;
  wire  \inst_dob_mux_b11/B0_28 ;
  wire  \inst_dob_mux_b11/B0_29 ;
  wire  \inst_dob_mux_b11/B0_3 ;
  wire  \inst_dob_mux_b11/B0_30 ;
  wire  \inst_dob_mux_b11/B0_31 ;
  wire  \inst_dob_mux_b11/B0_32 ;
  wire  \inst_dob_mux_b11/B0_33 ;
  wire  \inst_dob_mux_b11/B0_34 ;
  wire  \inst_dob_mux_b11/B0_35 ;
  wire  \inst_dob_mux_b11/B0_36 ;
  wire  \inst_dob_mux_b11/B0_37 ;
  wire  \inst_dob_mux_b11/B0_38 ;
  wire  \inst_dob_mux_b11/B0_39 ;
  wire  \inst_dob_mux_b11/B0_4 ;
  wire  \inst_dob_mux_b11/B0_40 ;
  wire  \inst_dob_mux_b11/B0_41 ;
  wire  \inst_dob_mux_b11/B0_42 ;
  wire  \inst_dob_mux_b11/B0_43 ;
  wire  \inst_dob_mux_b11/B0_44 ;
  wire  \inst_dob_mux_b11/B0_45 ;
  wire  \inst_dob_mux_b11/B0_46 ;
  wire  \inst_dob_mux_b11/B0_47 ;
  wire  \inst_dob_mux_b11/B0_48 ;
  wire  \inst_dob_mux_b11/B0_49 ;
  wire  \inst_dob_mux_b11/B0_5 ;
  wire  \inst_dob_mux_b11/B0_50 ;
  wire  \inst_dob_mux_b11/B0_51 ;
  wire  \inst_dob_mux_b11/B0_52 ;
  wire  \inst_dob_mux_b11/B0_53 ;
  wire  \inst_dob_mux_b11/B0_54 ;
  wire  \inst_dob_mux_b11/B0_55 ;
  wire  \inst_dob_mux_b11/B0_56 ;
  wire  \inst_dob_mux_b11/B0_57 ;
  wire  \inst_dob_mux_b11/B0_58 ;
  wire  \inst_dob_mux_b11/B0_59 ;
  wire  \inst_dob_mux_b11/B0_6 ;
  wire  \inst_dob_mux_b11/B0_60 ;
  wire  \inst_dob_mux_b11/B0_61 ;
  wire  \inst_dob_mux_b11/B0_62 ;
  wire  \inst_dob_mux_b11/B0_63 ;
  wire  \inst_dob_mux_b11/B0_7 ;
  wire  \inst_dob_mux_b11/B0_8 ;
  wire  \inst_dob_mux_b11/B0_9 ;
  wire  \inst_dob_mux_b11/B1_0 ;
  wire  \inst_dob_mux_b11/B1_1 ;
  wire  \inst_dob_mux_b11/B1_10 ;
  wire  \inst_dob_mux_b11/B1_11 ;
  wire  \inst_dob_mux_b11/B1_12 ;
  wire  \inst_dob_mux_b11/B1_13 ;
  wire  \inst_dob_mux_b11/B1_14 ;
  wire  \inst_dob_mux_b11/B1_15 ;
  wire  \inst_dob_mux_b11/B1_16 ;
  wire  \inst_dob_mux_b11/B1_17 ;
  wire  \inst_dob_mux_b11/B1_18 ;
  wire  \inst_dob_mux_b11/B1_19 ;
  wire  \inst_dob_mux_b11/B1_2 ;
  wire  \inst_dob_mux_b11/B1_20 ;
  wire  \inst_dob_mux_b11/B1_21 ;
  wire  \inst_dob_mux_b11/B1_22 ;
  wire  \inst_dob_mux_b11/B1_23 ;
  wire  \inst_dob_mux_b11/B1_24 ;
  wire  \inst_dob_mux_b11/B1_25 ;
  wire  \inst_dob_mux_b11/B1_26 ;
  wire  \inst_dob_mux_b11/B1_27 ;
  wire  \inst_dob_mux_b11/B1_28 ;
  wire  \inst_dob_mux_b11/B1_29 ;
  wire  \inst_dob_mux_b11/B1_3 ;
  wire  \inst_dob_mux_b11/B1_30 ;
  wire  \inst_dob_mux_b11/B1_31 ;
  wire  \inst_dob_mux_b11/B1_4 ;
  wire  \inst_dob_mux_b11/B1_5 ;
  wire  \inst_dob_mux_b11/B1_6 ;
  wire  \inst_dob_mux_b11/B1_7 ;
  wire  \inst_dob_mux_b11/B1_8 ;
  wire  \inst_dob_mux_b11/B1_9 ;
  wire  \inst_dob_mux_b11/B2_0 ;
  wire  \inst_dob_mux_b11/B2_1 ;
  wire  \inst_dob_mux_b11/B2_10 ;
  wire  \inst_dob_mux_b11/B2_11 ;
  wire  \inst_dob_mux_b11/B2_12 ;
  wire  \inst_dob_mux_b11/B2_13 ;
  wire  \inst_dob_mux_b11/B2_14 ;
  wire  \inst_dob_mux_b11/B2_15 ;
  wire  \inst_dob_mux_b11/B2_2 ;
  wire  \inst_dob_mux_b11/B2_3 ;
  wire  \inst_dob_mux_b11/B2_4 ;
  wire  \inst_dob_mux_b11/B2_5 ;
  wire  \inst_dob_mux_b11/B2_6 ;
  wire  \inst_dob_mux_b11/B2_7 ;
  wire  \inst_dob_mux_b11/B2_8 ;
  wire  \inst_dob_mux_b11/B2_9 ;
  wire  \inst_dob_mux_b11/B3_0 ;
  wire  \inst_dob_mux_b11/B3_1 ;
  wire  \inst_dob_mux_b11/B3_2 ;
  wire  \inst_dob_mux_b11/B3_3 ;
  wire  \inst_dob_mux_b11/B3_4 ;
  wire  \inst_dob_mux_b11/B3_5 ;
  wire  \inst_dob_mux_b11/B3_6 ;
  wire  \inst_dob_mux_b11/B3_7 ;
  wire  \inst_dob_mux_b11/B4_0 ;
  wire  \inst_dob_mux_b11/B4_1 ;
  wire  \inst_dob_mux_b11/B4_2 ;
  wire  \inst_dob_mux_b11/B4_3 ;
  wire  \inst_dob_mux_b11/B5_0 ;
  wire  \inst_dob_mux_b11/B5_1 ;
  wire  \inst_dob_mux_b12/B0_0 ;
  wire  \inst_dob_mux_b12/B0_1 ;
  wire  \inst_dob_mux_b12/B0_10 ;
  wire  \inst_dob_mux_b12/B0_11 ;
  wire  \inst_dob_mux_b12/B0_12 ;
  wire  \inst_dob_mux_b12/B0_13 ;
  wire  \inst_dob_mux_b12/B0_14 ;
  wire  \inst_dob_mux_b12/B0_15 ;
  wire  \inst_dob_mux_b12/B0_16 ;
  wire  \inst_dob_mux_b12/B0_17 ;
  wire  \inst_dob_mux_b12/B0_18 ;
  wire  \inst_dob_mux_b12/B0_19 ;
  wire  \inst_dob_mux_b12/B0_2 ;
  wire  \inst_dob_mux_b12/B0_20 ;
  wire  \inst_dob_mux_b12/B0_21 ;
  wire  \inst_dob_mux_b12/B0_22 ;
  wire  \inst_dob_mux_b12/B0_23 ;
  wire  \inst_dob_mux_b12/B0_24 ;
  wire  \inst_dob_mux_b12/B0_25 ;
  wire  \inst_dob_mux_b12/B0_26 ;
  wire  \inst_dob_mux_b12/B0_27 ;
  wire  \inst_dob_mux_b12/B0_28 ;
  wire  \inst_dob_mux_b12/B0_29 ;
  wire  \inst_dob_mux_b12/B0_3 ;
  wire  \inst_dob_mux_b12/B0_30 ;
  wire  \inst_dob_mux_b12/B0_31 ;
  wire  \inst_dob_mux_b12/B0_32 ;
  wire  \inst_dob_mux_b12/B0_33 ;
  wire  \inst_dob_mux_b12/B0_34 ;
  wire  \inst_dob_mux_b12/B0_35 ;
  wire  \inst_dob_mux_b12/B0_36 ;
  wire  \inst_dob_mux_b12/B0_37 ;
  wire  \inst_dob_mux_b12/B0_38 ;
  wire  \inst_dob_mux_b12/B0_39 ;
  wire  \inst_dob_mux_b12/B0_4 ;
  wire  \inst_dob_mux_b12/B0_40 ;
  wire  \inst_dob_mux_b12/B0_41 ;
  wire  \inst_dob_mux_b12/B0_42 ;
  wire  \inst_dob_mux_b12/B0_43 ;
  wire  \inst_dob_mux_b12/B0_44 ;
  wire  \inst_dob_mux_b12/B0_45 ;
  wire  \inst_dob_mux_b12/B0_46 ;
  wire  \inst_dob_mux_b12/B0_47 ;
  wire  \inst_dob_mux_b12/B0_48 ;
  wire  \inst_dob_mux_b12/B0_49 ;
  wire  \inst_dob_mux_b12/B0_5 ;
  wire  \inst_dob_mux_b12/B0_50 ;
  wire  \inst_dob_mux_b12/B0_51 ;
  wire  \inst_dob_mux_b12/B0_52 ;
  wire  \inst_dob_mux_b12/B0_53 ;
  wire  \inst_dob_mux_b12/B0_54 ;
  wire  \inst_dob_mux_b12/B0_55 ;
  wire  \inst_dob_mux_b12/B0_56 ;
  wire  \inst_dob_mux_b12/B0_57 ;
  wire  \inst_dob_mux_b12/B0_58 ;
  wire  \inst_dob_mux_b12/B0_59 ;
  wire  \inst_dob_mux_b12/B0_6 ;
  wire  \inst_dob_mux_b12/B0_60 ;
  wire  \inst_dob_mux_b12/B0_61 ;
  wire  \inst_dob_mux_b12/B0_62 ;
  wire  \inst_dob_mux_b12/B0_63 ;
  wire  \inst_dob_mux_b12/B0_7 ;
  wire  \inst_dob_mux_b12/B0_8 ;
  wire  \inst_dob_mux_b12/B0_9 ;
  wire  \inst_dob_mux_b12/B1_0 ;
  wire  \inst_dob_mux_b12/B1_1 ;
  wire  \inst_dob_mux_b12/B1_10 ;
  wire  \inst_dob_mux_b12/B1_11 ;
  wire  \inst_dob_mux_b12/B1_12 ;
  wire  \inst_dob_mux_b12/B1_13 ;
  wire  \inst_dob_mux_b12/B1_14 ;
  wire  \inst_dob_mux_b12/B1_15 ;
  wire  \inst_dob_mux_b12/B1_16 ;
  wire  \inst_dob_mux_b12/B1_17 ;
  wire  \inst_dob_mux_b12/B1_18 ;
  wire  \inst_dob_mux_b12/B1_19 ;
  wire  \inst_dob_mux_b12/B1_2 ;
  wire  \inst_dob_mux_b12/B1_20 ;
  wire  \inst_dob_mux_b12/B1_21 ;
  wire  \inst_dob_mux_b12/B1_22 ;
  wire  \inst_dob_mux_b12/B1_23 ;
  wire  \inst_dob_mux_b12/B1_24 ;
  wire  \inst_dob_mux_b12/B1_25 ;
  wire  \inst_dob_mux_b12/B1_26 ;
  wire  \inst_dob_mux_b12/B1_27 ;
  wire  \inst_dob_mux_b12/B1_28 ;
  wire  \inst_dob_mux_b12/B1_29 ;
  wire  \inst_dob_mux_b12/B1_3 ;
  wire  \inst_dob_mux_b12/B1_30 ;
  wire  \inst_dob_mux_b12/B1_31 ;
  wire  \inst_dob_mux_b12/B1_4 ;
  wire  \inst_dob_mux_b12/B1_5 ;
  wire  \inst_dob_mux_b12/B1_6 ;
  wire  \inst_dob_mux_b12/B1_7 ;
  wire  \inst_dob_mux_b12/B1_8 ;
  wire  \inst_dob_mux_b12/B1_9 ;
  wire  \inst_dob_mux_b12/B2_0 ;
  wire  \inst_dob_mux_b12/B2_1 ;
  wire  \inst_dob_mux_b12/B2_10 ;
  wire  \inst_dob_mux_b12/B2_11 ;
  wire  \inst_dob_mux_b12/B2_12 ;
  wire  \inst_dob_mux_b12/B2_13 ;
  wire  \inst_dob_mux_b12/B2_14 ;
  wire  \inst_dob_mux_b12/B2_15 ;
  wire  \inst_dob_mux_b12/B2_2 ;
  wire  \inst_dob_mux_b12/B2_3 ;
  wire  \inst_dob_mux_b12/B2_4 ;
  wire  \inst_dob_mux_b12/B2_5 ;
  wire  \inst_dob_mux_b12/B2_6 ;
  wire  \inst_dob_mux_b12/B2_7 ;
  wire  \inst_dob_mux_b12/B2_8 ;
  wire  \inst_dob_mux_b12/B2_9 ;
  wire  \inst_dob_mux_b12/B3_0 ;
  wire  \inst_dob_mux_b12/B3_1 ;
  wire  \inst_dob_mux_b12/B3_2 ;
  wire  \inst_dob_mux_b12/B3_3 ;
  wire  \inst_dob_mux_b12/B3_4 ;
  wire  \inst_dob_mux_b12/B3_5 ;
  wire  \inst_dob_mux_b12/B3_6 ;
  wire  \inst_dob_mux_b12/B3_7 ;
  wire  \inst_dob_mux_b12/B4_0 ;
  wire  \inst_dob_mux_b12/B4_1 ;
  wire  \inst_dob_mux_b12/B4_2 ;
  wire  \inst_dob_mux_b12/B4_3 ;
  wire  \inst_dob_mux_b12/B5_0 ;
  wire  \inst_dob_mux_b12/B5_1 ;
  wire  \inst_dob_mux_b13/B0_0 ;
  wire  \inst_dob_mux_b13/B0_1 ;
  wire  \inst_dob_mux_b13/B0_10 ;
  wire  \inst_dob_mux_b13/B0_11 ;
  wire  \inst_dob_mux_b13/B0_12 ;
  wire  \inst_dob_mux_b13/B0_13 ;
  wire  \inst_dob_mux_b13/B0_14 ;
  wire  \inst_dob_mux_b13/B0_15 ;
  wire  \inst_dob_mux_b13/B0_16 ;
  wire  \inst_dob_mux_b13/B0_17 ;
  wire  \inst_dob_mux_b13/B0_18 ;
  wire  \inst_dob_mux_b13/B0_19 ;
  wire  \inst_dob_mux_b13/B0_2 ;
  wire  \inst_dob_mux_b13/B0_20 ;
  wire  \inst_dob_mux_b13/B0_21 ;
  wire  \inst_dob_mux_b13/B0_22 ;
  wire  \inst_dob_mux_b13/B0_23 ;
  wire  \inst_dob_mux_b13/B0_24 ;
  wire  \inst_dob_mux_b13/B0_25 ;
  wire  \inst_dob_mux_b13/B0_26 ;
  wire  \inst_dob_mux_b13/B0_27 ;
  wire  \inst_dob_mux_b13/B0_28 ;
  wire  \inst_dob_mux_b13/B0_29 ;
  wire  \inst_dob_mux_b13/B0_3 ;
  wire  \inst_dob_mux_b13/B0_30 ;
  wire  \inst_dob_mux_b13/B0_31 ;
  wire  \inst_dob_mux_b13/B0_32 ;
  wire  \inst_dob_mux_b13/B0_33 ;
  wire  \inst_dob_mux_b13/B0_34 ;
  wire  \inst_dob_mux_b13/B0_35 ;
  wire  \inst_dob_mux_b13/B0_36 ;
  wire  \inst_dob_mux_b13/B0_37 ;
  wire  \inst_dob_mux_b13/B0_38 ;
  wire  \inst_dob_mux_b13/B0_39 ;
  wire  \inst_dob_mux_b13/B0_4 ;
  wire  \inst_dob_mux_b13/B0_40 ;
  wire  \inst_dob_mux_b13/B0_41 ;
  wire  \inst_dob_mux_b13/B0_42 ;
  wire  \inst_dob_mux_b13/B0_43 ;
  wire  \inst_dob_mux_b13/B0_44 ;
  wire  \inst_dob_mux_b13/B0_45 ;
  wire  \inst_dob_mux_b13/B0_46 ;
  wire  \inst_dob_mux_b13/B0_47 ;
  wire  \inst_dob_mux_b13/B0_48 ;
  wire  \inst_dob_mux_b13/B0_49 ;
  wire  \inst_dob_mux_b13/B0_5 ;
  wire  \inst_dob_mux_b13/B0_50 ;
  wire  \inst_dob_mux_b13/B0_51 ;
  wire  \inst_dob_mux_b13/B0_52 ;
  wire  \inst_dob_mux_b13/B0_53 ;
  wire  \inst_dob_mux_b13/B0_54 ;
  wire  \inst_dob_mux_b13/B0_55 ;
  wire  \inst_dob_mux_b13/B0_56 ;
  wire  \inst_dob_mux_b13/B0_57 ;
  wire  \inst_dob_mux_b13/B0_58 ;
  wire  \inst_dob_mux_b13/B0_59 ;
  wire  \inst_dob_mux_b13/B0_6 ;
  wire  \inst_dob_mux_b13/B0_60 ;
  wire  \inst_dob_mux_b13/B0_61 ;
  wire  \inst_dob_mux_b13/B0_62 ;
  wire  \inst_dob_mux_b13/B0_63 ;
  wire  \inst_dob_mux_b13/B0_7 ;
  wire  \inst_dob_mux_b13/B0_8 ;
  wire  \inst_dob_mux_b13/B0_9 ;
  wire  \inst_dob_mux_b13/B1_0 ;
  wire  \inst_dob_mux_b13/B1_1 ;
  wire  \inst_dob_mux_b13/B1_10 ;
  wire  \inst_dob_mux_b13/B1_11 ;
  wire  \inst_dob_mux_b13/B1_12 ;
  wire  \inst_dob_mux_b13/B1_13 ;
  wire  \inst_dob_mux_b13/B1_14 ;
  wire  \inst_dob_mux_b13/B1_15 ;
  wire  \inst_dob_mux_b13/B1_16 ;
  wire  \inst_dob_mux_b13/B1_17 ;
  wire  \inst_dob_mux_b13/B1_18 ;
  wire  \inst_dob_mux_b13/B1_19 ;
  wire  \inst_dob_mux_b13/B1_2 ;
  wire  \inst_dob_mux_b13/B1_20 ;
  wire  \inst_dob_mux_b13/B1_21 ;
  wire  \inst_dob_mux_b13/B1_22 ;
  wire  \inst_dob_mux_b13/B1_23 ;
  wire  \inst_dob_mux_b13/B1_24 ;
  wire  \inst_dob_mux_b13/B1_25 ;
  wire  \inst_dob_mux_b13/B1_26 ;
  wire  \inst_dob_mux_b13/B1_27 ;
  wire  \inst_dob_mux_b13/B1_28 ;
  wire  \inst_dob_mux_b13/B1_29 ;
  wire  \inst_dob_mux_b13/B1_3 ;
  wire  \inst_dob_mux_b13/B1_30 ;
  wire  \inst_dob_mux_b13/B1_31 ;
  wire  \inst_dob_mux_b13/B1_4 ;
  wire  \inst_dob_mux_b13/B1_5 ;
  wire  \inst_dob_mux_b13/B1_6 ;
  wire  \inst_dob_mux_b13/B1_7 ;
  wire  \inst_dob_mux_b13/B1_8 ;
  wire  \inst_dob_mux_b13/B1_9 ;
  wire  \inst_dob_mux_b13/B2_0 ;
  wire  \inst_dob_mux_b13/B2_1 ;
  wire  \inst_dob_mux_b13/B2_10 ;
  wire  \inst_dob_mux_b13/B2_11 ;
  wire  \inst_dob_mux_b13/B2_12 ;
  wire  \inst_dob_mux_b13/B2_13 ;
  wire  \inst_dob_mux_b13/B2_14 ;
  wire  \inst_dob_mux_b13/B2_15 ;
  wire  \inst_dob_mux_b13/B2_2 ;
  wire  \inst_dob_mux_b13/B2_3 ;
  wire  \inst_dob_mux_b13/B2_4 ;
  wire  \inst_dob_mux_b13/B2_5 ;
  wire  \inst_dob_mux_b13/B2_6 ;
  wire  \inst_dob_mux_b13/B2_7 ;
  wire  \inst_dob_mux_b13/B2_8 ;
  wire  \inst_dob_mux_b13/B2_9 ;
  wire  \inst_dob_mux_b13/B3_0 ;
  wire  \inst_dob_mux_b13/B3_1 ;
  wire  \inst_dob_mux_b13/B3_2 ;
  wire  \inst_dob_mux_b13/B3_3 ;
  wire  \inst_dob_mux_b13/B3_4 ;
  wire  \inst_dob_mux_b13/B3_5 ;
  wire  \inst_dob_mux_b13/B3_6 ;
  wire  \inst_dob_mux_b13/B3_7 ;
  wire  \inst_dob_mux_b13/B4_0 ;
  wire  \inst_dob_mux_b13/B4_1 ;
  wire  \inst_dob_mux_b13/B4_2 ;
  wire  \inst_dob_mux_b13/B4_3 ;
  wire  \inst_dob_mux_b13/B5_0 ;
  wire  \inst_dob_mux_b13/B5_1 ;
  wire  \inst_dob_mux_b14/B0_0 ;
  wire  \inst_dob_mux_b14/B0_1 ;
  wire  \inst_dob_mux_b14/B0_10 ;
  wire  \inst_dob_mux_b14/B0_11 ;
  wire  \inst_dob_mux_b14/B0_12 ;
  wire  \inst_dob_mux_b14/B0_13 ;
  wire  \inst_dob_mux_b14/B0_14 ;
  wire  \inst_dob_mux_b14/B0_15 ;
  wire  \inst_dob_mux_b14/B0_16 ;
  wire  \inst_dob_mux_b14/B0_17 ;
  wire  \inst_dob_mux_b14/B0_18 ;
  wire  \inst_dob_mux_b14/B0_19 ;
  wire  \inst_dob_mux_b14/B0_2 ;
  wire  \inst_dob_mux_b14/B0_20 ;
  wire  \inst_dob_mux_b14/B0_21 ;
  wire  \inst_dob_mux_b14/B0_22 ;
  wire  \inst_dob_mux_b14/B0_23 ;
  wire  \inst_dob_mux_b14/B0_24 ;
  wire  \inst_dob_mux_b14/B0_25 ;
  wire  \inst_dob_mux_b14/B0_26 ;
  wire  \inst_dob_mux_b14/B0_27 ;
  wire  \inst_dob_mux_b14/B0_28 ;
  wire  \inst_dob_mux_b14/B0_29 ;
  wire  \inst_dob_mux_b14/B0_3 ;
  wire  \inst_dob_mux_b14/B0_30 ;
  wire  \inst_dob_mux_b14/B0_31 ;
  wire  \inst_dob_mux_b14/B0_32 ;
  wire  \inst_dob_mux_b14/B0_33 ;
  wire  \inst_dob_mux_b14/B0_34 ;
  wire  \inst_dob_mux_b14/B0_35 ;
  wire  \inst_dob_mux_b14/B0_36 ;
  wire  \inst_dob_mux_b14/B0_37 ;
  wire  \inst_dob_mux_b14/B0_38 ;
  wire  \inst_dob_mux_b14/B0_39 ;
  wire  \inst_dob_mux_b14/B0_4 ;
  wire  \inst_dob_mux_b14/B0_40 ;
  wire  \inst_dob_mux_b14/B0_41 ;
  wire  \inst_dob_mux_b14/B0_42 ;
  wire  \inst_dob_mux_b14/B0_43 ;
  wire  \inst_dob_mux_b14/B0_44 ;
  wire  \inst_dob_mux_b14/B0_45 ;
  wire  \inst_dob_mux_b14/B0_46 ;
  wire  \inst_dob_mux_b14/B0_47 ;
  wire  \inst_dob_mux_b14/B0_48 ;
  wire  \inst_dob_mux_b14/B0_49 ;
  wire  \inst_dob_mux_b14/B0_5 ;
  wire  \inst_dob_mux_b14/B0_50 ;
  wire  \inst_dob_mux_b14/B0_51 ;
  wire  \inst_dob_mux_b14/B0_52 ;
  wire  \inst_dob_mux_b14/B0_53 ;
  wire  \inst_dob_mux_b14/B0_54 ;
  wire  \inst_dob_mux_b14/B0_55 ;
  wire  \inst_dob_mux_b14/B0_56 ;
  wire  \inst_dob_mux_b14/B0_57 ;
  wire  \inst_dob_mux_b14/B0_58 ;
  wire  \inst_dob_mux_b14/B0_59 ;
  wire  \inst_dob_mux_b14/B0_6 ;
  wire  \inst_dob_mux_b14/B0_60 ;
  wire  \inst_dob_mux_b14/B0_61 ;
  wire  \inst_dob_mux_b14/B0_62 ;
  wire  \inst_dob_mux_b14/B0_63 ;
  wire  \inst_dob_mux_b14/B0_7 ;
  wire  \inst_dob_mux_b14/B0_8 ;
  wire  \inst_dob_mux_b14/B0_9 ;
  wire  \inst_dob_mux_b14/B1_0 ;
  wire  \inst_dob_mux_b14/B1_1 ;
  wire  \inst_dob_mux_b14/B1_10 ;
  wire  \inst_dob_mux_b14/B1_11 ;
  wire  \inst_dob_mux_b14/B1_12 ;
  wire  \inst_dob_mux_b14/B1_13 ;
  wire  \inst_dob_mux_b14/B1_14 ;
  wire  \inst_dob_mux_b14/B1_15 ;
  wire  \inst_dob_mux_b14/B1_16 ;
  wire  \inst_dob_mux_b14/B1_17 ;
  wire  \inst_dob_mux_b14/B1_18 ;
  wire  \inst_dob_mux_b14/B1_19 ;
  wire  \inst_dob_mux_b14/B1_2 ;
  wire  \inst_dob_mux_b14/B1_20 ;
  wire  \inst_dob_mux_b14/B1_21 ;
  wire  \inst_dob_mux_b14/B1_22 ;
  wire  \inst_dob_mux_b14/B1_23 ;
  wire  \inst_dob_mux_b14/B1_24 ;
  wire  \inst_dob_mux_b14/B1_25 ;
  wire  \inst_dob_mux_b14/B1_26 ;
  wire  \inst_dob_mux_b14/B1_27 ;
  wire  \inst_dob_mux_b14/B1_28 ;
  wire  \inst_dob_mux_b14/B1_29 ;
  wire  \inst_dob_mux_b14/B1_3 ;
  wire  \inst_dob_mux_b14/B1_30 ;
  wire  \inst_dob_mux_b14/B1_31 ;
  wire  \inst_dob_mux_b14/B1_4 ;
  wire  \inst_dob_mux_b14/B1_5 ;
  wire  \inst_dob_mux_b14/B1_6 ;
  wire  \inst_dob_mux_b14/B1_7 ;
  wire  \inst_dob_mux_b14/B1_8 ;
  wire  \inst_dob_mux_b14/B1_9 ;
  wire  \inst_dob_mux_b14/B2_0 ;
  wire  \inst_dob_mux_b14/B2_1 ;
  wire  \inst_dob_mux_b14/B2_10 ;
  wire  \inst_dob_mux_b14/B2_11 ;
  wire  \inst_dob_mux_b14/B2_12 ;
  wire  \inst_dob_mux_b14/B2_13 ;
  wire  \inst_dob_mux_b14/B2_14 ;
  wire  \inst_dob_mux_b14/B2_15 ;
  wire  \inst_dob_mux_b14/B2_2 ;
  wire  \inst_dob_mux_b14/B2_3 ;
  wire  \inst_dob_mux_b14/B2_4 ;
  wire  \inst_dob_mux_b14/B2_5 ;
  wire  \inst_dob_mux_b14/B2_6 ;
  wire  \inst_dob_mux_b14/B2_7 ;
  wire  \inst_dob_mux_b14/B2_8 ;
  wire  \inst_dob_mux_b14/B2_9 ;
  wire  \inst_dob_mux_b14/B3_0 ;
  wire  \inst_dob_mux_b14/B3_1 ;
  wire  \inst_dob_mux_b14/B3_2 ;
  wire  \inst_dob_mux_b14/B3_3 ;
  wire  \inst_dob_mux_b14/B3_4 ;
  wire  \inst_dob_mux_b14/B3_5 ;
  wire  \inst_dob_mux_b14/B3_6 ;
  wire  \inst_dob_mux_b14/B3_7 ;
  wire  \inst_dob_mux_b14/B4_0 ;
  wire  \inst_dob_mux_b14/B4_1 ;
  wire  \inst_dob_mux_b14/B4_2 ;
  wire  \inst_dob_mux_b14/B4_3 ;
  wire  \inst_dob_mux_b14/B5_0 ;
  wire  \inst_dob_mux_b14/B5_1 ;
  wire  \inst_dob_mux_b15/B0_0 ;
  wire  \inst_dob_mux_b15/B0_1 ;
  wire  \inst_dob_mux_b15/B0_10 ;
  wire  \inst_dob_mux_b15/B0_11 ;
  wire  \inst_dob_mux_b15/B0_12 ;
  wire  \inst_dob_mux_b15/B0_13 ;
  wire  \inst_dob_mux_b15/B0_14 ;
  wire  \inst_dob_mux_b15/B0_15 ;
  wire  \inst_dob_mux_b15/B0_16 ;
  wire  \inst_dob_mux_b15/B0_17 ;
  wire  \inst_dob_mux_b15/B0_18 ;
  wire  \inst_dob_mux_b15/B0_19 ;
  wire  \inst_dob_mux_b15/B0_2 ;
  wire  \inst_dob_mux_b15/B0_20 ;
  wire  \inst_dob_mux_b15/B0_21 ;
  wire  \inst_dob_mux_b15/B0_22 ;
  wire  \inst_dob_mux_b15/B0_23 ;
  wire  \inst_dob_mux_b15/B0_24 ;
  wire  \inst_dob_mux_b15/B0_25 ;
  wire  \inst_dob_mux_b15/B0_26 ;
  wire  \inst_dob_mux_b15/B0_27 ;
  wire  \inst_dob_mux_b15/B0_28 ;
  wire  \inst_dob_mux_b15/B0_29 ;
  wire  \inst_dob_mux_b15/B0_3 ;
  wire  \inst_dob_mux_b15/B0_30 ;
  wire  \inst_dob_mux_b15/B0_31 ;
  wire  \inst_dob_mux_b15/B0_32 ;
  wire  \inst_dob_mux_b15/B0_33 ;
  wire  \inst_dob_mux_b15/B0_34 ;
  wire  \inst_dob_mux_b15/B0_35 ;
  wire  \inst_dob_mux_b15/B0_36 ;
  wire  \inst_dob_mux_b15/B0_37 ;
  wire  \inst_dob_mux_b15/B0_38 ;
  wire  \inst_dob_mux_b15/B0_39 ;
  wire  \inst_dob_mux_b15/B0_4 ;
  wire  \inst_dob_mux_b15/B0_40 ;
  wire  \inst_dob_mux_b15/B0_41 ;
  wire  \inst_dob_mux_b15/B0_42 ;
  wire  \inst_dob_mux_b15/B0_43 ;
  wire  \inst_dob_mux_b15/B0_44 ;
  wire  \inst_dob_mux_b15/B0_45 ;
  wire  \inst_dob_mux_b15/B0_46 ;
  wire  \inst_dob_mux_b15/B0_47 ;
  wire  \inst_dob_mux_b15/B0_48 ;
  wire  \inst_dob_mux_b15/B0_49 ;
  wire  \inst_dob_mux_b15/B0_5 ;
  wire  \inst_dob_mux_b15/B0_50 ;
  wire  \inst_dob_mux_b15/B0_51 ;
  wire  \inst_dob_mux_b15/B0_52 ;
  wire  \inst_dob_mux_b15/B0_53 ;
  wire  \inst_dob_mux_b15/B0_54 ;
  wire  \inst_dob_mux_b15/B0_55 ;
  wire  \inst_dob_mux_b15/B0_56 ;
  wire  \inst_dob_mux_b15/B0_57 ;
  wire  \inst_dob_mux_b15/B0_58 ;
  wire  \inst_dob_mux_b15/B0_59 ;
  wire  \inst_dob_mux_b15/B0_6 ;
  wire  \inst_dob_mux_b15/B0_60 ;
  wire  \inst_dob_mux_b15/B0_61 ;
  wire  \inst_dob_mux_b15/B0_62 ;
  wire  \inst_dob_mux_b15/B0_63 ;
  wire  \inst_dob_mux_b15/B0_7 ;
  wire  \inst_dob_mux_b15/B0_8 ;
  wire  \inst_dob_mux_b15/B0_9 ;
  wire  \inst_dob_mux_b15/B1_0 ;
  wire  \inst_dob_mux_b15/B1_1 ;
  wire  \inst_dob_mux_b15/B1_10 ;
  wire  \inst_dob_mux_b15/B1_11 ;
  wire  \inst_dob_mux_b15/B1_12 ;
  wire  \inst_dob_mux_b15/B1_13 ;
  wire  \inst_dob_mux_b15/B1_14 ;
  wire  \inst_dob_mux_b15/B1_15 ;
  wire  \inst_dob_mux_b15/B1_16 ;
  wire  \inst_dob_mux_b15/B1_17 ;
  wire  \inst_dob_mux_b15/B1_18 ;
  wire  \inst_dob_mux_b15/B1_19 ;
  wire  \inst_dob_mux_b15/B1_2 ;
  wire  \inst_dob_mux_b15/B1_20 ;
  wire  \inst_dob_mux_b15/B1_21 ;
  wire  \inst_dob_mux_b15/B1_22 ;
  wire  \inst_dob_mux_b15/B1_23 ;
  wire  \inst_dob_mux_b15/B1_24 ;
  wire  \inst_dob_mux_b15/B1_25 ;
  wire  \inst_dob_mux_b15/B1_26 ;
  wire  \inst_dob_mux_b15/B1_27 ;
  wire  \inst_dob_mux_b15/B1_28 ;
  wire  \inst_dob_mux_b15/B1_29 ;
  wire  \inst_dob_mux_b15/B1_3 ;
  wire  \inst_dob_mux_b15/B1_30 ;
  wire  \inst_dob_mux_b15/B1_31 ;
  wire  \inst_dob_mux_b15/B1_4 ;
  wire  \inst_dob_mux_b15/B1_5 ;
  wire  \inst_dob_mux_b15/B1_6 ;
  wire  \inst_dob_mux_b15/B1_7 ;
  wire  \inst_dob_mux_b15/B1_8 ;
  wire  \inst_dob_mux_b15/B1_9 ;
  wire  \inst_dob_mux_b15/B2_0 ;
  wire  \inst_dob_mux_b15/B2_1 ;
  wire  \inst_dob_mux_b15/B2_10 ;
  wire  \inst_dob_mux_b15/B2_11 ;
  wire  \inst_dob_mux_b15/B2_12 ;
  wire  \inst_dob_mux_b15/B2_13 ;
  wire  \inst_dob_mux_b15/B2_14 ;
  wire  \inst_dob_mux_b15/B2_15 ;
  wire  \inst_dob_mux_b15/B2_2 ;
  wire  \inst_dob_mux_b15/B2_3 ;
  wire  \inst_dob_mux_b15/B2_4 ;
  wire  \inst_dob_mux_b15/B2_5 ;
  wire  \inst_dob_mux_b15/B2_6 ;
  wire  \inst_dob_mux_b15/B2_7 ;
  wire  \inst_dob_mux_b15/B2_8 ;
  wire  \inst_dob_mux_b15/B2_9 ;
  wire  \inst_dob_mux_b15/B3_0 ;
  wire  \inst_dob_mux_b15/B3_1 ;
  wire  \inst_dob_mux_b15/B3_2 ;
  wire  \inst_dob_mux_b15/B3_3 ;
  wire  \inst_dob_mux_b15/B3_4 ;
  wire  \inst_dob_mux_b15/B3_5 ;
  wire  \inst_dob_mux_b15/B3_6 ;
  wire  \inst_dob_mux_b15/B3_7 ;
  wire  \inst_dob_mux_b15/B4_0 ;
  wire  \inst_dob_mux_b15/B4_1 ;
  wire  \inst_dob_mux_b15/B4_2 ;
  wire  \inst_dob_mux_b15/B4_3 ;
  wire  \inst_dob_mux_b15/B5_0 ;
  wire  \inst_dob_mux_b15/B5_1 ;
  wire  \inst_dob_mux_b2/B0_0 ;
  wire  \inst_dob_mux_b2/B0_1 ;
  wire  \inst_dob_mux_b2/B0_10 ;
  wire  \inst_dob_mux_b2/B0_11 ;
  wire  \inst_dob_mux_b2/B0_12 ;
  wire  \inst_dob_mux_b2/B0_13 ;
  wire  \inst_dob_mux_b2/B0_14 ;
  wire  \inst_dob_mux_b2/B0_15 ;
  wire  \inst_dob_mux_b2/B0_16 ;
  wire  \inst_dob_mux_b2/B0_17 ;
  wire  \inst_dob_mux_b2/B0_18 ;
  wire  \inst_dob_mux_b2/B0_19 ;
  wire  \inst_dob_mux_b2/B0_2 ;
  wire  \inst_dob_mux_b2/B0_20 ;
  wire  \inst_dob_mux_b2/B0_21 ;
  wire  \inst_dob_mux_b2/B0_22 ;
  wire  \inst_dob_mux_b2/B0_23 ;
  wire  \inst_dob_mux_b2/B0_24 ;
  wire  \inst_dob_mux_b2/B0_25 ;
  wire  \inst_dob_mux_b2/B0_26 ;
  wire  \inst_dob_mux_b2/B0_27 ;
  wire  \inst_dob_mux_b2/B0_28 ;
  wire  \inst_dob_mux_b2/B0_29 ;
  wire  \inst_dob_mux_b2/B0_3 ;
  wire  \inst_dob_mux_b2/B0_30 ;
  wire  \inst_dob_mux_b2/B0_31 ;
  wire  \inst_dob_mux_b2/B0_32 ;
  wire  \inst_dob_mux_b2/B0_33 ;
  wire  \inst_dob_mux_b2/B0_34 ;
  wire  \inst_dob_mux_b2/B0_35 ;
  wire  \inst_dob_mux_b2/B0_36 ;
  wire  \inst_dob_mux_b2/B0_37 ;
  wire  \inst_dob_mux_b2/B0_38 ;
  wire  \inst_dob_mux_b2/B0_39 ;
  wire  \inst_dob_mux_b2/B0_4 ;
  wire  \inst_dob_mux_b2/B0_40 ;
  wire  \inst_dob_mux_b2/B0_41 ;
  wire  \inst_dob_mux_b2/B0_42 ;
  wire  \inst_dob_mux_b2/B0_43 ;
  wire  \inst_dob_mux_b2/B0_44 ;
  wire  \inst_dob_mux_b2/B0_45 ;
  wire  \inst_dob_mux_b2/B0_46 ;
  wire  \inst_dob_mux_b2/B0_47 ;
  wire  \inst_dob_mux_b2/B0_48 ;
  wire  \inst_dob_mux_b2/B0_49 ;
  wire  \inst_dob_mux_b2/B0_5 ;
  wire  \inst_dob_mux_b2/B0_50 ;
  wire  \inst_dob_mux_b2/B0_51 ;
  wire  \inst_dob_mux_b2/B0_52 ;
  wire  \inst_dob_mux_b2/B0_53 ;
  wire  \inst_dob_mux_b2/B0_54 ;
  wire  \inst_dob_mux_b2/B0_55 ;
  wire  \inst_dob_mux_b2/B0_56 ;
  wire  \inst_dob_mux_b2/B0_57 ;
  wire  \inst_dob_mux_b2/B0_58 ;
  wire  \inst_dob_mux_b2/B0_59 ;
  wire  \inst_dob_mux_b2/B0_6 ;
  wire  \inst_dob_mux_b2/B0_60 ;
  wire  \inst_dob_mux_b2/B0_61 ;
  wire  \inst_dob_mux_b2/B0_62 ;
  wire  \inst_dob_mux_b2/B0_63 ;
  wire  \inst_dob_mux_b2/B0_7 ;
  wire  \inst_dob_mux_b2/B0_8 ;
  wire  \inst_dob_mux_b2/B0_9 ;
  wire  \inst_dob_mux_b2/B1_0 ;
  wire  \inst_dob_mux_b2/B1_1 ;
  wire  \inst_dob_mux_b2/B1_10 ;
  wire  \inst_dob_mux_b2/B1_11 ;
  wire  \inst_dob_mux_b2/B1_12 ;
  wire  \inst_dob_mux_b2/B1_13 ;
  wire  \inst_dob_mux_b2/B1_14 ;
  wire  \inst_dob_mux_b2/B1_15 ;
  wire  \inst_dob_mux_b2/B1_16 ;
  wire  \inst_dob_mux_b2/B1_17 ;
  wire  \inst_dob_mux_b2/B1_18 ;
  wire  \inst_dob_mux_b2/B1_19 ;
  wire  \inst_dob_mux_b2/B1_2 ;
  wire  \inst_dob_mux_b2/B1_20 ;
  wire  \inst_dob_mux_b2/B1_21 ;
  wire  \inst_dob_mux_b2/B1_22 ;
  wire  \inst_dob_mux_b2/B1_23 ;
  wire  \inst_dob_mux_b2/B1_24 ;
  wire  \inst_dob_mux_b2/B1_25 ;
  wire  \inst_dob_mux_b2/B1_26 ;
  wire  \inst_dob_mux_b2/B1_27 ;
  wire  \inst_dob_mux_b2/B1_28 ;
  wire  \inst_dob_mux_b2/B1_29 ;
  wire  \inst_dob_mux_b2/B1_3 ;
  wire  \inst_dob_mux_b2/B1_30 ;
  wire  \inst_dob_mux_b2/B1_31 ;
  wire  \inst_dob_mux_b2/B1_4 ;
  wire  \inst_dob_mux_b2/B1_5 ;
  wire  \inst_dob_mux_b2/B1_6 ;
  wire  \inst_dob_mux_b2/B1_7 ;
  wire  \inst_dob_mux_b2/B1_8 ;
  wire  \inst_dob_mux_b2/B1_9 ;
  wire  \inst_dob_mux_b2/B2_0 ;
  wire  \inst_dob_mux_b2/B2_1 ;
  wire  \inst_dob_mux_b2/B2_10 ;
  wire  \inst_dob_mux_b2/B2_11 ;
  wire  \inst_dob_mux_b2/B2_12 ;
  wire  \inst_dob_mux_b2/B2_13 ;
  wire  \inst_dob_mux_b2/B2_14 ;
  wire  \inst_dob_mux_b2/B2_15 ;
  wire  \inst_dob_mux_b2/B2_2 ;
  wire  \inst_dob_mux_b2/B2_3 ;
  wire  \inst_dob_mux_b2/B2_4 ;
  wire  \inst_dob_mux_b2/B2_5 ;
  wire  \inst_dob_mux_b2/B2_6 ;
  wire  \inst_dob_mux_b2/B2_7 ;
  wire  \inst_dob_mux_b2/B2_8 ;
  wire  \inst_dob_mux_b2/B2_9 ;
  wire  \inst_dob_mux_b2/B3_0 ;
  wire  \inst_dob_mux_b2/B3_1 ;
  wire  \inst_dob_mux_b2/B3_2 ;
  wire  \inst_dob_mux_b2/B3_3 ;
  wire  \inst_dob_mux_b2/B3_4 ;
  wire  \inst_dob_mux_b2/B3_5 ;
  wire  \inst_dob_mux_b2/B3_6 ;
  wire  \inst_dob_mux_b2/B3_7 ;
  wire  \inst_dob_mux_b2/B4_0 ;
  wire  \inst_dob_mux_b2/B4_1 ;
  wire  \inst_dob_mux_b2/B4_2 ;
  wire  \inst_dob_mux_b2/B4_3 ;
  wire  \inst_dob_mux_b2/B5_0 ;
  wire  \inst_dob_mux_b2/B5_1 ;
  wire  \inst_dob_mux_b3/B0_0 ;
  wire  \inst_dob_mux_b3/B0_1 ;
  wire  \inst_dob_mux_b3/B0_10 ;
  wire  \inst_dob_mux_b3/B0_11 ;
  wire  \inst_dob_mux_b3/B0_12 ;
  wire  \inst_dob_mux_b3/B0_13 ;
  wire  \inst_dob_mux_b3/B0_14 ;
  wire  \inst_dob_mux_b3/B0_15 ;
  wire  \inst_dob_mux_b3/B0_16 ;
  wire  \inst_dob_mux_b3/B0_17 ;
  wire  \inst_dob_mux_b3/B0_18 ;
  wire  \inst_dob_mux_b3/B0_19 ;
  wire  \inst_dob_mux_b3/B0_2 ;
  wire  \inst_dob_mux_b3/B0_20 ;
  wire  \inst_dob_mux_b3/B0_21 ;
  wire  \inst_dob_mux_b3/B0_22 ;
  wire  \inst_dob_mux_b3/B0_23 ;
  wire  \inst_dob_mux_b3/B0_24 ;
  wire  \inst_dob_mux_b3/B0_25 ;
  wire  \inst_dob_mux_b3/B0_26 ;
  wire  \inst_dob_mux_b3/B0_27 ;
  wire  \inst_dob_mux_b3/B0_28 ;
  wire  \inst_dob_mux_b3/B0_29 ;
  wire  \inst_dob_mux_b3/B0_3 ;
  wire  \inst_dob_mux_b3/B0_30 ;
  wire  \inst_dob_mux_b3/B0_31 ;
  wire  \inst_dob_mux_b3/B0_32 ;
  wire  \inst_dob_mux_b3/B0_33 ;
  wire  \inst_dob_mux_b3/B0_34 ;
  wire  \inst_dob_mux_b3/B0_35 ;
  wire  \inst_dob_mux_b3/B0_36 ;
  wire  \inst_dob_mux_b3/B0_37 ;
  wire  \inst_dob_mux_b3/B0_38 ;
  wire  \inst_dob_mux_b3/B0_39 ;
  wire  \inst_dob_mux_b3/B0_4 ;
  wire  \inst_dob_mux_b3/B0_40 ;
  wire  \inst_dob_mux_b3/B0_41 ;
  wire  \inst_dob_mux_b3/B0_42 ;
  wire  \inst_dob_mux_b3/B0_43 ;
  wire  \inst_dob_mux_b3/B0_44 ;
  wire  \inst_dob_mux_b3/B0_45 ;
  wire  \inst_dob_mux_b3/B0_46 ;
  wire  \inst_dob_mux_b3/B0_47 ;
  wire  \inst_dob_mux_b3/B0_48 ;
  wire  \inst_dob_mux_b3/B0_49 ;
  wire  \inst_dob_mux_b3/B0_5 ;
  wire  \inst_dob_mux_b3/B0_50 ;
  wire  \inst_dob_mux_b3/B0_51 ;
  wire  \inst_dob_mux_b3/B0_52 ;
  wire  \inst_dob_mux_b3/B0_53 ;
  wire  \inst_dob_mux_b3/B0_54 ;
  wire  \inst_dob_mux_b3/B0_55 ;
  wire  \inst_dob_mux_b3/B0_56 ;
  wire  \inst_dob_mux_b3/B0_57 ;
  wire  \inst_dob_mux_b3/B0_58 ;
  wire  \inst_dob_mux_b3/B0_59 ;
  wire  \inst_dob_mux_b3/B0_6 ;
  wire  \inst_dob_mux_b3/B0_60 ;
  wire  \inst_dob_mux_b3/B0_61 ;
  wire  \inst_dob_mux_b3/B0_62 ;
  wire  \inst_dob_mux_b3/B0_63 ;
  wire  \inst_dob_mux_b3/B0_7 ;
  wire  \inst_dob_mux_b3/B0_8 ;
  wire  \inst_dob_mux_b3/B0_9 ;
  wire  \inst_dob_mux_b3/B1_0 ;
  wire  \inst_dob_mux_b3/B1_1 ;
  wire  \inst_dob_mux_b3/B1_10 ;
  wire  \inst_dob_mux_b3/B1_11 ;
  wire  \inst_dob_mux_b3/B1_12 ;
  wire  \inst_dob_mux_b3/B1_13 ;
  wire  \inst_dob_mux_b3/B1_14 ;
  wire  \inst_dob_mux_b3/B1_15 ;
  wire  \inst_dob_mux_b3/B1_16 ;
  wire  \inst_dob_mux_b3/B1_17 ;
  wire  \inst_dob_mux_b3/B1_18 ;
  wire  \inst_dob_mux_b3/B1_19 ;
  wire  \inst_dob_mux_b3/B1_2 ;
  wire  \inst_dob_mux_b3/B1_20 ;
  wire  \inst_dob_mux_b3/B1_21 ;
  wire  \inst_dob_mux_b3/B1_22 ;
  wire  \inst_dob_mux_b3/B1_23 ;
  wire  \inst_dob_mux_b3/B1_24 ;
  wire  \inst_dob_mux_b3/B1_25 ;
  wire  \inst_dob_mux_b3/B1_26 ;
  wire  \inst_dob_mux_b3/B1_27 ;
  wire  \inst_dob_mux_b3/B1_28 ;
  wire  \inst_dob_mux_b3/B1_29 ;
  wire  \inst_dob_mux_b3/B1_3 ;
  wire  \inst_dob_mux_b3/B1_30 ;
  wire  \inst_dob_mux_b3/B1_31 ;
  wire  \inst_dob_mux_b3/B1_4 ;
  wire  \inst_dob_mux_b3/B1_5 ;
  wire  \inst_dob_mux_b3/B1_6 ;
  wire  \inst_dob_mux_b3/B1_7 ;
  wire  \inst_dob_mux_b3/B1_8 ;
  wire  \inst_dob_mux_b3/B1_9 ;
  wire  \inst_dob_mux_b3/B2_0 ;
  wire  \inst_dob_mux_b3/B2_1 ;
  wire  \inst_dob_mux_b3/B2_10 ;
  wire  \inst_dob_mux_b3/B2_11 ;
  wire  \inst_dob_mux_b3/B2_12 ;
  wire  \inst_dob_mux_b3/B2_13 ;
  wire  \inst_dob_mux_b3/B2_14 ;
  wire  \inst_dob_mux_b3/B2_15 ;
  wire  \inst_dob_mux_b3/B2_2 ;
  wire  \inst_dob_mux_b3/B2_3 ;
  wire  \inst_dob_mux_b3/B2_4 ;
  wire  \inst_dob_mux_b3/B2_5 ;
  wire  \inst_dob_mux_b3/B2_6 ;
  wire  \inst_dob_mux_b3/B2_7 ;
  wire  \inst_dob_mux_b3/B2_8 ;
  wire  \inst_dob_mux_b3/B2_9 ;
  wire  \inst_dob_mux_b3/B3_0 ;
  wire  \inst_dob_mux_b3/B3_1 ;
  wire  \inst_dob_mux_b3/B3_2 ;
  wire  \inst_dob_mux_b3/B3_3 ;
  wire  \inst_dob_mux_b3/B3_4 ;
  wire  \inst_dob_mux_b3/B3_5 ;
  wire  \inst_dob_mux_b3/B3_6 ;
  wire  \inst_dob_mux_b3/B3_7 ;
  wire  \inst_dob_mux_b3/B4_0 ;
  wire  \inst_dob_mux_b3/B4_1 ;
  wire  \inst_dob_mux_b3/B4_2 ;
  wire  \inst_dob_mux_b3/B4_3 ;
  wire  \inst_dob_mux_b3/B5_0 ;
  wire  \inst_dob_mux_b3/B5_1 ;
  wire  \inst_dob_mux_b4/B0_0 ;
  wire  \inst_dob_mux_b4/B0_1 ;
  wire  \inst_dob_mux_b4/B0_10 ;
  wire  \inst_dob_mux_b4/B0_11 ;
  wire  \inst_dob_mux_b4/B0_12 ;
  wire  \inst_dob_mux_b4/B0_13 ;
  wire  \inst_dob_mux_b4/B0_14 ;
  wire  \inst_dob_mux_b4/B0_15 ;
  wire  \inst_dob_mux_b4/B0_16 ;
  wire  \inst_dob_mux_b4/B0_17 ;
  wire  \inst_dob_mux_b4/B0_18 ;
  wire  \inst_dob_mux_b4/B0_19 ;
  wire  \inst_dob_mux_b4/B0_2 ;
  wire  \inst_dob_mux_b4/B0_20 ;
  wire  \inst_dob_mux_b4/B0_21 ;
  wire  \inst_dob_mux_b4/B0_22 ;
  wire  \inst_dob_mux_b4/B0_23 ;
  wire  \inst_dob_mux_b4/B0_24 ;
  wire  \inst_dob_mux_b4/B0_25 ;
  wire  \inst_dob_mux_b4/B0_26 ;
  wire  \inst_dob_mux_b4/B0_27 ;
  wire  \inst_dob_mux_b4/B0_28 ;
  wire  \inst_dob_mux_b4/B0_29 ;
  wire  \inst_dob_mux_b4/B0_3 ;
  wire  \inst_dob_mux_b4/B0_30 ;
  wire  \inst_dob_mux_b4/B0_31 ;
  wire  \inst_dob_mux_b4/B0_32 ;
  wire  \inst_dob_mux_b4/B0_33 ;
  wire  \inst_dob_mux_b4/B0_34 ;
  wire  \inst_dob_mux_b4/B0_35 ;
  wire  \inst_dob_mux_b4/B0_36 ;
  wire  \inst_dob_mux_b4/B0_37 ;
  wire  \inst_dob_mux_b4/B0_38 ;
  wire  \inst_dob_mux_b4/B0_39 ;
  wire  \inst_dob_mux_b4/B0_4 ;
  wire  \inst_dob_mux_b4/B0_40 ;
  wire  \inst_dob_mux_b4/B0_41 ;
  wire  \inst_dob_mux_b4/B0_42 ;
  wire  \inst_dob_mux_b4/B0_43 ;
  wire  \inst_dob_mux_b4/B0_44 ;
  wire  \inst_dob_mux_b4/B0_45 ;
  wire  \inst_dob_mux_b4/B0_46 ;
  wire  \inst_dob_mux_b4/B0_47 ;
  wire  \inst_dob_mux_b4/B0_48 ;
  wire  \inst_dob_mux_b4/B0_49 ;
  wire  \inst_dob_mux_b4/B0_5 ;
  wire  \inst_dob_mux_b4/B0_50 ;
  wire  \inst_dob_mux_b4/B0_51 ;
  wire  \inst_dob_mux_b4/B0_52 ;
  wire  \inst_dob_mux_b4/B0_53 ;
  wire  \inst_dob_mux_b4/B0_54 ;
  wire  \inst_dob_mux_b4/B0_55 ;
  wire  \inst_dob_mux_b4/B0_56 ;
  wire  \inst_dob_mux_b4/B0_57 ;
  wire  \inst_dob_mux_b4/B0_58 ;
  wire  \inst_dob_mux_b4/B0_59 ;
  wire  \inst_dob_mux_b4/B0_6 ;
  wire  \inst_dob_mux_b4/B0_60 ;
  wire  \inst_dob_mux_b4/B0_61 ;
  wire  \inst_dob_mux_b4/B0_62 ;
  wire  \inst_dob_mux_b4/B0_63 ;
  wire  \inst_dob_mux_b4/B0_7 ;
  wire  \inst_dob_mux_b4/B0_8 ;
  wire  \inst_dob_mux_b4/B0_9 ;
  wire  \inst_dob_mux_b4/B1_0 ;
  wire  \inst_dob_mux_b4/B1_1 ;
  wire  \inst_dob_mux_b4/B1_10 ;
  wire  \inst_dob_mux_b4/B1_11 ;
  wire  \inst_dob_mux_b4/B1_12 ;
  wire  \inst_dob_mux_b4/B1_13 ;
  wire  \inst_dob_mux_b4/B1_14 ;
  wire  \inst_dob_mux_b4/B1_15 ;
  wire  \inst_dob_mux_b4/B1_16 ;
  wire  \inst_dob_mux_b4/B1_17 ;
  wire  \inst_dob_mux_b4/B1_18 ;
  wire  \inst_dob_mux_b4/B1_19 ;
  wire  \inst_dob_mux_b4/B1_2 ;
  wire  \inst_dob_mux_b4/B1_20 ;
  wire  \inst_dob_mux_b4/B1_21 ;
  wire  \inst_dob_mux_b4/B1_22 ;
  wire  \inst_dob_mux_b4/B1_23 ;
  wire  \inst_dob_mux_b4/B1_24 ;
  wire  \inst_dob_mux_b4/B1_25 ;
  wire  \inst_dob_mux_b4/B1_26 ;
  wire  \inst_dob_mux_b4/B1_27 ;
  wire  \inst_dob_mux_b4/B1_28 ;
  wire  \inst_dob_mux_b4/B1_29 ;
  wire  \inst_dob_mux_b4/B1_3 ;
  wire  \inst_dob_mux_b4/B1_30 ;
  wire  \inst_dob_mux_b4/B1_31 ;
  wire  \inst_dob_mux_b4/B1_4 ;
  wire  \inst_dob_mux_b4/B1_5 ;
  wire  \inst_dob_mux_b4/B1_6 ;
  wire  \inst_dob_mux_b4/B1_7 ;
  wire  \inst_dob_mux_b4/B1_8 ;
  wire  \inst_dob_mux_b4/B1_9 ;
  wire  \inst_dob_mux_b4/B2_0 ;
  wire  \inst_dob_mux_b4/B2_1 ;
  wire  \inst_dob_mux_b4/B2_10 ;
  wire  \inst_dob_mux_b4/B2_11 ;
  wire  \inst_dob_mux_b4/B2_12 ;
  wire  \inst_dob_mux_b4/B2_13 ;
  wire  \inst_dob_mux_b4/B2_14 ;
  wire  \inst_dob_mux_b4/B2_15 ;
  wire  \inst_dob_mux_b4/B2_2 ;
  wire  \inst_dob_mux_b4/B2_3 ;
  wire  \inst_dob_mux_b4/B2_4 ;
  wire  \inst_dob_mux_b4/B2_5 ;
  wire  \inst_dob_mux_b4/B2_6 ;
  wire  \inst_dob_mux_b4/B2_7 ;
  wire  \inst_dob_mux_b4/B2_8 ;
  wire  \inst_dob_mux_b4/B2_9 ;
  wire  \inst_dob_mux_b4/B3_0 ;
  wire  \inst_dob_mux_b4/B3_1 ;
  wire  \inst_dob_mux_b4/B3_2 ;
  wire  \inst_dob_mux_b4/B3_3 ;
  wire  \inst_dob_mux_b4/B3_4 ;
  wire  \inst_dob_mux_b4/B3_5 ;
  wire  \inst_dob_mux_b4/B3_6 ;
  wire  \inst_dob_mux_b4/B3_7 ;
  wire  \inst_dob_mux_b4/B4_0 ;
  wire  \inst_dob_mux_b4/B4_1 ;
  wire  \inst_dob_mux_b4/B4_2 ;
  wire  \inst_dob_mux_b4/B4_3 ;
  wire  \inst_dob_mux_b4/B5_0 ;
  wire  \inst_dob_mux_b4/B5_1 ;
  wire  \inst_dob_mux_b5/B0_0 ;
  wire  \inst_dob_mux_b5/B0_1 ;
  wire  \inst_dob_mux_b5/B0_10 ;
  wire  \inst_dob_mux_b5/B0_11 ;
  wire  \inst_dob_mux_b5/B0_12 ;
  wire  \inst_dob_mux_b5/B0_13 ;
  wire  \inst_dob_mux_b5/B0_14 ;
  wire  \inst_dob_mux_b5/B0_15 ;
  wire  \inst_dob_mux_b5/B0_16 ;
  wire  \inst_dob_mux_b5/B0_17 ;
  wire  \inst_dob_mux_b5/B0_18 ;
  wire  \inst_dob_mux_b5/B0_19 ;
  wire  \inst_dob_mux_b5/B0_2 ;
  wire  \inst_dob_mux_b5/B0_20 ;
  wire  \inst_dob_mux_b5/B0_21 ;
  wire  \inst_dob_mux_b5/B0_22 ;
  wire  \inst_dob_mux_b5/B0_23 ;
  wire  \inst_dob_mux_b5/B0_24 ;
  wire  \inst_dob_mux_b5/B0_25 ;
  wire  \inst_dob_mux_b5/B0_26 ;
  wire  \inst_dob_mux_b5/B0_27 ;
  wire  \inst_dob_mux_b5/B0_28 ;
  wire  \inst_dob_mux_b5/B0_29 ;
  wire  \inst_dob_mux_b5/B0_3 ;
  wire  \inst_dob_mux_b5/B0_30 ;
  wire  \inst_dob_mux_b5/B0_31 ;
  wire  \inst_dob_mux_b5/B0_32 ;
  wire  \inst_dob_mux_b5/B0_33 ;
  wire  \inst_dob_mux_b5/B0_34 ;
  wire  \inst_dob_mux_b5/B0_35 ;
  wire  \inst_dob_mux_b5/B0_36 ;
  wire  \inst_dob_mux_b5/B0_37 ;
  wire  \inst_dob_mux_b5/B0_38 ;
  wire  \inst_dob_mux_b5/B0_39 ;
  wire  \inst_dob_mux_b5/B0_4 ;
  wire  \inst_dob_mux_b5/B0_40 ;
  wire  \inst_dob_mux_b5/B0_41 ;
  wire  \inst_dob_mux_b5/B0_42 ;
  wire  \inst_dob_mux_b5/B0_43 ;
  wire  \inst_dob_mux_b5/B0_44 ;
  wire  \inst_dob_mux_b5/B0_45 ;
  wire  \inst_dob_mux_b5/B0_46 ;
  wire  \inst_dob_mux_b5/B0_47 ;
  wire  \inst_dob_mux_b5/B0_48 ;
  wire  \inst_dob_mux_b5/B0_49 ;
  wire  \inst_dob_mux_b5/B0_5 ;
  wire  \inst_dob_mux_b5/B0_50 ;
  wire  \inst_dob_mux_b5/B0_51 ;
  wire  \inst_dob_mux_b5/B0_52 ;
  wire  \inst_dob_mux_b5/B0_53 ;
  wire  \inst_dob_mux_b5/B0_54 ;
  wire  \inst_dob_mux_b5/B0_55 ;
  wire  \inst_dob_mux_b5/B0_56 ;
  wire  \inst_dob_mux_b5/B0_57 ;
  wire  \inst_dob_mux_b5/B0_58 ;
  wire  \inst_dob_mux_b5/B0_59 ;
  wire  \inst_dob_mux_b5/B0_6 ;
  wire  \inst_dob_mux_b5/B0_60 ;
  wire  \inst_dob_mux_b5/B0_61 ;
  wire  \inst_dob_mux_b5/B0_62 ;
  wire  \inst_dob_mux_b5/B0_63 ;
  wire  \inst_dob_mux_b5/B0_7 ;
  wire  \inst_dob_mux_b5/B0_8 ;
  wire  \inst_dob_mux_b5/B0_9 ;
  wire  \inst_dob_mux_b5/B1_0 ;
  wire  \inst_dob_mux_b5/B1_1 ;
  wire  \inst_dob_mux_b5/B1_10 ;
  wire  \inst_dob_mux_b5/B1_11 ;
  wire  \inst_dob_mux_b5/B1_12 ;
  wire  \inst_dob_mux_b5/B1_13 ;
  wire  \inst_dob_mux_b5/B1_14 ;
  wire  \inst_dob_mux_b5/B1_15 ;
  wire  \inst_dob_mux_b5/B1_16 ;
  wire  \inst_dob_mux_b5/B1_17 ;
  wire  \inst_dob_mux_b5/B1_18 ;
  wire  \inst_dob_mux_b5/B1_19 ;
  wire  \inst_dob_mux_b5/B1_2 ;
  wire  \inst_dob_mux_b5/B1_20 ;
  wire  \inst_dob_mux_b5/B1_21 ;
  wire  \inst_dob_mux_b5/B1_22 ;
  wire  \inst_dob_mux_b5/B1_23 ;
  wire  \inst_dob_mux_b5/B1_24 ;
  wire  \inst_dob_mux_b5/B1_25 ;
  wire  \inst_dob_mux_b5/B1_26 ;
  wire  \inst_dob_mux_b5/B1_27 ;
  wire  \inst_dob_mux_b5/B1_28 ;
  wire  \inst_dob_mux_b5/B1_29 ;
  wire  \inst_dob_mux_b5/B1_3 ;
  wire  \inst_dob_mux_b5/B1_30 ;
  wire  \inst_dob_mux_b5/B1_31 ;
  wire  \inst_dob_mux_b5/B1_4 ;
  wire  \inst_dob_mux_b5/B1_5 ;
  wire  \inst_dob_mux_b5/B1_6 ;
  wire  \inst_dob_mux_b5/B1_7 ;
  wire  \inst_dob_mux_b5/B1_8 ;
  wire  \inst_dob_mux_b5/B1_9 ;
  wire  \inst_dob_mux_b5/B2_0 ;
  wire  \inst_dob_mux_b5/B2_1 ;
  wire  \inst_dob_mux_b5/B2_10 ;
  wire  \inst_dob_mux_b5/B2_11 ;
  wire  \inst_dob_mux_b5/B2_12 ;
  wire  \inst_dob_mux_b5/B2_13 ;
  wire  \inst_dob_mux_b5/B2_14 ;
  wire  \inst_dob_mux_b5/B2_15 ;
  wire  \inst_dob_mux_b5/B2_2 ;
  wire  \inst_dob_mux_b5/B2_3 ;
  wire  \inst_dob_mux_b5/B2_4 ;
  wire  \inst_dob_mux_b5/B2_5 ;
  wire  \inst_dob_mux_b5/B2_6 ;
  wire  \inst_dob_mux_b5/B2_7 ;
  wire  \inst_dob_mux_b5/B2_8 ;
  wire  \inst_dob_mux_b5/B2_9 ;
  wire  \inst_dob_mux_b5/B3_0 ;
  wire  \inst_dob_mux_b5/B3_1 ;
  wire  \inst_dob_mux_b5/B3_2 ;
  wire  \inst_dob_mux_b5/B3_3 ;
  wire  \inst_dob_mux_b5/B3_4 ;
  wire  \inst_dob_mux_b5/B3_5 ;
  wire  \inst_dob_mux_b5/B3_6 ;
  wire  \inst_dob_mux_b5/B3_7 ;
  wire  \inst_dob_mux_b5/B4_0 ;
  wire  \inst_dob_mux_b5/B4_1 ;
  wire  \inst_dob_mux_b5/B4_2 ;
  wire  \inst_dob_mux_b5/B4_3 ;
  wire  \inst_dob_mux_b5/B5_0 ;
  wire  \inst_dob_mux_b5/B5_1 ;
  wire  \inst_dob_mux_b6/B0_0 ;
  wire  \inst_dob_mux_b6/B0_1 ;
  wire  \inst_dob_mux_b6/B0_10 ;
  wire  \inst_dob_mux_b6/B0_11 ;
  wire  \inst_dob_mux_b6/B0_12 ;
  wire  \inst_dob_mux_b6/B0_13 ;
  wire  \inst_dob_mux_b6/B0_14 ;
  wire  \inst_dob_mux_b6/B0_15 ;
  wire  \inst_dob_mux_b6/B0_16 ;
  wire  \inst_dob_mux_b6/B0_17 ;
  wire  \inst_dob_mux_b6/B0_18 ;
  wire  \inst_dob_mux_b6/B0_19 ;
  wire  \inst_dob_mux_b6/B0_2 ;
  wire  \inst_dob_mux_b6/B0_20 ;
  wire  \inst_dob_mux_b6/B0_21 ;
  wire  \inst_dob_mux_b6/B0_22 ;
  wire  \inst_dob_mux_b6/B0_23 ;
  wire  \inst_dob_mux_b6/B0_24 ;
  wire  \inst_dob_mux_b6/B0_25 ;
  wire  \inst_dob_mux_b6/B0_26 ;
  wire  \inst_dob_mux_b6/B0_27 ;
  wire  \inst_dob_mux_b6/B0_28 ;
  wire  \inst_dob_mux_b6/B0_29 ;
  wire  \inst_dob_mux_b6/B0_3 ;
  wire  \inst_dob_mux_b6/B0_30 ;
  wire  \inst_dob_mux_b6/B0_31 ;
  wire  \inst_dob_mux_b6/B0_32 ;
  wire  \inst_dob_mux_b6/B0_33 ;
  wire  \inst_dob_mux_b6/B0_34 ;
  wire  \inst_dob_mux_b6/B0_35 ;
  wire  \inst_dob_mux_b6/B0_36 ;
  wire  \inst_dob_mux_b6/B0_37 ;
  wire  \inst_dob_mux_b6/B0_38 ;
  wire  \inst_dob_mux_b6/B0_39 ;
  wire  \inst_dob_mux_b6/B0_4 ;
  wire  \inst_dob_mux_b6/B0_40 ;
  wire  \inst_dob_mux_b6/B0_41 ;
  wire  \inst_dob_mux_b6/B0_42 ;
  wire  \inst_dob_mux_b6/B0_43 ;
  wire  \inst_dob_mux_b6/B0_44 ;
  wire  \inst_dob_mux_b6/B0_45 ;
  wire  \inst_dob_mux_b6/B0_46 ;
  wire  \inst_dob_mux_b6/B0_47 ;
  wire  \inst_dob_mux_b6/B0_48 ;
  wire  \inst_dob_mux_b6/B0_49 ;
  wire  \inst_dob_mux_b6/B0_5 ;
  wire  \inst_dob_mux_b6/B0_50 ;
  wire  \inst_dob_mux_b6/B0_51 ;
  wire  \inst_dob_mux_b6/B0_52 ;
  wire  \inst_dob_mux_b6/B0_53 ;
  wire  \inst_dob_mux_b6/B0_54 ;
  wire  \inst_dob_mux_b6/B0_55 ;
  wire  \inst_dob_mux_b6/B0_56 ;
  wire  \inst_dob_mux_b6/B0_57 ;
  wire  \inst_dob_mux_b6/B0_58 ;
  wire  \inst_dob_mux_b6/B0_59 ;
  wire  \inst_dob_mux_b6/B0_6 ;
  wire  \inst_dob_mux_b6/B0_60 ;
  wire  \inst_dob_mux_b6/B0_61 ;
  wire  \inst_dob_mux_b6/B0_62 ;
  wire  \inst_dob_mux_b6/B0_63 ;
  wire  \inst_dob_mux_b6/B0_7 ;
  wire  \inst_dob_mux_b6/B0_8 ;
  wire  \inst_dob_mux_b6/B0_9 ;
  wire  \inst_dob_mux_b6/B1_0 ;
  wire  \inst_dob_mux_b6/B1_1 ;
  wire  \inst_dob_mux_b6/B1_10 ;
  wire  \inst_dob_mux_b6/B1_11 ;
  wire  \inst_dob_mux_b6/B1_12 ;
  wire  \inst_dob_mux_b6/B1_13 ;
  wire  \inst_dob_mux_b6/B1_14 ;
  wire  \inst_dob_mux_b6/B1_15 ;
  wire  \inst_dob_mux_b6/B1_16 ;
  wire  \inst_dob_mux_b6/B1_17 ;
  wire  \inst_dob_mux_b6/B1_18 ;
  wire  \inst_dob_mux_b6/B1_19 ;
  wire  \inst_dob_mux_b6/B1_2 ;
  wire  \inst_dob_mux_b6/B1_20 ;
  wire  \inst_dob_mux_b6/B1_21 ;
  wire  \inst_dob_mux_b6/B1_22 ;
  wire  \inst_dob_mux_b6/B1_23 ;
  wire  \inst_dob_mux_b6/B1_24 ;
  wire  \inst_dob_mux_b6/B1_25 ;
  wire  \inst_dob_mux_b6/B1_26 ;
  wire  \inst_dob_mux_b6/B1_27 ;
  wire  \inst_dob_mux_b6/B1_28 ;
  wire  \inst_dob_mux_b6/B1_29 ;
  wire  \inst_dob_mux_b6/B1_3 ;
  wire  \inst_dob_mux_b6/B1_30 ;
  wire  \inst_dob_mux_b6/B1_31 ;
  wire  \inst_dob_mux_b6/B1_4 ;
  wire  \inst_dob_mux_b6/B1_5 ;
  wire  \inst_dob_mux_b6/B1_6 ;
  wire  \inst_dob_mux_b6/B1_7 ;
  wire  \inst_dob_mux_b6/B1_8 ;
  wire  \inst_dob_mux_b6/B1_9 ;
  wire  \inst_dob_mux_b6/B2_0 ;
  wire  \inst_dob_mux_b6/B2_1 ;
  wire  \inst_dob_mux_b6/B2_10 ;
  wire  \inst_dob_mux_b6/B2_11 ;
  wire  \inst_dob_mux_b6/B2_12 ;
  wire  \inst_dob_mux_b6/B2_13 ;
  wire  \inst_dob_mux_b6/B2_14 ;
  wire  \inst_dob_mux_b6/B2_15 ;
  wire  \inst_dob_mux_b6/B2_2 ;
  wire  \inst_dob_mux_b6/B2_3 ;
  wire  \inst_dob_mux_b6/B2_4 ;
  wire  \inst_dob_mux_b6/B2_5 ;
  wire  \inst_dob_mux_b6/B2_6 ;
  wire  \inst_dob_mux_b6/B2_7 ;
  wire  \inst_dob_mux_b6/B2_8 ;
  wire  \inst_dob_mux_b6/B2_9 ;
  wire  \inst_dob_mux_b6/B3_0 ;
  wire  \inst_dob_mux_b6/B3_1 ;
  wire  \inst_dob_mux_b6/B3_2 ;
  wire  \inst_dob_mux_b6/B3_3 ;
  wire  \inst_dob_mux_b6/B3_4 ;
  wire  \inst_dob_mux_b6/B3_5 ;
  wire  \inst_dob_mux_b6/B3_6 ;
  wire  \inst_dob_mux_b6/B3_7 ;
  wire  \inst_dob_mux_b6/B4_0 ;
  wire  \inst_dob_mux_b6/B4_1 ;
  wire  \inst_dob_mux_b6/B4_2 ;
  wire  \inst_dob_mux_b6/B4_3 ;
  wire  \inst_dob_mux_b6/B5_0 ;
  wire  \inst_dob_mux_b6/B5_1 ;
  wire  \inst_dob_mux_b7/B0_0 ;
  wire  \inst_dob_mux_b7/B0_1 ;
  wire  \inst_dob_mux_b7/B0_10 ;
  wire  \inst_dob_mux_b7/B0_11 ;
  wire  \inst_dob_mux_b7/B0_12 ;
  wire  \inst_dob_mux_b7/B0_13 ;
  wire  \inst_dob_mux_b7/B0_14 ;
  wire  \inst_dob_mux_b7/B0_15 ;
  wire  \inst_dob_mux_b7/B0_16 ;
  wire  \inst_dob_mux_b7/B0_17 ;
  wire  \inst_dob_mux_b7/B0_18 ;
  wire  \inst_dob_mux_b7/B0_19 ;
  wire  \inst_dob_mux_b7/B0_2 ;
  wire  \inst_dob_mux_b7/B0_20 ;
  wire  \inst_dob_mux_b7/B0_21 ;
  wire  \inst_dob_mux_b7/B0_22 ;
  wire  \inst_dob_mux_b7/B0_23 ;
  wire  \inst_dob_mux_b7/B0_24 ;
  wire  \inst_dob_mux_b7/B0_25 ;
  wire  \inst_dob_mux_b7/B0_26 ;
  wire  \inst_dob_mux_b7/B0_27 ;
  wire  \inst_dob_mux_b7/B0_28 ;
  wire  \inst_dob_mux_b7/B0_29 ;
  wire  \inst_dob_mux_b7/B0_3 ;
  wire  \inst_dob_mux_b7/B0_30 ;
  wire  \inst_dob_mux_b7/B0_31 ;
  wire  \inst_dob_mux_b7/B0_32 ;
  wire  \inst_dob_mux_b7/B0_33 ;
  wire  \inst_dob_mux_b7/B0_34 ;
  wire  \inst_dob_mux_b7/B0_35 ;
  wire  \inst_dob_mux_b7/B0_36 ;
  wire  \inst_dob_mux_b7/B0_37 ;
  wire  \inst_dob_mux_b7/B0_38 ;
  wire  \inst_dob_mux_b7/B0_39 ;
  wire  \inst_dob_mux_b7/B0_4 ;
  wire  \inst_dob_mux_b7/B0_40 ;
  wire  \inst_dob_mux_b7/B0_41 ;
  wire  \inst_dob_mux_b7/B0_42 ;
  wire  \inst_dob_mux_b7/B0_43 ;
  wire  \inst_dob_mux_b7/B0_44 ;
  wire  \inst_dob_mux_b7/B0_45 ;
  wire  \inst_dob_mux_b7/B0_46 ;
  wire  \inst_dob_mux_b7/B0_47 ;
  wire  \inst_dob_mux_b7/B0_48 ;
  wire  \inst_dob_mux_b7/B0_49 ;
  wire  \inst_dob_mux_b7/B0_5 ;
  wire  \inst_dob_mux_b7/B0_50 ;
  wire  \inst_dob_mux_b7/B0_51 ;
  wire  \inst_dob_mux_b7/B0_52 ;
  wire  \inst_dob_mux_b7/B0_53 ;
  wire  \inst_dob_mux_b7/B0_54 ;
  wire  \inst_dob_mux_b7/B0_55 ;
  wire  \inst_dob_mux_b7/B0_56 ;
  wire  \inst_dob_mux_b7/B0_57 ;
  wire  \inst_dob_mux_b7/B0_58 ;
  wire  \inst_dob_mux_b7/B0_59 ;
  wire  \inst_dob_mux_b7/B0_6 ;
  wire  \inst_dob_mux_b7/B0_60 ;
  wire  \inst_dob_mux_b7/B0_61 ;
  wire  \inst_dob_mux_b7/B0_62 ;
  wire  \inst_dob_mux_b7/B0_63 ;
  wire  \inst_dob_mux_b7/B0_7 ;
  wire  \inst_dob_mux_b7/B0_8 ;
  wire  \inst_dob_mux_b7/B0_9 ;
  wire  \inst_dob_mux_b7/B1_0 ;
  wire  \inst_dob_mux_b7/B1_1 ;
  wire  \inst_dob_mux_b7/B1_10 ;
  wire  \inst_dob_mux_b7/B1_11 ;
  wire  \inst_dob_mux_b7/B1_12 ;
  wire  \inst_dob_mux_b7/B1_13 ;
  wire  \inst_dob_mux_b7/B1_14 ;
  wire  \inst_dob_mux_b7/B1_15 ;
  wire  \inst_dob_mux_b7/B1_16 ;
  wire  \inst_dob_mux_b7/B1_17 ;
  wire  \inst_dob_mux_b7/B1_18 ;
  wire  \inst_dob_mux_b7/B1_19 ;
  wire  \inst_dob_mux_b7/B1_2 ;
  wire  \inst_dob_mux_b7/B1_20 ;
  wire  \inst_dob_mux_b7/B1_21 ;
  wire  \inst_dob_mux_b7/B1_22 ;
  wire  \inst_dob_mux_b7/B1_23 ;
  wire  \inst_dob_mux_b7/B1_24 ;
  wire  \inst_dob_mux_b7/B1_25 ;
  wire  \inst_dob_mux_b7/B1_26 ;
  wire  \inst_dob_mux_b7/B1_27 ;
  wire  \inst_dob_mux_b7/B1_28 ;
  wire  \inst_dob_mux_b7/B1_29 ;
  wire  \inst_dob_mux_b7/B1_3 ;
  wire  \inst_dob_mux_b7/B1_30 ;
  wire  \inst_dob_mux_b7/B1_31 ;
  wire  \inst_dob_mux_b7/B1_4 ;
  wire  \inst_dob_mux_b7/B1_5 ;
  wire  \inst_dob_mux_b7/B1_6 ;
  wire  \inst_dob_mux_b7/B1_7 ;
  wire  \inst_dob_mux_b7/B1_8 ;
  wire  \inst_dob_mux_b7/B1_9 ;
  wire  \inst_dob_mux_b7/B2_0 ;
  wire  \inst_dob_mux_b7/B2_1 ;
  wire  \inst_dob_mux_b7/B2_10 ;
  wire  \inst_dob_mux_b7/B2_11 ;
  wire  \inst_dob_mux_b7/B2_12 ;
  wire  \inst_dob_mux_b7/B2_13 ;
  wire  \inst_dob_mux_b7/B2_14 ;
  wire  \inst_dob_mux_b7/B2_15 ;
  wire  \inst_dob_mux_b7/B2_2 ;
  wire  \inst_dob_mux_b7/B2_3 ;
  wire  \inst_dob_mux_b7/B2_4 ;
  wire  \inst_dob_mux_b7/B2_5 ;
  wire  \inst_dob_mux_b7/B2_6 ;
  wire  \inst_dob_mux_b7/B2_7 ;
  wire  \inst_dob_mux_b7/B2_8 ;
  wire  \inst_dob_mux_b7/B2_9 ;
  wire  \inst_dob_mux_b7/B3_0 ;
  wire  \inst_dob_mux_b7/B3_1 ;
  wire  \inst_dob_mux_b7/B3_2 ;
  wire  \inst_dob_mux_b7/B3_3 ;
  wire  \inst_dob_mux_b7/B3_4 ;
  wire  \inst_dob_mux_b7/B3_5 ;
  wire  \inst_dob_mux_b7/B3_6 ;
  wire  \inst_dob_mux_b7/B3_7 ;
  wire  \inst_dob_mux_b7/B4_0 ;
  wire  \inst_dob_mux_b7/B4_1 ;
  wire  \inst_dob_mux_b7/B4_2 ;
  wire  \inst_dob_mux_b7/B4_3 ;
  wire  \inst_dob_mux_b7/B5_0 ;
  wire  \inst_dob_mux_b7/B5_1 ;
  wire  \inst_dob_mux_b8/B0_0 ;
  wire  \inst_dob_mux_b8/B0_1 ;
  wire  \inst_dob_mux_b8/B0_10 ;
  wire  \inst_dob_mux_b8/B0_11 ;
  wire  \inst_dob_mux_b8/B0_12 ;
  wire  \inst_dob_mux_b8/B0_13 ;
  wire  \inst_dob_mux_b8/B0_14 ;
  wire  \inst_dob_mux_b8/B0_15 ;
  wire  \inst_dob_mux_b8/B0_16 ;
  wire  \inst_dob_mux_b8/B0_17 ;
  wire  \inst_dob_mux_b8/B0_18 ;
  wire  \inst_dob_mux_b8/B0_19 ;
  wire  \inst_dob_mux_b8/B0_2 ;
  wire  \inst_dob_mux_b8/B0_20 ;
  wire  \inst_dob_mux_b8/B0_21 ;
  wire  \inst_dob_mux_b8/B0_22 ;
  wire  \inst_dob_mux_b8/B0_23 ;
  wire  \inst_dob_mux_b8/B0_24 ;
  wire  \inst_dob_mux_b8/B0_25 ;
  wire  \inst_dob_mux_b8/B0_26 ;
  wire  \inst_dob_mux_b8/B0_27 ;
  wire  \inst_dob_mux_b8/B0_28 ;
  wire  \inst_dob_mux_b8/B0_29 ;
  wire  \inst_dob_mux_b8/B0_3 ;
  wire  \inst_dob_mux_b8/B0_30 ;
  wire  \inst_dob_mux_b8/B0_31 ;
  wire  \inst_dob_mux_b8/B0_32 ;
  wire  \inst_dob_mux_b8/B0_33 ;
  wire  \inst_dob_mux_b8/B0_34 ;
  wire  \inst_dob_mux_b8/B0_35 ;
  wire  \inst_dob_mux_b8/B0_36 ;
  wire  \inst_dob_mux_b8/B0_37 ;
  wire  \inst_dob_mux_b8/B0_38 ;
  wire  \inst_dob_mux_b8/B0_39 ;
  wire  \inst_dob_mux_b8/B0_4 ;
  wire  \inst_dob_mux_b8/B0_40 ;
  wire  \inst_dob_mux_b8/B0_41 ;
  wire  \inst_dob_mux_b8/B0_42 ;
  wire  \inst_dob_mux_b8/B0_43 ;
  wire  \inst_dob_mux_b8/B0_44 ;
  wire  \inst_dob_mux_b8/B0_45 ;
  wire  \inst_dob_mux_b8/B0_46 ;
  wire  \inst_dob_mux_b8/B0_47 ;
  wire  \inst_dob_mux_b8/B0_48 ;
  wire  \inst_dob_mux_b8/B0_49 ;
  wire  \inst_dob_mux_b8/B0_5 ;
  wire  \inst_dob_mux_b8/B0_50 ;
  wire  \inst_dob_mux_b8/B0_51 ;
  wire  \inst_dob_mux_b8/B0_52 ;
  wire  \inst_dob_mux_b8/B0_53 ;
  wire  \inst_dob_mux_b8/B0_54 ;
  wire  \inst_dob_mux_b8/B0_55 ;
  wire  \inst_dob_mux_b8/B0_56 ;
  wire  \inst_dob_mux_b8/B0_57 ;
  wire  \inst_dob_mux_b8/B0_58 ;
  wire  \inst_dob_mux_b8/B0_59 ;
  wire  \inst_dob_mux_b8/B0_6 ;
  wire  \inst_dob_mux_b8/B0_60 ;
  wire  \inst_dob_mux_b8/B0_61 ;
  wire  \inst_dob_mux_b8/B0_62 ;
  wire  \inst_dob_mux_b8/B0_63 ;
  wire  \inst_dob_mux_b8/B0_7 ;
  wire  \inst_dob_mux_b8/B0_8 ;
  wire  \inst_dob_mux_b8/B0_9 ;
  wire  \inst_dob_mux_b8/B1_0 ;
  wire  \inst_dob_mux_b8/B1_1 ;
  wire  \inst_dob_mux_b8/B1_10 ;
  wire  \inst_dob_mux_b8/B1_11 ;
  wire  \inst_dob_mux_b8/B1_12 ;
  wire  \inst_dob_mux_b8/B1_13 ;
  wire  \inst_dob_mux_b8/B1_14 ;
  wire  \inst_dob_mux_b8/B1_15 ;
  wire  \inst_dob_mux_b8/B1_16 ;
  wire  \inst_dob_mux_b8/B1_17 ;
  wire  \inst_dob_mux_b8/B1_18 ;
  wire  \inst_dob_mux_b8/B1_19 ;
  wire  \inst_dob_mux_b8/B1_2 ;
  wire  \inst_dob_mux_b8/B1_20 ;
  wire  \inst_dob_mux_b8/B1_21 ;
  wire  \inst_dob_mux_b8/B1_22 ;
  wire  \inst_dob_mux_b8/B1_23 ;
  wire  \inst_dob_mux_b8/B1_24 ;
  wire  \inst_dob_mux_b8/B1_25 ;
  wire  \inst_dob_mux_b8/B1_26 ;
  wire  \inst_dob_mux_b8/B1_27 ;
  wire  \inst_dob_mux_b8/B1_28 ;
  wire  \inst_dob_mux_b8/B1_29 ;
  wire  \inst_dob_mux_b8/B1_3 ;
  wire  \inst_dob_mux_b8/B1_30 ;
  wire  \inst_dob_mux_b8/B1_31 ;
  wire  \inst_dob_mux_b8/B1_4 ;
  wire  \inst_dob_mux_b8/B1_5 ;
  wire  \inst_dob_mux_b8/B1_6 ;
  wire  \inst_dob_mux_b8/B1_7 ;
  wire  \inst_dob_mux_b8/B1_8 ;
  wire  \inst_dob_mux_b8/B1_9 ;
  wire  \inst_dob_mux_b8/B2_0 ;
  wire  \inst_dob_mux_b8/B2_1 ;
  wire  \inst_dob_mux_b8/B2_10 ;
  wire  \inst_dob_mux_b8/B2_11 ;
  wire  \inst_dob_mux_b8/B2_12 ;
  wire  \inst_dob_mux_b8/B2_13 ;
  wire  \inst_dob_mux_b8/B2_14 ;
  wire  \inst_dob_mux_b8/B2_15 ;
  wire  \inst_dob_mux_b8/B2_2 ;
  wire  \inst_dob_mux_b8/B2_3 ;
  wire  \inst_dob_mux_b8/B2_4 ;
  wire  \inst_dob_mux_b8/B2_5 ;
  wire  \inst_dob_mux_b8/B2_6 ;
  wire  \inst_dob_mux_b8/B2_7 ;
  wire  \inst_dob_mux_b8/B2_8 ;
  wire  \inst_dob_mux_b8/B2_9 ;
  wire  \inst_dob_mux_b8/B3_0 ;
  wire  \inst_dob_mux_b8/B3_1 ;
  wire  \inst_dob_mux_b8/B3_2 ;
  wire  \inst_dob_mux_b8/B3_3 ;
  wire  \inst_dob_mux_b8/B3_4 ;
  wire  \inst_dob_mux_b8/B3_5 ;
  wire  \inst_dob_mux_b8/B3_6 ;
  wire  \inst_dob_mux_b8/B3_7 ;
  wire  \inst_dob_mux_b8/B4_0 ;
  wire  \inst_dob_mux_b8/B4_1 ;
  wire  \inst_dob_mux_b8/B4_2 ;
  wire  \inst_dob_mux_b8/B4_3 ;
  wire  \inst_dob_mux_b8/B5_0 ;
  wire  \inst_dob_mux_b8/B5_1 ;
  wire  \inst_dob_mux_b9/B0_0 ;
  wire  \inst_dob_mux_b9/B0_1 ;
  wire  \inst_dob_mux_b9/B0_10 ;
  wire  \inst_dob_mux_b9/B0_11 ;
  wire  \inst_dob_mux_b9/B0_12 ;
  wire  \inst_dob_mux_b9/B0_13 ;
  wire  \inst_dob_mux_b9/B0_14 ;
  wire  \inst_dob_mux_b9/B0_15 ;
  wire  \inst_dob_mux_b9/B0_16 ;
  wire  \inst_dob_mux_b9/B0_17 ;
  wire  \inst_dob_mux_b9/B0_18 ;
  wire  \inst_dob_mux_b9/B0_19 ;
  wire  \inst_dob_mux_b9/B0_2 ;
  wire  \inst_dob_mux_b9/B0_20 ;
  wire  \inst_dob_mux_b9/B0_21 ;
  wire  \inst_dob_mux_b9/B0_22 ;
  wire  \inst_dob_mux_b9/B0_23 ;
  wire  \inst_dob_mux_b9/B0_24 ;
  wire  \inst_dob_mux_b9/B0_25 ;
  wire  \inst_dob_mux_b9/B0_26 ;
  wire  \inst_dob_mux_b9/B0_27 ;
  wire  \inst_dob_mux_b9/B0_28 ;
  wire  \inst_dob_mux_b9/B0_29 ;
  wire  \inst_dob_mux_b9/B0_3 ;
  wire  \inst_dob_mux_b9/B0_30 ;
  wire  \inst_dob_mux_b9/B0_31 ;
  wire  \inst_dob_mux_b9/B0_32 ;
  wire  \inst_dob_mux_b9/B0_33 ;
  wire  \inst_dob_mux_b9/B0_34 ;
  wire  \inst_dob_mux_b9/B0_35 ;
  wire  \inst_dob_mux_b9/B0_36 ;
  wire  \inst_dob_mux_b9/B0_37 ;
  wire  \inst_dob_mux_b9/B0_38 ;
  wire  \inst_dob_mux_b9/B0_39 ;
  wire  \inst_dob_mux_b9/B0_4 ;
  wire  \inst_dob_mux_b9/B0_40 ;
  wire  \inst_dob_mux_b9/B0_41 ;
  wire  \inst_dob_mux_b9/B0_42 ;
  wire  \inst_dob_mux_b9/B0_43 ;
  wire  \inst_dob_mux_b9/B0_44 ;
  wire  \inst_dob_mux_b9/B0_45 ;
  wire  \inst_dob_mux_b9/B0_46 ;
  wire  \inst_dob_mux_b9/B0_47 ;
  wire  \inst_dob_mux_b9/B0_48 ;
  wire  \inst_dob_mux_b9/B0_49 ;
  wire  \inst_dob_mux_b9/B0_5 ;
  wire  \inst_dob_mux_b9/B0_50 ;
  wire  \inst_dob_mux_b9/B0_51 ;
  wire  \inst_dob_mux_b9/B0_52 ;
  wire  \inst_dob_mux_b9/B0_53 ;
  wire  \inst_dob_mux_b9/B0_54 ;
  wire  \inst_dob_mux_b9/B0_55 ;
  wire  \inst_dob_mux_b9/B0_56 ;
  wire  \inst_dob_mux_b9/B0_57 ;
  wire  \inst_dob_mux_b9/B0_58 ;
  wire  \inst_dob_mux_b9/B0_59 ;
  wire  \inst_dob_mux_b9/B0_6 ;
  wire  \inst_dob_mux_b9/B0_60 ;
  wire  \inst_dob_mux_b9/B0_61 ;
  wire  \inst_dob_mux_b9/B0_62 ;
  wire  \inst_dob_mux_b9/B0_63 ;
  wire  \inst_dob_mux_b9/B0_7 ;
  wire  \inst_dob_mux_b9/B0_8 ;
  wire  \inst_dob_mux_b9/B0_9 ;
  wire  \inst_dob_mux_b9/B1_0 ;
  wire  \inst_dob_mux_b9/B1_1 ;
  wire  \inst_dob_mux_b9/B1_10 ;
  wire  \inst_dob_mux_b9/B1_11 ;
  wire  \inst_dob_mux_b9/B1_12 ;
  wire  \inst_dob_mux_b9/B1_13 ;
  wire  \inst_dob_mux_b9/B1_14 ;
  wire  \inst_dob_mux_b9/B1_15 ;
  wire  \inst_dob_mux_b9/B1_16 ;
  wire  \inst_dob_mux_b9/B1_17 ;
  wire  \inst_dob_mux_b9/B1_18 ;
  wire  \inst_dob_mux_b9/B1_19 ;
  wire  \inst_dob_mux_b9/B1_2 ;
  wire  \inst_dob_mux_b9/B1_20 ;
  wire  \inst_dob_mux_b9/B1_21 ;
  wire  \inst_dob_mux_b9/B1_22 ;
  wire  \inst_dob_mux_b9/B1_23 ;
  wire  \inst_dob_mux_b9/B1_24 ;
  wire  \inst_dob_mux_b9/B1_25 ;
  wire  \inst_dob_mux_b9/B1_26 ;
  wire  \inst_dob_mux_b9/B1_27 ;
  wire  \inst_dob_mux_b9/B1_28 ;
  wire  \inst_dob_mux_b9/B1_29 ;
  wire  \inst_dob_mux_b9/B1_3 ;
  wire  \inst_dob_mux_b9/B1_30 ;
  wire  \inst_dob_mux_b9/B1_31 ;
  wire  \inst_dob_mux_b9/B1_4 ;
  wire  \inst_dob_mux_b9/B1_5 ;
  wire  \inst_dob_mux_b9/B1_6 ;
  wire  \inst_dob_mux_b9/B1_7 ;
  wire  \inst_dob_mux_b9/B1_8 ;
  wire  \inst_dob_mux_b9/B1_9 ;
  wire  \inst_dob_mux_b9/B2_0 ;
  wire  \inst_dob_mux_b9/B2_1 ;
  wire  \inst_dob_mux_b9/B2_10 ;
  wire  \inst_dob_mux_b9/B2_11 ;
  wire  \inst_dob_mux_b9/B2_12 ;
  wire  \inst_dob_mux_b9/B2_13 ;
  wire  \inst_dob_mux_b9/B2_14 ;
  wire  \inst_dob_mux_b9/B2_15 ;
  wire  \inst_dob_mux_b9/B2_2 ;
  wire  \inst_dob_mux_b9/B2_3 ;
  wire  \inst_dob_mux_b9/B2_4 ;
  wire  \inst_dob_mux_b9/B2_5 ;
  wire  \inst_dob_mux_b9/B2_6 ;
  wire  \inst_dob_mux_b9/B2_7 ;
  wire  \inst_dob_mux_b9/B2_8 ;
  wire  \inst_dob_mux_b9/B2_9 ;
  wire  \inst_dob_mux_b9/B3_0 ;
  wire  \inst_dob_mux_b9/B3_1 ;
  wire  \inst_dob_mux_b9/B3_2 ;
  wire  \inst_dob_mux_b9/B3_3 ;
  wire  \inst_dob_mux_b9/B3_4 ;
  wire  \inst_dob_mux_b9/B3_5 ;
  wire  \inst_dob_mux_b9/B3_6 ;
  wire  \inst_dob_mux_b9/B3_7 ;
  wire  \inst_dob_mux_b9/B4_0 ;
  wire  \inst_dob_mux_b9/B4_1 ;
  wire  \inst_dob_mux_b9/B4_2 ;
  wire  \inst_dob_mux_b9/B4_3 ;
  wire  \inst_dob_mux_b9/B5_0 ;
  wire  \inst_dob_mux_b9/B5_1 ;
  wire \and_Naddra[11]_Naddr_o ;
  wire \and_Naddra[11]_Naddr_o_and_cea ;
  wire \and_Naddra[12]_Naddr_o ;
  wire \and_Naddra[12]_Naddr_o_al_n54 ;
  wire \and_Naddra[12]_addra_o ;
  wire \and_Naddra[12]_addra_o_al_n86 ;
  wire \and_Naddrb[11]_Naddr_o ;
  wire \and_Naddrb[11]_Naddr_o_and_ceb ;
  wire \and_Naddrb[12]_Naddr_o ;
  wire \and_Naddrb[12]_Naddr_o_al_n57 ;
  wire \and_Naddrb[12]_addrb_o ;
  wire \and_Naddrb[12]_addrb_o_al_n89 ;
  wire \and_addra[12]_Naddra_o ;
  wire \and_addra[12]_Naddra_o_al_n70 ;
  wire \and_addra[12]_addra[_o ;
  wire \and_addra[12]_addra[_o_al_n102 ;
  wire \and_addrb[12]_Naddrb_o ;
  wire \and_addrb[12]_Naddrb_o_al_n73 ;
  wire \and_addrb[12]_addrb[_o ;
  wire \and_addrb[12]_addrb[_o_al_n105 ;
  wire inst_dob_i0_000;
  wire inst_dob_i0_001;
  wire inst_dob_i0_002;
  wire inst_dob_i0_003;
  wire inst_dob_i0_004;
  wire inst_dob_i0_005;
  wire inst_dob_i0_006;
  wire inst_dob_i0_007;
  wire inst_dob_i0_008;
  wire inst_dob_i0_009;
  wire inst_dob_i0_010;
  wire inst_dob_i0_011;
  wire inst_dob_i0_012;
  wire inst_dob_i0_013;
  wire inst_dob_i0_014;
  wire inst_dob_i0_015;
  wire inst_dob_i10_000;
  wire inst_dob_i10_001;
  wire inst_dob_i10_002;
  wire inst_dob_i10_003;
  wire inst_dob_i10_004;
  wire inst_dob_i10_005;
  wire inst_dob_i10_006;
  wire inst_dob_i10_007;
  wire inst_dob_i10_008;
  wire inst_dob_i12_000;
  wire inst_dob_i12_001;
  wire inst_dob_i12_002;
  wire inst_dob_i12_003;
  wire inst_dob_i12_004;
  wire inst_dob_i12_005;
  wire inst_dob_i12_006;
  wire inst_dob_i12_007;
  wire inst_dob_i12_008;
  wire inst_dob_i14_000;
  wire inst_dob_i14_001;
  wire inst_dob_i14_002;
  wire inst_dob_i14_003;
  wire inst_dob_i14_004;
  wire inst_dob_i14_005;
  wire inst_dob_i14_006;
  wire inst_dob_i14_007;
  wire inst_dob_i14_008;
  wire inst_dob_i16_000;
  wire inst_dob_i16_001;
  wire inst_dob_i16_002;
  wire inst_dob_i16_003;
  wire inst_dob_i16_004;
  wire inst_dob_i16_005;
  wire inst_dob_i16_006;
  wire inst_dob_i16_007;
  wire inst_dob_i16_008;
  wire inst_dob_i16_009;
  wire inst_dob_i16_010;
  wire inst_dob_i16_011;
  wire inst_dob_i16_012;
  wire inst_dob_i16_013;
  wire inst_dob_i16_014;
  wire inst_dob_i16_015;
  wire inst_dob_i18_000;
  wire inst_dob_i18_001;
  wire inst_dob_i18_002;
  wire inst_dob_i18_003;
  wire inst_dob_i18_004;
  wire inst_dob_i18_005;
  wire inst_dob_i18_006;
  wire inst_dob_i18_007;
  wire inst_dob_i18_008;
  wire inst_dob_i20_000;
  wire inst_dob_i20_001;
  wire inst_dob_i20_002;
  wire inst_dob_i20_003;
  wire inst_dob_i20_004;
  wire inst_dob_i20_005;
  wire inst_dob_i20_006;
  wire inst_dob_i20_007;
  wire inst_dob_i20_008;
  wire inst_dob_i22_000;
  wire inst_dob_i22_001;
  wire inst_dob_i22_002;
  wire inst_dob_i22_003;
  wire inst_dob_i22_004;
  wire inst_dob_i22_005;
  wire inst_dob_i22_006;
  wire inst_dob_i22_007;
  wire inst_dob_i22_008;
  wire inst_dob_i24_000;
  wire inst_dob_i24_001;
  wire inst_dob_i24_002;
  wire inst_dob_i24_003;
  wire inst_dob_i24_004;
  wire inst_dob_i24_005;
  wire inst_dob_i24_006;
  wire inst_dob_i24_007;
  wire inst_dob_i24_008;
  wire inst_dob_i26_000;
  wire inst_dob_i26_001;
  wire inst_dob_i26_002;
  wire inst_dob_i26_003;
  wire inst_dob_i26_004;
  wire inst_dob_i26_005;
  wire inst_dob_i26_006;
  wire inst_dob_i26_007;
  wire inst_dob_i26_008;
  wire inst_dob_i28_000;
  wire inst_dob_i28_001;
  wire inst_dob_i28_002;
  wire inst_dob_i28_003;
  wire inst_dob_i28_004;
  wire inst_dob_i28_005;
  wire inst_dob_i28_006;
  wire inst_dob_i28_007;
  wire inst_dob_i28_008;
  wire inst_dob_i2_000;
  wire inst_dob_i2_001;
  wire inst_dob_i2_002;
  wire inst_dob_i2_003;
  wire inst_dob_i2_004;
  wire inst_dob_i2_005;
  wire inst_dob_i2_006;
  wire inst_dob_i2_007;
  wire inst_dob_i2_008;
  wire inst_dob_i30_000;
  wire inst_dob_i30_001;
  wire inst_dob_i30_002;
  wire inst_dob_i30_003;
  wire inst_dob_i30_004;
  wire inst_dob_i30_005;
  wire inst_dob_i30_006;
  wire inst_dob_i30_007;
  wire inst_dob_i30_008;
  wire inst_dob_i32_000;
  wire inst_dob_i32_001;
  wire inst_dob_i32_002;
  wire inst_dob_i32_003;
  wire inst_dob_i32_004;
  wire inst_dob_i32_005;
  wire inst_dob_i32_006;
  wire inst_dob_i32_007;
  wire inst_dob_i32_008;
  wire inst_dob_i32_009;
  wire inst_dob_i32_010;
  wire inst_dob_i32_011;
  wire inst_dob_i32_012;
  wire inst_dob_i32_013;
  wire inst_dob_i32_014;
  wire inst_dob_i32_015;
  wire inst_dob_i34_000;
  wire inst_dob_i34_001;
  wire inst_dob_i34_002;
  wire inst_dob_i34_003;
  wire inst_dob_i34_004;
  wire inst_dob_i34_005;
  wire inst_dob_i34_006;
  wire inst_dob_i34_007;
  wire inst_dob_i34_008;
  wire inst_dob_i36_000;
  wire inst_dob_i36_001;
  wire inst_dob_i36_002;
  wire inst_dob_i36_003;
  wire inst_dob_i36_004;
  wire inst_dob_i36_005;
  wire inst_dob_i36_006;
  wire inst_dob_i36_007;
  wire inst_dob_i36_008;
  wire inst_dob_i38_000;
  wire inst_dob_i38_001;
  wire inst_dob_i38_002;
  wire inst_dob_i38_003;
  wire inst_dob_i38_004;
  wire inst_dob_i38_005;
  wire inst_dob_i38_006;
  wire inst_dob_i38_007;
  wire inst_dob_i38_008;
  wire inst_dob_i40_000;
  wire inst_dob_i40_001;
  wire inst_dob_i40_002;
  wire inst_dob_i40_003;
  wire inst_dob_i40_004;
  wire inst_dob_i40_005;
  wire inst_dob_i40_006;
  wire inst_dob_i40_007;
  wire inst_dob_i40_008;
  wire inst_dob_i42_000;
  wire inst_dob_i42_001;
  wire inst_dob_i42_002;
  wire inst_dob_i42_003;
  wire inst_dob_i42_004;
  wire inst_dob_i42_005;
  wire inst_dob_i42_006;
  wire inst_dob_i42_007;
  wire inst_dob_i42_008;
  wire inst_dob_i44_000;
  wire inst_dob_i44_001;
  wire inst_dob_i44_002;
  wire inst_dob_i44_003;
  wire inst_dob_i44_004;
  wire inst_dob_i44_005;
  wire inst_dob_i44_006;
  wire inst_dob_i44_007;
  wire inst_dob_i44_008;
  wire inst_dob_i46_000;
  wire inst_dob_i46_001;
  wire inst_dob_i46_002;
  wire inst_dob_i46_003;
  wire inst_dob_i46_004;
  wire inst_dob_i46_005;
  wire inst_dob_i46_006;
  wire inst_dob_i46_007;
  wire inst_dob_i46_008;
  wire inst_dob_i48_000;
  wire inst_dob_i48_001;
  wire inst_dob_i48_002;
  wire inst_dob_i48_003;
  wire inst_dob_i48_004;
  wire inst_dob_i48_005;
  wire inst_dob_i48_006;
  wire inst_dob_i48_007;
  wire inst_dob_i48_008;
  wire inst_dob_i48_009;
  wire inst_dob_i48_010;
  wire inst_dob_i48_011;
  wire inst_dob_i48_012;
  wire inst_dob_i48_013;
  wire inst_dob_i48_014;
  wire inst_dob_i48_015;
  wire inst_dob_i4_000;
  wire inst_dob_i4_001;
  wire inst_dob_i4_002;
  wire inst_dob_i4_003;
  wire inst_dob_i4_004;
  wire inst_dob_i4_005;
  wire inst_dob_i4_006;
  wire inst_dob_i4_007;
  wire inst_dob_i4_008;
  wire inst_dob_i50_000;
  wire inst_dob_i50_001;
  wire inst_dob_i50_002;
  wire inst_dob_i50_003;
  wire inst_dob_i50_004;
  wire inst_dob_i50_005;
  wire inst_dob_i50_006;
  wire inst_dob_i50_007;
  wire inst_dob_i50_008;
  wire inst_dob_i52_000;
  wire inst_dob_i52_001;
  wire inst_dob_i52_002;
  wire inst_dob_i52_003;
  wire inst_dob_i52_004;
  wire inst_dob_i52_005;
  wire inst_dob_i52_006;
  wire inst_dob_i52_007;
  wire inst_dob_i52_008;
  wire inst_dob_i54_000;
  wire inst_dob_i54_001;
  wire inst_dob_i54_002;
  wire inst_dob_i54_003;
  wire inst_dob_i54_004;
  wire inst_dob_i54_005;
  wire inst_dob_i54_006;
  wire inst_dob_i54_007;
  wire inst_dob_i54_008;
  wire inst_dob_i56_000;
  wire inst_dob_i56_001;
  wire inst_dob_i56_002;
  wire inst_dob_i56_003;
  wire inst_dob_i56_004;
  wire inst_dob_i56_005;
  wire inst_dob_i56_006;
  wire inst_dob_i56_007;
  wire inst_dob_i56_008;
  wire inst_dob_i58_000;
  wire inst_dob_i58_001;
  wire inst_dob_i58_002;
  wire inst_dob_i58_003;
  wire inst_dob_i58_004;
  wire inst_dob_i58_005;
  wire inst_dob_i58_006;
  wire inst_dob_i58_007;
  wire inst_dob_i58_008;
  wire inst_dob_i60_000;
  wire inst_dob_i60_001;
  wire inst_dob_i60_002;
  wire inst_dob_i60_003;
  wire inst_dob_i60_004;
  wire inst_dob_i60_005;
  wire inst_dob_i60_006;
  wire inst_dob_i60_007;
  wire inst_dob_i60_008;
  wire inst_dob_i62_000;
  wire inst_dob_i62_001;
  wire inst_dob_i62_002;
  wire inst_dob_i62_003;
  wire inst_dob_i62_004;
  wire inst_dob_i62_005;
  wire inst_dob_i62_006;
  wire inst_dob_i62_007;
  wire inst_dob_i62_008;
  wire inst_dob_i64_000;
  wire inst_dob_i64_001;
  wire inst_dob_i64_002;
  wire inst_dob_i64_003;
  wire inst_dob_i64_004;
  wire inst_dob_i64_005;
  wire inst_dob_i64_006;
  wire inst_dob_i64_007;
  wire inst_dob_i64_008;
  wire inst_dob_i64_009;
  wire inst_dob_i64_010;
  wire inst_dob_i64_011;
  wire inst_dob_i64_012;
  wire inst_dob_i64_013;
  wire inst_dob_i64_014;
  wire inst_dob_i64_015;
  wire inst_dob_i6_000;
  wire inst_dob_i6_001;
  wire inst_dob_i6_002;
  wire inst_dob_i6_003;
  wire inst_dob_i6_004;
  wire inst_dob_i6_005;
  wire inst_dob_i6_006;
  wire inst_dob_i6_007;
  wire inst_dob_i6_008;
  wire inst_dob_i8_000;
  wire inst_dob_i8_001;
  wire inst_dob_i8_002;
  wire inst_dob_i8_003;
  wire inst_dob_i8_004;
  wire inst_dob_i8_005;
  wire inst_dob_i8_006;
  wire inst_dob_i8_007;
  wire inst_dob_i8_008;

  reg_sr_as_w1 addrb_pipe_b0 (
    .clk(clkb),
    .d(addrb[9]),
    .en(ceb),
    .reset(rstb),
    .set(1'b0),
    .q(addrb_piped[0]));
  reg_sr_as_w1 addrb_pipe_b1 (
    .clk(clkb),
    .d(addrb[10]),
    .en(ceb),
    .reset(rstb),
    .set(1'b0),
    .q(addrb_piped[1]));
  reg_sr_as_w1 addrb_pipe_b2 (
    .clk(clkb),
    .d(addrb[11]),
    .en(ceb),
    .reset(rstb),
    .set(1'b0),
    .q(addrb_piped[2]));
  reg_sr_as_w1 addrb_pipe_b3 (
    .clk(clkb),
    .d(addrb[12]),
    .en(ceb),
    .reset(rstb),
    .set(1'b0),
    .q(addrb_piped[3]));
  reg_sr_as_w1 addrb_pipe_b4 (
    .clk(clkb),
    .d(addrb[13]),
    .en(ceb),
    .reset(rstb),
    .set(1'b0),
    .q(addrb_piped[4]));
  reg_sr_as_w1 addrb_pipe_b5 (
    .clk(clkb),
    .d(addrb[14]),
    .en(ceb),
    .reset(rstb),
    .set(1'b0),
    .q(addrb_piped[5]));
  reg_sr_as_w1 addrb_pipe_b6 (
    .clk(clkb),
    .d(addrb[15]),
    .en(ceb),
    .reset(rstb),
    .set(1'b0),
    .q(addrb_piped[6]));
  reg_sr_as_w1 addrb_piped_pipe_b0 (
    .clk(clkb),
    .d(addrb_piped[0]),
    .en(ceb),
    .reset(rstb),
    .set(1'b0),
    .q(addrb_piped_piped[0]));
  reg_sr_as_w1 addrb_piped_pipe_b1 (
    .clk(clkb),
    .d(addrb_piped[1]),
    .en(ceb),
    .reset(rstb),
    .set(1'b0),
    .q(addrb_piped_piped[1]));
  reg_sr_as_w1 addrb_piped_pipe_b2 (
    .clk(clkb),
    .d(addrb_piped[2]),
    .en(ceb),
    .reset(rstb),
    .set(1'b0),
    .q(addrb_piped_piped[2]));
  reg_sr_as_w1 addrb_piped_pipe_b3 (
    .clk(clkb),
    .d(addrb_piped[3]),
    .en(ceb),
    .reset(rstb),
    .set(1'b0),
    .q(addrb_piped_piped[3]));
  reg_sr_as_w1 addrb_piped_pipe_b4 (
    .clk(clkb),
    .d(addrb_piped[4]),
    .en(ceb),
    .reset(rstb),
    .set(1'b0),
    .q(addrb_piped_piped[4]));
  reg_sr_as_w1 addrb_piped_pipe_b5 (
    .clk(clkb),
    .d(addrb_piped[5]),
    .en(ceb),
    .reset(rstb),
    .set(1'b0),
    .q(addrb_piped_piped[5]));
  reg_sr_as_w1 addrb_piped_pipe_b6 (
    .clk(clkb),
    .d(addrb_piped[6]),
    .en(ceb),
    .reset(rstb),
    .set(1'b0),
    .q(addrb_piped_piped[6]));
  and \and_Naddra[11]_Naddr  (\and_Naddra[11]_Naddr_o , ~addra[11], ~addra[12], ~addra[13], ~addra[14], addra[15]);
  and \and_Naddra[11]_Naddr_o_and_cea_i  (\and_Naddra[11]_Naddr_o_and_cea , \and_Naddra[11]_Naddr_o , cea);
  and \and_Naddra[12]_Naddr  (\and_Naddra[12]_Naddr_o , ~addra[12], ~addra[13], ~addra[14], ~addra[15]);
  and \and_Naddra[12]_Naddr_al_u54  (\and_Naddra[12]_Naddr_o_al_n54 , ~addra[12], ~addra[13], addra[14], ~addra[15]);
  and \and_Naddra[12]_addra  (\and_Naddra[12]_addra_o , ~addra[12], addra[13], ~addra[14], ~addra[15]);
  and \and_Naddra[12]_addra_al_u86  (\and_Naddra[12]_addra_o_al_n86 , ~addra[12], addra[13], addra[14], ~addra[15]);
  and \and_Naddrb[11]_Naddr  (\and_Naddrb[11]_Naddr_o , ~addrb[11], ~addrb[12], ~addrb[13], ~addrb[14], addrb[15]);
  and \and_Naddrb[11]_Naddr_o_and_ceb_i  (\and_Naddrb[11]_Naddr_o_and_ceb , \and_Naddrb[11]_Naddr_o , ceb);
  and \and_Naddrb[12]_Naddr  (\and_Naddrb[12]_Naddr_o , ~addrb[12], ~addrb[13], ~addrb[14], ~addrb[15]);
  and \and_Naddrb[12]_Naddr_al_u57  (\and_Naddrb[12]_Naddr_o_al_n57 , ~addrb[12], ~addrb[13], addrb[14], ~addrb[15]);
  and \and_Naddrb[12]_addrb  (\and_Naddrb[12]_addrb_o , ~addrb[12], addrb[13], ~addrb[14], ~addrb[15]);
  and \and_Naddrb[12]_addrb_al_u89  (\and_Naddrb[12]_addrb_o_al_n89 , ~addrb[12], addrb[13], addrb[14], ~addrb[15]);
  and \and_addra[12]_Naddra  (\and_addra[12]_Naddra_o , addra[12], ~addra[13], ~addra[14], ~addra[15]);
  and \and_addra[12]_Naddra_al_u70  (\and_addra[12]_Naddra_o_al_n70 , addra[12], ~addra[13], addra[14], ~addra[15]);
  and \and_addra[12]_addra[  (\and_addra[12]_addra[_o , addra[12], addra[13], ~addra[14], ~addra[15]);
  and \and_addra[12]_addra[_al_u102  (\and_addra[12]_addra[_o_al_n102 , addra[12], addra[13], addra[14], ~addra[15]);
  and \and_addrb[12]_Naddrb  (\and_addrb[12]_Naddrb_o , addrb[12], ~addrb[13], ~addrb[14], ~addrb[15]);
  and \and_addrb[12]_Naddrb_al_u73  (\and_addrb[12]_Naddrb_o_al_n73 , addrb[12], ~addrb[13], addrb[14], ~addrb[15]);
  and \and_addrb[12]_addrb[  (\and_addrb[12]_addrb[_o , addrb[12], addrb[13], ~addrb[14], ~addrb[15]);
  and \and_addrb[12]_addrb[_al_u105  (\and_addrb[12]_addrb[_o_al_n105 , addrb[12], addrb[13], addrb[14], ~addrb[15]);
  EG_PHY_CONFIG #(
    .DONE_PERSISTN("ENABLE"),
    .INIT_PERSISTN("ENABLE"),
    .JTAG_PERSISTN("DISABLE"),
    .PROGRAMN_PERSISTN("DISABLE"))
    config_inst ();
  // address_offset=0;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("INV"),
    .CSB1("INV"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_000000_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa({\and_Naddra[12]_Naddr_o ,addra[11:10]}),
    .csb({\and_Naddrb[12]_Naddr_o ,addrb[11:10]}),
    .dia(dia[8:0]),
    .rstb(rstb),
    .dob({inst_dob_i0_008,inst_dob_i0_007,inst_dob_i0_006,inst_dob_i0_005,inst_dob_i0_004,inst_dob_i0_003,inst_dob_i0_002,inst_dob_i0_001,inst_dob_i0_000}));
  // address_offset=0;data_offset=9;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("INV"),
    .CSB1("INV"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_000000_009 (
    .addra(addra[12:0]),
    .addrb(addrb[12:0]),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[15:13]),
    .csb(addrb[15:13]),
    .dia({open_n70,open_n71,open_n72,open_n73,open_n74,open_n75,open_n76,dia[9],open_n77}),
    .rstb(rstb),
    .dob({open_n101,open_n102,open_n103,open_n104,open_n105,open_n106,open_n107,open_n108,inst_dob_i0_009}));
  // address_offset=0;data_offset=10;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("INV"),
    .CSB1("INV"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_000000_010 (
    .addra(addra[12:0]),
    .addrb(addrb[12:0]),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[15:13]),
    .csb(addrb[15:13]),
    .dia({open_n109,open_n110,open_n111,open_n112,open_n113,open_n114,open_n115,dia[10],open_n116}),
    .rstb(rstb),
    .dob({open_n140,open_n141,open_n142,open_n143,open_n144,open_n145,open_n146,open_n147,inst_dob_i0_010}));
  // address_offset=0;data_offset=11;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("INV"),
    .CSB1("INV"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_000000_011 (
    .addra(addra[12:0]),
    .addrb(addrb[12:0]),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[15:13]),
    .csb(addrb[15:13]),
    .dia({open_n148,open_n149,open_n150,open_n151,open_n152,open_n153,open_n154,dia[11],open_n155}),
    .rstb(rstb),
    .dob({open_n179,open_n180,open_n181,open_n182,open_n183,open_n184,open_n185,open_n186,inst_dob_i0_011}));
  // address_offset=0;data_offset=12;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("INV"),
    .CSB1("INV"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_000000_012 (
    .addra(addra[12:0]),
    .addrb(addrb[12:0]),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[15:13]),
    .csb(addrb[15:13]),
    .dia({open_n187,open_n188,open_n189,open_n190,open_n191,open_n192,open_n193,dia[12],open_n194}),
    .rstb(rstb),
    .dob({open_n218,open_n219,open_n220,open_n221,open_n222,open_n223,open_n224,open_n225,inst_dob_i0_012}));
  // address_offset=0;data_offset=13;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("INV"),
    .CSB1("INV"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_000000_013 (
    .addra(addra[12:0]),
    .addrb(addrb[12:0]),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[15:13]),
    .csb(addrb[15:13]),
    .dia({open_n226,open_n227,open_n228,open_n229,open_n230,open_n231,open_n232,dia[13],open_n233}),
    .rstb(rstb),
    .dob({open_n257,open_n258,open_n259,open_n260,open_n261,open_n262,open_n263,open_n264,inst_dob_i0_013}));
  // address_offset=0;data_offset=14;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("INV"),
    .CSB1("INV"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_000000_014 (
    .addra(addra[12:0]),
    .addrb(addrb[12:0]),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[15:13]),
    .csb(addrb[15:13]),
    .dia({open_n265,open_n266,open_n267,open_n268,open_n269,open_n270,open_n271,dia[14],open_n272}),
    .rstb(rstb),
    .dob({open_n296,open_n297,open_n298,open_n299,open_n300,open_n301,open_n302,open_n303,inst_dob_i0_014}));
  // address_offset=0;data_offset=15;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("INV"),
    .CSB1("INV"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_000000_015 (
    .addra(addra[12:0]),
    .addrb(addrb[12:0]),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[15:13]),
    .csb(addrb[15:13]),
    .dia({open_n304,open_n305,open_n306,open_n307,open_n308,open_n309,open_n310,dia[15],open_n311}),
    .rstb(rstb),
    .dob({open_n335,open_n336,open_n337,open_n338,open_n339,open_n340,open_n341,open_n342,inst_dob_i0_015}));
  // address_offset=1024;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("SIG"),
    .CSB1("INV"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_001024_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa({\and_Naddra[12]_Naddr_o ,addra[11:10]}),
    .csb({\and_Naddrb[12]_Naddr_o ,addrb[11:10]}),
    .dia(dia[8:0]),
    .rstb(rstb),
    .dob({inst_dob_i2_008,inst_dob_i2_007,inst_dob_i2_006,inst_dob_i2_005,inst_dob_i2_004,inst_dob_i2_003,inst_dob_i2_002,inst_dob_i2_001,inst_dob_i2_000}));
  // address_offset=2048;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("INV"),
    .CSB1("SIG"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_002048_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa({\and_Naddra[12]_Naddr_o ,addra[11:10]}),
    .csb({\and_Naddrb[12]_Naddr_o ,addrb[11:10]}),
    .dia(dia[8:0]),
    .rstb(rstb),
    .dob({inst_dob_i4_008,inst_dob_i4_007,inst_dob_i4_006,inst_dob_i4_005,inst_dob_i4_004,inst_dob_i4_003,inst_dob_i4_002,inst_dob_i4_001,inst_dob_i4_000}));
  // address_offset=3072;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("SIG"),
    .CSB1("SIG"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_003072_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa({\and_Naddra[12]_Naddr_o ,addra[11:10]}),
    .csb({\and_Naddrb[12]_Naddr_o ,addrb[11:10]}),
    .dia(dia[8:0]),
    .rstb(rstb),
    .dob({inst_dob_i6_008,inst_dob_i6_007,inst_dob_i6_006,inst_dob_i6_005,inst_dob_i6_004,inst_dob_i6_003,inst_dob_i6_002,inst_dob_i6_001,inst_dob_i6_000}));
  // address_offset=4096;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("INV"),
    .CSB1("INV"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_004096_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa({\and_addra[12]_Naddra_o ,addra[11:10]}),
    .csb({\and_addrb[12]_Naddrb_o ,addrb[11:10]}),
    .dia(dia[8:0]),
    .rstb(rstb),
    .dob({inst_dob_i8_008,inst_dob_i8_007,inst_dob_i8_006,inst_dob_i8_005,inst_dob_i8_004,inst_dob_i8_003,inst_dob_i8_002,inst_dob_i8_001,inst_dob_i8_000}));
  // address_offset=5120;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("SIG"),
    .CSB1("INV"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_005120_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa({\and_addra[12]_Naddra_o ,addra[11:10]}),
    .csb({\and_addrb[12]_Naddrb_o ,addrb[11:10]}),
    .dia(dia[8:0]),
    .rstb(rstb),
    .dob({inst_dob_i10_008,inst_dob_i10_007,inst_dob_i10_006,inst_dob_i10_005,inst_dob_i10_004,inst_dob_i10_003,inst_dob_i10_002,inst_dob_i10_001,inst_dob_i10_000}));
  // address_offset=6144;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("INV"),
    .CSB1("SIG"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_006144_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa({\and_addra[12]_Naddra_o ,addra[11:10]}),
    .csb({\and_addrb[12]_Naddrb_o ,addrb[11:10]}),
    .dia(dia[8:0]),
    .rstb(rstb),
    .dob({inst_dob_i12_008,inst_dob_i12_007,inst_dob_i12_006,inst_dob_i12_005,inst_dob_i12_004,inst_dob_i12_003,inst_dob_i12_002,inst_dob_i12_001,inst_dob_i12_000}));
  // address_offset=7168;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("SIG"),
    .CSB1("SIG"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_007168_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa({\and_addra[12]_Naddra_o ,addra[11:10]}),
    .csb({\and_addrb[12]_Naddrb_o ,addrb[11:10]}),
    .dia(dia[8:0]),
    .rstb(rstb),
    .dob({inst_dob_i14_008,inst_dob_i14_007,inst_dob_i14_006,inst_dob_i14_005,inst_dob_i14_004,inst_dob_i14_003,inst_dob_i14_002,inst_dob_i14_001,inst_dob_i14_000}));
  // address_offset=8192;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("INV"),
    .CSB1("INV"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_008192_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa({\and_Naddra[12]_addra_o ,addra[11:10]}),
    .csb({\and_Naddrb[12]_addrb_o ,addrb[11:10]}),
    .dia(dia[8:0]),
    .rstb(rstb),
    .dob({inst_dob_i16_008,inst_dob_i16_007,inst_dob_i16_006,inst_dob_i16_005,inst_dob_i16_004,inst_dob_i16_003,inst_dob_i16_002,inst_dob_i16_001,inst_dob_i16_000}));
  // address_offset=8192;data_offset=9;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("SIG"),
    .CSB1("INV"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_008192_009 (
    .addra(addra[12:0]),
    .addrb(addrb[12:0]),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[15:13]),
    .csb(addrb[15:13]),
    .dia({open_n527,open_n528,open_n529,open_n530,open_n531,open_n532,open_n533,dia[9],open_n534}),
    .rstb(rstb),
    .dob({open_n558,open_n559,open_n560,open_n561,open_n562,open_n563,open_n564,open_n565,inst_dob_i16_009}));
  // address_offset=8192;data_offset=10;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("SIG"),
    .CSB1("INV"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_008192_010 (
    .addra(addra[12:0]),
    .addrb(addrb[12:0]),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[15:13]),
    .csb(addrb[15:13]),
    .dia({open_n566,open_n567,open_n568,open_n569,open_n570,open_n571,open_n572,dia[10],open_n573}),
    .rstb(rstb),
    .dob({open_n597,open_n598,open_n599,open_n600,open_n601,open_n602,open_n603,open_n604,inst_dob_i16_010}));
  // address_offset=8192;data_offset=11;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("SIG"),
    .CSB1("INV"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_008192_011 (
    .addra(addra[12:0]),
    .addrb(addrb[12:0]),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[15:13]),
    .csb(addrb[15:13]),
    .dia({open_n605,open_n606,open_n607,open_n608,open_n609,open_n610,open_n611,dia[11],open_n612}),
    .rstb(rstb),
    .dob({open_n636,open_n637,open_n638,open_n639,open_n640,open_n641,open_n642,open_n643,inst_dob_i16_011}));
  // address_offset=8192;data_offset=12;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("SIG"),
    .CSB1("INV"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_008192_012 (
    .addra(addra[12:0]),
    .addrb(addrb[12:0]),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[15:13]),
    .csb(addrb[15:13]),
    .dia({open_n644,open_n645,open_n646,open_n647,open_n648,open_n649,open_n650,dia[12],open_n651}),
    .rstb(rstb),
    .dob({open_n675,open_n676,open_n677,open_n678,open_n679,open_n680,open_n681,open_n682,inst_dob_i16_012}));
  // address_offset=8192;data_offset=13;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("SIG"),
    .CSB1("INV"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_008192_013 (
    .addra(addra[12:0]),
    .addrb(addrb[12:0]),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[15:13]),
    .csb(addrb[15:13]),
    .dia({open_n683,open_n684,open_n685,open_n686,open_n687,open_n688,open_n689,dia[13],open_n690}),
    .rstb(rstb),
    .dob({open_n714,open_n715,open_n716,open_n717,open_n718,open_n719,open_n720,open_n721,inst_dob_i16_013}));
  // address_offset=8192;data_offset=14;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("SIG"),
    .CSB1("INV"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_008192_014 (
    .addra(addra[12:0]),
    .addrb(addrb[12:0]),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[15:13]),
    .csb(addrb[15:13]),
    .dia({open_n722,open_n723,open_n724,open_n725,open_n726,open_n727,open_n728,dia[14],open_n729}),
    .rstb(rstb),
    .dob({open_n753,open_n754,open_n755,open_n756,open_n757,open_n758,open_n759,open_n760,inst_dob_i16_014}));
  // address_offset=8192;data_offset=15;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("SIG"),
    .CSB1("INV"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_008192_015 (
    .addra(addra[12:0]),
    .addrb(addrb[12:0]),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[15:13]),
    .csb(addrb[15:13]),
    .dia({open_n761,open_n762,open_n763,open_n764,open_n765,open_n766,open_n767,dia[15],open_n768}),
    .rstb(rstb),
    .dob({open_n792,open_n793,open_n794,open_n795,open_n796,open_n797,open_n798,open_n799,inst_dob_i16_015}));
  // address_offset=9216;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("SIG"),
    .CSB1("INV"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_009216_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa({\and_Naddra[12]_addra_o ,addra[11:10]}),
    .csb({\and_Naddrb[12]_addrb_o ,addrb[11:10]}),
    .dia(dia[8:0]),
    .rstb(rstb),
    .dob({inst_dob_i18_008,inst_dob_i18_007,inst_dob_i18_006,inst_dob_i18_005,inst_dob_i18_004,inst_dob_i18_003,inst_dob_i18_002,inst_dob_i18_001,inst_dob_i18_000}));
  // address_offset=10240;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("INV"),
    .CSB1("SIG"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_010240_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa({\and_Naddra[12]_addra_o ,addra[11:10]}),
    .csb({\and_Naddrb[12]_addrb_o ,addrb[11:10]}),
    .dia(dia[8:0]),
    .rstb(rstb),
    .dob({inst_dob_i20_008,inst_dob_i20_007,inst_dob_i20_006,inst_dob_i20_005,inst_dob_i20_004,inst_dob_i20_003,inst_dob_i20_002,inst_dob_i20_001,inst_dob_i20_000}));
  // address_offset=11264;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("SIG"),
    .CSB1("SIG"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_011264_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa({\and_Naddra[12]_addra_o ,addra[11:10]}),
    .csb({\and_Naddrb[12]_addrb_o ,addrb[11:10]}),
    .dia(dia[8:0]),
    .rstb(rstb),
    .dob({inst_dob_i22_008,inst_dob_i22_007,inst_dob_i22_006,inst_dob_i22_005,inst_dob_i22_004,inst_dob_i22_003,inst_dob_i22_002,inst_dob_i22_001,inst_dob_i22_000}));
  // address_offset=12288;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("INV"),
    .CSB1("INV"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_012288_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa({\and_addra[12]_addra[_o ,addra[11:10]}),
    .csb({\and_addrb[12]_addrb[_o ,addrb[11:10]}),
    .dia(dia[8:0]),
    .rstb(rstb),
    .dob({inst_dob_i24_008,inst_dob_i24_007,inst_dob_i24_006,inst_dob_i24_005,inst_dob_i24_004,inst_dob_i24_003,inst_dob_i24_002,inst_dob_i24_001,inst_dob_i24_000}));
  // address_offset=13312;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("SIG"),
    .CSB1("INV"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_013312_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa({\and_addra[12]_addra[_o ,addra[11:10]}),
    .csb({\and_addrb[12]_addrb[_o ,addrb[11:10]}),
    .dia(dia[8:0]),
    .rstb(rstb),
    .dob({inst_dob_i26_008,inst_dob_i26_007,inst_dob_i26_006,inst_dob_i26_005,inst_dob_i26_004,inst_dob_i26_003,inst_dob_i26_002,inst_dob_i26_001,inst_dob_i26_000}));
  // address_offset=14336;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("INV"),
    .CSB1("SIG"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_014336_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa({\and_addra[12]_addra[_o ,addra[11:10]}),
    .csb({\and_addrb[12]_addrb[_o ,addrb[11:10]}),
    .dia(dia[8:0]),
    .rstb(rstb),
    .dob({inst_dob_i28_008,inst_dob_i28_007,inst_dob_i28_006,inst_dob_i28_005,inst_dob_i28_004,inst_dob_i28_003,inst_dob_i28_002,inst_dob_i28_001,inst_dob_i28_000}));
  // address_offset=15360;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("SIG"),
    .CSB1("SIG"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_015360_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa({\and_addra[12]_addra[_o ,addra[11:10]}),
    .csb({\and_addrb[12]_addrb[_o ,addrb[11:10]}),
    .dia(dia[8:0]),
    .rstb(rstb),
    .dob({inst_dob_i30_008,inst_dob_i30_007,inst_dob_i30_006,inst_dob_i30_005,inst_dob_i30_004,inst_dob_i30_003,inst_dob_i30_002,inst_dob_i30_001,inst_dob_i30_000}));
  // address_offset=16384;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("INV"),
    .CSB1("INV"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_016384_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa({\and_Naddra[12]_Naddr_o_al_n54 ,addra[11:10]}),
    .csb({\and_Naddrb[12]_Naddr_o_al_n57 ,addrb[11:10]}),
    .dia(dia[8:0]),
    .rstb(rstb),
    .dob({inst_dob_i32_008,inst_dob_i32_007,inst_dob_i32_006,inst_dob_i32_005,inst_dob_i32_004,inst_dob_i32_003,inst_dob_i32_002,inst_dob_i32_001,inst_dob_i32_000}));
  // address_offset=16384;data_offset=9;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("INV"),
    .CSB1("SIG"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_016384_009 (
    .addra(addra[12:0]),
    .addrb(addrb[12:0]),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[15:13]),
    .csb(addrb[15:13]),
    .dia({open_n984,open_n985,open_n986,open_n987,open_n988,open_n989,open_n990,dia[9],open_n991}),
    .rstb(rstb),
    .dob({open_n1015,open_n1016,open_n1017,open_n1018,open_n1019,open_n1020,open_n1021,open_n1022,inst_dob_i32_009}));
  // address_offset=16384;data_offset=10;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("INV"),
    .CSB1("SIG"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_016384_010 (
    .addra(addra[12:0]),
    .addrb(addrb[12:0]),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[15:13]),
    .csb(addrb[15:13]),
    .dia({open_n1023,open_n1024,open_n1025,open_n1026,open_n1027,open_n1028,open_n1029,dia[10],open_n1030}),
    .rstb(rstb),
    .dob({open_n1054,open_n1055,open_n1056,open_n1057,open_n1058,open_n1059,open_n1060,open_n1061,inst_dob_i32_010}));
  // address_offset=16384;data_offset=11;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("INV"),
    .CSB1("SIG"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_016384_011 (
    .addra(addra[12:0]),
    .addrb(addrb[12:0]),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[15:13]),
    .csb(addrb[15:13]),
    .dia({open_n1062,open_n1063,open_n1064,open_n1065,open_n1066,open_n1067,open_n1068,dia[11],open_n1069}),
    .rstb(rstb),
    .dob({open_n1093,open_n1094,open_n1095,open_n1096,open_n1097,open_n1098,open_n1099,open_n1100,inst_dob_i32_011}));
  // address_offset=16384;data_offset=12;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("INV"),
    .CSB1("SIG"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_016384_012 (
    .addra(addra[12:0]),
    .addrb(addrb[12:0]),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[15:13]),
    .csb(addrb[15:13]),
    .dia({open_n1101,open_n1102,open_n1103,open_n1104,open_n1105,open_n1106,open_n1107,dia[12],open_n1108}),
    .rstb(rstb),
    .dob({open_n1132,open_n1133,open_n1134,open_n1135,open_n1136,open_n1137,open_n1138,open_n1139,inst_dob_i32_012}));
  // address_offset=16384;data_offset=13;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("INV"),
    .CSB1("SIG"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_016384_013 (
    .addra(addra[12:0]),
    .addrb(addrb[12:0]),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[15:13]),
    .csb(addrb[15:13]),
    .dia({open_n1140,open_n1141,open_n1142,open_n1143,open_n1144,open_n1145,open_n1146,dia[13],open_n1147}),
    .rstb(rstb),
    .dob({open_n1171,open_n1172,open_n1173,open_n1174,open_n1175,open_n1176,open_n1177,open_n1178,inst_dob_i32_013}));
  // address_offset=16384;data_offset=14;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("INV"),
    .CSB1("SIG"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_016384_014 (
    .addra(addra[12:0]),
    .addrb(addrb[12:0]),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[15:13]),
    .csb(addrb[15:13]),
    .dia({open_n1179,open_n1180,open_n1181,open_n1182,open_n1183,open_n1184,open_n1185,dia[14],open_n1186}),
    .rstb(rstb),
    .dob({open_n1210,open_n1211,open_n1212,open_n1213,open_n1214,open_n1215,open_n1216,open_n1217,inst_dob_i32_014}));
  // address_offset=16384;data_offset=15;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("INV"),
    .CSB1("SIG"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_016384_015 (
    .addra(addra[12:0]),
    .addrb(addrb[12:0]),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[15:13]),
    .csb(addrb[15:13]),
    .dia({open_n1218,open_n1219,open_n1220,open_n1221,open_n1222,open_n1223,open_n1224,dia[15],open_n1225}),
    .rstb(rstb),
    .dob({open_n1249,open_n1250,open_n1251,open_n1252,open_n1253,open_n1254,open_n1255,open_n1256,inst_dob_i32_015}));
  // address_offset=17408;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("SIG"),
    .CSB1("INV"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_017408_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa({\and_Naddra[12]_Naddr_o_al_n54 ,addra[11:10]}),
    .csb({\and_Naddrb[12]_Naddr_o_al_n57 ,addrb[11:10]}),
    .dia(dia[8:0]),
    .rstb(rstb),
    .dob({inst_dob_i34_008,inst_dob_i34_007,inst_dob_i34_006,inst_dob_i34_005,inst_dob_i34_004,inst_dob_i34_003,inst_dob_i34_002,inst_dob_i34_001,inst_dob_i34_000}));
  // address_offset=18432;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("INV"),
    .CSB1("SIG"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_018432_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa({\and_Naddra[12]_Naddr_o_al_n54 ,addra[11:10]}),
    .csb({\and_Naddrb[12]_Naddr_o_al_n57 ,addrb[11:10]}),
    .dia(dia[8:0]),
    .rstb(rstb),
    .dob({inst_dob_i36_008,inst_dob_i36_007,inst_dob_i36_006,inst_dob_i36_005,inst_dob_i36_004,inst_dob_i36_003,inst_dob_i36_002,inst_dob_i36_001,inst_dob_i36_000}));
  // address_offset=19456;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("SIG"),
    .CSB1("SIG"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_019456_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa({\and_Naddra[12]_Naddr_o_al_n54 ,addra[11:10]}),
    .csb({\and_Naddrb[12]_Naddr_o_al_n57 ,addrb[11:10]}),
    .dia(dia[8:0]),
    .rstb(rstb),
    .dob({inst_dob_i38_008,inst_dob_i38_007,inst_dob_i38_006,inst_dob_i38_005,inst_dob_i38_004,inst_dob_i38_003,inst_dob_i38_002,inst_dob_i38_001,inst_dob_i38_000}));
  // address_offset=20480;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("INV"),
    .CSB1("INV"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_020480_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa({\and_addra[12]_Naddra_o_al_n70 ,addra[11:10]}),
    .csb({\and_addrb[12]_Naddrb_o_al_n73 ,addrb[11:10]}),
    .dia(dia[8:0]),
    .rstb(rstb),
    .dob({inst_dob_i40_008,inst_dob_i40_007,inst_dob_i40_006,inst_dob_i40_005,inst_dob_i40_004,inst_dob_i40_003,inst_dob_i40_002,inst_dob_i40_001,inst_dob_i40_000}));
  // address_offset=21504;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("SIG"),
    .CSB1("INV"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_021504_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa({\and_addra[12]_Naddra_o_al_n70 ,addra[11:10]}),
    .csb({\and_addrb[12]_Naddrb_o_al_n73 ,addrb[11:10]}),
    .dia(dia[8:0]),
    .rstb(rstb),
    .dob({inst_dob_i42_008,inst_dob_i42_007,inst_dob_i42_006,inst_dob_i42_005,inst_dob_i42_004,inst_dob_i42_003,inst_dob_i42_002,inst_dob_i42_001,inst_dob_i42_000}));
  // address_offset=22528;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("INV"),
    .CSB1("SIG"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_022528_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa({\and_addra[12]_Naddra_o_al_n70 ,addra[11:10]}),
    .csb({\and_addrb[12]_Naddrb_o_al_n73 ,addrb[11:10]}),
    .dia(dia[8:0]),
    .rstb(rstb),
    .dob({inst_dob_i44_008,inst_dob_i44_007,inst_dob_i44_006,inst_dob_i44_005,inst_dob_i44_004,inst_dob_i44_003,inst_dob_i44_002,inst_dob_i44_001,inst_dob_i44_000}));
  // address_offset=23552;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("SIG"),
    .CSB1("SIG"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_023552_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa({\and_addra[12]_Naddra_o_al_n70 ,addra[11:10]}),
    .csb({\and_addrb[12]_Naddrb_o_al_n73 ,addrb[11:10]}),
    .dia(dia[8:0]),
    .rstb(rstb),
    .dob({inst_dob_i46_008,inst_dob_i46_007,inst_dob_i46_006,inst_dob_i46_005,inst_dob_i46_004,inst_dob_i46_003,inst_dob_i46_002,inst_dob_i46_001,inst_dob_i46_000}));
  // address_offset=24576;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("INV"),
    .CSB1("INV"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_024576_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa({\and_Naddra[12]_addra_o_al_n86 ,addra[11:10]}),
    .csb({\and_Naddrb[12]_addrb_o_al_n89 ,addrb[11:10]}),
    .dia(dia[8:0]),
    .rstb(rstb),
    .dob({inst_dob_i48_008,inst_dob_i48_007,inst_dob_i48_006,inst_dob_i48_005,inst_dob_i48_004,inst_dob_i48_003,inst_dob_i48_002,inst_dob_i48_001,inst_dob_i48_000}));
  // address_offset=24576;data_offset=9;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("SIG"),
    .CSB1("SIG"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_024576_009 (
    .addra(addra[12:0]),
    .addrb(addrb[12:0]),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[15:13]),
    .csb(addrb[15:13]),
    .dia({open_n1441,open_n1442,open_n1443,open_n1444,open_n1445,open_n1446,open_n1447,dia[9],open_n1448}),
    .rstb(rstb),
    .dob({open_n1472,open_n1473,open_n1474,open_n1475,open_n1476,open_n1477,open_n1478,open_n1479,inst_dob_i48_009}));
  // address_offset=24576;data_offset=10;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("SIG"),
    .CSB1("SIG"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_024576_010 (
    .addra(addra[12:0]),
    .addrb(addrb[12:0]),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[15:13]),
    .csb(addrb[15:13]),
    .dia({open_n1480,open_n1481,open_n1482,open_n1483,open_n1484,open_n1485,open_n1486,dia[10],open_n1487}),
    .rstb(rstb),
    .dob({open_n1511,open_n1512,open_n1513,open_n1514,open_n1515,open_n1516,open_n1517,open_n1518,inst_dob_i48_010}));
  // address_offset=24576;data_offset=11;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("SIG"),
    .CSB1("SIG"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_024576_011 (
    .addra(addra[12:0]),
    .addrb(addrb[12:0]),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[15:13]),
    .csb(addrb[15:13]),
    .dia({open_n1519,open_n1520,open_n1521,open_n1522,open_n1523,open_n1524,open_n1525,dia[11],open_n1526}),
    .rstb(rstb),
    .dob({open_n1550,open_n1551,open_n1552,open_n1553,open_n1554,open_n1555,open_n1556,open_n1557,inst_dob_i48_011}));
  // address_offset=24576;data_offset=12;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("SIG"),
    .CSB1("SIG"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_024576_012 (
    .addra(addra[12:0]),
    .addrb(addrb[12:0]),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[15:13]),
    .csb(addrb[15:13]),
    .dia({open_n1558,open_n1559,open_n1560,open_n1561,open_n1562,open_n1563,open_n1564,dia[12],open_n1565}),
    .rstb(rstb),
    .dob({open_n1589,open_n1590,open_n1591,open_n1592,open_n1593,open_n1594,open_n1595,open_n1596,inst_dob_i48_012}));
  // address_offset=24576;data_offset=13;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("SIG"),
    .CSB1("SIG"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_024576_013 (
    .addra(addra[12:0]),
    .addrb(addrb[12:0]),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[15:13]),
    .csb(addrb[15:13]),
    .dia({open_n1597,open_n1598,open_n1599,open_n1600,open_n1601,open_n1602,open_n1603,dia[13],open_n1604}),
    .rstb(rstb),
    .dob({open_n1628,open_n1629,open_n1630,open_n1631,open_n1632,open_n1633,open_n1634,open_n1635,inst_dob_i48_013}));
  // address_offset=24576;data_offset=14;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("SIG"),
    .CSB1("SIG"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_024576_014 (
    .addra(addra[12:0]),
    .addrb(addrb[12:0]),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[15:13]),
    .csb(addrb[15:13]),
    .dia({open_n1636,open_n1637,open_n1638,open_n1639,open_n1640,open_n1641,open_n1642,dia[14],open_n1643}),
    .rstb(rstb),
    .dob({open_n1667,open_n1668,open_n1669,open_n1670,open_n1671,open_n1672,open_n1673,open_n1674,inst_dob_i48_014}));
  // address_offset=24576;data_offset=15;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("SIG"),
    .CSB1("SIG"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_024576_015 (
    .addra(addra[12:0]),
    .addrb(addrb[12:0]),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[15:13]),
    .csb(addrb[15:13]),
    .dia({open_n1675,open_n1676,open_n1677,open_n1678,open_n1679,open_n1680,open_n1681,dia[15],open_n1682}),
    .rstb(rstb),
    .dob({open_n1706,open_n1707,open_n1708,open_n1709,open_n1710,open_n1711,open_n1712,open_n1713,inst_dob_i48_015}));
  // address_offset=25600;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("SIG"),
    .CSB1("INV"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_025600_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa({\and_Naddra[12]_addra_o_al_n86 ,addra[11:10]}),
    .csb({\and_Naddrb[12]_addrb_o_al_n89 ,addrb[11:10]}),
    .dia(dia[8:0]),
    .rstb(rstb),
    .dob({inst_dob_i50_008,inst_dob_i50_007,inst_dob_i50_006,inst_dob_i50_005,inst_dob_i50_004,inst_dob_i50_003,inst_dob_i50_002,inst_dob_i50_001,inst_dob_i50_000}));
  // address_offset=26624;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("INV"),
    .CSB1("SIG"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_026624_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa({\and_Naddra[12]_addra_o_al_n86 ,addra[11:10]}),
    .csb({\and_Naddrb[12]_addrb_o_al_n89 ,addrb[11:10]}),
    .dia(dia[8:0]),
    .rstb(rstb),
    .dob({inst_dob_i52_008,inst_dob_i52_007,inst_dob_i52_006,inst_dob_i52_005,inst_dob_i52_004,inst_dob_i52_003,inst_dob_i52_002,inst_dob_i52_001,inst_dob_i52_000}));
  // address_offset=27648;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("SIG"),
    .CSB1("SIG"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_027648_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa({\and_Naddra[12]_addra_o_al_n86 ,addra[11:10]}),
    .csb({\and_Naddrb[12]_addrb_o_al_n89 ,addrb[11:10]}),
    .dia(dia[8:0]),
    .rstb(rstb),
    .dob({inst_dob_i54_008,inst_dob_i54_007,inst_dob_i54_006,inst_dob_i54_005,inst_dob_i54_004,inst_dob_i54_003,inst_dob_i54_002,inst_dob_i54_001,inst_dob_i54_000}));
  // address_offset=28672;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("INV"),
    .CSB1("INV"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_028672_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa({\and_addra[12]_addra[_o_al_n102 ,addra[11:10]}),
    .csb({\and_addrb[12]_addrb[_o_al_n105 ,addrb[11:10]}),
    .dia(dia[8:0]),
    .rstb(rstb),
    .dob({inst_dob_i56_008,inst_dob_i56_007,inst_dob_i56_006,inst_dob_i56_005,inst_dob_i56_004,inst_dob_i56_003,inst_dob_i56_002,inst_dob_i56_001,inst_dob_i56_000}));
  // address_offset=29696;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("SIG"),
    .CSB1("INV"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_029696_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa({\and_addra[12]_addra[_o_al_n102 ,addra[11:10]}),
    .csb({\and_addrb[12]_addrb[_o_al_n105 ,addrb[11:10]}),
    .dia(dia[8:0]),
    .rstb(rstb),
    .dob({inst_dob_i58_008,inst_dob_i58_007,inst_dob_i58_006,inst_dob_i58_005,inst_dob_i58_004,inst_dob_i58_003,inst_dob_i58_002,inst_dob_i58_001,inst_dob_i58_000}));
  // address_offset=30720;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("INV"),
    .CSB1("SIG"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_030720_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa({\and_addra[12]_addra[_o_al_n102 ,addra[11:10]}),
    .csb({\and_addrb[12]_addrb[_o_al_n105 ,addrb[11:10]}),
    .dia(dia[8:0]),
    .rstb(rstb),
    .dob({inst_dob_i60_008,inst_dob_i60_007,inst_dob_i60_006,inst_dob_i60_005,inst_dob_i60_004,inst_dob_i60_003,inst_dob_i60_002,inst_dob_i60_001,inst_dob_i60_000}));
  // address_offset=31744;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("SIG"),
    .CSB1("SIG"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_031744_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa({\and_addra[12]_addra[_o_al_n102 ,addra[11:10]}),
    .csb({\and_addrb[12]_addrb[_o_al_n105 ,addrb[11:10]}),
    .dia(dia[8:0]),
    .rstb(rstb),
    .dob({inst_dob_i62_008,inst_dob_i62_007,inst_dob_i62_006,inst_dob_i62_005,inst_dob_i62_004,inst_dob_i62_003,inst_dob_i62_002,inst_dob_i62_001,inst_dob_i62_000}));
  // address_offset=32768;data_offset=0;depth=32;width=16;num_section=1;width_per_section=16;section_size=16;working_depth=512;working_width=18;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("1"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("INV"),
    .CSB1("INV"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("18"),
    .DATA_WIDTH_B("18"),
    .MODE("PDPW8K"),
    .OCEAMUX("1"),
    .OCEBMUX("1"),
    .REGMODE_A("OUTREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_032768_000 (
    .addra({addra[8:0],4'b1111}),
    .addrb({addrb[8:0],4'b1111}),
    .clka(clka),
    .clkb(clkb),
    .csa({\and_Naddra[11]_Naddr_o_and_cea ,addra[10:9]}),
    .csb({\and_Naddrb[11]_Naddr_o_and_ceb ,addrb[10:9]}),
    .dia(dia[8:0]),
    .dib({open_n1877,open_n1878,dia[15:9]}),
    .rstb(rstb),
    .doa({inst_dob_i64_008,inst_dob_i64_007,inst_dob_i64_006,inst_dob_i64_005,inst_dob_i64_004,inst_dob_i64_003,inst_dob_i64_002,inst_dob_i64_001,inst_dob_i64_000}),
    .dob({open_n1884,open_n1885,inst_dob_i64_015,inst_dob_i64_014,inst_dob_i64_013,inst_dob_i64_012,inst_dob_i64_011,inst_dob_i64_010,inst_dob_i64_009}));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_0  (
    .i0(inst_dob_i0_000),
    .i1(inst_dob_i0_000),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b0/B0_0 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_1  (
    .i0(inst_dob_i2_000),
    .i1(inst_dob_i2_000),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b0/B0_1 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_10  (
    .i0(inst_dob_i20_000),
    .i1(inst_dob_i20_000),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b0/B0_10 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_11  (
    .i0(inst_dob_i22_000),
    .i1(inst_dob_i22_000),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b0/B0_11 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_12  (
    .i0(inst_dob_i24_000),
    .i1(inst_dob_i24_000),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b0/B0_12 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_13  (
    .i0(inst_dob_i26_000),
    .i1(inst_dob_i26_000),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b0/B0_13 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_14  (
    .i0(inst_dob_i28_000),
    .i1(inst_dob_i28_000),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b0/B0_14 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_15  (
    .i0(inst_dob_i30_000),
    .i1(inst_dob_i30_000),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b0/B0_15 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_16  (
    .i0(inst_dob_i32_000),
    .i1(inst_dob_i32_000),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b0/B0_16 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_17  (
    .i0(inst_dob_i34_000),
    .i1(inst_dob_i34_000),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b0/B0_17 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_18  (
    .i0(inst_dob_i36_000),
    .i1(inst_dob_i36_000),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b0/B0_18 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_19  (
    .i0(inst_dob_i38_000),
    .i1(inst_dob_i38_000),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b0/B0_19 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_2  (
    .i0(inst_dob_i4_000),
    .i1(inst_dob_i4_000),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b0/B0_2 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_20  (
    .i0(inst_dob_i40_000),
    .i1(inst_dob_i40_000),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b0/B0_20 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_21  (
    .i0(inst_dob_i42_000),
    .i1(inst_dob_i42_000),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b0/B0_21 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_22  (
    .i0(inst_dob_i44_000),
    .i1(inst_dob_i44_000),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b0/B0_22 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_23  (
    .i0(inst_dob_i46_000),
    .i1(inst_dob_i46_000),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b0/B0_23 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_24  (
    .i0(inst_dob_i48_000),
    .i1(inst_dob_i48_000),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b0/B0_24 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_25  (
    .i0(inst_dob_i50_000),
    .i1(inst_dob_i50_000),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b0/B0_25 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_26  (
    .i0(inst_dob_i52_000),
    .i1(inst_dob_i52_000),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b0/B0_26 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_27  (
    .i0(inst_dob_i54_000),
    .i1(inst_dob_i54_000),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b0/B0_27 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_28  (
    .i0(inst_dob_i56_000),
    .i1(inst_dob_i56_000),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b0/B0_28 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_29  (
    .i0(inst_dob_i58_000),
    .i1(inst_dob_i58_000),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b0/B0_29 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_3  (
    .i0(inst_dob_i6_000),
    .i1(inst_dob_i6_000),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b0/B0_3 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_30  (
    .i0(inst_dob_i60_000),
    .i1(inst_dob_i60_000),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b0/B0_30 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_31  (
    .i0(inst_dob_i62_000),
    .i1(inst_dob_i62_000),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b0/B0_31 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_32  (
    .i0(inst_dob_i64_000),
    .i1(inst_dob_i64_000),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b0/B0_32 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_33  (
    .i0(inst_dob_i64_000),
    .i1(inst_dob_i64_000),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b0/B0_33 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_34  (
    .i0(inst_dob_i64_000),
    .i1(inst_dob_i64_000),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b0/B0_34 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_35  (
    .i0(inst_dob_i64_000),
    .i1(inst_dob_i64_000),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b0/B0_35 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_36  (
    .i0(inst_dob_i64_000),
    .i1(inst_dob_i64_000),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b0/B0_36 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_37  (
    .i0(inst_dob_i64_000),
    .i1(inst_dob_i64_000),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b0/B0_37 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_38  (
    .i0(inst_dob_i64_000),
    .i1(inst_dob_i64_000),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b0/B0_38 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_39  (
    .i0(inst_dob_i64_000),
    .i1(inst_dob_i64_000),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b0/B0_39 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_4  (
    .i0(inst_dob_i8_000),
    .i1(inst_dob_i8_000),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b0/B0_4 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_40  (
    .i0(inst_dob_i64_000),
    .i1(inst_dob_i64_000),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b0/B0_40 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_41  (
    .i0(inst_dob_i64_000),
    .i1(inst_dob_i64_000),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b0/B0_41 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_42  (
    .i0(inst_dob_i64_000),
    .i1(inst_dob_i64_000),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b0/B0_42 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_43  (
    .i0(inst_dob_i64_000),
    .i1(inst_dob_i64_000),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b0/B0_43 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_44  (
    .i0(inst_dob_i64_000),
    .i1(inst_dob_i64_000),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b0/B0_44 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_45  (
    .i0(inst_dob_i64_000),
    .i1(inst_dob_i64_000),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b0/B0_45 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_46  (
    .i0(inst_dob_i64_000),
    .i1(inst_dob_i64_000),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b0/B0_46 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_47  (
    .i0(inst_dob_i64_000),
    .i1(inst_dob_i64_000),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b0/B0_47 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_48  (
    .i0(inst_dob_i64_000),
    .i1(inst_dob_i64_000),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b0/B0_48 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_49  (
    .i0(inst_dob_i64_000),
    .i1(inst_dob_i64_000),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b0/B0_49 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_5  (
    .i0(inst_dob_i10_000),
    .i1(inst_dob_i10_000),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b0/B0_5 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_50  (
    .i0(inst_dob_i64_000),
    .i1(inst_dob_i64_000),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b0/B0_50 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_51  (
    .i0(inst_dob_i64_000),
    .i1(inst_dob_i64_000),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b0/B0_51 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_52  (
    .i0(inst_dob_i64_000),
    .i1(inst_dob_i64_000),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b0/B0_52 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_53  (
    .i0(inst_dob_i64_000),
    .i1(inst_dob_i64_000),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b0/B0_53 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_54  (
    .i0(inst_dob_i64_000),
    .i1(inst_dob_i64_000),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b0/B0_54 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_55  (
    .i0(inst_dob_i64_000),
    .i1(inst_dob_i64_000),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b0/B0_55 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_56  (
    .i0(inst_dob_i64_000),
    .i1(inst_dob_i64_000),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b0/B0_56 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_57  (
    .i0(inst_dob_i64_000),
    .i1(inst_dob_i64_000),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b0/B0_57 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_58  (
    .i0(inst_dob_i64_000),
    .i1(inst_dob_i64_000),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b0/B0_58 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_59  (
    .i0(inst_dob_i64_000),
    .i1(inst_dob_i64_000),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b0/B0_59 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_6  (
    .i0(inst_dob_i12_000),
    .i1(inst_dob_i12_000),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b0/B0_6 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_60  (
    .i0(inst_dob_i64_000),
    .i1(inst_dob_i64_000),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b0/B0_60 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_61  (
    .i0(inst_dob_i64_000),
    .i1(inst_dob_i64_000),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b0/B0_61 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_62  (
    .i0(inst_dob_i64_000),
    .i1(inst_dob_i64_000),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b0/B0_62 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_63  (
    .i0(inst_dob_i64_000),
    .i1(inst_dob_i64_000),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b0/B0_63 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_7  (
    .i0(inst_dob_i14_000),
    .i1(inst_dob_i14_000),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b0/B0_7 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_8  (
    .i0(inst_dob_i16_000),
    .i1(inst_dob_i16_000),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b0/B0_8 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_9  (
    .i0(inst_dob_i18_000),
    .i1(inst_dob_i18_000),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b0/B0_9 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_1_0  (
    .i0(\inst_dob_mux_b0/B0_0 ),
    .i1(\inst_dob_mux_b0/B0_1 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b0/B1_0 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_1_1  (
    .i0(\inst_dob_mux_b0/B0_2 ),
    .i1(\inst_dob_mux_b0/B0_3 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b0/B1_1 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_1_10  (
    .i0(\inst_dob_mux_b0/B0_20 ),
    .i1(\inst_dob_mux_b0/B0_21 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b0/B1_10 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_1_11  (
    .i0(\inst_dob_mux_b0/B0_22 ),
    .i1(\inst_dob_mux_b0/B0_23 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b0/B1_11 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_1_12  (
    .i0(\inst_dob_mux_b0/B0_24 ),
    .i1(\inst_dob_mux_b0/B0_25 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b0/B1_12 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_1_13  (
    .i0(\inst_dob_mux_b0/B0_26 ),
    .i1(\inst_dob_mux_b0/B0_27 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b0/B1_13 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_1_14  (
    .i0(\inst_dob_mux_b0/B0_28 ),
    .i1(\inst_dob_mux_b0/B0_29 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b0/B1_14 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_1_15  (
    .i0(\inst_dob_mux_b0/B0_30 ),
    .i1(\inst_dob_mux_b0/B0_31 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b0/B1_15 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_1_16  (
    .i0(\inst_dob_mux_b0/B0_32 ),
    .i1(\inst_dob_mux_b0/B0_33 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b0/B1_16 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_1_17  (
    .i0(\inst_dob_mux_b0/B0_34 ),
    .i1(\inst_dob_mux_b0/B0_35 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b0/B1_17 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_1_18  (
    .i0(\inst_dob_mux_b0/B0_36 ),
    .i1(\inst_dob_mux_b0/B0_37 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b0/B1_18 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_1_19  (
    .i0(\inst_dob_mux_b0/B0_38 ),
    .i1(\inst_dob_mux_b0/B0_39 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b0/B1_19 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_1_2  (
    .i0(\inst_dob_mux_b0/B0_4 ),
    .i1(\inst_dob_mux_b0/B0_5 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b0/B1_2 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_1_20  (
    .i0(\inst_dob_mux_b0/B0_40 ),
    .i1(\inst_dob_mux_b0/B0_41 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b0/B1_20 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_1_21  (
    .i0(\inst_dob_mux_b0/B0_42 ),
    .i1(\inst_dob_mux_b0/B0_43 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b0/B1_21 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_1_22  (
    .i0(\inst_dob_mux_b0/B0_44 ),
    .i1(\inst_dob_mux_b0/B0_45 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b0/B1_22 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_1_23  (
    .i0(\inst_dob_mux_b0/B0_46 ),
    .i1(\inst_dob_mux_b0/B0_47 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b0/B1_23 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_1_24  (
    .i0(\inst_dob_mux_b0/B0_48 ),
    .i1(\inst_dob_mux_b0/B0_49 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b0/B1_24 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_1_25  (
    .i0(\inst_dob_mux_b0/B0_50 ),
    .i1(\inst_dob_mux_b0/B0_51 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b0/B1_25 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_1_26  (
    .i0(\inst_dob_mux_b0/B0_52 ),
    .i1(\inst_dob_mux_b0/B0_53 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b0/B1_26 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_1_27  (
    .i0(\inst_dob_mux_b0/B0_54 ),
    .i1(\inst_dob_mux_b0/B0_55 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b0/B1_27 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_1_28  (
    .i0(\inst_dob_mux_b0/B0_56 ),
    .i1(\inst_dob_mux_b0/B0_57 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b0/B1_28 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_1_29  (
    .i0(\inst_dob_mux_b0/B0_58 ),
    .i1(\inst_dob_mux_b0/B0_59 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b0/B1_29 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_1_3  (
    .i0(\inst_dob_mux_b0/B0_6 ),
    .i1(\inst_dob_mux_b0/B0_7 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b0/B1_3 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_1_30  (
    .i0(\inst_dob_mux_b0/B0_60 ),
    .i1(\inst_dob_mux_b0/B0_61 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b0/B1_30 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_1_31  (
    .i0(\inst_dob_mux_b0/B0_62 ),
    .i1(\inst_dob_mux_b0/B0_63 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b0/B1_31 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_1_4  (
    .i0(\inst_dob_mux_b0/B0_8 ),
    .i1(\inst_dob_mux_b0/B0_9 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b0/B1_4 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_1_5  (
    .i0(\inst_dob_mux_b0/B0_10 ),
    .i1(\inst_dob_mux_b0/B0_11 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b0/B1_5 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_1_6  (
    .i0(\inst_dob_mux_b0/B0_12 ),
    .i1(\inst_dob_mux_b0/B0_13 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b0/B1_6 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_1_7  (
    .i0(\inst_dob_mux_b0/B0_14 ),
    .i1(\inst_dob_mux_b0/B0_15 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b0/B1_7 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_1_8  (
    .i0(\inst_dob_mux_b0/B0_16 ),
    .i1(\inst_dob_mux_b0/B0_17 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b0/B1_8 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_1_9  (
    .i0(\inst_dob_mux_b0/B0_18 ),
    .i1(\inst_dob_mux_b0/B0_19 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b0/B1_9 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_2_0  (
    .i0(\inst_dob_mux_b0/B1_0 ),
    .i1(\inst_dob_mux_b0/B1_1 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b0/B2_0 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_2_1  (
    .i0(\inst_dob_mux_b0/B1_2 ),
    .i1(\inst_dob_mux_b0/B1_3 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b0/B2_1 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_2_10  (
    .i0(\inst_dob_mux_b0/B1_20 ),
    .i1(\inst_dob_mux_b0/B1_21 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b0/B2_10 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_2_11  (
    .i0(\inst_dob_mux_b0/B1_22 ),
    .i1(\inst_dob_mux_b0/B1_23 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b0/B2_11 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_2_12  (
    .i0(\inst_dob_mux_b0/B1_24 ),
    .i1(\inst_dob_mux_b0/B1_25 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b0/B2_12 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_2_13  (
    .i0(\inst_dob_mux_b0/B1_26 ),
    .i1(\inst_dob_mux_b0/B1_27 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b0/B2_13 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_2_14  (
    .i0(\inst_dob_mux_b0/B1_28 ),
    .i1(\inst_dob_mux_b0/B1_29 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b0/B2_14 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_2_15  (
    .i0(\inst_dob_mux_b0/B1_30 ),
    .i1(\inst_dob_mux_b0/B1_31 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b0/B2_15 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_2_2  (
    .i0(\inst_dob_mux_b0/B1_4 ),
    .i1(\inst_dob_mux_b0/B1_5 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b0/B2_2 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_2_3  (
    .i0(\inst_dob_mux_b0/B1_6 ),
    .i1(\inst_dob_mux_b0/B1_7 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b0/B2_3 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_2_4  (
    .i0(\inst_dob_mux_b0/B1_8 ),
    .i1(\inst_dob_mux_b0/B1_9 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b0/B2_4 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_2_5  (
    .i0(\inst_dob_mux_b0/B1_10 ),
    .i1(\inst_dob_mux_b0/B1_11 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b0/B2_5 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_2_6  (
    .i0(\inst_dob_mux_b0/B1_12 ),
    .i1(\inst_dob_mux_b0/B1_13 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b0/B2_6 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_2_7  (
    .i0(\inst_dob_mux_b0/B1_14 ),
    .i1(\inst_dob_mux_b0/B1_15 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b0/B2_7 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_2_8  (
    .i0(\inst_dob_mux_b0/B1_16 ),
    .i1(\inst_dob_mux_b0/B1_17 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b0/B2_8 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_2_9  (
    .i0(\inst_dob_mux_b0/B1_18 ),
    .i1(\inst_dob_mux_b0/B1_19 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b0/B2_9 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_3_0  (
    .i0(\inst_dob_mux_b0/B2_0 ),
    .i1(\inst_dob_mux_b0/B2_1 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b0/B3_0 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_3_1  (
    .i0(\inst_dob_mux_b0/B2_2 ),
    .i1(\inst_dob_mux_b0/B2_3 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b0/B3_1 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_3_2  (
    .i0(\inst_dob_mux_b0/B2_4 ),
    .i1(\inst_dob_mux_b0/B2_5 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b0/B3_2 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_3_3  (
    .i0(\inst_dob_mux_b0/B2_6 ),
    .i1(\inst_dob_mux_b0/B2_7 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b0/B3_3 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_3_4  (
    .i0(\inst_dob_mux_b0/B2_8 ),
    .i1(\inst_dob_mux_b0/B2_9 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b0/B3_4 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_3_5  (
    .i0(\inst_dob_mux_b0/B2_10 ),
    .i1(\inst_dob_mux_b0/B2_11 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b0/B3_5 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_3_6  (
    .i0(\inst_dob_mux_b0/B2_12 ),
    .i1(\inst_dob_mux_b0/B2_13 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b0/B3_6 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_3_7  (
    .i0(\inst_dob_mux_b0/B2_14 ),
    .i1(\inst_dob_mux_b0/B2_15 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b0/B3_7 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_4_0  (
    .i0(\inst_dob_mux_b0/B3_0 ),
    .i1(\inst_dob_mux_b0/B3_1 ),
    .sel(addrb_piped_piped[4]),
    .o(\inst_dob_mux_b0/B4_0 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_4_1  (
    .i0(\inst_dob_mux_b0/B3_2 ),
    .i1(\inst_dob_mux_b0/B3_3 ),
    .sel(addrb_piped_piped[4]),
    .o(\inst_dob_mux_b0/B4_1 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_4_2  (
    .i0(\inst_dob_mux_b0/B3_4 ),
    .i1(\inst_dob_mux_b0/B3_5 ),
    .sel(addrb_piped_piped[4]),
    .o(\inst_dob_mux_b0/B4_2 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_4_3  (
    .i0(\inst_dob_mux_b0/B3_6 ),
    .i1(\inst_dob_mux_b0/B3_7 ),
    .sel(addrb_piped_piped[4]),
    .o(\inst_dob_mux_b0/B4_3 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_5_0  (
    .i0(\inst_dob_mux_b0/B4_0 ),
    .i1(\inst_dob_mux_b0/B4_1 ),
    .sel(addrb_piped_piped[5]),
    .o(\inst_dob_mux_b0/B5_0 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_5_1  (
    .i0(\inst_dob_mux_b0/B4_2 ),
    .i1(\inst_dob_mux_b0/B4_3 ),
    .sel(addrb_piped_piped[5]),
    .o(\inst_dob_mux_b0/B5_1 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_6_0  (
    .i0(\inst_dob_mux_b0/B5_0 ),
    .i1(\inst_dob_mux_b0/B5_1 ),
    .sel(addrb_piped_piped[6]),
    .o(dob[0]));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_0  (
    .i0(inst_dob_i0_001),
    .i1(inst_dob_i0_001),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b1/B0_0 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_1  (
    .i0(inst_dob_i2_001),
    .i1(inst_dob_i2_001),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b1/B0_1 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_10  (
    .i0(inst_dob_i20_001),
    .i1(inst_dob_i20_001),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b1/B0_10 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_11  (
    .i0(inst_dob_i22_001),
    .i1(inst_dob_i22_001),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b1/B0_11 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_12  (
    .i0(inst_dob_i24_001),
    .i1(inst_dob_i24_001),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b1/B0_12 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_13  (
    .i0(inst_dob_i26_001),
    .i1(inst_dob_i26_001),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b1/B0_13 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_14  (
    .i0(inst_dob_i28_001),
    .i1(inst_dob_i28_001),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b1/B0_14 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_15  (
    .i0(inst_dob_i30_001),
    .i1(inst_dob_i30_001),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b1/B0_15 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_16  (
    .i0(inst_dob_i32_001),
    .i1(inst_dob_i32_001),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b1/B0_16 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_17  (
    .i0(inst_dob_i34_001),
    .i1(inst_dob_i34_001),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b1/B0_17 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_18  (
    .i0(inst_dob_i36_001),
    .i1(inst_dob_i36_001),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b1/B0_18 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_19  (
    .i0(inst_dob_i38_001),
    .i1(inst_dob_i38_001),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b1/B0_19 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_2  (
    .i0(inst_dob_i4_001),
    .i1(inst_dob_i4_001),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b1/B0_2 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_20  (
    .i0(inst_dob_i40_001),
    .i1(inst_dob_i40_001),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b1/B0_20 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_21  (
    .i0(inst_dob_i42_001),
    .i1(inst_dob_i42_001),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b1/B0_21 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_22  (
    .i0(inst_dob_i44_001),
    .i1(inst_dob_i44_001),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b1/B0_22 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_23  (
    .i0(inst_dob_i46_001),
    .i1(inst_dob_i46_001),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b1/B0_23 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_24  (
    .i0(inst_dob_i48_001),
    .i1(inst_dob_i48_001),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b1/B0_24 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_25  (
    .i0(inst_dob_i50_001),
    .i1(inst_dob_i50_001),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b1/B0_25 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_26  (
    .i0(inst_dob_i52_001),
    .i1(inst_dob_i52_001),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b1/B0_26 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_27  (
    .i0(inst_dob_i54_001),
    .i1(inst_dob_i54_001),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b1/B0_27 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_28  (
    .i0(inst_dob_i56_001),
    .i1(inst_dob_i56_001),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b1/B0_28 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_29  (
    .i0(inst_dob_i58_001),
    .i1(inst_dob_i58_001),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b1/B0_29 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_3  (
    .i0(inst_dob_i6_001),
    .i1(inst_dob_i6_001),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b1/B0_3 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_30  (
    .i0(inst_dob_i60_001),
    .i1(inst_dob_i60_001),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b1/B0_30 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_31  (
    .i0(inst_dob_i62_001),
    .i1(inst_dob_i62_001),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b1/B0_31 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_32  (
    .i0(inst_dob_i64_001),
    .i1(inst_dob_i64_001),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b1/B0_32 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_33  (
    .i0(inst_dob_i64_001),
    .i1(inst_dob_i64_001),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b1/B0_33 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_34  (
    .i0(inst_dob_i64_001),
    .i1(inst_dob_i64_001),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b1/B0_34 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_35  (
    .i0(inst_dob_i64_001),
    .i1(inst_dob_i64_001),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b1/B0_35 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_36  (
    .i0(inst_dob_i64_001),
    .i1(inst_dob_i64_001),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b1/B0_36 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_37  (
    .i0(inst_dob_i64_001),
    .i1(inst_dob_i64_001),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b1/B0_37 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_38  (
    .i0(inst_dob_i64_001),
    .i1(inst_dob_i64_001),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b1/B0_38 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_39  (
    .i0(inst_dob_i64_001),
    .i1(inst_dob_i64_001),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b1/B0_39 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_4  (
    .i0(inst_dob_i8_001),
    .i1(inst_dob_i8_001),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b1/B0_4 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_40  (
    .i0(inst_dob_i64_001),
    .i1(inst_dob_i64_001),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b1/B0_40 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_41  (
    .i0(inst_dob_i64_001),
    .i1(inst_dob_i64_001),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b1/B0_41 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_42  (
    .i0(inst_dob_i64_001),
    .i1(inst_dob_i64_001),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b1/B0_42 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_43  (
    .i0(inst_dob_i64_001),
    .i1(inst_dob_i64_001),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b1/B0_43 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_44  (
    .i0(inst_dob_i64_001),
    .i1(inst_dob_i64_001),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b1/B0_44 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_45  (
    .i0(inst_dob_i64_001),
    .i1(inst_dob_i64_001),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b1/B0_45 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_46  (
    .i0(inst_dob_i64_001),
    .i1(inst_dob_i64_001),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b1/B0_46 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_47  (
    .i0(inst_dob_i64_001),
    .i1(inst_dob_i64_001),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b1/B0_47 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_48  (
    .i0(inst_dob_i64_001),
    .i1(inst_dob_i64_001),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b1/B0_48 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_49  (
    .i0(inst_dob_i64_001),
    .i1(inst_dob_i64_001),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b1/B0_49 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_5  (
    .i0(inst_dob_i10_001),
    .i1(inst_dob_i10_001),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b1/B0_5 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_50  (
    .i0(inst_dob_i64_001),
    .i1(inst_dob_i64_001),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b1/B0_50 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_51  (
    .i0(inst_dob_i64_001),
    .i1(inst_dob_i64_001),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b1/B0_51 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_52  (
    .i0(inst_dob_i64_001),
    .i1(inst_dob_i64_001),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b1/B0_52 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_53  (
    .i0(inst_dob_i64_001),
    .i1(inst_dob_i64_001),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b1/B0_53 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_54  (
    .i0(inst_dob_i64_001),
    .i1(inst_dob_i64_001),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b1/B0_54 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_55  (
    .i0(inst_dob_i64_001),
    .i1(inst_dob_i64_001),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b1/B0_55 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_56  (
    .i0(inst_dob_i64_001),
    .i1(inst_dob_i64_001),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b1/B0_56 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_57  (
    .i0(inst_dob_i64_001),
    .i1(inst_dob_i64_001),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b1/B0_57 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_58  (
    .i0(inst_dob_i64_001),
    .i1(inst_dob_i64_001),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b1/B0_58 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_59  (
    .i0(inst_dob_i64_001),
    .i1(inst_dob_i64_001),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b1/B0_59 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_6  (
    .i0(inst_dob_i12_001),
    .i1(inst_dob_i12_001),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b1/B0_6 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_60  (
    .i0(inst_dob_i64_001),
    .i1(inst_dob_i64_001),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b1/B0_60 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_61  (
    .i0(inst_dob_i64_001),
    .i1(inst_dob_i64_001),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b1/B0_61 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_62  (
    .i0(inst_dob_i64_001),
    .i1(inst_dob_i64_001),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b1/B0_62 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_63  (
    .i0(inst_dob_i64_001),
    .i1(inst_dob_i64_001),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b1/B0_63 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_7  (
    .i0(inst_dob_i14_001),
    .i1(inst_dob_i14_001),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b1/B0_7 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_8  (
    .i0(inst_dob_i16_001),
    .i1(inst_dob_i16_001),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b1/B0_8 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_9  (
    .i0(inst_dob_i18_001),
    .i1(inst_dob_i18_001),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b1/B0_9 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_1_0  (
    .i0(\inst_dob_mux_b1/B0_0 ),
    .i1(\inst_dob_mux_b1/B0_1 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b1/B1_0 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_1_1  (
    .i0(\inst_dob_mux_b1/B0_2 ),
    .i1(\inst_dob_mux_b1/B0_3 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b1/B1_1 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_1_10  (
    .i0(\inst_dob_mux_b1/B0_20 ),
    .i1(\inst_dob_mux_b1/B0_21 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b1/B1_10 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_1_11  (
    .i0(\inst_dob_mux_b1/B0_22 ),
    .i1(\inst_dob_mux_b1/B0_23 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b1/B1_11 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_1_12  (
    .i0(\inst_dob_mux_b1/B0_24 ),
    .i1(\inst_dob_mux_b1/B0_25 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b1/B1_12 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_1_13  (
    .i0(\inst_dob_mux_b1/B0_26 ),
    .i1(\inst_dob_mux_b1/B0_27 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b1/B1_13 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_1_14  (
    .i0(\inst_dob_mux_b1/B0_28 ),
    .i1(\inst_dob_mux_b1/B0_29 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b1/B1_14 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_1_15  (
    .i0(\inst_dob_mux_b1/B0_30 ),
    .i1(\inst_dob_mux_b1/B0_31 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b1/B1_15 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_1_16  (
    .i0(\inst_dob_mux_b1/B0_32 ),
    .i1(\inst_dob_mux_b1/B0_33 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b1/B1_16 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_1_17  (
    .i0(\inst_dob_mux_b1/B0_34 ),
    .i1(\inst_dob_mux_b1/B0_35 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b1/B1_17 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_1_18  (
    .i0(\inst_dob_mux_b1/B0_36 ),
    .i1(\inst_dob_mux_b1/B0_37 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b1/B1_18 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_1_19  (
    .i0(\inst_dob_mux_b1/B0_38 ),
    .i1(\inst_dob_mux_b1/B0_39 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b1/B1_19 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_1_2  (
    .i0(\inst_dob_mux_b1/B0_4 ),
    .i1(\inst_dob_mux_b1/B0_5 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b1/B1_2 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_1_20  (
    .i0(\inst_dob_mux_b1/B0_40 ),
    .i1(\inst_dob_mux_b1/B0_41 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b1/B1_20 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_1_21  (
    .i0(\inst_dob_mux_b1/B0_42 ),
    .i1(\inst_dob_mux_b1/B0_43 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b1/B1_21 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_1_22  (
    .i0(\inst_dob_mux_b1/B0_44 ),
    .i1(\inst_dob_mux_b1/B0_45 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b1/B1_22 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_1_23  (
    .i0(\inst_dob_mux_b1/B0_46 ),
    .i1(\inst_dob_mux_b1/B0_47 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b1/B1_23 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_1_24  (
    .i0(\inst_dob_mux_b1/B0_48 ),
    .i1(\inst_dob_mux_b1/B0_49 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b1/B1_24 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_1_25  (
    .i0(\inst_dob_mux_b1/B0_50 ),
    .i1(\inst_dob_mux_b1/B0_51 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b1/B1_25 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_1_26  (
    .i0(\inst_dob_mux_b1/B0_52 ),
    .i1(\inst_dob_mux_b1/B0_53 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b1/B1_26 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_1_27  (
    .i0(\inst_dob_mux_b1/B0_54 ),
    .i1(\inst_dob_mux_b1/B0_55 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b1/B1_27 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_1_28  (
    .i0(\inst_dob_mux_b1/B0_56 ),
    .i1(\inst_dob_mux_b1/B0_57 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b1/B1_28 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_1_29  (
    .i0(\inst_dob_mux_b1/B0_58 ),
    .i1(\inst_dob_mux_b1/B0_59 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b1/B1_29 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_1_3  (
    .i0(\inst_dob_mux_b1/B0_6 ),
    .i1(\inst_dob_mux_b1/B0_7 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b1/B1_3 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_1_30  (
    .i0(\inst_dob_mux_b1/B0_60 ),
    .i1(\inst_dob_mux_b1/B0_61 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b1/B1_30 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_1_31  (
    .i0(\inst_dob_mux_b1/B0_62 ),
    .i1(\inst_dob_mux_b1/B0_63 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b1/B1_31 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_1_4  (
    .i0(\inst_dob_mux_b1/B0_8 ),
    .i1(\inst_dob_mux_b1/B0_9 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b1/B1_4 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_1_5  (
    .i0(\inst_dob_mux_b1/B0_10 ),
    .i1(\inst_dob_mux_b1/B0_11 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b1/B1_5 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_1_6  (
    .i0(\inst_dob_mux_b1/B0_12 ),
    .i1(\inst_dob_mux_b1/B0_13 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b1/B1_6 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_1_7  (
    .i0(\inst_dob_mux_b1/B0_14 ),
    .i1(\inst_dob_mux_b1/B0_15 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b1/B1_7 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_1_8  (
    .i0(\inst_dob_mux_b1/B0_16 ),
    .i1(\inst_dob_mux_b1/B0_17 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b1/B1_8 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_1_9  (
    .i0(\inst_dob_mux_b1/B0_18 ),
    .i1(\inst_dob_mux_b1/B0_19 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b1/B1_9 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_2_0  (
    .i0(\inst_dob_mux_b1/B1_0 ),
    .i1(\inst_dob_mux_b1/B1_1 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b1/B2_0 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_2_1  (
    .i0(\inst_dob_mux_b1/B1_2 ),
    .i1(\inst_dob_mux_b1/B1_3 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b1/B2_1 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_2_10  (
    .i0(\inst_dob_mux_b1/B1_20 ),
    .i1(\inst_dob_mux_b1/B1_21 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b1/B2_10 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_2_11  (
    .i0(\inst_dob_mux_b1/B1_22 ),
    .i1(\inst_dob_mux_b1/B1_23 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b1/B2_11 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_2_12  (
    .i0(\inst_dob_mux_b1/B1_24 ),
    .i1(\inst_dob_mux_b1/B1_25 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b1/B2_12 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_2_13  (
    .i0(\inst_dob_mux_b1/B1_26 ),
    .i1(\inst_dob_mux_b1/B1_27 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b1/B2_13 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_2_14  (
    .i0(\inst_dob_mux_b1/B1_28 ),
    .i1(\inst_dob_mux_b1/B1_29 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b1/B2_14 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_2_15  (
    .i0(\inst_dob_mux_b1/B1_30 ),
    .i1(\inst_dob_mux_b1/B1_31 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b1/B2_15 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_2_2  (
    .i0(\inst_dob_mux_b1/B1_4 ),
    .i1(\inst_dob_mux_b1/B1_5 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b1/B2_2 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_2_3  (
    .i0(\inst_dob_mux_b1/B1_6 ),
    .i1(\inst_dob_mux_b1/B1_7 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b1/B2_3 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_2_4  (
    .i0(\inst_dob_mux_b1/B1_8 ),
    .i1(\inst_dob_mux_b1/B1_9 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b1/B2_4 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_2_5  (
    .i0(\inst_dob_mux_b1/B1_10 ),
    .i1(\inst_dob_mux_b1/B1_11 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b1/B2_5 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_2_6  (
    .i0(\inst_dob_mux_b1/B1_12 ),
    .i1(\inst_dob_mux_b1/B1_13 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b1/B2_6 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_2_7  (
    .i0(\inst_dob_mux_b1/B1_14 ),
    .i1(\inst_dob_mux_b1/B1_15 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b1/B2_7 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_2_8  (
    .i0(\inst_dob_mux_b1/B1_16 ),
    .i1(\inst_dob_mux_b1/B1_17 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b1/B2_8 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_2_9  (
    .i0(\inst_dob_mux_b1/B1_18 ),
    .i1(\inst_dob_mux_b1/B1_19 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b1/B2_9 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_3_0  (
    .i0(\inst_dob_mux_b1/B2_0 ),
    .i1(\inst_dob_mux_b1/B2_1 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b1/B3_0 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_3_1  (
    .i0(\inst_dob_mux_b1/B2_2 ),
    .i1(\inst_dob_mux_b1/B2_3 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b1/B3_1 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_3_2  (
    .i0(\inst_dob_mux_b1/B2_4 ),
    .i1(\inst_dob_mux_b1/B2_5 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b1/B3_2 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_3_3  (
    .i0(\inst_dob_mux_b1/B2_6 ),
    .i1(\inst_dob_mux_b1/B2_7 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b1/B3_3 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_3_4  (
    .i0(\inst_dob_mux_b1/B2_8 ),
    .i1(\inst_dob_mux_b1/B2_9 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b1/B3_4 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_3_5  (
    .i0(\inst_dob_mux_b1/B2_10 ),
    .i1(\inst_dob_mux_b1/B2_11 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b1/B3_5 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_3_6  (
    .i0(\inst_dob_mux_b1/B2_12 ),
    .i1(\inst_dob_mux_b1/B2_13 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b1/B3_6 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_3_7  (
    .i0(\inst_dob_mux_b1/B2_14 ),
    .i1(\inst_dob_mux_b1/B2_15 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b1/B3_7 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_4_0  (
    .i0(\inst_dob_mux_b1/B3_0 ),
    .i1(\inst_dob_mux_b1/B3_1 ),
    .sel(addrb_piped_piped[4]),
    .o(\inst_dob_mux_b1/B4_0 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_4_1  (
    .i0(\inst_dob_mux_b1/B3_2 ),
    .i1(\inst_dob_mux_b1/B3_3 ),
    .sel(addrb_piped_piped[4]),
    .o(\inst_dob_mux_b1/B4_1 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_4_2  (
    .i0(\inst_dob_mux_b1/B3_4 ),
    .i1(\inst_dob_mux_b1/B3_5 ),
    .sel(addrb_piped_piped[4]),
    .o(\inst_dob_mux_b1/B4_2 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_4_3  (
    .i0(\inst_dob_mux_b1/B3_6 ),
    .i1(\inst_dob_mux_b1/B3_7 ),
    .sel(addrb_piped_piped[4]),
    .o(\inst_dob_mux_b1/B4_3 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_5_0  (
    .i0(\inst_dob_mux_b1/B4_0 ),
    .i1(\inst_dob_mux_b1/B4_1 ),
    .sel(addrb_piped_piped[5]),
    .o(\inst_dob_mux_b1/B5_0 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_5_1  (
    .i0(\inst_dob_mux_b1/B4_2 ),
    .i1(\inst_dob_mux_b1/B4_3 ),
    .sel(addrb_piped_piped[5]),
    .o(\inst_dob_mux_b1/B5_1 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_6_0  (
    .i0(\inst_dob_mux_b1/B5_0 ),
    .i1(\inst_dob_mux_b1/B5_1 ),
    .sel(addrb_piped_piped[6]),
    .o(dob[1]));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_0  (
    .i0(inst_dob_i0_010),
    .i1(inst_dob_i0_010),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b10/B0_0 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_1  (
    .i0(inst_dob_i0_010),
    .i1(inst_dob_i0_010),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b10/B0_1 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_10  (
    .i0(inst_dob_i16_010),
    .i1(inst_dob_i16_010),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b10/B0_10 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_11  (
    .i0(inst_dob_i16_010),
    .i1(inst_dob_i16_010),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b10/B0_11 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_12  (
    .i0(inst_dob_i16_010),
    .i1(inst_dob_i16_010),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b10/B0_12 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_13  (
    .i0(inst_dob_i16_010),
    .i1(inst_dob_i16_010),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b10/B0_13 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_14  (
    .i0(inst_dob_i16_010),
    .i1(inst_dob_i16_010),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b10/B0_14 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_15  (
    .i0(inst_dob_i16_010),
    .i1(inst_dob_i16_010),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b10/B0_15 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_16  (
    .i0(inst_dob_i32_010),
    .i1(inst_dob_i32_010),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b10/B0_16 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_17  (
    .i0(inst_dob_i32_010),
    .i1(inst_dob_i32_010),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b10/B0_17 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_18  (
    .i0(inst_dob_i32_010),
    .i1(inst_dob_i32_010),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b10/B0_18 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_19  (
    .i0(inst_dob_i32_010),
    .i1(inst_dob_i32_010),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b10/B0_19 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_2  (
    .i0(inst_dob_i0_010),
    .i1(inst_dob_i0_010),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b10/B0_2 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_20  (
    .i0(inst_dob_i32_010),
    .i1(inst_dob_i32_010),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b10/B0_20 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_21  (
    .i0(inst_dob_i32_010),
    .i1(inst_dob_i32_010),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b10/B0_21 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_22  (
    .i0(inst_dob_i32_010),
    .i1(inst_dob_i32_010),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b10/B0_22 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_23  (
    .i0(inst_dob_i32_010),
    .i1(inst_dob_i32_010),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b10/B0_23 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_24  (
    .i0(inst_dob_i48_010),
    .i1(inst_dob_i48_010),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b10/B0_24 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_25  (
    .i0(inst_dob_i48_010),
    .i1(inst_dob_i48_010),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b10/B0_25 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_26  (
    .i0(inst_dob_i48_010),
    .i1(inst_dob_i48_010),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b10/B0_26 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_27  (
    .i0(inst_dob_i48_010),
    .i1(inst_dob_i48_010),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b10/B0_27 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_28  (
    .i0(inst_dob_i48_010),
    .i1(inst_dob_i48_010),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b10/B0_28 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_29  (
    .i0(inst_dob_i48_010),
    .i1(inst_dob_i48_010),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b10/B0_29 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_3  (
    .i0(inst_dob_i0_010),
    .i1(inst_dob_i0_010),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b10/B0_3 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_30  (
    .i0(inst_dob_i48_010),
    .i1(inst_dob_i48_010),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b10/B0_30 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_31  (
    .i0(inst_dob_i48_010),
    .i1(inst_dob_i48_010),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b10/B0_31 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_32  (
    .i0(inst_dob_i64_010),
    .i1(inst_dob_i64_010),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b10/B0_32 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_33  (
    .i0(inst_dob_i64_010),
    .i1(inst_dob_i64_010),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b10/B0_33 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_34  (
    .i0(inst_dob_i64_010),
    .i1(inst_dob_i64_010),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b10/B0_34 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_35  (
    .i0(inst_dob_i64_010),
    .i1(inst_dob_i64_010),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b10/B0_35 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_36  (
    .i0(inst_dob_i64_010),
    .i1(inst_dob_i64_010),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b10/B0_36 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_37  (
    .i0(inst_dob_i64_010),
    .i1(inst_dob_i64_010),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b10/B0_37 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_38  (
    .i0(inst_dob_i64_010),
    .i1(inst_dob_i64_010),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b10/B0_38 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_39  (
    .i0(inst_dob_i64_010),
    .i1(inst_dob_i64_010),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b10/B0_39 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_4  (
    .i0(inst_dob_i0_010),
    .i1(inst_dob_i0_010),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b10/B0_4 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_40  (
    .i0(inst_dob_i64_010),
    .i1(inst_dob_i64_010),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b10/B0_40 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_41  (
    .i0(inst_dob_i64_010),
    .i1(inst_dob_i64_010),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b10/B0_41 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_42  (
    .i0(inst_dob_i64_010),
    .i1(inst_dob_i64_010),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b10/B0_42 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_43  (
    .i0(inst_dob_i64_010),
    .i1(inst_dob_i64_010),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b10/B0_43 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_44  (
    .i0(inst_dob_i64_010),
    .i1(inst_dob_i64_010),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b10/B0_44 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_45  (
    .i0(inst_dob_i64_010),
    .i1(inst_dob_i64_010),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b10/B0_45 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_46  (
    .i0(inst_dob_i64_010),
    .i1(inst_dob_i64_010),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b10/B0_46 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_47  (
    .i0(inst_dob_i64_010),
    .i1(inst_dob_i64_010),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b10/B0_47 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_48  (
    .i0(inst_dob_i64_010),
    .i1(inst_dob_i64_010),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b10/B0_48 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_49  (
    .i0(inst_dob_i64_010),
    .i1(inst_dob_i64_010),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b10/B0_49 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_5  (
    .i0(inst_dob_i0_010),
    .i1(inst_dob_i0_010),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b10/B0_5 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_50  (
    .i0(inst_dob_i64_010),
    .i1(inst_dob_i64_010),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b10/B0_50 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_51  (
    .i0(inst_dob_i64_010),
    .i1(inst_dob_i64_010),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b10/B0_51 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_52  (
    .i0(inst_dob_i64_010),
    .i1(inst_dob_i64_010),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b10/B0_52 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_53  (
    .i0(inst_dob_i64_010),
    .i1(inst_dob_i64_010),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b10/B0_53 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_54  (
    .i0(inst_dob_i64_010),
    .i1(inst_dob_i64_010),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b10/B0_54 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_55  (
    .i0(inst_dob_i64_010),
    .i1(inst_dob_i64_010),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b10/B0_55 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_56  (
    .i0(inst_dob_i64_010),
    .i1(inst_dob_i64_010),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b10/B0_56 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_57  (
    .i0(inst_dob_i64_010),
    .i1(inst_dob_i64_010),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b10/B0_57 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_58  (
    .i0(inst_dob_i64_010),
    .i1(inst_dob_i64_010),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b10/B0_58 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_59  (
    .i0(inst_dob_i64_010),
    .i1(inst_dob_i64_010),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b10/B0_59 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_6  (
    .i0(inst_dob_i0_010),
    .i1(inst_dob_i0_010),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b10/B0_6 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_60  (
    .i0(inst_dob_i64_010),
    .i1(inst_dob_i64_010),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b10/B0_60 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_61  (
    .i0(inst_dob_i64_010),
    .i1(inst_dob_i64_010),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b10/B0_61 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_62  (
    .i0(inst_dob_i64_010),
    .i1(inst_dob_i64_010),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b10/B0_62 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_63  (
    .i0(inst_dob_i64_010),
    .i1(inst_dob_i64_010),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b10/B0_63 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_7  (
    .i0(inst_dob_i0_010),
    .i1(inst_dob_i0_010),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b10/B0_7 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_8  (
    .i0(inst_dob_i16_010),
    .i1(inst_dob_i16_010),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b10/B0_8 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_9  (
    .i0(inst_dob_i16_010),
    .i1(inst_dob_i16_010),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b10/B0_9 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_1_0  (
    .i0(\inst_dob_mux_b10/B0_0 ),
    .i1(\inst_dob_mux_b10/B0_1 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b10/B1_0 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_1_1  (
    .i0(\inst_dob_mux_b10/B0_2 ),
    .i1(\inst_dob_mux_b10/B0_3 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b10/B1_1 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_1_10  (
    .i0(\inst_dob_mux_b10/B0_20 ),
    .i1(\inst_dob_mux_b10/B0_21 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b10/B1_10 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_1_11  (
    .i0(\inst_dob_mux_b10/B0_22 ),
    .i1(\inst_dob_mux_b10/B0_23 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b10/B1_11 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_1_12  (
    .i0(\inst_dob_mux_b10/B0_24 ),
    .i1(\inst_dob_mux_b10/B0_25 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b10/B1_12 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_1_13  (
    .i0(\inst_dob_mux_b10/B0_26 ),
    .i1(\inst_dob_mux_b10/B0_27 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b10/B1_13 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_1_14  (
    .i0(\inst_dob_mux_b10/B0_28 ),
    .i1(\inst_dob_mux_b10/B0_29 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b10/B1_14 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_1_15  (
    .i0(\inst_dob_mux_b10/B0_30 ),
    .i1(\inst_dob_mux_b10/B0_31 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b10/B1_15 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_1_16  (
    .i0(\inst_dob_mux_b10/B0_32 ),
    .i1(\inst_dob_mux_b10/B0_33 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b10/B1_16 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_1_17  (
    .i0(\inst_dob_mux_b10/B0_34 ),
    .i1(\inst_dob_mux_b10/B0_35 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b10/B1_17 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_1_18  (
    .i0(\inst_dob_mux_b10/B0_36 ),
    .i1(\inst_dob_mux_b10/B0_37 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b10/B1_18 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_1_19  (
    .i0(\inst_dob_mux_b10/B0_38 ),
    .i1(\inst_dob_mux_b10/B0_39 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b10/B1_19 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_1_2  (
    .i0(\inst_dob_mux_b10/B0_4 ),
    .i1(\inst_dob_mux_b10/B0_5 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b10/B1_2 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_1_20  (
    .i0(\inst_dob_mux_b10/B0_40 ),
    .i1(\inst_dob_mux_b10/B0_41 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b10/B1_20 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_1_21  (
    .i0(\inst_dob_mux_b10/B0_42 ),
    .i1(\inst_dob_mux_b10/B0_43 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b10/B1_21 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_1_22  (
    .i0(\inst_dob_mux_b10/B0_44 ),
    .i1(\inst_dob_mux_b10/B0_45 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b10/B1_22 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_1_23  (
    .i0(\inst_dob_mux_b10/B0_46 ),
    .i1(\inst_dob_mux_b10/B0_47 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b10/B1_23 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_1_24  (
    .i0(\inst_dob_mux_b10/B0_48 ),
    .i1(\inst_dob_mux_b10/B0_49 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b10/B1_24 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_1_25  (
    .i0(\inst_dob_mux_b10/B0_50 ),
    .i1(\inst_dob_mux_b10/B0_51 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b10/B1_25 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_1_26  (
    .i0(\inst_dob_mux_b10/B0_52 ),
    .i1(\inst_dob_mux_b10/B0_53 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b10/B1_26 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_1_27  (
    .i0(\inst_dob_mux_b10/B0_54 ),
    .i1(\inst_dob_mux_b10/B0_55 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b10/B1_27 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_1_28  (
    .i0(\inst_dob_mux_b10/B0_56 ),
    .i1(\inst_dob_mux_b10/B0_57 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b10/B1_28 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_1_29  (
    .i0(\inst_dob_mux_b10/B0_58 ),
    .i1(\inst_dob_mux_b10/B0_59 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b10/B1_29 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_1_3  (
    .i0(\inst_dob_mux_b10/B0_6 ),
    .i1(\inst_dob_mux_b10/B0_7 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b10/B1_3 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_1_30  (
    .i0(\inst_dob_mux_b10/B0_60 ),
    .i1(\inst_dob_mux_b10/B0_61 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b10/B1_30 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_1_31  (
    .i0(\inst_dob_mux_b10/B0_62 ),
    .i1(\inst_dob_mux_b10/B0_63 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b10/B1_31 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_1_4  (
    .i0(\inst_dob_mux_b10/B0_8 ),
    .i1(\inst_dob_mux_b10/B0_9 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b10/B1_4 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_1_5  (
    .i0(\inst_dob_mux_b10/B0_10 ),
    .i1(\inst_dob_mux_b10/B0_11 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b10/B1_5 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_1_6  (
    .i0(\inst_dob_mux_b10/B0_12 ),
    .i1(\inst_dob_mux_b10/B0_13 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b10/B1_6 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_1_7  (
    .i0(\inst_dob_mux_b10/B0_14 ),
    .i1(\inst_dob_mux_b10/B0_15 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b10/B1_7 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_1_8  (
    .i0(\inst_dob_mux_b10/B0_16 ),
    .i1(\inst_dob_mux_b10/B0_17 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b10/B1_8 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_1_9  (
    .i0(\inst_dob_mux_b10/B0_18 ),
    .i1(\inst_dob_mux_b10/B0_19 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b10/B1_9 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_2_0  (
    .i0(\inst_dob_mux_b10/B1_0 ),
    .i1(\inst_dob_mux_b10/B1_1 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b10/B2_0 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_2_1  (
    .i0(\inst_dob_mux_b10/B1_2 ),
    .i1(\inst_dob_mux_b10/B1_3 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b10/B2_1 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_2_10  (
    .i0(\inst_dob_mux_b10/B1_20 ),
    .i1(\inst_dob_mux_b10/B1_21 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b10/B2_10 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_2_11  (
    .i0(\inst_dob_mux_b10/B1_22 ),
    .i1(\inst_dob_mux_b10/B1_23 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b10/B2_11 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_2_12  (
    .i0(\inst_dob_mux_b10/B1_24 ),
    .i1(\inst_dob_mux_b10/B1_25 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b10/B2_12 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_2_13  (
    .i0(\inst_dob_mux_b10/B1_26 ),
    .i1(\inst_dob_mux_b10/B1_27 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b10/B2_13 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_2_14  (
    .i0(\inst_dob_mux_b10/B1_28 ),
    .i1(\inst_dob_mux_b10/B1_29 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b10/B2_14 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_2_15  (
    .i0(\inst_dob_mux_b10/B1_30 ),
    .i1(\inst_dob_mux_b10/B1_31 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b10/B2_15 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_2_2  (
    .i0(\inst_dob_mux_b10/B1_4 ),
    .i1(\inst_dob_mux_b10/B1_5 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b10/B2_2 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_2_3  (
    .i0(\inst_dob_mux_b10/B1_6 ),
    .i1(\inst_dob_mux_b10/B1_7 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b10/B2_3 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_2_4  (
    .i0(\inst_dob_mux_b10/B1_8 ),
    .i1(\inst_dob_mux_b10/B1_9 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b10/B2_4 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_2_5  (
    .i0(\inst_dob_mux_b10/B1_10 ),
    .i1(\inst_dob_mux_b10/B1_11 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b10/B2_5 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_2_6  (
    .i0(\inst_dob_mux_b10/B1_12 ),
    .i1(\inst_dob_mux_b10/B1_13 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b10/B2_6 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_2_7  (
    .i0(\inst_dob_mux_b10/B1_14 ),
    .i1(\inst_dob_mux_b10/B1_15 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b10/B2_7 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_2_8  (
    .i0(\inst_dob_mux_b10/B1_16 ),
    .i1(\inst_dob_mux_b10/B1_17 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b10/B2_8 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_2_9  (
    .i0(\inst_dob_mux_b10/B1_18 ),
    .i1(\inst_dob_mux_b10/B1_19 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b10/B2_9 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_3_0  (
    .i0(\inst_dob_mux_b10/B2_0 ),
    .i1(\inst_dob_mux_b10/B2_1 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b10/B3_0 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_3_1  (
    .i0(\inst_dob_mux_b10/B2_2 ),
    .i1(\inst_dob_mux_b10/B2_3 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b10/B3_1 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_3_2  (
    .i0(\inst_dob_mux_b10/B2_4 ),
    .i1(\inst_dob_mux_b10/B2_5 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b10/B3_2 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_3_3  (
    .i0(\inst_dob_mux_b10/B2_6 ),
    .i1(\inst_dob_mux_b10/B2_7 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b10/B3_3 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_3_4  (
    .i0(\inst_dob_mux_b10/B2_8 ),
    .i1(\inst_dob_mux_b10/B2_9 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b10/B3_4 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_3_5  (
    .i0(\inst_dob_mux_b10/B2_10 ),
    .i1(\inst_dob_mux_b10/B2_11 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b10/B3_5 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_3_6  (
    .i0(\inst_dob_mux_b10/B2_12 ),
    .i1(\inst_dob_mux_b10/B2_13 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b10/B3_6 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_3_7  (
    .i0(\inst_dob_mux_b10/B2_14 ),
    .i1(\inst_dob_mux_b10/B2_15 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b10/B3_7 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_4_0  (
    .i0(\inst_dob_mux_b10/B3_0 ),
    .i1(\inst_dob_mux_b10/B3_1 ),
    .sel(addrb_piped_piped[4]),
    .o(\inst_dob_mux_b10/B4_0 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_4_1  (
    .i0(\inst_dob_mux_b10/B3_2 ),
    .i1(\inst_dob_mux_b10/B3_3 ),
    .sel(addrb_piped_piped[4]),
    .o(\inst_dob_mux_b10/B4_1 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_4_2  (
    .i0(\inst_dob_mux_b10/B3_4 ),
    .i1(\inst_dob_mux_b10/B3_5 ),
    .sel(addrb_piped_piped[4]),
    .o(\inst_dob_mux_b10/B4_2 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_4_3  (
    .i0(\inst_dob_mux_b10/B3_6 ),
    .i1(\inst_dob_mux_b10/B3_7 ),
    .sel(addrb_piped_piped[4]),
    .o(\inst_dob_mux_b10/B4_3 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_5_0  (
    .i0(\inst_dob_mux_b10/B4_0 ),
    .i1(\inst_dob_mux_b10/B4_1 ),
    .sel(addrb_piped_piped[5]),
    .o(\inst_dob_mux_b10/B5_0 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_5_1  (
    .i0(\inst_dob_mux_b10/B4_2 ),
    .i1(\inst_dob_mux_b10/B4_3 ),
    .sel(addrb_piped_piped[5]),
    .o(\inst_dob_mux_b10/B5_1 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_6_0  (
    .i0(\inst_dob_mux_b10/B5_0 ),
    .i1(\inst_dob_mux_b10/B5_1 ),
    .sel(addrb_piped_piped[6]),
    .o(dob[10]));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_0  (
    .i0(inst_dob_i0_011),
    .i1(inst_dob_i0_011),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b11/B0_0 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_1  (
    .i0(inst_dob_i0_011),
    .i1(inst_dob_i0_011),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b11/B0_1 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_10  (
    .i0(inst_dob_i16_011),
    .i1(inst_dob_i16_011),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b11/B0_10 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_11  (
    .i0(inst_dob_i16_011),
    .i1(inst_dob_i16_011),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b11/B0_11 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_12  (
    .i0(inst_dob_i16_011),
    .i1(inst_dob_i16_011),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b11/B0_12 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_13  (
    .i0(inst_dob_i16_011),
    .i1(inst_dob_i16_011),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b11/B0_13 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_14  (
    .i0(inst_dob_i16_011),
    .i1(inst_dob_i16_011),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b11/B0_14 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_15  (
    .i0(inst_dob_i16_011),
    .i1(inst_dob_i16_011),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b11/B0_15 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_16  (
    .i0(inst_dob_i32_011),
    .i1(inst_dob_i32_011),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b11/B0_16 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_17  (
    .i0(inst_dob_i32_011),
    .i1(inst_dob_i32_011),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b11/B0_17 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_18  (
    .i0(inst_dob_i32_011),
    .i1(inst_dob_i32_011),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b11/B0_18 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_19  (
    .i0(inst_dob_i32_011),
    .i1(inst_dob_i32_011),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b11/B0_19 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_2  (
    .i0(inst_dob_i0_011),
    .i1(inst_dob_i0_011),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b11/B0_2 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_20  (
    .i0(inst_dob_i32_011),
    .i1(inst_dob_i32_011),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b11/B0_20 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_21  (
    .i0(inst_dob_i32_011),
    .i1(inst_dob_i32_011),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b11/B0_21 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_22  (
    .i0(inst_dob_i32_011),
    .i1(inst_dob_i32_011),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b11/B0_22 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_23  (
    .i0(inst_dob_i32_011),
    .i1(inst_dob_i32_011),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b11/B0_23 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_24  (
    .i0(inst_dob_i48_011),
    .i1(inst_dob_i48_011),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b11/B0_24 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_25  (
    .i0(inst_dob_i48_011),
    .i1(inst_dob_i48_011),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b11/B0_25 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_26  (
    .i0(inst_dob_i48_011),
    .i1(inst_dob_i48_011),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b11/B0_26 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_27  (
    .i0(inst_dob_i48_011),
    .i1(inst_dob_i48_011),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b11/B0_27 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_28  (
    .i0(inst_dob_i48_011),
    .i1(inst_dob_i48_011),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b11/B0_28 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_29  (
    .i0(inst_dob_i48_011),
    .i1(inst_dob_i48_011),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b11/B0_29 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_3  (
    .i0(inst_dob_i0_011),
    .i1(inst_dob_i0_011),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b11/B0_3 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_30  (
    .i0(inst_dob_i48_011),
    .i1(inst_dob_i48_011),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b11/B0_30 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_31  (
    .i0(inst_dob_i48_011),
    .i1(inst_dob_i48_011),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b11/B0_31 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_32  (
    .i0(inst_dob_i64_011),
    .i1(inst_dob_i64_011),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b11/B0_32 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_33  (
    .i0(inst_dob_i64_011),
    .i1(inst_dob_i64_011),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b11/B0_33 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_34  (
    .i0(inst_dob_i64_011),
    .i1(inst_dob_i64_011),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b11/B0_34 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_35  (
    .i0(inst_dob_i64_011),
    .i1(inst_dob_i64_011),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b11/B0_35 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_36  (
    .i0(inst_dob_i64_011),
    .i1(inst_dob_i64_011),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b11/B0_36 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_37  (
    .i0(inst_dob_i64_011),
    .i1(inst_dob_i64_011),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b11/B0_37 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_38  (
    .i0(inst_dob_i64_011),
    .i1(inst_dob_i64_011),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b11/B0_38 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_39  (
    .i0(inst_dob_i64_011),
    .i1(inst_dob_i64_011),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b11/B0_39 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_4  (
    .i0(inst_dob_i0_011),
    .i1(inst_dob_i0_011),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b11/B0_4 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_40  (
    .i0(inst_dob_i64_011),
    .i1(inst_dob_i64_011),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b11/B0_40 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_41  (
    .i0(inst_dob_i64_011),
    .i1(inst_dob_i64_011),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b11/B0_41 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_42  (
    .i0(inst_dob_i64_011),
    .i1(inst_dob_i64_011),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b11/B0_42 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_43  (
    .i0(inst_dob_i64_011),
    .i1(inst_dob_i64_011),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b11/B0_43 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_44  (
    .i0(inst_dob_i64_011),
    .i1(inst_dob_i64_011),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b11/B0_44 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_45  (
    .i0(inst_dob_i64_011),
    .i1(inst_dob_i64_011),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b11/B0_45 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_46  (
    .i0(inst_dob_i64_011),
    .i1(inst_dob_i64_011),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b11/B0_46 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_47  (
    .i0(inst_dob_i64_011),
    .i1(inst_dob_i64_011),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b11/B0_47 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_48  (
    .i0(inst_dob_i64_011),
    .i1(inst_dob_i64_011),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b11/B0_48 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_49  (
    .i0(inst_dob_i64_011),
    .i1(inst_dob_i64_011),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b11/B0_49 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_5  (
    .i0(inst_dob_i0_011),
    .i1(inst_dob_i0_011),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b11/B0_5 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_50  (
    .i0(inst_dob_i64_011),
    .i1(inst_dob_i64_011),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b11/B0_50 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_51  (
    .i0(inst_dob_i64_011),
    .i1(inst_dob_i64_011),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b11/B0_51 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_52  (
    .i0(inst_dob_i64_011),
    .i1(inst_dob_i64_011),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b11/B0_52 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_53  (
    .i0(inst_dob_i64_011),
    .i1(inst_dob_i64_011),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b11/B0_53 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_54  (
    .i0(inst_dob_i64_011),
    .i1(inst_dob_i64_011),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b11/B0_54 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_55  (
    .i0(inst_dob_i64_011),
    .i1(inst_dob_i64_011),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b11/B0_55 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_56  (
    .i0(inst_dob_i64_011),
    .i1(inst_dob_i64_011),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b11/B0_56 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_57  (
    .i0(inst_dob_i64_011),
    .i1(inst_dob_i64_011),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b11/B0_57 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_58  (
    .i0(inst_dob_i64_011),
    .i1(inst_dob_i64_011),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b11/B0_58 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_59  (
    .i0(inst_dob_i64_011),
    .i1(inst_dob_i64_011),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b11/B0_59 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_6  (
    .i0(inst_dob_i0_011),
    .i1(inst_dob_i0_011),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b11/B0_6 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_60  (
    .i0(inst_dob_i64_011),
    .i1(inst_dob_i64_011),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b11/B0_60 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_61  (
    .i0(inst_dob_i64_011),
    .i1(inst_dob_i64_011),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b11/B0_61 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_62  (
    .i0(inst_dob_i64_011),
    .i1(inst_dob_i64_011),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b11/B0_62 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_63  (
    .i0(inst_dob_i64_011),
    .i1(inst_dob_i64_011),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b11/B0_63 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_7  (
    .i0(inst_dob_i0_011),
    .i1(inst_dob_i0_011),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b11/B0_7 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_8  (
    .i0(inst_dob_i16_011),
    .i1(inst_dob_i16_011),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b11/B0_8 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_9  (
    .i0(inst_dob_i16_011),
    .i1(inst_dob_i16_011),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b11/B0_9 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_1_0  (
    .i0(\inst_dob_mux_b11/B0_0 ),
    .i1(\inst_dob_mux_b11/B0_1 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b11/B1_0 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_1_1  (
    .i0(\inst_dob_mux_b11/B0_2 ),
    .i1(\inst_dob_mux_b11/B0_3 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b11/B1_1 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_1_10  (
    .i0(\inst_dob_mux_b11/B0_20 ),
    .i1(\inst_dob_mux_b11/B0_21 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b11/B1_10 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_1_11  (
    .i0(\inst_dob_mux_b11/B0_22 ),
    .i1(\inst_dob_mux_b11/B0_23 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b11/B1_11 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_1_12  (
    .i0(\inst_dob_mux_b11/B0_24 ),
    .i1(\inst_dob_mux_b11/B0_25 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b11/B1_12 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_1_13  (
    .i0(\inst_dob_mux_b11/B0_26 ),
    .i1(\inst_dob_mux_b11/B0_27 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b11/B1_13 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_1_14  (
    .i0(\inst_dob_mux_b11/B0_28 ),
    .i1(\inst_dob_mux_b11/B0_29 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b11/B1_14 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_1_15  (
    .i0(\inst_dob_mux_b11/B0_30 ),
    .i1(\inst_dob_mux_b11/B0_31 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b11/B1_15 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_1_16  (
    .i0(\inst_dob_mux_b11/B0_32 ),
    .i1(\inst_dob_mux_b11/B0_33 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b11/B1_16 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_1_17  (
    .i0(\inst_dob_mux_b11/B0_34 ),
    .i1(\inst_dob_mux_b11/B0_35 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b11/B1_17 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_1_18  (
    .i0(\inst_dob_mux_b11/B0_36 ),
    .i1(\inst_dob_mux_b11/B0_37 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b11/B1_18 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_1_19  (
    .i0(\inst_dob_mux_b11/B0_38 ),
    .i1(\inst_dob_mux_b11/B0_39 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b11/B1_19 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_1_2  (
    .i0(\inst_dob_mux_b11/B0_4 ),
    .i1(\inst_dob_mux_b11/B0_5 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b11/B1_2 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_1_20  (
    .i0(\inst_dob_mux_b11/B0_40 ),
    .i1(\inst_dob_mux_b11/B0_41 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b11/B1_20 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_1_21  (
    .i0(\inst_dob_mux_b11/B0_42 ),
    .i1(\inst_dob_mux_b11/B0_43 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b11/B1_21 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_1_22  (
    .i0(\inst_dob_mux_b11/B0_44 ),
    .i1(\inst_dob_mux_b11/B0_45 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b11/B1_22 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_1_23  (
    .i0(\inst_dob_mux_b11/B0_46 ),
    .i1(\inst_dob_mux_b11/B0_47 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b11/B1_23 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_1_24  (
    .i0(\inst_dob_mux_b11/B0_48 ),
    .i1(\inst_dob_mux_b11/B0_49 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b11/B1_24 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_1_25  (
    .i0(\inst_dob_mux_b11/B0_50 ),
    .i1(\inst_dob_mux_b11/B0_51 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b11/B1_25 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_1_26  (
    .i0(\inst_dob_mux_b11/B0_52 ),
    .i1(\inst_dob_mux_b11/B0_53 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b11/B1_26 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_1_27  (
    .i0(\inst_dob_mux_b11/B0_54 ),
    .i1(\inst_dob_mux_b11/B0_55 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b11/B1_27 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_1_28  (
    .i0(\inst_dob_mux_b11/B0_56 ),
    .i1(\inst_dob_mux_b11/B0_57 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b11/B1_28 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_1_29  (
    .i0(\inst_dob_mux_b11/B0_58 ),
    .i1(\inst_dob_mux_b11/B0_59 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b11/B1_29 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_1_3  (
    .i0(\inst_dob_mux_b11/B0_6 ),
    .i1(\inst_dob_mux_b11/B0_7 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b11/B1_3 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_1_30  (
    .i0(\inst_dob_mux_b11/B0_60 ),
    .i1(\inst_dob_mux_b11/B0_61 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b11/B1_30 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_1_31  (
    .i0(\inst_dob_mux_b11/B0_62 ),
    .i1(\inst_dob_mux_b11/B0_63 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b11/B1_31 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_1_4  (
    .i0(\inst_dob_mux_b11/B0_8 ),
    .i1(\inst_dob_mux_b11/B0_9 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b11/B1_4 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_1_5  (
    .i0(\inst_dob_mux_b11/B0_10 ),
    .i1(\inst_dob_mux_b11/B0_11 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b11/B1_5 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_1_6  (
    .i0(\inst_dob_mux_b11/B0_12 ),
    .i1(\inst_dob_mux_b11/B0_13 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b11/B1_6 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_1_7  (
    .i0(\inst_dob_mux_b11/B0_14 ),
    .i1(\inst_dob_mux_b11/B0_15 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b11/B1_7 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_1_8  (
    .i0(\inst_dob_mux_b11/B0_16 ),
    .i1(\inst_dob_mux_b11/B0_17 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b11/B1_8 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_1_9  (
    .i0(\inst_dob_mux_b11/B0_18 ),
    .i1(\inst_dob_mux_b11/B0_19 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b11/B1_9 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_2_0  (
    .i0(\inst_dob_mux_b11/B1_0 ),
    .i1(\inst_dob_mux_b11/B1_1 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b11/B2_0 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_2_1  (
    .i0(\inst_dob_mux_b11/B1_2 ),
    .i1(\inst_dob_mux_b11/B1_3 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b11/B2_1 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_2_10  (
    .i0(\inst_dob_mux_b11/B1_20 ),
    .i1(\inst_dob_mux_b11/B1_21 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b11/B2_10 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_2_11  (
    .i0(\inst_dob_mux_b11/B1_22 ),
    .i1(\inst_dob_mux_b11/B1_23 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b11/B2_11 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_2_12  (
    .i0(\inst_dob_mux_b11/B1_24 ),
    .i1(\inst_dob_mux_b11/B1_25 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b11/B2_12 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_2_13  (
    .i0(\inst_dob_mux_b11/B1_26 ),
    .i1(\inst_dob_mux_b11/B1_27 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b11/B2_13 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_2_14  (
    .i0(\inst_dob_mux_b11/B1_28 ),
    .i1(\inst_dob_mux_b11/B1_29 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b11/B2_14 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_2_15  (
    .i0(\inst_dob_mux_b11/B1_30 ),
    .i1(\inst_dob_mux_b11/B1_31 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b11/B2_15 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_2_2  (
    .i0(\inst_dob_mux_b11/B1_4 ),
    .i1(\inst_dob_mux_b11/B1_5 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b11/B2_2 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_2_3  (
    .i0(\inst_dob_mux_b11/B1_6 ),
    .i1(\inst_dob_mux_b11/B1_7 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b11/B2_3 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_2_4  (
    .i0(\inst_dob_mux_b11/B1_8 ),
    .i1(\inst_dob_mux_b11/B1_9 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b11/B2_4 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_2_5  (
    .i0(\inst_dob_mux_b11/B1_10 ),
    .i1(\inst_dob_mux_b11/B1_11 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b11/B2_5 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_2_6  (
    .i0(\inst_dob_mux_b11/B1_12 ),
    .i1(\inst_dob_mux_b11/B1_13 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b11/B2_6 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_2_7  (
    .i0(\inst_dob_mux_b11/B1_14 ),
    .i1(\inst_dob_mux_b11/B1_15 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b11/B2_7 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_2_8  (
    .i0(\inst_dob_mux_b11/B1_16 ),
    .i1(\inst_dob_mux_b11/B1_17 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b11/B2_8 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_2_9  (
    .i0(\inst_dob_mux_b11/B1_18 ),
    .i1(\inst_dob_mux_b11/B1_19 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b11/B2_9 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_3_0  (
    .i0(\inst_dob_mux_b11/B2_0 ),
    .i1(\inst_dob_mux_b11/B2_1 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b11/B3_0 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_3_1  (
    .i0(\inst_dob_mux_b11/B2_2 ),
    .i1(\inst_dob_mux_b11/B2_3 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b11/B3_1 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_3_2  (
    .i0(\inst_dob_mux_b11/B2_4 ),
    .i1(\inst_dob_mux_b11/B2_5 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b11/B3_2 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_3_3  (
    .i0(\inst_dob_mux_b11/B2_6 ),
    .i1(\inst_dob_mux_b11/B2_7 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b11/B3_3 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_3_4  (
    .i0(\inst_dob_mux_b11/B2_8 ),
    .i1(\inst_dob_mux_b11/B2_9 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b11/B3_4 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_3_5  (
    .i0(\inst_dob_mux_b11/B2_10 ),
    .i1(\inst_dob_mux_b11/B2_11 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b11/B3_5 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_3_6  (
    .i0(\inst_dob_mux_b11/B2_12 ),
    .i1(\inst_dob_mux_b11/B2_13 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b11/B3_6 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_3_7  (
    .i0(\inst_dob_mux_b11/B2_14 ),
    .i1(\inst_dob_mux_b11/B2_15 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b11/B3_7 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_4_0  (
    .i0(\inst_dob_mux_b11/B3_0 ),
    .i1(\inst_dob_mux_b11/B3_1 ),
    .sel(addrb_piped_piped[4]),
    .o(\inst_dob_mux_b11/B4_0 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_4_1  (
    .i0(\inst_dob_mux_b11/B3_2 ),
    .i1(\inst_dob_mux_b11/B3_3 ),
    .sel(addrb_piped_piped[4]),
    .o(\inst_dob_mux_b11/B4_1 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_4_2  (
    .i0(\inst_dob_mux_b11/B3_4 ),
    .i1(\inst_dob_mux_b11/B3_5 ),
    .sel(addrb_piped_piped[4]),
    .o(\inst_dob_mux_b11/B4_2 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_4_3  (
    .i0(\inst_dob_mux_b11/B3_6 ),
    .i1(\inst_dob_mux_b11/B3_7 ),
    .sel(addrb_piped_piped[4]),
    .o(\inst_dob_mux_b11/B4_3 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_5_0  (
    .i0(\inst_dob_mux_b11/B4_0 ),
    .i1(\inst_dob_mux_b11/B4_1 ),
    .sel(addrb_piped_piped[5]),
    .o(\inst_dob_mux_b11/B5_0 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_5_1  (
    .i0(\inst_dob_mux_b11/B4_2 ),
    .i1(\inst_dob_mux_b11/B4_3 ),
    .sel(addrb_piped_piped[5]),
    .o(\inst_dob_mux_b11/B5_1 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_6_0  (
    .i0(\inst_dob_mux_b11/B5_0 ),
    .i1(\inst_dob_mux_b11/B5_1 ),
    .sel(addrb_piped_piped[6]),
    .o(dob[11]));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_0  (
    .i0(inst_dob_i0_012),
    .i1(inst_dob_i0_012),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b12/B0_0 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_1  (
    .i0(inst_dob_i0_012),
    .i1(inst_dob_i0_012),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b12/B0_1 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_10  (
    .i0(inst_dob_i16_012),
    .i1(inst_dob_i16_012),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b12/B0_10 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_11  (
    .i0(inst_dob_i16_012),
    .i1(inst_dob_i16_012),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b12/B0_11 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_12  (
    .i0(inst_dob_i16_012),
    .i1(inst_dob_i16_012),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b12/B0_12 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_13  (
    .i0(inst_dob_i16_012),
    .i1(inst_dob_i16_012),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b12/B0_13 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_14  (
    .i0(inst_dob_i16_012),
    .i1(inst_dob_i16_012),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b12/B0_14 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_15  (
    .i0(inst_dob_i16_012),
    .i1(inst_dob_i16_012),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b12/B0_15 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_16  (
    .i0(inst_dob_i32_012),
    .i1(inst_dob_i32_012),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b12/B0_16 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_17  (
    .i0(inst_dob_i32_012),
    .i1(inst_dob_i32_012),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b12/B0_17 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_18  (
    .i0(inst_dob_i32_012),
    .i1(inst_dob_i32_012),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b12/B0_18 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_19  (
    .i0(inst_dob_i32_012),
    .i1(inst_dob_i32_012),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b12/B0_19 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_2  (
    .i0(inst_dob_i0_012),
    .i1(inst_dob_i0_012),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b12/B0_2 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_20  (
    .i0(inst_dob_i32_012),
    .i1(inst_dob_i32_012),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b12/B0_20 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_21  (
    .i0(inst_dob_i32_012),
    .i1(inst_dob_i32_012),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b12/B0_21 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_22  (
    .i0(inst_dob_i32_012),
    .i1(inst_dob_i32_012),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b12/B0_22 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_23  (
    .i0(inst_dob_i32_012),
    .i1(inst_dob_i32_012),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b12/B0_23 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_24  (
    .i0(inst_dob_i48_012),
    .i1(inst_dob_i48_012),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b12/B0_24 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_25  (
    .i0(inst_dob_i48_012),
    .i1(inst_dob_i48_012),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b12/B0_25 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_26  (
    .i0(inst_dob_i48_012),
    .i1(inst_dob_i48_012),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b12/B0_26 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_27  (
    .i0(inst_dob_i48_012),
    .i1(inst_dob_i48_012),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b12/B0_27 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_28  (
    .i0(inst_dob_i48_012),
    .i1(inst_dob_i48_012),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b12/B0_28 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_29  (
    .i0(inst_dob_i48_012),
    .i1(inst_dob_i48_012),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b12/B0_29 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_3  (
    .i0(inst_dob_i0_012),
    .i1(inst_dob_i0_012),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b12/B0_3 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_30  (
    .i0(inst_dob_i48_012),
    .i1(inst_dob_i48_012),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b12/B0_30 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_31  (
    .i0(inst_dob_i48_012),
    .i1(inst_dob_i48_012),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b12/B0_31 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_32  (
    .i0(inst_dob_i64_012),
    .i1(inst_dob_i64_012),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b12/B0_32 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_33  (
    .i0(inst_dob_i64_012),
    .i1(inst_dob_i64_012),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b12/B0_33 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_34  (
    .i0(inst_dob_i64_012),
    .i1(inst_dob_i64_012),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b12/B0_34 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_35  (
    .i0(inst_dob_i64_012),
    .i1(inst_dob_i64_012),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b12/B0_35 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_36  (
    .i0(inst_dob_i64_012),
    .i1(inst_dob_i64_012),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b12/B0_36 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_37  (
    .i0(inst_dob_i64_012),
    .i1(inst_dob_i64_012),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b12/B0_37 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_38  (
    .i0(inst_dob_i64_012),
    .i1(inst_dob_i64_012),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b12/B0_38 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_39  (
    .i0(inst_dob_i64_012),
    .i1(inst_dob_i64_012),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b12/B0_39 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_4  (
    .i0(inst_dob_i0_012),
    .i1(inst_dob_i0_012),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b12/B0_4 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_40  (
    .i0(inst_dob_i64_012),
    .i1(inst_dob_i64_012),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b12/B0_40 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_41  (
    .i0(inst_dob_i64_012),
    .i1(inst_dob_i64_012),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b12/B0_41 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_42  (
    .i0(inst_dob_i64_012),
    .i1(inst_dob_i64_012),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b12/B0_42 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_43  (
    .i0(inst_dob_i64_012),
    .i1(inst_dob_i64_012),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b12/B0_43 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_44  (
    .i0(inst_dob_i64_012),
    .i1(inst_dob_i64_012),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b12/B0_44 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_45  (
    .i0(inst_dob_i64_012),
    .i1(inst_dob_i64_012),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b12/B0_45 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_46  (
    .i0(inst_dob_i64_012),
    .i1(inst_dob_i64_012),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b12/B0_46 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_47  (
    .i0(inst_dob_i64_012),
    .i1(inst_dob_i64_012),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b12/B0_47 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_48  (
    .i0(inst_dob_i64_012),
    .i1(inst_dob_i64_012),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b12/B0_48 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_49  (
    .i0(inst_dob_i64_012),
    .i1(inst_dob_i64_012),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b12/B0_49 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_5  (
    .i0(inst_dob_i0_012),
    .i1(inst_dob_i0_012),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b12/B0_5 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_50  (
    .i0(inst_dob_i64_012),
    .i1(inst_dob_i64_012),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b12/B0_50 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_51  (
    .i0(inst_dob_i64_012),
    .i1(inst_dob_i64_012),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b12/B0_51 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_52  (
    .i0(inst_dob_i64_012),
    .i1(inst_dob_i64_012),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b12/B0_52 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_53  (
    .i0(inst_dob_i64_012),
    .i1(inst_dob_i64_012),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b12/B0_53 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_54  (
    .i0(inst_dob_i64_012),
    .i1(inst_dob_i64_012),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b12/B0_54 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_55  (
    .i0(inst_dob_i64_012),
    .i1(inst_dob_i64_012),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b12/B0_55 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_56  (
    .i0(inst_dob_i64_012),
    .i1(inst_dob_i64_012),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b12/B0_56 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_57  (
    .i0(inst_dob_i64_012),
    .i1(inst_dob_i64_012),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b12/B0_57 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_58  (
    .i0(inst_dob_i64_012),
    .i1(inst_dob_i64_012),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b12/B0_58 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_59  (
    .i0(inst_dob_i64_012),
    .i1(inst_dob_i64_012),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b12/B0_59 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_6  (
    .i0(inst_dob_i0_012),
    .i1(inst_dob_i0_012),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b12/B0_6 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_60  (
    .i0(inst_dob_i64_012),
    .i1(inst_dob_i64_012),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b12/B0_60 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_61  (
    .i0(inst_dob_i64_012),
    .i1(inst_dob_i64_012),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b12/B0_61 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_62  (
    .i0(inst_dob_i64_012),
    .i1(inst_dob_i64_012),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b12/B0_62 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_63  (
    .i0(inst_dob_i64_012),
    .i1(inst_dob_i64_012),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b12/B0_63 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_7  (
    .i0(inst_dob_i0_012),
    .i1(inst_dob_i0_012),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b12/B0_7 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_8  (
    .i0(inst_dob_i16_012),
    .i1(inst_dob_i16_012),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b12/B0_8 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_9  (
    .i0(inst_dob_i16_012),
    .i1(inst_dob_i16_012),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b12/B0_9 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_1_0  (
    .i0(\inst_dob_mux_b12/B0_0 ),
    .i1(\inst_dob_mux_b12/B0_1 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b12/B1_0 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_1_1  (
    .i0(\inst_dob_mux_b12/B0_2 ),
    .i1(\inst_dob_mux_b12/B0_3 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b12/B1_1 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_1_10  (
    .i0(\inst_dob_mux_b12/B0_20 ),
    .i1(\inst_dob_mux_b12/B0_21 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b12/B1_10 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_1_11  (
    .i0(\inst_dob_mux_b12/B0_22 ),
    .i1(\inst_dob_mux_b12/B0_23 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b12/B1_11 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_1_12  (
    .i0(\inst_dob_mux_b12/B0_24 ),
    .i1(\inst_dob_mux_b12/B0_25 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b12/B1_12 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_1_13  (
    .i0(\inst_dob_mux_b12/B0_26 ),
    .i1(\inst_dob_mux_b12/B0_27 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b12/B1_13 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_1_14  (
    .i0(\inst_dob_mux_b12/B0_28 ),
    .i1(\inst_dob_mux_b12/B0_29 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b12/B1_14 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_1_15  (
    .i0(\inst_dob_mux_b12/B0_30 ),
    .i1(\inst_dob_mux_b12/B0_31 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b12/B1_15 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_1_16  (
    .i0(\inst_dob_mux_b12/B0_32 ),
    .i1(\inst_dob_mux_b12/B0_33 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b12/B1_16 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_1_17  (
    .i0(\inst_dob_mux_b12/B0_34 ),
    .i1(\inst_dob_mux_b12/B0_35 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b12/B1_17 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_1_18  (
    .i0(\inst_dob_mux_b12/B0_36 ),
    .i1(\inst_dob_mux_b12/B0_37 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b12/B1_18 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_1_19  (
    .i0(\inst_dob_mux_b12/B0_38 ),
    .i1(\inst_dob_mux_b12/B0_39 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b12/B1_19 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_1_2  (
    .i0(\inst_dob_mux_b12/B0_4 ),
    .i1(\inst_dob_mux_b12/B0_5 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b12/B1_2 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_1_20  (
    .i0(\inst_dob_mux_b12/B0_40 ),
    .i1(\inst_dob_mux_b12/B0_41 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b12/B1_20 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_1_21  (
    .i0(\inst_dob_mux_b12/B0_42 ),
    .i1(\inst_dob_mux_b12/B0_43 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b12/B1_21 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_1_22  (
    .i0(\inst_dob_mux_b12/B0_44 ),
    .i1(\inst_dob_mux_b12/B0_45 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b12/B1_22 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_1_23  (
    .i0(\inst_dob_mux_b12/B0_46 ),
    .i1(\inst_dob_mux_b12/B0_47 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b12/B1_23 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_1_24  (
    .i0(\inst_dob_mux_b12/B0_48 ),
    .i1(\inst_dob_mux_b12/B0_49 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b12/B1_24 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_1_25  (
    .i0(\inst_dob_mux_b12/B0_50 ),
    .i1(\inst_dob_mux_b12/B0_51 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b12/B1_25 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_1_26  (
    .i0(\inst_dob_mux_b12/B0_52 ),
    .i1(\inst_dob_mux_b12/B0_53 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b12/B1_26 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_1_27  (
    .i0(\inst_dob_mux_b12/B0_54 ),
    .i1(\inst_dob_mux_b12/B0_55 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b12/B1_27 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_1_28  (
    .i0(\inst_dob_mux_b12/B0_56 ),
    .i1(\inst_dob_mux_b12/B0_57 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b12/B1_28 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_1_29  (
    .i0(\inst_dob_mux_b12/B0_58 ),
    .i1(\inst_dob_mux_b12/B0_59 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b12/B1_29 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_1_3  (
    .i0(\inst_dob_mux_b12/B0_6 ),
    .i1(\inst_dob_mux_b12/B0_7 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b12/B1_3 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_1_30  (
    .i0(\inst_dob_mux_b12/B0_60 ),
    .i1(\inst_dob_mux_b12/B0_61 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b12/B1_30 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_1_31  (
    .i0(\inst_dob_mux_b12/B0_62 ),
    .i1(\inst_dob_mux_b12/B0_63 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b12/B1_31 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_1_4  (
    .i0(\inst_dob_mux_b12/B0_8 ),
    .i1(\inst_dob_mux_b12/B0_9 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b12/B1_4 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_1_5  (
    .i0(\inst_dob_mux_b12/B0_10 ),
    .i1(\inst_dob_mux_b12/B0_11 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b12/B1_5 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_1_6  (
    .i0(\inst_dob_mux_b12/B0_12 ),
    .i1(\inst_dob_mux_b12/B0_13 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b12/B1_6 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_1_7  (
    .i0(\inst_dob_mux_b12/B0_14 ),
    .i1(\inst_dob_mux_b12/B0_15 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b12/B1_7 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_1_8  (
    .i0(\inst_dob_mux_b12/B0_16 ),
    .i1(\inst_dob_mux_b12/B0_17 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b12/B1_8 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_1_9  (
    .i0(\inst_dob_mux_b12/B0_18 ),
    .i1(\inst_dob_mux_b12/B0_19 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b12/B1_9 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_2_0  (
    .i0(\inst_dob_mux_b12/B1_0 ),
    .i1(\inst_dob_mux_b12/B1_1 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b12/B2_0 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_2_1  (
    .i0(\inst_dob_mux_b12/B1_2 ),
    .i1(\inst_dob_mux_b12/B1_3 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b12/B2_1 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_2_10  (
    .i0(\inst_dob_mux_b12/B1_20 ),
    .i1(\inst_dob_mux_b12/B1_21 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b12/B2_10 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_2_11  (
    .i0(\inst_dob_mux_b12/B1_22 ),
    .i1(\inst_dob_mux_b12/B1_23 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b12/B2_11 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_2_12  (
    .i0(\inst_dob_mux_b12/B1_24 ),
    .i1(\inst_dob_mux_b12/B1_25 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b12/B2_12 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_2_13  (
    .i0(\inst_dob_mux_b12/B1_26 ),
    .i1(\inst_dob_mux_b12/B1_27 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b12/B2_13 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_2_14  (
    .i0(\inst_dob_mux_b12/B1_28 ),
    .i1(\inst_dob_mux_b12/B1_29 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b12/B2_14 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_2_15  (
    .i0(\inst_dob_mux_b12/B1_30 ),
    .i1(\inst_dob_mux_b12/B1_31 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b12/B2_15 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_2_2  (
    .i0(\inst_dob_mux_b12/B1_4 ),
    .i1(\inst_dob_mux_b12/B1_5 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b12/B2_2 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_2_3  (
    .i0(\inst_dob_mux_b12/B1_6 ),
    .i1(\inst_dob_mux_b12/B1_7 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b12/B2_3 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_2_4  (
    .i0(\inst_dob_mux_b12/B1_8 ),
    .i1(\inst_dob_mux_b12/B1_9 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b12/B2_4 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_2_5  (
    .i0(\inst_dob_mux_b12/B1_10 ),
    .i1(\inst_dob_mux_b12/B1_11 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b12/B2_5 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_2_6  (
    .i0(\inst_dob_mux_b12/B1_12 ),
    .i1(\inst_dob_mux_b12/B1_13 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b12/B2_6 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_2_7  (
    .i0(\inst_dob_mux_b12/B1_14 ),
    .i1(\inst_dob_mux_b12/B1_15 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b12/B2_7 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_2_8  (
    .i0(\inst_dob_mux_b12/B1_16 ),
    .i1(\inst_dob_mux_b12/B1_17 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b12/B2_8 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_2_9  (
    .i0(\inst_dob_mux_b12/B1_18 ),
    .i1(\inst_dob_mux_b12/B1_19 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b12/B2_9 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_3_0  (
    .i0(\inst_dob_mux_b12/B2_0 ),
    .i1(\inst_dob_mux_b12/B2_1 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b12/B3_0 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_3_1  (
    .i0(\inst_dob_mux_b12/B2_2 ),
    .i1(\inst_dob_mux_b12/B2_3 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b12/B3_1 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_3_2  (
    .i0(\inst_dob_mux_b12/B2_4 ),
    .i1(\inst_dob_mux_b12/B2_5 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b12/B3_2 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_3_3  (
    .i0(\inst_dob_mux_b12/B2_6 ),
    .i1(\inst_dob_mux_b12/B2_7 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b12/B3_3 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_3_4  (
    .i0(\inst_dob_mux_b12/B2_8 ),
    .i1(\inst_dob_mux_b12/B2_9 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b12/B3_4 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_3_5  (
    .i0(\inst_dob_mux_b12/B2_10 ),
    .i1(\inst_dob_mux_b12/B2_11 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b12/B3_5 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_3_6  (
    .i0(\inst_dob_mux_b12/B2_12 ),
    .i1(\inst_dob_mux_b12/B2_13 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b12/B3_6 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_3_7  (
    .i0(\inst_dob_mux_b12/B2_14 ),
    .i1(\inst_dob_mux_b12/B2_15 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b12/B3_7 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_4_0  (
    .i0(\inst_dob_mux_b12/B3_0 ),
    .i1(\inst_dob_mux_b12/B3_1 ),
    .sel(addrb_piped_piped[4]),
    .o(\inst_dob_mux_b12/B4_0 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_4_1  (
    .i0(\inst_dob_mux_b12/B3_2 ),
    .i1(\inst_dob_mux_b12/B3_3 ),
    .sel(addrb_piped_piped[4]),
    .o(\inst_dob_mux_b12/B4_1 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_4_2  (
    .i0(\inst_dob_mux_b12/B3_4 ),
    .i1(\inst_dob_mux_b12/B3_5 ),
    .sel(addrb_piped_piped[4]),
    .o(\inst_dob_mux_b12/B4_2 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_4_3  (
    .i0(\inst_dob_mux_b12/B3_6 ),
    .i1(\inst_dob_mux_b12/B3_7 ),
    .sel(addrb_piped_piped[4]),
    .o(\inst_dob_mux_b12/B4_3 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_5_0  (
    .i0(\inst_dob_mux_b12/B4_0 ),
    .i1(\inst_dob_mux_b12/B4_1 ),
    .sel(addrb_piped_piped[5]),
    .o(\inst_dob_mux_b12/B5_0 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_5_1  (
    .i0(\inst_dob_mux_b12/B4_2 ),
    .i1(\inst_dob_mux_b12/B4_3 ),
    .sel(addrb_piped_piped[5]),
    .o(\inst_dob_mux_b12/B5_1 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_6_0  (
    .i0(\inst_dob_mux_b12/B5_0 ),
    .i1(\inst_dob_mux_b12/B5_1 ),
    .sel(addrb_piped_piped[6]),
    .o(dob[12]));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_0  (
    .i0(inst_dob_i0_013),
    .i1(inst_dob_i0_013),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b13/B0_0 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_1  (
    .i0(inst_dob_i0_013),
    .i1(inst_dob_i0_013),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b13/B0_1 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_10  (
    .i0(inst_dob_i16_013),
    .i1(inst_dob_i16_013),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b13/B0_10 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_11  (
    .i0(inst_dob_i16_013),
    .i1(inst_dob_i16_013),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b13/B0_11 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_12  (
    .i0(inst_dob_i16_013),
    .i1(inst_dob_i16_013),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b13/B0_12 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_13  (
    .i0(inst_dob_i16_013),
    .i1(inst_dob_i16_013),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b13/B0_13 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_14  (
    .i0(inst_dob_i16_013),
    .i1(inst_dob_i16_013),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b13/B0_14 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_15  (
    .i0(inst_dob_i16_013),
    .i1(inst_dob_i16_013),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b13/B0_15 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_16  (
    .i0(inst_dob_i32_013),
    .i1(inst_dob_i32_013),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b13/B0_16 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_17  (
    .i0(inst_dob_i32_013),
    .i1(inst_dob_i32_013),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b13/B0_17 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_18  (
    .i0(inst_dob_i32_013),
    .i1(inst_dob_i32_013),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b13/B0_18 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_19  (
    .i0(inst_dob_i32_013),
    .i1(inst_dob_i32_013),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b13/B0_19 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_2  (
    .i0(inst_dob_i0_013),
    .i1(inst_dob_i0_013),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b13/B0_2 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_20  (
    .i0(inst_dob_i32_013),
    .i1(inst_dob_i32_013),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b13/B0_20 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_21  (
    .i0(inst_dob_i32_013),
    .i1(inst_dob_i32_013),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b13/B0_21 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_22  (
    .i0(inst_dob_i32_013),
    .i1(inst_dob_i32_013),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b13/B0_22 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_23  (
    .i0(inst_dob_i32_013),
    .i1(inst_dob_i32_013),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b13/B0_23 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_24  (
    .i0(inst_dob_i48_013),
    .i1(inst_dob_i48_013),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b13/B0_24 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_25  (
    .i0(inst_dob_i48_013),
    .i1(inst_dob_i48_013),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b13/B0_25 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_26  (
    .i0(inst_dob_i48_013),
    .i1(inst_dob_i48_013),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b13/B0_26 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_27  (
    .i0(inst_dob_i48_013),
    .i1(inst_dob_i48_013),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b13/B0_27 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_28  (
    .i0(inst_dob_i48_013),
    .i1(inst_dob_i48_013),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b13/B0_28 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_29  (
    .i0(inst_dob_i48_013),
    .i1(inst_dob_i48_013),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b13/B0_29 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_3  (
    .i0(inst_dob_i0_013),
    .i1(inst_dob_i0_013),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b13/B0_3 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_30  (
    .i0(inst_dob_i48_013),
    .i1(inst_dob_i48_013),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b13/B0_30 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_31  (
    .i0(inst_dob_i48_013),
    .i1(inst_dob_i48_013),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b13/B0_31 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_32  (
    .i0(inst_dob_i64_013),
    .i1(inst_dob_i64_013),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b13/B0_32 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_33  (
    .i0(inst_dob_i64_013),
    .i1(inst_dob_i64_013),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b13/B0_33 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_34  (
    .i0(inst_dob_i64_013),
    .i1(inst_dob_i64_013),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b13/B0_34 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_35  (
    .i0(inst_dob_i64_013),
    .i1(inst_dob_i64_013),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b13/B0_35 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_36  (
    .i0(inst_dob_i64_013),
    .i1(inst_dob_i64_013),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b13/B0_36 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_37  (
    .i0(inst_dob_i64_013),
    .i1(inst_dob_i64_013),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b13/B0_37 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_38  (
    .i0(inst_dob_i64_013),
    .i1(inst_dob_i64_013),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b13/B0_38 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_39  (
    .i0(inst_dob_i64_013),
    .i1(inst_dob_i64_013),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b13/B0_39 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_4  (
    .i0(inst_dob_i0_013),
    .i1(inst_dob_i0_013),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b13/B0_4 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_40  (
    .i0(inst_dob_i64_013),
    .i1(inst_dob_i64_013),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b13/B0_40 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_41  (
    .i0(inst_dob_i64_013),
    .i1(inst_dob_i64_013),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b13/B0_41 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_42  (
    .i0(inst_dob_i64_013),
    .i1(inst_dob_i64_013),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b13/B0_42 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_43  (
    .i0(inst_dob_i64_013),
    .i1(inst_dob_i64_013),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b13/B0_43 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_44  (
    .i0(inst_dob_i64_013),
    .i1(inst_dob_i64_013),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b13/B0_44 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_45  (
    .i0(inst_dob_i64_013),
    .i1(inst_dob_i64_013),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b13/B0_45 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_46  (
    .i0(inst_dob_i64_013),
    .i1(inst_dob_i64_013),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b13/B0_46 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_47  (
    .i0(inst_dob_i64_013),
    .i1(inst_dob_i64_013),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b13/B0_47 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_48  (
    .i0(inst_dob_i64_013),
    .i1(inst_dob_i64_013),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b13/B0_48 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_49  (
    .i0(inst_dob_i64_013),
    .i1(inst_dob_i64_013),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b13/B0_49 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_5  (
    .i0(inst_dob_i0_013),
    .i1(inst_dob_i0_013),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b13/B0_5 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_50  (
    .i0(inst_dob_i64_013),
    .i1(inst_dob_i64_013),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b13/B0_50 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_51  (
    .i0(inst_dob_i64_013),
    .i1(inst_dob_i64_013),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b13/B0_51 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_52  (
    .i0(inst_dob_i64_013),
    .i1(inst_dob_i64_013),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b13/B0_52 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_53  (
    .i0(inst_dob_i64_013),
    .i1(inst_dob_i64_013),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b13/B0_53 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_54  (
    .i0(inst_dob_i64_013),
    .i1(inst_dob_i64_013),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b13/B0_54 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_55  (
    .i0(inst_dob_i64_013),
    .i1(inst_dob_i64_013),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b13/B0_55 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_56  (
    .i0(inst_dob_i64_013),
    .i1(inst_dob_i64_013),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b13/B0_56 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_57  (
    .i0(inst_dob_i64_013),
    .i1(inst_dob_i64_013),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b13/B0_57 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_58  (
    .i0(inst_dob_i64_013),
    .i1(inst_dob_i64_013),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b13/B0_58 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_59  (
    .i0(inst_dob_i64_013),
    .i1(inst_dob_i64_013),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b13/B0_59 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_6  (
    .i0(inst_dob_i0_013),
    .i1(inst_dob_i0_013),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b13/B0_6 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_60  (
    .i0(inst_dob_i64_013),
    .i1(inst_dob_i64_013),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b13/B0_60 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_61  (
    .i0(inst_dob_i64_013),
    .i1(inst_dob_i64_013),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b13/B0_61 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_62  (
    .i0(inst_dob_i64_013),
    .i1(inst_dob_i64_013),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b13/B0_62 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_63  (
    .i0(inst_dob_i64_013),
    .i1(inst_dob_i64_013),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b13/B0_63 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_7  (
    .i0(inst_dob_i0_013),
    .i1(inst_dob_i0_013),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b13/B0_7 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_8  (
    .i0(inst_dob_i16_013),
    .i1(inst_dob_i16_013),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b13/B0_8 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_9  (
    .i0(inst_dob_i16_013),
    .i1(inst_dob_i16_013),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b13/B0_9 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_1_0  (
    .i0(\inst_dob_mux_b13/B0_0 ),
    .i1(\inst_dob_mux_b13/B0_1 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b13/B1_0 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_1_1  (
    .i0(\inst_dob_mux_b13/B0_2 ),
    .i1(\inst_dob_mux_b13/B0_3 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b13/B1_1 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_1_10  (
    .i0(\inst_dob_mux_b13/B0_20 ),
    .i1(\inst_dob_mux_b13/B0_21 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b13/B1_10 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_1_11  (
    .i0(\inst_dob_mux_b13/B0_22 ),
    .i1(\inst_dob_mux_b13/B0_23 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b13/B1_11 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_1_12  (
    .i0(\inst_dob_mux_b13/B0_24 ),
    .i1(\inst_dob_mux_b13/B0_25 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b13/B1_12 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_1_13  (
    .i0(\inst_dob_mux_b13/B0_26 ),
    .i1(\inst_dob_mux_b13/B0_27 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b13/B1_13 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_1_14  (
    .i0(\inst_dob_mux_b13/B0_28 ),
    .i1(\inst_dob_mux_b13/B0_29 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b13/B1_14 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_1_15  (
    .i0(\inst_dob_mux_b13/B0_30 ),
    .i1(\inst_dob_mux_b13/B0_31 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b13/B1_15 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_1_16  (
    .i0(\inst_dob_mux_b13/B0_32 ),
    .i1(\inst_dob_mux_b13/B0_33 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b13/B1_16 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_1_17  (
    .i0(\inst_dob_mux_b13/B0_34 ),
    .i1(\inst_dob_mux_b13/B0_35 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b13/B1_17 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_1_18  (
    .i0(\inst_dob_mux_b13/B0_36 ),
    .i1(\inst_dob_mux_b13/B0_37 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b13/B1_18 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_1_19  (
    .i0(\inst_dob_mux_b13/B0_38 ),
    .i1(\inst_dob_mux_b13/B0_39 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b13/B1_19 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_1_2  (
    .i0(\inst_dob_mux_b13/B0_4 ),
    .i1(\inst_dob_mux_b13/B0_5 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b13/B1_2 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_1_20  (
    .i0(\inst_dob_mux_b13/B0_40 ),
    .i1(\inst_dob_mux_b13/B0_41 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b13/B1_20 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_1_21  (
    .i0(\inst_dob_mux_b13/B0_42 ),
    .i1(\inst_dob_mux_b13/B0_43 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b13/B1_21 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_1_22  (
    .i0(\inst_dob_mux_b13/B0_44 ),
    .i1(\inst_dob_mux_b13/B0_45 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b13/B1_22 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_1_23  (
    .i0(\inst_dob_mux_b13/B0_46 ),
    .i1(\inst_dob_mux_b13/B0_47 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b13/B1_23 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_1_24  (
    .i0(\inst_dob_mux_b13/B0_48 ),
    .i1(\inst_dob_mux_b13/B0_49 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b13/B1_24 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_1_25  (
    .i0(\inst_dob_mux_b13/B0_50 ),
    .i1(\inst_dob_mux_b13/B0_51 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b13/B1_25 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_1_26  (
    .i0(\inst_dob_mux_b13/B0_52 ),
    .i1(\inst_dob_mux_b13/B0_53 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b13/B1_26 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_1_27  (
    .i0(\inst_dob_mux_b13/B0_54 ),
    .i1(\inst_dob_mux_b13/B0_55 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b13/B1_27 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_1_28  (
    .i0(\inst_dob_mux_b13/B0_56 ),
    .i1(\inst_dob_mux_b13/B0_57 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b13/B1_28 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_1_29  (
    .i0(\inst_dob_mux_b13/B0_58 ),
    .i1(\inst_dob_mux_b13/B0_59 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b13/B1_29 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_1_3  (
    .i0(\inst_dob_mux_b13/B0_6 ),
    .i1(\inst_dob_mux_b13/B0_7 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b13/B1_3 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_1_30  (
    .i0(\inst_dob_mux_b13/B0_60 ),
    .i1(\inst_dob_mux_b13/B0_61 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b13/B1_30 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_1_31  (
    .i0(\inst_dob_mux_b13/B0_62 ),
    .i1(\inst_dob_mux_b13/B0_63 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b13/B1_31 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_1_4  (
    .i0(\inst_dob_mux_b13/B0_8 ),
    .i1(\inst_dob_mux_b13/B0_9 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b13/B1_4 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_1_5  (
    .i0(\inst_dob_mux_b13/B0_10 ),
    .i1(\inst_dob_mux_b13/B0_11 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b13/B1_5 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_1_6  (
    .i0(\inst_dob_mux_b13/B0_12 ),
    .i1(\inst_dob_mux_b13/B0_13 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b13/B1_6 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_1_7  (
    .i0(\inst_dob_mux_b13/B0_14 ),
    .i1(\inst_dob_mux_b13/B0_15 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b13/B1_7 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_1_8  (
    .i0(\inst_dob_mux_b13/B0_16 ),
    .i1(\inst_dob_mux_b13/B0_17 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b13/B1_8 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_1_9  (
    .i0(\inst_dob_mux_b13/B0_18 ),
    .i1(\inst_dob_mux_b13/B0_19 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b13/B1_9 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_2_0  (
    .i0(\inst_dob_mux_b13/B1_0 ),
    .i1(\inst_dob_mux_b13/B1_1 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b13/B2_0 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_2_1  (
    .i0(\inst_dob_mux_b13/B1_2 ),
    .i1(\inst_dob_mux_b13/B1_3 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b13/B2_1 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_2_10  (
    .i0(\inst_dob_mux_b13/B1_20 ),
    .i1(\inst_dob_mux_b13/B1_21 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b13/B2_10 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_2_11  (
    .i0(\inst_dob_mux_b13/B1_22 ),
    .i1(\inst_dob_mux_b13/B1_23 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b13/B2_11 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_2_12  (
    .i0(\inst_dob_mux_b13/B1_24 ),
    .i1(\inst_dob_mux_b13/B1_25 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b13/B2_12 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_2_13  (
    .i0(\inst_dob_mux_b13/B1_26 ),
    .i1(\inst_dob_mux_b13/B1_27 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b13/B2_13 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_2_14  (
    .i0(\inst_dob_mux_b13/B1_28 ),
    .i1(\inst_dob_mux_b13/B1_29 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b13/B2_14 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_2_15  (
    .i0(\inst_dob_mux_b13/B1_30 ),
    .i1(\inst_dob_mux_b13/B1_31 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b13/B2_15 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_2_2  (
    .i0(\inst_dob_mux_b13/B1_4 ),
    .i1(\inst_dob_mux_b13/B1_5 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b13/B2_2 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_2_3  (
    .i0(\inst_dob_mux_b13/B1_6 ),
    .i1(\inst_dob_mux_b13/B1_7 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b13/B2_3 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_2_4  (
    .i0(\inst_dob_mux_b13/B1_8 ),
    .i1(\inst_dob_mux_b13/B1_9 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b13/B2_4 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_2_5  (
    .i0(\inst_dob_mux_b13/B1_10 ),
    .i1(\inst_dob_mux_b13/B1_11 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b13/B2_5 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_2_6  (
    .i0(\inst_dob_mux_b13/B1_12 ),
    .i1(\inst_dob_mux_b13/B1_13 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b13/B2_6 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_2_7  (
    .i0(\inst_dob_mux_b13/B1_14 ),
    .i1(\inst_dob_mux_b13/B1_15 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b13/B2_7 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_2_8  (
    .i0(\inst_dob_mux_b13/B1_16 ),
    .i1(\inst_dob_mux_b13/B1_17 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b13/B2_8 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_2_9  (
    .i0(\inst_dob_mux_b13/B1_18 ),
    .i1(\inst_dob_mux_b13/B1_19 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b13/B2_9 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_3_0  (
    .i0(\inst_dob_mux_b13/B2_0 ),
    .i1(\inst_dob_mux_b13/B2_1 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b13/B3_0 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_3_1  (
    .i0(\inst_dob_mux_b13/B2_2 ),
    .i1(\inst_dob_mux_b13/B2_3 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b13/B3_1 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_3_2  (
    .i0(\inst_dob_mux_b13/B2_4 ),
    .i1(\inst_dob_mux_b13/B2_5 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b13/B3_2 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_3_3  (
    .i0(\inst_dob_mux_b13/B2_6 ),
    .i1(\inst_dob_mux_b13/B2_7 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b13/B3_3 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_3_4  (
    .i0(\inst_dob_mux_b13/B2_8 ),
    .i1(\inst_dob_mux_b13/B2_9 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b13/B3_4 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_3_5  (
    .i0(\inst_dob_mux_b13/B2_10 ),
    .i1(\inst_dob_mux_b13/B2_11 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b13/B3_5 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_3_6  (
    .i0(\inst_dob_mux_b13/B2_12 ),
    .i1(\inst_dob_mux_b13/B2_13 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b13/B3_6 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_3_7  (
    .i0(\inst_dob_mux_b13/B2_14 ),
    .i1(\inst_dob_mux_b13/B2_15 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b13/B3_7 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_4_0  (
    .i0(\inst_dob_mux_b13/B3_0 ),
    .i1(\inst_dob_mux_b13/B3_1 ),
    .sel(addrb_piped_piped[4]),
    .o(\inst_dob_mux_b13/B4_0 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_4_1  (
    .i0(\inst_dob_mux_b13/B3_2 ),
    .i1(\inst_dob_mux_b13/B3_3 ),
    .sel(addrb_piped_piped[4]),
    .o(\inst_dob_mux_b13/B4_1 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_4_2  (
    .i0(\inst_dob_mux_b13/B3_4 ),
    .i1(\inst_dob_mux_b13/B3_5 ),
    .sel(addrb_piped_piped[4]),
    .o(\inst_dob_mux_b13/B4_2 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_4_3  (
    .i0(\inst_dob_mux_b13/B3_6 ),
    .i1(\inst_dob_mux_b13/B3_7 ),
    .sel(addrb_piped_piped[4]),
    .o(\inst_dob_mux_b13/B4_3 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_5_0  (
    .i0(\inst_dob_mux_b13/B4_0 ),
    .i1(\inst_dob_mux_b13/B4_1 ),
    .sel(addrb_piped_piped[5]),
    .o(\inst_dob_mux_b13/B5_0 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_5_1  (
    .i0(\inst_dob_mux_b13/B4_2 ),
    .i1(\inst_dob_mux_b13/B4_3 ),
    .sel(addrb_piped_piped[5]),
    .o(\inst_dob_mux_b13/B5_1 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_6_0  (
    .i0(\inst_dob_mux_b13/B5_0 ),
    .i1(\inst_dob_mux_b13/B5_1 ),
    .sel(addrb_piped_piped[6]),
    .o(dob[13]));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_0  (
    .i0(inst_dob_i0_014),
    .i1(inst_dob_i0_014),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b14/B0_0 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_1  (
    .i0(inst_dob_i0_014),
    .i1(inst_dob_i0_014),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b14/B0_1 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_10  (
    .i0(inst_dob_i16_014),
    .i1(inst_dob_i16_014),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b14/B0_10 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_11  (
    .i0(inst_dob_i16_014),
    .i1(inst_dob_i16_014),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b14/B0_11 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_12  (
    .i0(inst_dob_i16_014),
    .i1(inst_dob_i16_014),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b14/B0_12 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_13  (
    .i0(inst_dob_i16_014),
    .i1(inst_dob_i16_014),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b14/B0_13 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_14  (
    .i0(inst_dob_i16_014),
    .i1(inst_dob_i16_014),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b14/B0_14 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_15  (
    .i0(inst_dob_i16_014),
    .i1(inst_dob_i16_014),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b14/B0_15 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_16  (
    .i0(inst_dob_i32_014),
    .i1(inst_dob_i32_014),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b14/B0_16 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_17  (
    .i0(inst_dob_i32_014),
    .i1(inst_dob_i32_014),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b14/B0_17 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_18  (
    .i0(inst_dob_i32_014),
    .i1(inst_dob_i32_014),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b14/B0_18 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_19  (
    .i0(inst_dob_i32_014),
    .i1(inst_dob_i32_014),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b14/B0_19 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_2  (
    .i0(inst_dob_i0_014),
    .i1(inst_dob_i0_014),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b14/B0_2 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_20  (
    .i0(inst_dob_i32_014),
    .i1(inst_dob_i32_014),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b14/B0_20 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_21  (
    .i0(inst_dob_i32_014),
    .i1(inst_dob_i32_014),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b14/B0_21 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_22  (
    .i0(inst_dob_i32_014),
    .i1(inst_dob_i32_014),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b14/B0_22 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_23  (
    .i0(inst_dob_i32_014),
    .i1(inst_dob_i32_014),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b14/B0_23 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_24  (
    .i0(inst_dob_i48_014),
    .i1(inst_dob_i48_014),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b14/B0_24 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_25  (
    .i0(inst_dob_i48_014),
    .i1(inst_dob_i48_014),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b14/B0_25 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_26  (
    .i0(inst_dob_i48_014),
    .i1(inst_dob_i48_014),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b14/B0_26 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_27  (
    .i0(inst_dob_i48_014),
    .i1(inst_dob_i48_014),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b14/B0_27 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_28  (
    .i0(inst_dob_i48_014),
    .i1(inst_dob_i48_014),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b14/B0_28 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_29  (
    .i0(inst_dob_i48_014),
    .i1(inst_dob_i48_014),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b14/B0_29 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_3  (
    .i0(inst_dob_i0_014),
    .i1(inst_dob_i0_014),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b14/B0_3 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_30  (
    .i0(inst_dob_i48_014),
    .i1(inst_dob_i48_014),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b14/B0_30 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_31  (
    .i0(inst_dob_i48_014),
    .i1(inst_dob_i48_014),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b14/B0_31 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_32  (
    .i0(inst_dob_i64_014),
    .i1(inst_dob_i64_014),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b14/B0_32 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_33  (
    .i0(inst_dob_i64_014),
    .i1(inst_dob_i64_014),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b14/B0_33 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_34  (
    .i0(inst_dob_i64_014),
    .i1(inst_dob_i64_014),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b14/B0_34 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_35  (
    .i0(inst_dob_i64_014),
    .i1(inst_dob_i64_014),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b14/B0_35 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_36  (
    .i0(inst_dob_i64_014),
    .i1(inst_dob_i64_014),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b14/B0_36 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_37  (
    .i0(inst_dob_i64_014),
    .i1(inst_dob_i64_014),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b14/B0_37 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_38  (
    .i0(inst_dob_i64_014),
    .i1(inst_dob_i64_014),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b14/B0_38 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_39  (
    .i0(inst_dob_i64_014),
    .i1(inst_dob_i64_014),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b14/B0_39 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_4  (
    .i0(inst_dob_i0_014),
    .i1(inst_dob_i0_014),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b14/B0_4 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_40  (
    .i0(inst_dob_i64_014),
    .i1(inst_dob_i64_014),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b14/B0_40 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_41  (
    .i0(inst_dob_i64_014),
    .i1(inst_dob_i64_014),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b14/B0_41 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_42  (
    .i0(inst_dob_i64_014),
    .i1(inst_dob_i64_014),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b14/B0_42 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_43  (
    .i0(inst_dob_i64_014),
    .i1(inst_dob_i64_014),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b14/B0_43 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_44  (
    .i0(inst_dob_i64_014),
    .i1(inst_dob_i64_014),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b14/B0_44 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_45  (
    .i0(inst_dob_i64_014),
    .i1(inst_dob_i64_014),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b14/B0_45 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_46  (
    .i0(inst_dob_i64_014),
    .i1(inst_dob_i64_014),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b14/B0_46 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_47  (
    .i0(inst_dob_i64_014),
    .i1(inst_dob_i64_014),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b14/B0_47 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_48  (
    .i0(inst_dob_i64_014),
    .i1(inst_dob_i64_014),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b14/B0_48 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_49  (
    .i0(inst_dob_i64_014),
    .i1(inst_dob_i64_014),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b14/B0_49 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_5  (
    .i0(inst_dob_i0_014),
    .i1(inst_dob_i0_014),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b14/B0_5 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_50  (
    .i0(inst_dob_i64_014),
    .i1(inst_dob_i64_014),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b14/B0_50 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_51  (
    .i0(inst_dob_i64_014),
    .i1(inst_dob_i64_014),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b14/B0_51 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_52  (
    .i0(inst_dob_i64_014),
    .i1(inst_dob_i64_014),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b14/B0_52 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_53  (
    .i0(inst_dob_i64_014),
    .i1(inst_dob_i64_014),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b14/B0_53 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_54  (
    .i0(inst_dob_i64_014),
    .i1(inst_dob_i64_014),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b14/B0_54 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_55  (
    .i0(inst_dob_i64_014),
    .i1(inst_dob_i64_014),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b14/B0_55 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_56  (
    .i0(inst_dob_i64_014),
    .i1(inst_dob_i64_014),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b14/B0_56 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_57  (
    .i0(inst_dob_i64_014),
    .i1(inst_dob_i64_014),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b14/B0_57 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_58  (
    .i0(inst_dob_i64_014),
    .i1(inst_dob_i64_014),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b14/B0_58 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_59  (
    .i0(inst_dob_i64_014),
    .i1(inst_dob_i64_014),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b14/B0_59 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_6  (
    .i0(inst_dob_i0_014),
    .i1(inst_dob_i0_014),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b14/B0_6 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_60  (
    .i0(inst_dob_i64_014),
    .i1(inst_dob_i64_014),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b14/B0_60 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_61  (
    .i0(inst_dob_i64_014),
    .i1(inst_dob_i64_014),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b14/B0_61 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_62  (
    .i0(inst_dob_i64_014),
    .i1(inst_dob_i64_014),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b14/B0_62 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_63  (
    .i0(inst_dob_i64_014),
    .i1(inst_dob_i64_014),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b14/B0_63 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_7  (
    .i0(inst_dob_i0_014),
    .i1(inst_dob_i0_014),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b14/B0_7 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_8  (
    .i0(inst_dob_i16_014),
    .i1(inst_dob_i16_014),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b14/B0_8 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_9  (
    .i0(inst_dob_i16_014),
    .i1(inst_dob_i16_014),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b14/B0_9 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_1_0  (
    .i0(\inst_dob_mux_b14/B0_0 ),
    .i1(\inst_dob_mux_b14/B0_1 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b14/B1_0 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_1_1  (
    .i0(\inst_dob_mux_b14/B0_2 ),
    .i1(\inst_dob_mux_b14/B0_3 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b14/B1_1 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_1_10  (
    .i0(\inst_dob_mux_b14/B0_20 ),
    .i1(\inst_dob_mux_b14/B0_21 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b14/B1_10 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_1_11  (
    .i0(\inst_dob_mux_b14/B0_22 ),
    .i1(\inst_dob_mux_b14/B0_23 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b14/B1_11 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_1_12  (
    .i0(\inst_dob_mux_b14/B0_24 ),
    .i1(\inst_dob_mux_b14/B0_25 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b14/B1_12 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_1_13  (
    .i0(\inst_dob_mux_b14/B0_26 ),
    .i1(\inst_dob_mux_b14/B0_27 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b14/B1_13 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_1_14  (
    .i0(\inst_dob_mux_b14/B0_28 ),
    .i1(\inst_dob_mux_b14/B0_29 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b14/B1_14 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_1_15  (
    .i0(\inst_dob_mux_b14/B0_30 ),
    .i1(\inst_dob_mux_b14/B0_31 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b14/B1_15 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_1_16  (
    .i0(\inst_dob_mux_b14/B0_32 ),
    .i1(\inst_dob_mux_b14/B0_33 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b14/B1_16 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_1_17  (
    .i0(\inst_dob_mux_b14/B0_34 ),
    .i1(\inst_dob_mux_b14/B0_35 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b14/B1_17 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_1_18  (
    .i0(\inst_dob_mux_b14/B0_36 ),
    .i1(\inst_dob_mux_b14/B0_37 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b14/B1_18 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_1_19  (
    .i0(\inst_dob_mux_b14/B0_38 ),
    .i1(\inst_dob_mux_b14/B0_39 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b14/B1_19 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_1_2  (
    .i0(\inst_dob_mux_b14/B0_4 ),
    .i1(\inst_dob_mux_b14/B0_5 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b14/B1_2 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_1_20  (
    .i0(\inst_dob_mux_b14/B0_40 ),
    .i1(\inst_dob_mux_b14/B0_41 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b14/B1_20 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_1_21  (
    .i0(\inst_dob_mux_b14/B0_42 ),
    .i1(\inst_dob_mux_b14/B0_43 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b14/B1_21 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_1_22  (
    .i0(\inst_dob_mux_b14/B0_44 ),
    .i1(\inst_dob_mux_b14/B0_45 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b14/B1_22 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_1_23  (
    .i0(\inst_dob_mux_b14/B0_46 ),
    .i1(\inst_dob_mux_b14/B0_47 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b14/B1_23 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_1_24  (
    .i0(\inst_dob_mux_b14/B0_48 ),
    .i1(\inst_dob_mux_b14/B0_49 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b14/B1_24 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_1_25  (
    .i0(\inst_dob_mux_b14/B0_50 ),
    .i1(\inst_dob_mux_b14/B0_51 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b14/B1_25 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_1_26  (
    .i0(\inst_dob_mux_b14/B0_52 ),
    .i1(\inst_dob_mux_b14/B0_53 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b14/B1_26 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_1_27  (
    .i0(\inst_dob_mux_b14/B0_54 ),
    .i1(\inst_dob_mux_b14/B0_55 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b14/B1_27 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_1_28  (
    .i0(\inst_dob_mux_b14/B0_56 ),
    .i1(\inst_dob_mux_b14/B0_57 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b14/B1_28 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_1_29  (
    .i0(\inst_dob_mux_b14/B0_58 ),
    .i1(\inst_dob_mux_b14/B0_59 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b14/B1_29 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_1_3  (
    .i0(\inst_dob_mux_b14/B0_6 ),
    .i1(\inst_dob_mux_b14/B0_7 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b14/B1_3 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_1_30  (
    .i0(\inst_dob_mux_b14/B0_60 ),
    .i1(\inst_dob_mux_b14/B0_61 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b14/B1_30 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_1_31  (
    .i0(\inst_dob_mux_b14/B0_62 ),
    .i1(\inst_dob_mux_b14/B0_63 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b14/B1_31 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_1_4  (
    .i0(\inst_dob_mux_b14/B0_8 ),
    .i1(\inst_dob_mux_b14/B0_9 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b14/B1_4 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_1_5  (
    .i0(\inst_dob_mux_b14/B0_10 ),
    .i1(\inst_dob_mux_b14/B0_11 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b14/B1_5 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_1_6  (
    .i0(\inst_dob_mux_b14/B0_12 ),
    .i1(\inst_dob_mux_b14/B0_13 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b14/B1_6 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_1_7  (
    .i0(\inst_dob_mux_b14/B0_14 ),
    .i1(\inst_dob_mux_b14/B0_15 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b14/B1_7 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_1_8  (
    .i0(\inst_dob_mux_b14/B0_16 ),
    .i1(\inst_dob_mux_b14/B0_17 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b14/B1_8 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_1_9  (
    .i0(\inst_dob_mux_b14/B0_18 ),
    .i1(\inst_dob_mux_b14/B0_19 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b14/B1_9 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_2_0  (
    .i0(\inst_dob_mux_b14/B1_0 ),
    .i1(\inst_dob_mux_b14/B1_1 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b14/B2_0 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_2_1  (
    .i0(\inst_dob_mux_b14/B1_2 ),
    .i1(\inst_dob_mux_b14/B1_3 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b14/B2_1 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_2_10  (
    .i0(\inst_dob_mux_b14/B1_20 ),
    .i1(\inst_dob_mux_b14/B1_21 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b14/B2_10 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_2_11  (
    .i0(\inst_dob_mux_b14/B1_22 ),
    .i1(\inst_dob_mux_b14/B1_23 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b14/B2_11 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_2_12  (
    .i0(\inst_dob_mux_b14/B1_24 ),
    .i1(\inst_dob_mux_b14/B1_25 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b14/B2_12 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_2_13  (
    .i0(\inst_dob_mux_b14/B1_26 ),
    .i1(\inst_dob_mux_b14/B1_27 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b14/B2_13 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_2_14  (
    .i0(\inst_dob_mux_b14/B1_28 ),
    .i1(\inst_dob_mux_b14/B1_29 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b14/B2_14 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_2_15  (
    .i0(\inst_dob_mux_b14/B1_30 ),
    .i1(\inst_dob_mux_b14/B1_31 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b14/B2_15 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_2_2  (
    .i0(\inst_dob_mux_b14/B1_4 ),
    .i1(\inst_dob_mux_b14/B1_5 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b14/B2_2 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_2_3  (
    .i0(\inst_dob_mux_b14/B1_6 ),
    .i1(\inst_dob_mux_b14/B1_7 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b14/B2_3 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_2_4  (
    .i0(\inst_dob_mux_b14/B1_8 ),
    .i1(\inst_dob_mux_b14/B1_9 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b14/B2_4 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_2_5  (
    .i0(\inst_dob_mux_b14/B1_10 ),
    .i1(\inst_dob_mux_b14/B1_11 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b14/B2_5 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_2_6  (
    .i0(\inst_dob_mux_b14/B1_12 ),
    .i1(\inst_dob_mux_b14/B1_13 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b14/B2_6 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_2_7  (
    .i0(\inst_dob_mux_b14/B1_14 ),
    .i1(\inst_dob_mux_b14/B1_15 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b14/B2_7 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_2_8  (
    .i0(\inst_dob_mux_b14/B1_16 ),
    .i1(\inst_dob_mux_b14/B1_17 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b14/B2_8 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_2_9  (
    .i0(\inst_dob_mux_b14/B1_18 ),
    .i1(\inst_dob_mux_b14/B1_19 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b14/B2_9 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_3_0  (
    .i0(\inst_dob_mux_b14/B2_0 ),
    .i1(\inst_dob_mux_b14/B2_1 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b14/B3_0 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_3_1  (
    .i0(\inst_dob_mux_b14/B2_2 ),
    .i1(\inst_dob_mux_b14/B2_3 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b14/B3_1 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_3_2  (
    .i0(\inst_dob_mux_b14/B2_4 ),
    .i1(\inst_dob_mux_b14/B2_5 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b14/B3_2 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_3_3  (
    .i0(\inst_dob_mux_b14/B2_6 ),
    .i1(\inst_dob_mux_b14/B2_7 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b14/B3_3 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_3_4  (
    .i0(\inst_dob_mux_b14/B2_8 ),
    .i1(\inst_dob_mux_b14/B2_9 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b14/B3_4 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_3_5  (
    .i0(\inst_dob_mux_b14/B2_10 ),
    .i1(\inst_dob_mux_b14/B2_11 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b14/B3_5 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_3_6  (
    .i0(\inst_dob_mux_b14/B2_12 ),
    .i1(\inst_dob_mux_b14/B2_13 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b14/B3_6 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_3_7  (
    .i0(\inst_dob_mux_b14/B2_14 ),
    .i1(\inst_dob_mux_b14/B2_15 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b14/B3_7 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_4_0  (
    .i0(\inst_dob_mux_b14/B3_0 ),
    .i1(\inst_dob_mux_b14/B3_1 ),
    .sel(addrb_piped_piped[4]),
    .o(\inst_dob_mux_b14/B4_0 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_4_1  (
    .i0(\inst_dob_mux_b14/B3_2 ),
    .i1(\inst_dob_mux_b14/B3_3 ),
    .sel(addrb_piped_piped[4]),
    .o(\inst_dob_mux_b14/B4_1 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_4_2  (
    .i0(\inst_dob_mux_b14/B3_4 ),
    .i1(\inst_dob_mux_b14/B3_5 ),
    .sel(addrb_piped_piped[4]),
    .o(\inst_dob_mux_b14/B4_2 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_4_3  (
    .i0(\inst_dob_mux_b14/B3_6 ),
    .i1(\inst_dob_mux_b14/B3_7 ),
    .sel(addrb_piped_piped[4]),
    .o(\inst_dob_mux_b14/B4_3 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_5_0  (
    .i0(\inst_dob_mux_b14/B4_0 ),
    .i1(\inst_dob_mux_b14/B4_1 ),
    .sel(addrb_piped_piped[5]),
    .o(\inst_dob_mux_b14/B5_0 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_5_1  (
    .i0(\inst_dob_mux_b14/B4_2 ),
    .i1(\inst_dob_mux_b14/B4_3 ),
    .sel(addrb_piped_piped[5]),
    .o(\inst_dob_mux_b14/B5_1 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_6_0  (
    .i0(\inst_dob_mux_b14/B5_0 ),
    .i1(\inst_dob_mux_b14/B5_1 ),
    .sel(addrb_piped_piped[6]),
    .o(dob[14]));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_0  (
    .i0(inst_dob_i0_015),
    .i1(inst_dob_i0_015),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b15/B0_0 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_1  (
    .i0(inst_dob_i0_015),
    .i1(inst_dob_i0_015),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b15/B0_1 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_10  (
    .i0(inst_dob_i16_015),
    .i1(inst_dob_i16_015),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b15/B0_10 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_11  (
    .i0(inst_dob_i16_015),
    .i1(inst_dob_i16_015),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b15/B0_11 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_12  (
    .i0(inst_dob_i16_015),
    .i1(inst_dob_i16_015),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b15/B0_12 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_13  (
    .i0(inst_dob_i16_015),
    .i1(inst_dob_i16_015),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b15/B0_13 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_14  (
    .i0(inst_dob_i16_015),
    .i1(inst_dob_i16_015),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b15/B0_14 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_15  (
    .i0(inst_dob_i16_015),
    .i1(inst_dob_i16_015),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b15/B0_15 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_16  (
    .i0(inst_dob_i32_015),
    .i1(inst_dob_i32_015),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b15/B0_16 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_17  (
    .i0(inst_dob_i32_015),
    .i1(inst_dob_i32_015),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b15/B0_17 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_18  (
    .i0(inst_dob_i32_015),
    .i1(inst_dob_i32_015),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b15/B0_18 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_19  (
    .i0(inst_dob_i32_015),
    .i1(inst_dob_i32_015),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b15/B0_19 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_2  (
    .i0(inst_dob_i0_015),
    .i1(inst_dob_i0_015),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b15/B0_2 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_20  (
    .i0(inst_dob_i32_015),
    .i1(inst_dob_i32_015),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b15/B0_20 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_21  (
    .i0(inst_dob_i32_015),
    .i1(inst_dob_i32_015),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b15/B0_21 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_22  (
    .i0(inst_dob_i32_015),
    .i1(inst_dob_i32_015),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b15/B0_22 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_23  (
    .i0(inst_dob_i32_015),
    .i1(inst_dob_i32_015),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b15/B0_23 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_24  (
    .i0(inst_dob_i48_015),
    .i1(inst_dob_i48_015),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b15/B0_24 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_25  (
    .i0(inst_dob_i48_015),
    .i1(inst_dob_i48_015),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b15/B0_25 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_26  (
    .i0(inst_dob_i48_015),
    .i1(inst_dob_i48_015),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b15/B0_26 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_27  (
    .i0(inst_dob_i48_015),
    .i1(inst_dob_i48_015),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b15/B0_27 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_28  (
    .i0(inst_dob_i48_015),
    .i1(inst_dob_i48_015),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b15/B0_28 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_29  (
    .i0(inst_dob_i48_015),
    .i1(inst_dob_i48_015),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b15/B0_29 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_3  (
    .i0(inst_dob_i0_015),
    .i1(inst_dob_i0_015),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b15/B0_3 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_30  (
    .i0(inst_dob_i48_015),
    .i1(inst_dob_i48_015),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b15/B0_30 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_31  (
    .i0(inst_dob_i48_015),
    .i1(inst_dob_i48_015),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b15/B0_31 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_32  (
    .i0(inst_dob_i64_015),
    .i1(inst_dob_i64_015),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b15/B0_32 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_33  (
    .i0(inst_dob_i64_015),
    .i1(inst_dob_i64_015),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b15/B0_33 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_34  (
    .i0(inst_dob_i64_015),
    .i1(inst_dob_i64_015),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b15/B0_34 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_35  (
    .i0(inst_dob_i64_015),
    .i1(inst_dob_i64_015),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b15/B0_35 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_36  (
    .i0(inst_dob_i64_015),
    .i1(inst_dob_i64_015),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b15/B0_36 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_37  (
    .i0(inst_dob_i64_015),
    .i1(inst_dob_i64_015),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b15/B0_37 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_38  (
    .i0(inst_dob_i64_015),
    .i1(inst_dob_i64_015),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b15/B0_38 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_39  (
    .i0(inst_dob_i64_015),
    .i1(inst_dob_i64_015),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b15/B0_39 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_4  (
    .i0(inst_dob_i0_015),
    .i1(inst_dob_i0_015),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b15/B0_4 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_40  (
    .i0(inst_dob_i64_015),
    .i1(inst_dob_i64_015),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b15/B0_40 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_41  (
    .i0(inst_dob_i64_015),
    .i1(inst_dob_i64_015),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b15/B0_41 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_42  (
    .i0(inst_dob_i64_015),
    .i1(inst_dob_i64_015),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b15/B0_42 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_43  (
    .i0(inst_dob_i64_015),
    .i1(inst_dob_i64_015),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b15/B0_43 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_44  (
    .i0(inst_dob_i64_015),
    .i1(inst_dob_i64_015),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b15/B0_44 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_45  (
    .i0(inst_dob_i64_015),
    .i1(inst_dob_i64_015),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b15/B0_45 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_46  (
    .i0(inst_dob_i64_015),
    .i1(inst_dob_i64_015),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b15/B0_46 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_47  (
    .i0(inst_dob_i64_015),
    .i1(inst_dob_i64_015),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b15/B0_47 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_48  (
    .i0(inst_dob_i64_015),
    .i1(inst_dob_i64_015),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b15/B0_48 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_49  (
    .i0(inst_dob_i64_015),
    .i1(inst_dob_i64_015),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b15/B0_49 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_5  (
    .i0(inst_dob_i0_015),
    .i1(inst_dob_i0_015),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b15/B0_5 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_50  (
    .i0(inst_dob_i64_015),
    .i1(inst_dob_i64_015),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b15/B0_50 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_51  (
    .i0(inst_dob_i64_015),
    .i1(inst_dob_i64_015),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b15/B0_51 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_52  (
    .i0(inst_dob_i64_015),
    .i1(inst_dob_i64_015),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b15/B0_52 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_53  (
    .i0(inst_dob_i64_015),
    .i1(inst_dob_i64_015),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b15/B0_53 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_54  (
    .i0(inst_dob_i64_015),
    .i1(inst_dob_i64_015),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b15/B0_54 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_55  (
    .i0(inst_dob_i64_015),
    .i1(inst_dob_i64_015),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b15/B0_55 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_56  (
    .i0(inst_dob_i64_015),
    .i1(inst_dob_i64_015),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b15/B0_56 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_57  (
    .i0(inst_dob_i64_015),
    .i1(inst_dob_i64_015),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b15/B0_57 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_58  (
    .i0(inst_dob_i64_015),
    .i1(inst_dob_i64_015),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b15/B0_58 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_59  (
    .i0(inst_dob_i64_015),
    .i1(inst_dob_i64_015),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b15/B0_59 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_6  (
    .i0(inst_dob_i0_015),
    .i1(inst_dob_i0_015),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b15/B0_6 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_60  (
    .i0(inst_dob_i64_015),
    .i1(inst_dob_i64_015),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b15/B0_60 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_61  (
    .i0(inst_dob_i64_015),
    .i1(inst_dob_i64_015),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b15/B0_61 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_62  (
    .i0(inst_dob_i64_015),
    .i1(inst_dob_i64_015),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b15/B0_62 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_63  (
    .i0(inst_dob_i64_015),
    .i1(inst_dob_i64_015),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b15/B0_63 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_7  (
    .i0(inst_dob_i0_015),
    .i1(inst_dob_i0_015),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b15/B0_7 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_8  (
    .i0(inst_dob_i16_015),
    .i1(inst_dob_i16_015),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b15/B0_8 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_9  (
    .i0(inst_dob_i16_015),
    .i1(inst_dob_i16_015),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b15/B0_9 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_1_0  (
    .i0(\inst_dob_mux_b15/B0_0 ),
    .i1(\inst_dob_mux_b15/B0_1 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b15/B1_0 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_1_1  (
    .i0(\inst_dob_mux_b15/B0_2 ),
    .i1(\inst_dob_mux_b15/B0_3 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b15/B1_1 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_1_10  (
    .i0(\inst_dob_mux_b15/B0_20 ),
    .i1(\inst_dob_mux_b15/B0_21 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b15/B1_10 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_1_11  (
    .i0(\inst_dob_mux_b15/B0_22 ),
    .i1(\inst_dob_mux_b15/B0_23 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b15/B1_11 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_1_12  (
    .i0(\inst_dob_mux_b15/B0_24 ),
    .i1(\inst_dob_mux_b15/B0_25 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b15/B1_12 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_1_13  (
    .i0(\inst_dob_mux_b15/B0_26 ),
    .i1(\inst_dob_mux_b15/B0_27 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b15/B1_13 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_1_14  (
    .i0(\inst_dob_mux_b15/B0_28 ),
    .i1(\inst_dob_mux_b15/B0_29 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b15/B1_14 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_1_15  (
    .i0(\inst_dob_mux_b15/B0_30 ),
    .i1(\inst_dob_mux_b15/B0_31 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b15/B1_15 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_1_16  (
    .i0(\inst_dob_mux_b15/B0_32 ),
    .i1(\inst_dob_mux_b15/B0_33 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b15/B1_16 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_1_17  (
    .i0(\inst_dob_mux_b15/B0_34 ),
    .i1(\inst_dob_mux_b15/B0_35 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b15/B1_17 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_1_18  (
    .i0(\inst_dob_mux_b15/B0_36 ),
    .i1(\inst_dob_mux_b15/B0_37 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b15/B1_18 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_1_19  (
    .i0(\inst_dob_mux_b15/B0_38 ),
    .i1(\inst_dob_mux_b15/B0_39 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b15/B1_19 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_1_2  (
    .i0(\inst_dob_mux_b15/B0_4 ),
    .i1(\inst_dob_mux_b15/B0_5 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b15/B1_2 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_1_20  (
    .i0(\inst_dob_mux_b15/B0_40 ),
    .i1(\inst_dob_mux_b15/B0_41 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b15/B1_20 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_1_21  (
    .i0(\inst_dob_mux_b15/B0_42 ),
    .i1(\inst_dob_mux_b15/B0_43 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b15/B1_21 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_1_22  (
    .i0(\inst_dob_mux_b15/B0_44 ),
    .i1(\inst_dob_mux_b15/B0_45 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b15/B1_22 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_1_23  (
    .i0(\inst_dob_mux_b15/B0_46 ),
    .i1(\inst_dob_mux_b15/B0_47 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b15/B1_23 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_1_24  (
    .i0(\inst_dob_mux_b15/B0_48 ),
    .i1(\inst_dob_mux_b15/B0_49 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b15/B1_24 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_1_25  (
    .i0(\inst_dob_mux_b15/B0_50 ),
    .i1(\inst_dob_mux_b15/B0_51 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b15/B1_25 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_1_26  (
    .i0(\inst_dob_mux_b15/B0_52 ),
    .i1(\inst_dob_mux_b15/B0_53 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b15/B1_26 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_1_27  (
    .i0(\inst_dob_mux_b15/B0_54 ),
    .i1(\inst_dob_mux_b15/B0_55 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b15/B1_27 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_1_28  (
    .i0(\inst_dob_mux_b15/B0_56 ),
    .i1(\inst_dob_mux_b15/B0_57 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b15/B1_28 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_1_29  (
    .i0(\inst_dob_mux_b15/B0_58 ),
    .i1(\inst_dob_mux_b15/B0_59 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b15/B1_29 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_1_3  (
    .i0(\inst_dob_mux_b15/B0_6 ),
    .i1(\inst_dob_mux_b15/B0_7 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b15/B1_3 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_1_30  (
    .i0(\inst_dob_mux_b15/B0_60 ),
    .i1(\inst_dob_mux_b15/B0_61 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b15/B1_30 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_1_31  (
    .i0(\inst_dob_mux_b15/B0_62 ),
    .i1(\inst_dob_mux_b15/B0_63 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b15/B1_31 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_1_4  (
    .i0(\inst_dob_mux_b15/B0_8 ),
    .i1(\inst_dob_mux_b15/B0_9 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b15/B1_4 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_1_5  (
    .i0(\inst_dob_mux_b15/B0_10 ),
    .i1(\inst_dob_mux_b15/B0_11 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b15/B1_5 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_1_6  (
    .i0(\inst_dob_mux_b15/B0_12 ),
    .i1(\inst_dob_mux_b15/B0_13 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b15/B1_6 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_1_7  (
    .i0(\inst_dob_mux_b15/B0_14 ),
    .i1(\inst_dob_mux_b15/B0_15 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b15/B1_7 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_1_8  (
    .i0(\inst_dob_mux_b15/B0_16 ),
    .i1(\inst_dob_mux_b15/B0_17 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b15/B1_8 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_1_9  (
    .i0(\inst_dob_mux_b15/B0_18 ),
    .i1(\inst_dob_mux_b15/B0_19 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b15/B1_9 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_2_0  (
    .i0(\inst_dob_mux_b15/B1_0 ),
    .i1(\inst_dob_mux_b15/B1_1 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b15/B2_0 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_2_1  (
    .i0(\inst_dob_mux_b15/B1_2 ),
    .i1(\inst_dob_mux_b15/B1_3 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b15/B2_1 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_2_10  (
    .i0(\inst_dob_mux_b15/B1_20 ),
    .i1(\inst_dob_mux_b15/B1_21 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b15/B2_10 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_2_11  (
    .i0(\inst_dob_mux_b15/B1_22 ),
    .i1(\inst_dob_mux_b15/B1_23 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b15/B2_11 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_2_12  (
    .i0(\inst_dob_mux_b15/B1_24 ),
    .i1(\inst_dob_mux_b15/B1_25 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b15/B2_12 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_2_13  (
    .i0(\inst_dob_mux_b15/B1_26 ),
    .i1(\inst_dob_mux_b15/B1_27 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b15/B2_13 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_2_14  (
    .i0(\inst_dob_mux_b15/B1_28 ),
    .i1(\inst_dob_mux_b15/B1_29 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b15/B2_14 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_2_15  (
    .i0(\inst_dob_mux_b15/B1_30 ),
    .i1(\inst_dob_mux_b15/B1_31 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b15/B2_15 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_2_2  (
    .i0(\inst_dob_mux_b15/B1_4 ),
    .i1(\inst_dob_mux_b15/B1_5 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b15/B2_2 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_2_3  (
    .i0(\inst_dob_mux_b15/B1_6 ),
    .i1(\inst_dob_mux_b15/B1_7 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b15/B2_3 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_2_4  (
    .i0(\inst_dob_mux_b15/B1_8 ),
    .i1(\inst_dob_mux_b15/B1_9 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b15/B2_4 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_2_5  (
    .i0(\inst_dob_mux_b15/B1_10 ),
    .i1(\inst_dob_mux_b15/B1_11 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b15/B2_5 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_2_6  (
    .i0(\inst_dob_mux_b15/B1_12 ),
    .i1(\inst_dob_mux_b15/B1_13 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b15/B2_6 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_2_7  (
    .i0(\inst_dob_mux_b15/B1_14 ),
    .i1(\inst_dob_mux_b15/B1_15 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b15/B2_7 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_2_8  (
    .i0(\inst_dob_mux_b15/B1_16 ),
    .i1(\inst_dob_mux_b15/B1_17 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b15/B2_8 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_2_9  (
    .i0(\inst_dob_mux_b15/B1_18 ),
    .i1(\inst_dob_mux_b15/B1_19 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b15/B2_9 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_3_0  (
    .i0(\inst_dob_mux_b15/B2_0 ),
    .i1(\inst_dob_mux_b15/B2_1 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b15/B3_0 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_3_1  (
    .i0(\inst_dob_mux_b15/B2_2 ),
    .i1(\inst_dob_mux_b15/B2_3 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b15/B3_1 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_3_2  (
    .i0(\inst_dob_mux_b15/B2_4 ),
    .i1(\inst_dob_mux_b15/B2_5 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b15/B3_2 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_3_3  (
    .i0(\inst_dob_mux_b15/B2_6 ),
    .i1(\inst_dob_mux_b15/B2_7 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b15/B3_3 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_3_4  (
    .i0(\inst_dob_mux_b15/B2_8 ),
    .i1(\inst_dob_mux_b15/B2_9 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b15/B3_4 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_3_5  (
    .i0(\inst_dob_mux_b15/B2_10 ),
    .i1(\inst_dob_mux_b15/B2_11 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b15/B3_5 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_3_6  (
    .i0(\inst_dob_mux_b15/B2_12 ),
    .i1(\inst_dob_mux_b15/B2_13 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b15/B3_6 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_3_7  (
    .i0(\inst_dob_mux_b15/B2_14 ),
    .i1(\inst_dob_mux_b15/B2_15 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b15/B3_7 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_4_0  (
    .i0(\inst_dob_mux_b15/B3_0 ),
    .i1(\inst_dob_mux_b15/B3_1 ),
    .sel(addrb_piped_piped[4]),
    .o(\inst_dob_mux_b15/B4_0 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_4_1  (
    .i0(\inst_dob_mux_b15/B3_2 ),
    .i1(\inst_dob_mux_b15/B3_3 ),
    .sel(addrb_piped_piped[4]),
    .o(\inst_dob_mux_b15/B4_1 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_4_2  (
    .i0(\inst_dob_mux_b15/B3_4 ),
    .i1(\inst_dob_mux_b15/B3_5 ),
    .sel(addrb_piped_piped[4]),
    .o(\inst_dob_mux_b15/B4_2 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_4_3  (
    .i0(\inst_dob_mux_b15/B3_6 ),
    .i1(\inst_dob_mux_b15/B3_7 ),
    .sel(addrb_piped_piped[4]),
    .o(\inst_dob_mux_b15/B4_3 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_5_0  (
    .i0(\inst_dob_mux_b15/B4_0 ),
    .i1(\inst_dob_mux_b15/B4_1 ),
    .sel(addrb_piped_piped[5]),
    .o(\inst_dob_mux_b15/B5_0 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_5_1  (
    .i0(\inst_dob_mux_b15/B4_2 ),
    .i1(\inst_dob_mux_b15/B4_3 ),
    .sel(addrb_piped_piped[5]),
    .o(\inst_dob_mux_b15/B5_1 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_6_0  (
    .i0(\inst_dob_mux_b15/B5_0 ),
    .i1(\inst_dob_mux_b15/B5_1 ),
    .sel(addrb_piped_piped[6]),
    .o(dob[15]));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_0  (
    .i0(inst_dob_i0_002),
    .i1(inst_dob_i0_002),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b2/B0_0 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_1  (
    .i0(inst_dob_i2_002),
    .i1(inst_dob_i2_002),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b2/B0_1 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_10  (
    .i0(inst_dob_i20_002),
    .i1(inst_dob_i20_002),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b2/B0_10 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_11  (
    .i0(inst_dob_i22_002),
    .i1(inst_dob_i22_002),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b2/B0_11 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_12  (
    .i0(inst_dob_i24_002),
    .i1(inst_dob_i24_002),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b2/B0_12 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_13  (
    .i0(inst_dob_i26_002),
    .i1(inst_dob_i26_002),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b2/B0_13 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_14  (
    .i0(inst_dob_i28_002),
    .i1(inst_dob_i28_002),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b2/B0_14 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_15  (
    .i0(inst_dob_i30_002),
    .i1(inst_dob_i30_002),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b2/B0_15 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_16  (
    .i0(inst_dob_i32_002),
    .i1(inst_dob_i32_002),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b2/B0_16 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_17  (
    .i0(inst_dob_i34_002),
    .i1(inst_dob_i34_002),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b2/B0_17 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_18  (
    .i0(inst_dob_i36_002),
    .i1(inst_dob_i36_002),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b2/B0_18 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_19  (
    .i0(inst_dob_i38_002),
    .i1(inst_dob_i38_002),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b2/B0_19 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_2  (
    .i0(inst_dob_i4_002),
    .i1(inst_dob_i4_002),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b2/B0_2 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_20  (
    .i0(inst_dob_i40_002),
    .i1(inst_dob_i40_002),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b2/B0_20 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_21  (
    .i0(inst_dob_i42_002),
    .i1(inst_dob_i42_002),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b2/B0_21 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_22  (
    .i0(inst_dob_i44_002),
    .i1(inst_dob_i44_002),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b2/B0_22 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_23  (
    .i0(inst_dob_i46_002),
    .i1(inst_dob_i46_002),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b2/B0_23 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_24  (
    .i0(inst_dob_i48_002),
    .i1(inst_dob_i48_002),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b2/B0_24 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_25  (
    .i0(inst_dob_i50_002),
    .i1(inst_dob_i50_002),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b2/B0_25 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_26  (
    .i0(inst_dob_i52_002),
    .i1(inst_dob_i52_002),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b2/B0_26 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_27  (
    .i0(inst_dob_i54_002),
    .i1(inst_dob_i54_002),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b2/B0_27 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_28  (
    .i0(inst_dob_i56_002),
    .i1(inst_dob_i56_002),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b2/B0_28 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_29  (
    .i0(inst_dob_i58_002),
    .i1(inst_dob_i58_002),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b2/B0_29 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_3  (
    .i0(inst_dob_i6_002),
    .i1(inst_dob_i6_002),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b2/B0_3 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_30  (
    .i0(inst_dob_i60_002),
    .i1(inst_dob_i60_002),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b2/B0_30 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_31  (
    .i0(inst_dob_i62_002),
    .i1(inst_dob_i62_002),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b2/B0_31 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_32  (
    .i0(inst_dob_i64_002),
    .i1(inst_dob_i64_002),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b2/B0_32 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_33  (
    .i0(inst_dob_i64_002),
    .i1(inst_dob_i64_002),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b2/B0_33 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_34  (
    .i0(inst_dob_i64_002),
    .i1(inst_dob_i64_002),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b2/B0_34 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_35  (
    .i0(inst_dob_i64_002),
    .i1(inst_dob_i64_002),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b2/B0_35 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_36  (
    .i0(inst_dob_i64_002),
    .i1(inst_dob_i64_002),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b2/B0_36 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_37  (
    .i0(inst_dob_i64_002),
    .i1(inst_dob_i64_002),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b2/B0_37 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_38  (
    .i0(inst_dob_i64_002),
    .i1(inst_dob_i64_002),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b2/B0_38 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_39  (
    .i0(inst_dob_i64_002),
    .i1(inst_dob_i64_002),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b2/B0_39 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_4  (
    .i0(inst_dob_i8_002),
    .i1(inst_dob_i8_002),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b2/B0_4 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_40  (
    .i0(inst_dob_i64_002),
    .i1(inst_dob_i64_002),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b2/B0_40 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_41  (
    .i0(inst_dob_i64_002),
    .i1(inst_dob_i64_002),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b2/B0_41 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_42  (
    .i0(inst_dob_i64_002),
    .i1(inst_dob_i64_002),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b2/B0_42 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_43  (
    .i0(inst_dob_i64_002),
    .i1(inst_dob_i64_002),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b2/B0_43 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_44  (
    .i0(inst_dob_i64_002),
    .i1(inst_dob_i64_002),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b2/B0_44 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_45  (
    .i0(inst_dob_i64_002),
    .i1(inst_dob_i64_002),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b2/B0_45 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_46  (
    .i0(inst_dob_i64_002),
    .i1(inst_dob_i64_002),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b2/B0_46 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_47  (
    .i0(inst_dob_i64_002),
    .i1(inst_dob_i64_002),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b2/B0_47 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_48  (
    .i0(inst_dob_i64_002),
    .i1(inst_dob_i64_002),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b2/B0_48 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_49  (
    .i0(inst_dob_i64_002),
    .i1(inst_dob_i64_002),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b2/B0_49 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_5  (
    .i0(inst_dob_i10_002),
    .i1(inst_dob_i10_002),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b2/B0_5 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_50  (
    .i0(inst_dob_i64_002),
    .i1(inst_dob_i64_002),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b2/B0_50 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_51  (
    .i0(inst_dob_i64_002),
    .i1(inst_dob_i64_002),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b2/B0_51 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_52  (
    .i0(inst_dob_i64_002),
    .i1(inst_dob_i64_002),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b2/B0_52 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_53  (
    .i0(inst_dob_i64_002),
    .i1(inst_dob_i64_002),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b2/B0_53 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_54  (
    .i0(inst_dob_i64_002),
    .i1(inst_dob_i64_002),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b2/B0_54 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_55  (
    .i0(inst_dob_i64_002),
    .i1(inst_dob_i64_002),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b2/B0_55 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_56  (
    .i0(inst_dob_i64_002),
    .i1(inst_dob_i64_002),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b2/B0_56 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_57  (
    .i0(inst_dob_i64_002),
    .i1(inst_dob_i64_002),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b2/B0_57 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_58  (
    .i0(inst_dob_i64_002),
    .i1(inst_dob_i64_002),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b2/B0_58 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_59  (
    .i0(inst_dob_i64_002),
    .i1(inst_dob_i64_002),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b2/B0_59 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_6  (
    .i0(inst_dob_i12_002),
    .i1(inst_dob_i12_002),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b2/B0_6 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_60  (
    .i0(inst_dob_i64_002),
    .i1(inst_dob_i64_002),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b2/B0_60 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_61  (
    .i0(inst_dob_i64_002),
    .i1(inst_dob_i64_002),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b2/B0_61 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_62  (
    .i0(inst_dob_i64_002),
    .i1(inst_dob_i64_002),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b2/B0_62 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_63  (
    .i0(inst_dob_i64_002),
    .i1(inst_dob_i64_002),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b2/B0_63 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_7  (
    .i0(inst_dob_i14_002),
    .i1(inst_dob_i14_002),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b2/B0_7 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_8  (
    .i0(inst_dob_i16_002),
    .i1(inst_dob_i16_002),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b2/B0_8 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_9  (
    .i0(inst_dob_i18_002),
    .i1(inst_dob_i18_002),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b2/B0_9 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_1_0  (
    .i0(\inst_dob_mux_b2/B0_0 ),
    .i1(\inst_dob_mux_b2/B0_1 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b2/B1_0 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_1_1  (
    .i0(\inst_dob_mux_b2/B0_2 ),
    .i1(\inst_dob_mux_b2/B0_3 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b2/B1_1 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_1_10  (
    .i0(\inst_dob_mux_b2/B0_20 ),
    .i1(\inst_dob_mux_b2/B0_21 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b2/B1_10 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_1_11  (
    .i0(\inst_dob_mux_b2/B0_22 ),
    .i1(\inst_dob_mux_b2/B0_23 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b2/B1_11 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_1_12  (
    .i0(\inst_dob_mux_b2/B0_24 ),
    .i1(\inst_dob_mux_b2/B0_25 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b2/B1_12 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_1_13  (
    .i0(\inst_dob_mux_b2/B0_26 ),
    .i1(\inst_dob_mux_b2/B0_27 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b2/B1_13 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_1_14  (
    .i0(\inst_dob_mux_b2/B0_28 ),
    .i1(\inst_dob_mux_b2/B0_29 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b2/B1_14 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_1_15  (
    .i0(\inst_dob_mux_b2/B0_30 ),
    .i1(\inst_dob_mux_b2/B0_31 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b2/B1_15 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_1_16  (
    .i0(\inst_dob_mux_b2/B0_32 ),
    .i1(\inst_dob_mux_b2/B0_33 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b2/B1_16 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_1_17  (
    .i0(\inst_dob_mux_b2/B0_34 ),
    .i1(\inst_dob_mux_b2/B0_35 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b2/B1_17 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_1_18  (
    .i0(\inst_dob_mux_b2/B0_36 ),
    .i1(\inst_dob_mux_b2/B0_37 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b2/B1_18 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_1_19  (
    .i0(\inst_dob_mux_b2/B0_38 ),
    .i1(\inst_dob_mux_b2/B0_39 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b2/B1_19 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_1_2  (
    .i0(\inst_dob_mux_b2/B0_4 ),
    .i1(\inst_dob_mux_b2/B0_5 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b2/B1_2 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_1_20  (
    .i0(\inst_dob_mux_b2/B0_40 ),
    .i1(\inst_dob_mux_b2/B0_41 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b2/B1_20 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_1_21  (
    .i0(\inst_dob_mux_b2/B0_42 ),
    .i1(\inst_dob_mux_b2/B0_43 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b2/B1_21 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_1_22  (
    .i0(\inst_dob_mux_b2/B0_44 ),
    .i1(\inst_dob_mux_b2/B0_45 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b2/B1_22 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_1_23  (
    .i0(\inst_dob_mux_b2/B0_46 ),
    .i1(\inst_dob_mux_b2/B0_47 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b2/B1_23 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_1_24  (
    .i0(\inst_dob_mux_b2/B0_48 ),
    .i1(\inst_dob_mux_b2/B0_49 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b2/B1_24 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_1_25  (
    .i0(\inst_dob_mux_b2/B0_50 ),
    .i1(\inst_dob_mux_b2/B0_51 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b2/B1_25 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_1_26  (
    .i0(\inst_dob_mux_b2/B0_52 ),
    .i1(\inst_dob_mux_b2/B0_53 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b2/B1_26 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_1_27  (
    .i0(\inst_dob_mux_b2/B0_54 ),
    .i1(\inst_dob_mux_b2/B0_55 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b2/B1_27 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_1_28  (
    .i0(\inst_dob_mux_b2/B0_56 ),
    .i1(\inst_dob_mux_b2/B0_57 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b2/B1_28 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_1_29  (
    .i0(\inst_dob_mux_b2/B0_58 ),
    .i1(\inst_dob_mux_b2/B0_59 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b2/B1_29 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_1_3  (
    .i0(\inst_dob_mux_b2/B0_6 ),
    .i1(\inst_dob_mux_b2/B0_7 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b2/B1_3 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_1_30  (
    .i0(\inst_dob_mux_b2/B0_60 ),
    .i1(\inst_dob_mux_b2/B0_61 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b2/B1_30 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_1_31  (
    .i0(\inst_dob_mux_b2/B0_62 ),
    .i1(\inst_dob_mux_b2/B0_63 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b2/B1_31 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_1_4  (
    .i0(\inst_dob_mux_b2/B0_8 ),
    .i1(\inst_dob_mux_b2/B0_9 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b2/B1_4 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_1_5  (
    .i0(\inst_dob_mux_b2/B0_10 ),
    .i1(\inst_dob_mux_b2/B0_11 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b2/B1_5 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_1_6  (
    .i0(\inst_dob_mux_b2/B0_12 ),
    .i1(\inst_dob_mux_b2/B0_13 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b2/B1_6 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_1_7  (
    .i0(\inst_dob_mux_b2/B0_14 ),
    .i1(\inst_dob_mux_b2/B0_15 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b2/B1_7 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_1_8  (
    .i0(\inst_dob_mux_b2/B0_16 ),
    .i1(\inst_dob_mux_b2/B0_17 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b2/B1_8 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_1_9  (
    .i0(\inst_dob_mux_b2/B0_18 ),
    .i1(\inst_dob_mux_b2/B0_19 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b2/B1_9 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_2_0  (
    .i0(\inst_dob_mux_b2/B1_0 ),
    .i1(\inst_dob_mux_b2/B1_1 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b2/B2_0 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_2_1  (
    .i0(\inst_dob_mux_b2/B1_2 ),
    .i1(\inst_dob_mux_b2/B1_3 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b2/B2_1 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_2_10  (
    .i0(\inst_dob_mux_b2/B1_20 ),
    .i1(\inst_dob_mux_b2/B1_21 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b2/B2_10 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_2_11  (
    .i0(\inst_dob_mux_b2/B1_22 ),
    .i1(\inst_dob_mux_b2/B1_23 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b2/B2_11 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_2_12  (
    .i0(\inst_dob_mux_b2/B1_24 ),
    .i1(\inst_dob_mux_b2/B1_25 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b2/B2_12 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_2_13  (
    .i0(\inst_dob_mux_b2/B1_26 ),
    .i1(\inst_dob_mux_b2/B1_27 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b2/B2_13 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_2_14  (
    .i0(\inst_dob_mux_b2/B1_28 ),
    .i1(\inst_dob_mux_b2/B1_29 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b2/B2_14 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_2_15  (
    .i0(\inst_dob_mux_b2/B1_30 ),
    .i1(\inst_dob_mux_b2/B1_31 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b2/B2_15 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_2_2  (
    .i0(\inst_dob_mux_b2/B1_4 ),
    .i1(\inst_dob_mux_b2/B1_5 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b2/B2_2 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_2_3  (
    .i0(\inst_dob_mux_b2/B1_6 ),
    .i1(\inst_dob_mux_b2/B1_7 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b2/B2_3 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_2_4  (
    .i0(\inst_dob_mux_b2/B1_8 ),
    .i1(\inst_dob_mux_b2/B1_9 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b2/B2_4 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_2_5  (
    .i0(\inst_dob_mux_b2/B1_10 ),
    .i1(\inst_dob_mux_b2/B1_11 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b2/B2_5 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_2_6  (
    .i0(\inst_dob_mux_b2/B1_12 ),
    .i1(\inst_dob_mux_b2/B1_13 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b2/B2_6 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_2_7  (
    .i0(\inst_dob_mux_b2/B1_14 ),
    .i1(\inst_dob_mux_b2/B1_15 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b2/B2_7 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_2_8  (
    .i0(\inst_dob_mux_b2/B1_16 ),
    .i1(\inst_dob_mux_b2/B1_17 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b2/B2_8 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_2_9  (
    .i0(\inst_dob_mux_b2/B1_18 ),
    .i1(\inst_dob_mux_b2/B1_19 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b2/B2_9 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_3_0  (
    .i0(\inst_dob_mux_b2/B2_0 ),
    .i1(\inst_dob_mux_b2/B2_1 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b2/B3_0 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_3_1  (
    .i0(\inst_dob_mux_b2/B2_2 ),
    .i1(\inst_dob_mux_b2/B2_3 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b2/B3_1 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_3_2  (
    .i0(\inst_dob_mux_b2/B2_4 ),
    .i1(\inst_dob_mux_b2/B2_5 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b2/B3_2 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_3_3  (
    .i0(\inst_dob_mux_b2/B2_6 ),
    .i1(\inst_dob_mux_b2/B2_7 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b2/B3_3 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_3_4  (
    .i0(\inst_dob_mux_b2/B2_8 ),
    .i1(\inst_dob_mux_b2/B2_9 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b2/B3_4 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_3_5  (
    .i0(\inst_dob_mux_b2/B2_10 ),
    .i1(\inst_dob_mux_b2/B2_11 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b2/B3_5 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_3_6  (
    .i0(\inst_dob_mux_b2/B2_12 ),
    .i1(\inst_dob_mux_b2/B2_13 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b2/B3_6 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_3_7  (
    .i0(\inst_dob_mux_b2/B2_14 ),
    .i1(\inst_dob_mux_b2/B2_15 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b2/B3_7 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_4_0  (
    .i0(\inst_dob_mux_b2/B3_0 ),
    .i1(\inst_dob_mux_b2/B3_1 ),
    .sel(addrb_piped_piped[4]),
    .o(\inst_dob_mux_b2/B4_0 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_4_1  (
    .i0(\inst_dob_mux_b2/B3_2 ),
    .i1(\inst_dob_mux_b2/B3_3 ),
    .sel(addrb_piped_piped[4]),
    .o(\inst_dob_mux_b2/B4_1 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_4_2  (
    .i0(\inst_dob_mux_b2/B3_4 ),
    .i1(\inst_dob_mux_b2/B3_5 ),
    .sel(addrb_piped_piped[4]),
    .o(\inst_dob_mux_b2/B4_2 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_4_3  (
    .i0(\inst_dob_mux_b2/B3_6 ),
    .i1(\inst_dob_mux_b2/B3_7 ),
    .sel(addrb_piped_piped[4]),
    .o(\inst_dob_mux_b2/B4_3 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_5_0  (
    .i0(\inst_dob_mux_b2/B4_0 ),
    .i1(\inst_dob_mux_b2/B4_1 ),
    .sel(addrb_piped_piped[5]),
    .o(\inst_dob_mux_b2/B5_0 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_5_1  (
    .i0(\inst_dob_mux_b2/B4_2 ),
    .i1(\inst_dob_mux_b2/B4_3 ),
    .sel(addrb_piped_piped[5]),
    .o(\inst_dob_mux_b2/B5_1 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_6_0  (
    .i0(\inst_dob_mux_b2/B5_0 ),
    .i1(\inst_dob_mux_b2/B5_1 ),
    .sel(addrb_piped_piped[6]),
    .o(dob[2]));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_0  (
    .i0(inst_dob_i0_003),
    .i1(inst_dob_i0_003),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b3/B0_0 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_1  (
    .i0(inst_dob_i2_003),
    .i1(inst_dob_i2_003),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b3/B0_1 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_10  (
    .i0(inst_dob_i20_003),
    .i1(inst_dob_i20_003),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b3/B0_10 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_11  (
    .i0(inst_dob_i22_003),
    .i1(inst_dob_i22_003),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b3/B0_11 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_12  (
    .i0(inst_dob_i24_003),
    .i1(inst_dob_i24_003),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b3/B0_12 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_13  (
    .i0(inst_dob_i26_003),
    .i1(inst_dob_i26_003),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b3/B0_13 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_14  (
    .i0(inst_dob_i28_003),
    .i1(inst_dob_i28_003),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b3/B0_14 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_15  (
    .i0(inst_dob_i30_003),
    .i1(inst_dob_i30_003),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b3/B0_15 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_16  (
    .i0(inst_dob_i32_003),
    .i1(inst_dob_i32_003),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b3/B0_16 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_17  (
    .i0(inst_dob_i34_003),
    .i1(inst_dob_i34_003),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b3/B0_17 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_18  (
    .i0(inst_dob_i36_003),
    .i1(inst_dob_i36_003),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b3/B0_18 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_19  (
    .i0(inst_dob_i38_003),
    .i1(inst_dob_i38_003),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b3/B0_19 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_2  (
    .i0(inst_dob_i4_003),
    .i1(inst_dob_i4_003),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b3/B0_2 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_20  (
    .i0(inst_dob_i40_003),
    .i1(inst_dob_i40_003),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b3/B0_20 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_21  (
    .i0(inst_dob_i42_003),
    .i1(inst_dob_i42_003),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b3/B0_21 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_22  (
    .i0(inst_dob_i44_003),
    .i1(inst_dob_i44_003),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b3/B0_22 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_23  (
    .i0(inst_dob_i46_003),
    .i1(inst_dob_i46_003),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b3/B0_23 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_24  (
    .i0(inst_dob_i48_003),
    .i1(inst_dob_i48_003),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b3/B0_24 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_25  (
    .i0(inst_dob_i50_003),
    .i1(inst_dob_i50_003),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b3/B0_25 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_26  (
    .i0(inst_dob_i52_003),
    .i1(inst_dob_i52_003),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b3/B0_26 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_27  (
    .i0(inst_dob_i54_003),
    .i1(inst_dob_i54_003),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b3/B0_27 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_28  (
    .i0(inst_dob_i56_003),
    .i1(inst_dob_i56_003),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b3/B0_28 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_29  (
    .i0(inst_dob_i58_003),
    .i1(inst_dob_i58_003),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b3/B0_29 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_3  (
    .i0(inst_dob_i6_003),
    .i1(inst_dob_i6_003),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b3/B0_3 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_30  (
    .i0(inst_dob_i60_003),
    .i1(inst_dob_i60_003),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b3/B0_30 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_31  (
    .i0(inst_dob_i62_003),
    .i1(inst_dob_i62_003),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b3/B0_31 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_32  (
    .i0(inst_dob_i64_003),
    .i1(inst_dob_i64_003),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b3/B0_32 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_33  (
    .i0(inst_dob_i64_003),
    .i1(inst_dob_i64_003),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b3/B0_33 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_34  (
    .i0(inst_dob_i64_003),
    .i1(inst_dob_i64_003),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b3/B0_34 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_35  (
    .i0(inst_dob_i64_003),
    .i1(inst_dob_i64_003),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b3/B0_35 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_36  (
    .i0(inst_dob_i64_003),
    .i1(inst_dob_i64_003),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b3/B0_36 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_37  (
    .i0(inst_dob_i64_003),
    .i1(inst_dob_i64_003),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b3/B0_37 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_38  (
    .i0(inst_dob_i64_003),
    .i1(inst_dob_i64_003),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b3/B0_38 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_39  (
    .i0(inst_dob_i64_003),
    .i1(inst_dob_i64_003),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b3/B0_39 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_4  (
    .i0(inst_dob_i8_003),
    .i1(inst_dob_i8_003),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b3/B0_4 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_40  (
    .i0(inst_dob_i64_003),
    .i1(inst_dob_i64_003),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b3/B0_40 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_41  (
    .i0(inst_dob_i64_003),
    .i1(inst_dob_i64_003),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b3/B0_41 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_42  (
    .i0(inst_dob_i64_003),
    .i1(inst_dob_i64_003),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b3/B0_42 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_43  (
    .i0(inst_dob_i64_003),
    .i1(inst_dob_i64_003),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b3/B0_43 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_44  (
    .i0(inst_dob_i64_003),
    .i1(inst_dob_i64_003),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b3/B0_44 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_45  (
    .i0(inst_dob_i64_003),
    .i1(inst_dob_i64_003),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b3/B0_45 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_46  (
    .i0(inst_dob_i64_003),
    .i1(inst_dob_i64_003),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b3/B0_46 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_47  (
    .i0(inst_dob_i64_003),
    .i1(inst_dob_i64_003),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b3/B0_47 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_48  (
    .i0(inst_dob_i64_003),
    .i1(inst_dob_i64_003),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b3/B0_48 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_49  (
    .i0(inst_dob_i64_003),
    .i1(inst_dob_i64_003),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b3/B0_49 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_5  (
    .i0(inst_dob_i10_003),
    .i1(inst_dob_i10_003),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b3/B0_5 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_50  (
    .i0(inst_dob_i64_003),
    .i1(inst_dob_i64_003),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b3/B0_50 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_51  (
    .i0(inst_dob_i64_003),
    .i1(inst_dob_i64_003),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b3/B0_51 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_52  (
    .i0(inst_dob_i64_003),
    .i1(inst_dob_i64_003),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b3/B0_52 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_53  (
    .i0(inst_dob_i64_003),
    .i1(inst_dob_i64_003),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b3/B0_53 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_54  (
    .i0(inst_dob_i64_003),
    .i1(inst_dob_i64_003),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b3/B0_54 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_55  (
    .i0(inst_dob_i64_003),
    .i1(inst_dob_i64_003),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b3/B0_55 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_56  (
    .i0(inst_dob_i64_003),
    .i1(inst_dob_i64_003),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b3/B0_56 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_57  (
    .i0(inst_dob_i64_003),
    .i1(inst_dob_i64_003),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b3/B0_57 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_58  (
    .i0(inst_dob_i64_003),
    .i1(inst_dob_i64_003),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b3/B0_58 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_59  (
    .i0(inst_dob_i64_003),
    .i1(inst_dob_i64_003),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b3/B0_59 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_6  (
    .i0(inst_dob_i12_003),
    .i1(inst_dob_i12_003),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b3/B0_6 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_60  (
    .i0(inst_dob_i64_003),
    .i1(inst_dob_i64_003),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b3/B0_60 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_61  (
    .i0(inst_dob_i64_003),
    .i1(inst_dob_i64_003),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b3/B0_61 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_62  (
    .i0(inst_dob_i64_003),
    .i1(inst_dob_i64_003),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b3/B0_62 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_63  (
    .i0(inst_dob_i64_003),
    .i1(inst_dob_i64_003),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b3/B0_63 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_7  (
    .i0(inst_dob_i14_003),
    .i1(inst_dob_i14_003),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b3/B0_7 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_8  (
    .i0(inst_dob_i16_003),
    .i1(inst_dob_i16_003),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b3/B0_8 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_9  (
    .i0(inst_dob_i18_003),
    .i1(inst_dob_i18_003),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b3/B0_9 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_1_0  (
    .i0(\inst_dob_mux_b3/B0_0 ),
    .i1(\inst_dob_mux_b3/B0_1 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b3/B1_0 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_1_1  (
    .i0(\inst_dob_mux_b3/B0_2 ),
    .i1(\inst_dob_mux_b3/B0_3 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b3/B1_1 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_1_10  (
    .i0(\inst_dob_mux_b3/B0_20 ),
    .i1(\inst_dob_mux_b3/B0_21 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b3/B1_10 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_1_11  (
    .i0(\inst_dob_mux_b3/B0_22 ),
    .i1(\inst_dob_mux_b3/B0_23 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b3/B1_11 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_1_12  (
    .i0(\inst_dob_mux_b3/B0_24 ),
    .i1(\inst_dob_mux_b3/B0_25 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b3/B1_12 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_1_13  (
    .i0(\inst_dob_mux_b3/B0_26 ),
    .i1(\inst_dob_mux_b3/B0_27 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b3/B1_13 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_1_14  (
    .i0(\inst_dob_mux_b3/B0_28 ),
    .i1(\inst_dob_mux_b3/B0_29 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b3/B1_14 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_1_15  (
    .i0(\inst_dob_mux_b3/B0_30 ),
    .i1(\inst_dob_mux_b3/B0_31 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b3/B1_15 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_1_16  (
    .i0(\inst_dob_mux_b3/B0_32 ),
    .i1(\inst_dob_mux_b3/B0_33 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b3/B1_16 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_1_17  (
    .i0(\inst_dob_mux_b3/B0_34 ),
    .i1(\inst_dob_mux_b3/B0_35 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b3/B1_17 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_1_18  (
    .i0(\inst_dob_mux_b3/B0_36 ),
    .i1(\inst_dob_mux_b3/B0_37 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b3/B1_18 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_1_19  (
    .i0(\inst_dob_mux_b3/B0_38 ),
    .i1(\inst_dob_mux_b3/B0_39 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b3/B1_19 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_1_2  (
    .i0(\inst_dob_mux_b3/B0_4 ),
    .i1(\inst_dob_mux_b3/B0_5 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b3/B1_2 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_1_20  (
    .i0(\inst_dob_mux_b3/B0_40 ),
    .i1(\inst_dob_mux_b3/B0_41 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b3/B1_20 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_1_21  (
    .i0(\inst_dob_mux_b3/B0_42 ),
    .i1(\inst_dob_mux_b3/B0_43 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b3/B1_21 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_1_22  (
    .i0(\inst_dob_mux_b3/B0_44 ),
    .i1(\inst_dob_mux_b3/B0_45 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b3/B1_22 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_1_23  (
    .i0(\inst_dob_mux_b3/B0_46 ),
    .i1(\inst_dob_mux_b3/B0_47 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b3/B1_23 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_1_24  (
    .i0(\inst_dob_mux_b3/B0_48 ),
    .i1(\inst_dob_mux_b3/B0_49 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b3/B1_24 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_1_25  (
    .i0(\inst_dob_mux_b3/B0_50 ),
    .i1(\inst_dob_mux_b3/B0_51 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b3/B1_25 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_1_26  (
    .i0(\inst_dob_mux_b3/B0_52 ),
    .i1(\inst_dob_mux_b3/B0_53 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b3/B1_26 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_1_27  (
    .i0(\inst_dob_mux_b3/B0_54 ),
    .i1(\inst_dob_mux_b3/B0_55 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b3/B1_27 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_1_28  (
    .i0(\inst_dob_mux_b3/B0_56 ),
    .i1(\inst_dob_mux_b3/B0_57 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b3/B1_28 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_1_29  (
    .i0(\inst_dob_mux_b3/B0_58 ),
    .i1(\inst_dob_mux_b3/B0_59 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b3/B1_29 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_1_3  (
    .i0(\inst_dob_mux_b3/B0_6 ),
    .i1(\inst_dob_mux_b3/B0_7 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b3/B1_3 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_1_30  (
    .i0(\inst_dob_mux_b3/B0_60 ),
    .i1(\inst_dob_mux_b3/B0_61 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b3/B1_30 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_1_31  (
    .i0(\inst_dob_mux_b3/B0_62 ),
    .i1(\inst_dob_mux_b3/B0_63 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b3/B1_31 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_1_4  (
    .i0(\inst_dob_mux_b3/B0_8 ),
    .i1(\inst_dob_mux_b3/B0_9 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b3/B1_4 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_1_5  (
    .i0(\inst_dob_mux_b3/B0_10 ),
    .i1(\inst_dob_mux_b3/B0_11 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b3/B1_5 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_1_6  (
    .i0(\inst_dob_mux_b3/B0_12 ),
    .i1(\inst_dob_mux_b3/B0_13 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b3/B1_6 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_1_7  (
    .i0(\inst_dob_mux_b3/B0_14 ),
    .i1(\inst_dob_mux_b3/B0_15 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b3/B1_7 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_1_8  (
    .i0(\inst_dob_mux_b3/B0_16 ),
    .i1(\inst_dob_mux_b3/B0_17 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b3/B1_8 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_1_9  (
    .i0(\inst_dob_mux_b3/B0_18 ),
    .i1(\inst_dob_mux_b3/B0_19 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b3/B1_9 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_2_0  (
    .i0(\inst_dob_mux_b3/B1_0 ),
    .i1(\inst_dob_mux_b3/B1_1 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b3/B2_0 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_2_1  (
    .i0(\inst_dob_mux_b3/B1_2 ),
    .i1(\inst_dob_mux_b3/B1_3 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b3/B2_1 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_2_10  (
    .i0(\inst_dob_mux_b3/B1_20 ),
    .i1(\inst_dob_mux_b3/B1_21 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b3/B2_10 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_2_11  (
    .i0(\inst_dob_mux_b3/B1_22 ),
    .i1(\inst_dob_mux_b3/B1_23 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b3/B2_11 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_2_12  (
    .i0(\inst_dob_mux_b3/B1_24 ),
    .i1(\inst_dob_mux_b3/B1_25 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b3/B2_12 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_2_13  (
    .i0(\inst_dob_mux_b3/B1_26 ),
    .i1(\inst_dob_mux_b3/B1_27 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b3/B2_13 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_2_14  (
    .i0(\inst_dob_mux_b3/B1_28 ),
    .i1(\inst_dob_mux_b3/B1_29 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b3/B2_14 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_2_15  (
    .i0(\inst_dob_mux_b3/B1_30 ),
    .i1(\inst_dob_mux_b3/B1_31 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b3/B2_15 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_2_2  (
    .i0(\inst_dob_mux_b3/B1_4 ),
    .i1(\inst_dob_mux_b3/B1_5 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b3/B2_2 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_2_3  (
    .i0(\inst_dob_mux_b3/B1_6 ),
    .i1(\inst_dob_mux_b3/B1_7 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b3/B2_3 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_2_4  (
    .i0(\inst_dob_mux_b3/B1_8 ),
    .i1(\inst_dob_mux_b3/B1_9 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b3/B2_4 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_2_5  (
    .i0(\inst_dob_mux_b3/B1_10 ),
    .i1(\inst_dob_mux_b3/B1_11 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b3/B2_5 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_2_6  (
    .i0(\inst_dob_mux_b3/B1_12 ),
    .i1(\inst_dob_mux_b3/B1_13 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b3/B2_6 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_2_7  (
    .i0(\inst_dob_mux_b3/B1_14 ),
    .i1(\inst_dob_mux_b3/B1_15 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b3/B2_7 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_2_8  (
    .i0(\inst_dob_mux_b3/B1_16 ),
    .i1(\inst_dob_mux_b3/B1_17 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b3/B2_8 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_2_9  (
    .i0(\inst_dob_mux_b3/B1_18 ),
    .i1(\inst_dob_mux_b3/B1_19 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b3/B2_9 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_3_0  (
    .i0(\inst_dob_mux_b3/B2_0 ),
    .i1(\inst_dob_mux_b3/B2_1 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b3/B3_0 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_3_1  (
    .i0(\inst_dob_mux_b3/B2_2 ),
    .i1(\inst_dob_mux_b3/B2_3 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b3/B3_1 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_3_2  (
    .i0(\inst_dob_mux_b3/B2_4 ),
    .i1(\inst_dob_mux_b3/B2_5 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b3/B3_2 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_3_3  (
    .i0(\inst_dob_mux_b3/B2_6 ),
    .i1(\inst_dob_mux_b3/B2_7 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b3/B3_3 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_3_4  (
    .i0(\inst_dob_mux_b3/B2_8 ),
    .i1(\inst_dob_mux_b3/B2_9 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b3/B3_4 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_3_5  (
    .i0(\inst_dob_mux_b3/B2_10 ),
    .i1(\inst_dob_mux_b3/B2_11 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b3/B3_5 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_3_6  (
    .i0(\inst_dob_mux_b3/B2_12 ),
    .i1(\inst_dob_mux_b3/B2_13 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b3/B3_6 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_3_7  (
    .i0(\inst_dob_mux_b3/B2_14 ),
    .i1(\inst_dob_mux_b3/B2_15 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b3/B3_7 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_4_0  (
    .i0(\inst_dob_mux_b3/B3_0 ),
    .i1(\inst_dob_mux_b3/B3_1 ),
    .sel(addrb_piped_piped[4]),
    .o(\inst_dob_mux_b3/B4_0 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_4_1  (
    .i0(\inst_dob_mux_b3/B3_2 ),
    .i1(\inst_dob_mux_b3/B3_3 ),
    .sel(addrb_piped_piped[4]),
    .o(\inst_dob_mux_b3/B4_1 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_4_2  (
    .i0(\inst_dob_mux_b3/B3_4 ),
    .i1(\inst_dob_mux_b3/B3_5 ),
    .sel(addrb_piped_piped[4]),
    .o(\inst_dob_mux_b3/B4_2 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_4_3  (
    .i0(\inst_dob_mux_b3/B3_6 ),
    .i1(\inst_dob_mux_b3/B3_7 ),
    .sel(addrb_piped_piped[4]),
    .o(\inst_dob_mux_b3/B4_3 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_5_0  (
    .i0(\inst_dob_mux_b3/B4_0 ),
    .i1(\inst_dob_mux_b3/B4_1 ),
    .sel(addrb_piped_piped[5]),
    .o(\inst_dob_mux_b3/B5_0 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_5_1  (
    .i0(\inst_dob_mux_b3/B4_2 ),
    .i1(\inst_dob_mux_b3/B4_3 ),
    .sel(addrb_piped_piped[5]),
    .o(\inst_dob_mux_b3/B5_1 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_6_0  (
    .i0(\inst_dob_mux_b3/B5_0 ),
    .i1(\inst_dob_mux_b3/B5_1 ),
    .sel(addrb_piped_piped[6]),
    .o(dob[3]));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_0  (
    .i0(inst_dob_i0_004),
    .i1(inst_dob_i0_004),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b4/B0_0 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_1  (
    .i0(inst_dob_i2_004),
    .i1(inst_dob_i2_004),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b4/B0_1 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_10  (
    .i0(inst_dob_i20_004),
    .i1(inst_dob_i20_004),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b4/B0_10 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_11  (
    .i0(inst_dob_i22_004),
    .i1(inst_dob_i22_004),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b4/B0_11 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_12  (
    .i0(inst_dob_i24_004),
    .i1(inst_dob_i24_004),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b4/B0_12 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_13  (
    .i0(inst_dob_i26_004),
    .i1(inst_dob_i26_004),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b4/B0_13 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_14  (
    .i0(inst_dob_i28_004),
    .i1(inst_dob_i28_004),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b4/B0_14 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_15  (
    .i0(inst_dob_i30_004),
    .i1(inst_dob_i30_004),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b4/B0_15 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_16  (
    .i0(inst_dob_i32_004),
    .i1(inst_dob_i32_004),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b4/B0_16 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_17  (
    .i0(inst_dob_i34_004),
    .i1(inst_dob_i34_004),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b4/B0_17 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_18  (
    .i0(inst_dob_i36_004),
    .i1(inst_dob_i36_004),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b4/B0_18 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_19  (
    .i0(inst_dob_i38_004),
    .i1(inst_dob_i38_004),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b4/B0_19 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_2  (
    .i0(inst_dob_i4_004),
    .i1(inst_dob_i4_004),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b4/B0_2 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_20  (
    .i0(inst_dob_i40_004),
    .i1(inst_dob_i40_004),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b4/B0_20 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_21  (
    .i0(inst_dob_i42_004),
    .i1(inst_dob_i42_004),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b4/B0_21 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_22  (
    .i0(inst_dob_i44_004),
    .i1(inst_dob_i44_004),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b4/B0_22 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_23  (
    .i0(inst_dob_i46_004),
    .i1(inst_dob_i46_004),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b4/B0_23 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_24  (
    .i0(inst_dob_i48_004),
    .i1(inst_dob_i48_004),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b4/B0_24 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_25  (
    .i0(inst_dob_i50_004),
    .i1(inst_dob_i50_004),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b4/B0_25 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_26  (
    .i0(inst_dob_i52_004),
    .i1(inst_dob_i52_004),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b4/B0_26 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_27  (
    .i0(inst_dob_i54_004),
    .i1(inst_dob_i54_004),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b4/B0_27 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_28  (
    .i0(inst_dob_i56_004),
    .i1(inst_dob_i56_004),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b4/B0_28 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_29  (
    .i0(inst_dob_i58_004),
    .i1(inst_dob_i58_004),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b4/B0_29 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_3  (
    .i0(inst_dob_i6_004),
    .i1(inst_dob_i6_004),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b4/B0_3 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_30  (
    .i0(inst_dob_i60_004),
    .i1(inst_dob_i60_004),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b4/B0_30 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_31  (
    .i0(inst_dob_i62_004),
    .i1(inst_dob_i62_004),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b4/B0_31 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_32  (
    .i0(inst_dob_i64_004),
    .i1(inst_dob_i64_004),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b4/B0_32 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_33  (
    .i0(inst_dob_i64_004),
    .i1(inst_dob_i64_004),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b4/B0_33 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_34  (
    .i0(inst_dob_i64_004),
    .i1(inst_dob_i64_004),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b4/B0_34 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_35  (
    .i0(inst_dob_i64_004),
    .i1(inst_dob_i64_004),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b4/B0_35 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_36  (
    .i0(inst_dob_i64_004),
    .i1(inst_dob_i64_004),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b4/B0_36 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_37  (
    .i0(inst_dob_i64_004),
    .i1(inst_dob_i64_004),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b4/B0_37 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_38  (
    .i0(inst_dob_i64_004),
    .i1(inst_dob_i64_004),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b4/B0_38 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_39  (
    .i0(inst_dob_i64_004),
    .i1(inst_dob_i64_004),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b4/B0_39 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_4  (
    .i0(inst_dob_i8_004),
    .i1(inst_dob_i8_004),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b4/B0_4 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_40  (
    .i0(inst_dob_i64_004),
    .i1(inst_dob_i64_004),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b4/B0_40 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_41  (
    .i0(inst_dob_i64_004),
    .i1(inst_dob_i64_004),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b4/B0_41 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_42  (
    .i0(inst_dob_i64_004),
    .i1(inst_dob_i64_004),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b4/B0_42 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_43  (
    .i0(inst_dob_i64_004),
    .i1(inst_dob_i64_004),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b4/B0_43 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_44  (
    .i0(inst_dob_i64_004),
    .i1(inst_dob_i64_004),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b4/B0_44 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_45  (
    .i0(inst_dob_i64_004),
    .i1(inst_dob_i64_004),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b4/B0_45 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_46  (
    .i0(inst_dob_i64_004),
    .i1(inst_dob_i64_004),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b4/B0_46 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_47  (
    .i0(inst_dob_i64_004),
    .i1(inst_dob_i64_004),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b4/B0_47 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_48  (
    .i0(inst_dob_i64_004),
    .i1(inst_dob_i64_004),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b4/B0_48 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_49  (
    .i0(inst_dob_i64_004),
    .i1(inst_dob_i64_004),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b4/B0_49 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_5  (
    .i0(inst_dob_i10_004),
    .i1(inst_dob_i10_004),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b4/B0_5 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_50  (
    .i0(inst_dob_i64_004),
    .i1(inst_dob_i64_004),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b4/B0_50 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_51  (
    .i0(inst_dob_i64_004),
    .i1(inst_dob_i64_004),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b4/B0_51 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_52  (
    .i0(inst_dob_i64_004),
    .i1(inst_dob_i64_004),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b4/B0_52 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_53  (
    .i0(inst_dob_i64_004),
    .i1(inst_dob_i64_004),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b4/B0_53 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_54  (
    .i0(inst_dob_i64_004),
    .i1(inst_dob_i64_004),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b4/B0_54 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_55  (
    .i0(inst_dob_i64_004),
    .i1(inst_dob_i64_004),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b4/B0_55 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_56  (
    .i0(inst_dob_i64_004),
    .i1(inst_dob_i64_004),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b4/B0_56 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_57  (
    .i0(inst_dob_i64_004),
    .i1(inst_dob_i64_004),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b4/B0_57 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_58  (
    .i0(inst_dob_i64_004),
    .i1(inst_dob_i64_004),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b4/B0_58 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_59  (
    .i0(inst_dob_i64_004),
    .i1(inst_dob_i64_004),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b4/B0_59 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_6  (
    .i0(inst_dob_i12_004),
    .i1(inst_dob_i12_004),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b4/B0_6 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_60  (
    .i0(inst_dob_i64_004),
    .i1(inst_dob_i64_004),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b4/B0_60 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_61  (
    .i0(inst_dob_i64_004),
    .i1(inst_dob_i64_004),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b4/B0_61 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_62  (
    .i0(inst_dob_i64_004),
    .i1(inst_dob_i64_004),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b4/B0_62 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_63  (
    .i0(inst_dob_i64_004),
    .i1(inst_dob_i64_004),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b4/B0_63 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_7  (
    .i0(inst_dob_i14_004),
    .i1(inst_dob_i14_004),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b4/B0_7 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_8  (
    .i0(inst_dob_i16_004),
    .i1(inst_dob_i16_004),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b4/B0_8 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_9  (
    .i0(inst_dob_i18_004),
    .i1(inst_dob_i18_004),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b4/B0_9 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_1_0  (
    .i0(\inst_dob_mux_b4/B0_0 ),
    .i1(\inst_dob_mux_b4/B0_1 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b4/B1_0 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_1_1  (
    .i0(\inst_dob_mux_b4/B0_2 ),
    .i1(\inst_dob_mux_b4/B0_3 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b4/B1_1 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_1_10  (
    .i0(\inst_dob_mux_b4/B0_20 ),
    .i1(\inst_dob_mux_b4/B0_21 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b4/B1_10 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_1_11  (
    .i0(\inst_dob_mux_b4/B0_22 ),
    .i1(\inst_dob_mux_b4/B0_23 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b4/B1_11 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_1_12  (
    .i0(\inst_dob_mux_b4/B0_24 ),
    .i1(\inst_dob_mux_b4/B0_25 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b4/B1_12 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_1_13  (
    .i0(\inst_dob_mux_b4/B0_26 ),
    .i1(\inst_dob_mux_b4/B0_27 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b4/B1_13 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_1_14  (
    .i0(\inst_dob_mux_b4/B0_28 ),
    .i1(\inst_dob_mux_b4/B0_29 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b4/B1_14 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_1_15  (
    .i0(\inst_dob_mux_b4/B0_30 ),
    .i1(\inst_dob_mux_b4/B0_31 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b4/B1_15 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_1_16  (
    .i0(\inst_dob_mux_b4/B0_32 ),
    .i1(\inst_dob_mux_b4/B0_33 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b4/B1_16 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_1_17  (
    .i0(\inst_dob_mux_b4/B0_34 ),
    .i1(\inst_dob_mux_b4/B0_35 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b4/B1_17 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_1_18  (
    .i0(\inst_dob_mux_b4/B0_36 ),
    .i1(\inst_dob_mux_b4/B0_37 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b4/B1_18 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_1_19  (
    .i0(\inst_dob_mux_b4/B0_38 ),
    .i1(\inst_dob_mux_b4/B0_39 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b4/B1_19 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_1_2  (
    .i0(\inst_dob_mux_b4/B0_4 ),
    .i1(\inst_dob_mux_b4/B0_5 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b4/B1_2 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_1_20  (
    .i0(\inst_dob_mux_b4/B0_40 ),
    .i1(\inst_dob_mux_b4/B0_41 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b4/B1_20 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_1_21  (
    .i0(\inst_dob_mux_b4/B0_42 ),
    .i1(\inst_dob_mux_b4/B0_43 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b4/B1_21 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_1_22  (
    .i0(\inst_dob_mux_b4/B0_44 ),
    .i1(\inst_dob_mux_b4/B0_45 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b4/B1_22 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_1_23  (
    .i0(\inst_dob_mux_b4/B0_46 ),
    .i1(\inst_dob_mux_b4/B0_47 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b4/B1_23 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_1_24  (
    .i0(\inst_dob_mux_b4/B0_48 ),
    .i1(\inst_dob_mux_b4/B0_49 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b4/B1_24 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_1_25  (
    .i0(\inst_dob_mux_b4/B0_50 ),
    .i1(\inst_dob_mux_b4/B0_51 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b4/B1_25 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_1_26  (
    .i0(\inst_dob_mux_b4/B0_52 ),
    .i1(\inst_dob_mux_b4/B0_53 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b4/B1_26 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_1_27  (
    .i0(\inst_dob_mux_b4/B0_54 ),
    .i1(\inst_dob_mux_b4/B0_55 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b4/B1_27 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_1_28  (
    .i0(\inst_dob_mux_b4/B0_56 ),
    .i1(\inst_dob_mux_b4/B0_57 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b4/B1_28 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_1_29  (
    .i0(\inst_dob_mux_b4/B0_58 ),
    .i1(\inst_dob_mux_b4/B0_59 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b4/B1_29 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_1_3  (
    .i0(\inst_dob_mux_b4/B0_6 ),
    .i1(\inst_dob_mux_b4/B0_7 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b4/B1_3 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_1_30  (
    .i0(\inst_dob_mux_b4/B0_60 ),
    .i1(\inst_dob_mux_b4/B0_61 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b4/B1_30 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_1_31  (
    .i0(\inst_dob_mux_b4/B0_62 ),
    .i1(\inst_dob_mux_b4/B0_63 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b4/B1_31 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_1_4  (
    .i0(\inst_dob_mux_b4/B0_8 ),
    .i1(\inst_dob_mux_b4/B0_9 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b4/B1_4 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_1_5  (
    .i0(\inst_dob_mux_b4/B0_10 ),
    .i1(\inst_dob_mux_b4/B0_11 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b4/B1_5 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_1_6  (
    .i0(\inst_dob_mux_b4/B0_12 ),
    .i1(\inst_dob_mux_b4/B0_13 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b4/B1_6 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_1_7  (
    .i0(\inst_dob_mux_b4/B0_14 ),
    .i1(\inst_dob_mux_b4/B0_15 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b4/B1_7 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_1_8  (
    .i0(\inst_dob_mux_b4/B0_16 ),
    .i1(\inst_dob_mux_b4/B0_17 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b4/B1_8 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_1_9  (
    .i0(\inst_dob_mux_b4/B0_18 ),
    .i1(\inst_dob_mux_b4/B0_19 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b4/B1_9 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_2_0  (
    .i0(\inst_dob_mux_b4/B1_0 ),
    .i1(\inst_dob_mux_b4/B1_1 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b4/B2_0 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_2_1  (
    .i0(\inst_dob_mux_b4/B1_2 ),
    .i1(\inst_dob_mux_b4/B1_3 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b4/B2_1 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_2_10  (
    .i0(\inst_dob_mux_b4/B1_20 ),
    .i1(\inst_dob_mux_b4/B1_21 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b4/B2_10 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_2_11  (
    .i0(\inst_dob_mux_b4/B1_22 ),
    .i1(\inst_dob_mux_b4/B1_23 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b4/B2_11 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_2_12  (
    .i0(\inst_dob_mux_b4/B1_24 ),
    .i1(\inst_dob_mux_b4/B1_25 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b4/B2_12 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_2_13  (
    .i0(\inst_dob_mux_b4/B1_26 ),
    .i1(\inst_dob_mux_b4/B1_27 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b4/B2_13 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_2_14  (
    .i0(\inst_dob_mux_b4/B1_28 ),
    .i1(\inst_dob_mux_b4/B1_29 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b4/B2_14 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_2_15  (
    .i0(\inst_dob_mux_b4/B1_30 ),
    .i1(\inst_dob_mux_b4/B1_31 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b4/B2_15 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_2_2  (
    .i0(\inst_dob_mux_b4/B1_4 ),
    .i1(\inst_dob_mux_b4/B1_5 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b4/B2_2 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_2_3  (
    .i0(\inst_dob_mux_b4/B1_6 ),
    .i1(\inst_dob_mux_b4/B1_7 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b4/B2_3 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_2_4  (
    .i0(\inst_dob_mux_b4/B1_8 ),
    .i1(\inst_dob_mux_b4/B1_9 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b4/B2_4 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_2_5  (
    .i0(\inst_dob_mux_b4/B1_10 ),
    .i1(\inst_dob_mux_b4/B1_11 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b4/B2_5 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_2_6  (
    .i0(\inst_dob_mux_b4/B1_12 ),
    .i1(\inst_dob_mux_b4/B1_13 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b4/B2_6 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_2_7  (
    .i0(\inst_dob_mux_b4/B1_14 ),
    .i1(\inst_dob_mux_b4/B1_15 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b4/B2_7 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_2_8  (
    .i0(\inst_dob_mux_b4/B1_16 ),
    .i1(\inst_dob_mux_b4/B1_17 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b4/B2_8 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_2_9  (
    .i0(\inst_dob_mux_b4/B1_18 ),
    .i1(\inst_dob_mux_b4/B1_19 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b4/B2_9 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_3_0  (
    .i0(\inst_dob_mux_b4/B2_0 ),
    .i1(\inst_dob_mux_b4/B2_1 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b4/B3_0 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_3_1  (
    .i0(\inst_dob_mux_b4/B2_2 ),
    .i1(\inst_dob_mux_b4/B2_3 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b4/B3_1 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_3_2  (
    .i0(\inst_dob_mux_b4/B2_4 ),
    .i1(\inst_dob_mux_b4/B2_5 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b4/B3_2 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_3_3  (
    .i0(\inst_dob_mux_b4/B2_6 ),
    .i1(\inst_dob_mux_b4/B2_7 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b4/B3_3 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_3_4  (
    .i0(\inst_dob_mux_b4/B2_8 ),
    .i1(\inst_dob_mux_b4/B2_9 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b4/B3_4 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_3_5  (
    .i0(\inst_dob_mux_b4/B2_10 ),
    .i1(\inst_dob_mux_b4/B2_11 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b4/B3_5 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_3_6  (
    .i0(\inst_dob_mux_b4/B2_12 ),
    .i1(\inst_dob_mux_b4/B2_13 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b4/B3_6 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_3_7  (
    .i0(\inst_dob_mux_b4/B2_14 ),
    .i1(\inst_dob_mux_b4/B2_15 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b4/B3_7 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_4_0  (
    .i0(\inst_dob_mux_b4/B3_0 ),
    .i1(\inst_dob_mux_b4/B3_1 ),
    .sel(addrb_piped_piped[4]),
    .o(\inst_dob_mux_b4/B4_0 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_4_1  (
    .i0(\inst_dob_mux_b4/B3_2 ),
    .i1(\inst_dob_mux_b4/B3_3 ),
    .sel(addrb_piped_piped[4]),
    .o(\inst_dob_mux_b4/B4_1 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_4_2  (
    .i0(\inst_dob_mux_b4/B3_4 ),
    .i1(\inst_dob_mux_b4/B3_5 ),
    .sel(addrb_piped_piped[4]),
    .o(\inst_dob_mux_b4/B4_2 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_4_3  (
    .i0(\inst_dob_mux_b4/B3_6 ),
    .i1(\inst_dob_mux_b4/B3_7 ),
    .sel(addrb_piped_piped[4]),
    .o(\inst_dob_mux_b4/B4_3 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_5_0  (
    .i0(\inst_dob_mux_b4/B4_0 ),
    .i1(\inst_dob_mux_b4/B4_1 ),
    .sel(addrb_piped_piped[5]),
    .o(\inst_dob_mux_b4/B5_0 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_5_1  (
    .i0(\inst_dob_mux_b4/B4_2 ),
    .i1(\inst_dob_mux_b4/B4_3 ),
    .sel(addrb_piped_piped[5]),
    .o(\inst_dob_mux_b4/B5_1 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_6_0  (
    .i0(\inst_dob_mux_b4/B5_0 ),
    .i1(\inst_dob_mux_b4/B5_1 ),
    .sel(addrb_piped_piped[6]),
    .o(dob[4]));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_0  (
    .i0(inst_dob_i0_005),
    .i1(inst_dob_i0_005),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b5/B0_0 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_1  (
    .i0(inst_dob_i2_005),
    .i1(inst_dob_i2_005),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b5/B0_1 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_10  (
    .i0(inst_dob_i20_005),
    .i1(inst_dob_i20_005),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b5/B0_10 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_11  (
    .i0(inst_dob_i22_005),
    .i1(inst_dob_i22_005),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b5/B0_11 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_12  (
    .i0(inst_dob_i24_005),
    .i1(inst_dob_i24_005),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b5/B0_12 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_13  (
    .i0(inst_dob_i26_005),
    .i1(inst_dob_i26_005),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b5/B0_13 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_14  (
    .i0(inst_dob_i28_005),
    .i1(inst_dob_i28_005),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b5/B0_14 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_15  (
    .i0(inst_dob_i30_005),
    .i1(inst_dob_i30_005),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b5/B0_15 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_16  (
    .i0(inst_dob_i32_005),
    .i1(inst_dob_i32_005),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b5/B0_16 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_17  (
    .i0(inst_dob_i34_005),
    .i1(inst_dob_i34_005),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b5/B0_17 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_18  (
    .i0(inst_dob_i36_005),
    .i1(inst_dob_i36_005),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b5/B0_18 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_19  (
    .i0(inst_dob_i38_005),
    .i1(inst_dob_i38_005),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b5/B0_19 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_2  (
    .i0(inst_dob_i4_005),
    .i1(inst_dob_i4_005),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b5/B0_2 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_20  (
    .i0(inst_dob_i40_005),
    .i1(inst_dob_i40_005),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b5/B0_20 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_21  (
    .i0(inst_dob_i42_005),
    .i1(inst_dob_i42_005),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b5/B0_21 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_22  (
    .i0(inst_dob_i44_005),
    .i1(inst_dob_i44_005),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b5/B0_22 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_23  (
    .i0(inst_dob_i46_005),
    .i1(inst_dob_i46_005),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b5/B0_23 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_24  (
    .i0(inst_dob_i48_005),
    .i1(inst_dob_i48_005),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b5/B0_24 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_25  (
    .i0(inst_dob_i50_005),
    .i1(inst_dob_i50_005),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b5/B0_25 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_26  (
    .i0(inst_dob_i52_005),
    .i1(inst_dob_i52_005),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b5/B0_26 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_27  (
    .i0(inst_dob_i54_005),
    .i1(inst_dob_i54_005),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b5/B0_27 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_28  (
    .i0(inst_dob_i56_005),
    .i1(inst_dob_i56_005),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b5/B0_28 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_29  (
    .i0(inst_dob_i58_005),
    .i1(inst_dob_i58_005),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b5/B0_29 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_3  (
    .i0(inst_dob_i6_005),
    .i1(inst_dob_i6_005),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b5/B0_3 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_30  (
    .i0(inst_dob_i60_005),
    .i1(inst_dob_i60_005),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b5/B0_30 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_31  (
    .i0(inst_dob_i62_005),
    .i1(inst_dob_i62_005),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b5/B0_31 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_32  (
    .i0(inst_dob_i64_005),
    .i1(inst_dob_i64_005),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b5/B0_32 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_33  (
    .i0(inst_dob_i64_005),
    .i1(inst_dob_i64_005),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b5/B0_33 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_34  (
    .i0(inst_dob_i64_005),
    .i1(inst_dob_i64_005),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b5/B0_34 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_35  (
    .i0(inst_dob_i64_005),
    .i1(inst_dob_i64_005),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b5/B0_35 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_36  (
    .i0(inst_dob_i64_005),
    .i1(inst_dob_i64_005),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b5/B0_36 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_37  (
    .i0(inst_dob_i64_005),
    .i1(inst_dob_i64_005),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b5/B0_37 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_38  (
    .i0(inst_dob_i64_005),
    .i1(inst_dob_i64_005),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b5/B0_38 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_39  (
    .i0(inst_dob_i64_005),
    .i1(inst_dob_i64_005),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b5/B0_39 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_4  (
    .i0(inst_dob_i8_005),
    .i1(inst_dob_i8_005),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b5/B0_4 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_40  (
    .i0(inst_dob_i64_005),
    .i1(inst_dob_i64_005),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b5/B0_40 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_41  (
    .i0(inst_dob_i64_005),
    .i1(inst_dob_i64_005),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b5/B0_41 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_42  (
    .i0(inst_dob_i64_005),
    .i1(inst_dob_i64_005),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b5/B0_42 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_43  (
    .i0(inst_dob_i64_005),
    .i1(inst_dob_i64_005),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b5/B0_43 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_44  (
    .i0(inst_dob_i64_005),
    .i1(inst_dob_i64_005),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b5/B0_44 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_45  (
    .i0(inst_dob_i64_005),
    .i1(inst_dob_i64_005),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b5/B0_45 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_46  (
    .i0(inst_dob_i64_005),
    .i1(inst_dob_i64_005),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b5/B0_46 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_47  (
    .i0(inst_dob_i64_005),
    .i1(inst_dob_i64_005),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b5/B0_47 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_48  (
    .i0(inst_dob_i64_005),
    .i1(inst_dob_i64_005),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b5/B0_48 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_49  (
    .i0(inst_dob_i64_005),
    .i1(inst_dob_i64_005),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b5/B0_49 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_5  (
    .i0(inst_dob_i10_005),
    .i1(inst_dob_i10_005),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b5/B0_5 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_50  (
    .i0(inst_dob_i64_005),
    .i1(inst_dob_i64_005),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b5/B0_50 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_51  (
    .i0(inst_dob_i64_005),
    .i1(inst_dob_i64_005),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b5/B0_51 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_52  (
    .i0(inst_dob_i64_005),
    .i1(inst_dob_i64_005),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b5/B0_52 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_53  (
    .i0(inst_dob_i64_005),
    .i1(inst_dob_i64_005),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b5/B0_53 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_54  (
    .i0(inst_dob_i64_005),
    .i1(inst_dob_i64_005),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b5/B0_54 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_55  (
    .i0(inst_dob_i64_005),
    .i1(inst_dob_i64_005),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b5/B0_55 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_56  (
    .i0(inst_dob_i64_005),
    .i1(inst_dob_i64_005),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b5/B0_56 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_57  (
    .i0(inst_dob_i64_005),
    .i1(inst_dob_i64_005),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b5/B0_57 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_58  (
    .i0(inst_dob_i64_005),
    .i1(inst_dob_i64_005),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b5/B0_58 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_59  (
    .i0(inst_dob_i64_005),
    .i1(inst_dob_i64_005),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b5/B0_59 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_6  (
    .i0(inst_dob_i12_005),
    .i1(inst_dob_i12_005),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b5/B0_6 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_60  (
    .i0(inst_dob_i64_005),
    .i1(inst_dob_i64_005),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b5/B0_60 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_61  (
    .i0(inst_dob_i64_005),
    .i1(inst_dob_i64_005),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b5/B0_61 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_62  (
    .i0(inst_dob_i64_005),
    .i1(inst_dob_i64_005),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b5/B0_62 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_63  (
    .i0(inst_dob_i64_005),
    .i1(inst_dob_i64_005),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b5/B0_63 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_7  (
    .i0(inst_dob_i14_005),
    .i1(inst_dob_i14_005),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b5/B0_7 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_8  (
    .i0(inst_dob_i16_005),
    .i1(inst_dob_i16_005),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b5/B0_8 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_9  (
    .i0(inst_dob_i18_005),
    .i1(inst_dob_i18_005),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b5/B0_9 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_1_0  (
    .i0(\inst_dob_mux_b5/B0_0 ),
    .i1(\inst_dob_mux_b5/B0_1 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b5/B1_0 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_1_1  (
    .i0(\inst_dob_mux_b5/B0_2 ),
    .i1(\inst_dob_mux_b5/B0_3 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b5/B1_1 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_1_10  (
    .i0(\inst_dob_mux_b5/B0_20 ),
    .i1(\inst_dob_mux_b5/B0_21 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b5/B1_10 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_1_11  (
    .i0(\inst_dob_mux_b5/B0_22 ),
    .i1(\inst_dob_mux_b5/B0_23 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b5/B1_11 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_1_12  (
    .i0(\inst_dob_mux_b5/B0_24 ),
    .i1(\inst_dob_mux_b5/B0_25 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b5/B1_12 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_1_13  (
    .i0(\inst_dob_mux_b5/B0_26 ),
    .i1(\inst_dob_mux_b5/B0_27 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b5/B1_13 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_1_14  (
    .i0(\inst_dob_mux_b5/B0_28 ),
    .i1(\inst_dob_mux_b5/B0_29 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b5/B1_14 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_1_15  (
    .i0(\inst_dob_mux_b5/B0_30 ),
    .i1(\inst_dob_mux_b5/B0_31 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b5/B1_15 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_1_16  (
    .i0(\inst_dob_mux_b5/B0_32 ),
    .i1(\inst_dob_mux_b5/B0_33 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b5/B1_16 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_1_17  (
    .i0(\inst_dob_mux_b5/B0_34 ),
    .i1(\inst_dob_mux_b5/B0_35 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b5/B1_17 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_1_18  (
    .i0(\inst_dob_mux_b5/B0_36 ),
    .i1(\inst_dob_mux_b5/B0_37 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b5/B1_18 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_1_19  (
    .i0(\inst_dob_mux_b5/B0_38 ),
    .i1(\inst_dob_mux_b5/B0_39 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b5/B1_19 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_1_2  (
    .i0(\inst_dob_mux_b5/B0_4 ),
    .i1(\inst_dob_mux_b5/B0_5 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b5/B1_2 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_1_20  (
    .i0(\inst_dob_mux_b5/B0_40 ),
    .i1(\inst_dob_mux_b5/B0_41 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b5/B1_20 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_1_21  (
    .i0(\inst_dob_mux_b5/B0_42 ),
    .i1(\inst_dob_mux_b5/B0_43 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b5/B1_21 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_1_22  (
    .i0(\inst_dob_mux_b5/B0_44 ),
    .i1(\inst_dob_mux_b5/B0_45 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b5/B1_22 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_1_23  (
    .i0(\inst_dob_mux_b5/B0_46 ),
    .i1(\inst_dob_mux_b5/B0_47 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b5/B1_23 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_1_24  (
    .i0(\inst_dob_mux_b5/B0_48 ),
    .i1(\inst_dob_mux_b5/B0_49 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b5/B1_24 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_1_25  (
    .i0(\inst_dob_mux_b5/B0_50 ),
    .i1(\inst_dob_mux_b5/B0_51 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b5/B1_25 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_1_26  (
    .i0(\inst_dob_mux_b5/B0_52 ),
    .i1(\inst_dob_mux_b5/B0_53 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b5/B1_26 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_1_27  (
    .i0(\inst_dob_mux_b5/B0_54 ),
    .i1(\inst_dob_mux_b5/B0_55 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b5/B1_27 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_1_28  (
    .i0(\inst_dob_mux_b5/B0_56 ),
    .i1(\inst_dob_mux_b5/B0_57 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b5/B1_28 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_1_29  (
    .i0(\inst_dob_mux_b5/B0_58 ),
    .i1(\inst_dob_mux_b5/B0_59 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b5/B1_29 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_1_3  (
    .i0(\inst_dob_mux_b5/B0_6 ),
    .i1(\inst_dob_mux_b5/B0_7 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b5/B1_3 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_1_30  (
    .i0(\inst_dob_mux_b5/B0_60 ),
    .i1(\inst_dob_mux_b5/B0_61 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b5/B1_30 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_1_31  (
    .i0(\inst_dob_mux_b5/B0_62 ),
    .i1(\inst_dob_mux_b5/B0_63 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b5/B1_31 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_1_4  (
    .i0(\inst_dob_mux_b5/B0_8 ),
    .i1(\inst_dob_mux_b5/B0_9 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b5/B1_4 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_1_5  (
    .i0(\inst_dob_mux_b5/B0_10 ),
    .i1(\inst_dob_mux_b5/B0_11 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b5/B1_5 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_1_6  (
    .i0(\inst_dob_mux_b5/B0_12 ),
    .i1(\inst_dob_mux_b5/B0_13 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b5/B1_6 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_1_7  (
    .i0(\inst_dob_mux_b5/B0_14 ),
    .i1(\inst_dob_mux_b5/B0_15 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b5/B1_7 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_1_8  (
    .i0(\inst_dob_mux_b5/B0_16 ),
    .i1(\inst_dob_mux_b5/B0_17 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b5/B1_8 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_1_9  (
    .i0(\inst_dob_mux_b5/B0_18 ),
    .i1(\inst_dob_mux_b5/B0_19 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b5/B1_9 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_2_0  (
    .i0(\inst_dob_mux_b5/B1_0 ),
    .i1(\inst_dob_mux_b5/B1_1 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b5/B2_0 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_2_1  (
    .i0(\inst_dob_mux_b5/B1_2 ),
    .i1(\inst_dob_mux_b5/B1_3 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b5/B2_1 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_2_10  (
    .i0(\inst_dob_mux_b5/B1_20 ),
    .i1(\inst_dob_mux_b5/B1_21 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b5/B2_10 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_2_11  (
    .i0(\inst_dob_mux_b5/B1_22 ),
    .i1(\inst_dob_mux_b5/B1_23 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b5/B2_11 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_2_12  (
    .i0(\inst_dob_mux_b5/B1_24 ),
    .i1(\inst_dob_mux_b5/B1_25 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b5/B2_12 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_2_13  (
    .i0(\inst_dob_mux_b5/B1_26 ),
    .i1(\inst_dob_mux_b5/B1_27 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b5/B2_13 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_2_14  (
    .i0(\inst_dob_mux_b5/B1_28 ),
    .i1(\inst_dob_mux_b5/B1_29 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b5/B2_14 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_2_15  (
    .i0(\inst_dob_mux_b5/B1_30 ),
    .i1(\inst_dob_mux_b5/B1_31 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b5/B2_15 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_2_2  (
    .i0(\inst_dob_mux_b5/B1_4 ),
    .i1(\inst_dob_mux_b5/B1_5 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b5/B2_2 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_2_3  (
    .i0(\inst_dob_mux_b5/B1_6 ),
    .i1(\inst_dob_mux_b5/B1_7 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b5/B2_3 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_2_4  (
    .i0(\inst_dob_mux_b5/B1_8 ),
    .i1(\inst_dob_mux_b5/B1_9 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b5/B2_4 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_2_5  (
    .i0(\inst_dob_mux_b5/B1_10 ),
    .i1(\inst_dob_mux_b5/B1_11 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b5/B2_5 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_2_6  (
    .i0(\inst_dob_mux_b5/B1_12 ),
    .i1(\inst_dob_mux_b5/B1_13 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b5/B2_6 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_2_7  (
    .i0(\inst_dob_mux_b5/B1_14 ),
    .i1(\inst_dob_mux_b5/B1_15 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b5/B2_7 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_2_8  (
    .i0(\inst_dob_mux_b5/B1_16 ),
    .i1(\inst_dob_mux_b5/B1_17 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b5/B2_8 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_2_9  (
    .i0(\inst_dob_mux_b5/B1_18 ),
    .i1(\inst_dob_mux_b5/B1_19 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b5/B2_9 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_3_0  (
    .i0(\inst_dob_mux_b5/B2_0 ),
    .i1(\inst_dob_mux_b5/B2_1 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b5/B3_0 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_3_1  (
    .i0(\inst_dob_mux_b5/B2_2 ),
    .i1(\inst_dob_mux_b5/B2_3 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b5/B3_1 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_3_2  (
    .i0(\inst_dob_mux_b5/B2_4 ),
    .i1(\inst_dob_mux_b5/B2_5 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b5/B3_2 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_3_3  (
    .i0(\inst_dob_mux_b5/B2_6 ),
    .i1(\inst_dob_mux_b5/B2_7 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b5/B3_3 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_3_4  (
    .i0(\inst_dob_mux_b5/B2_8 ),
    .i1(\inst_dob_mux_b5/B2_9 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b5/B3_4 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_3_5  (
    .i0(\inst_dob_mux_b5/B2_10 ),
    .i1(\inst_dob_mux_b5/B2_11 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b5/B3_5 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_3_6  (
    .i0(\inst_dob_mux_b5/B2_12 ),
    .i1(\inst_dob_mux_b5/B2_13 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b5/B3_6 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_3_7  (
    .i0(\inst_dob_mux_b5/B2_14 ),
    .i1(\inst_dob_mux_b5/B2_15 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b5/B3_7 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_4_0  (
    .i0(\inst_dob_mux_b5/B3_0 ),
    .i1(\inst_dob_mux_b5/B3_1 ),
    .sel(addrb_piped_piped[4]),
    .o(\inst_dob_mux_b5/B4_0 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_4_1  (
    .i0(\inst_dob_mux_b5/B3_2 ),
    .i1(\inst_dob_mux_b5/B3_3 ),
    .sel(addrb_piped_piped[4]),
    .o(\inst_dob_mux_b5/B4_1 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_4_2  (
    .i0(\inst_dob_mux_b5/B3_4 ),
    .i1(\inst_dob_mux_b5/B3_5 ),
    .sel(addrb_piped_piped[4]),
    .o(\inst_dob_mux_b5/B4_2 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_4_3  (
    .i0(\inst_dob_mux_b5/B3_6 ),
    .i1(\inst_dob_mux_b5/B3_7 ),
    .sel(addrb_piped_piped[4]),
    .o(\inst_dob_mux_b5/B4_3 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_5_0  (
    .i0(\inst_dob_mux_b5/B4_0 ),
    .i1(\inst_dob_mux_b5/B4_1 ),
    .sel(addrb_piped_piped[5]),
    .o(\inst_dob_mux_b5/B5_0 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_5_1  (
    .i0(\inst_dob_mux_b5/B4_2 ),
    .i1(\inst_dob_mux_b5/B4_3 ),
    .sel(addrb_piped_piped[5]),
    .o(\inst_dob_mux_b5/B5_1 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_6_0  (
    .i0(\inst_dob_mux_b5/B5_0 ),
    .i1(\inst_dob_mux_b5/B5_1 ),
    .sel(addrb_piped_piped[6]),
    .o(dob[5]));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_0  (
    .i0(inst_dob_i0_006),
    .i1(inst_dob_i0_006),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b6/B0_0 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_1  (
    .i0(inst_dob_i2_006),
    .i1(inst_dob_i2_006),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b6/B0_1 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_10  (
    .i0(inst_dob_i20_006),
    .i1(inst_dob_i20_006),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b6/B0_10 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_11  (
    .i0(inst_dob_i22_006),
    .i1(inst_dob_i22_006),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b6/B0_11 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_12  (
    .i0(inst_dob_i24_006),
    .i1(inst_dob_i24_006),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b6/B0_12 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_13  (
    .i0(inst_dob_i26_006),
    .i1(inst_dob_i26_006),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b6/B0_13 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_14  (
    .i0(inst_dob_i28_006),
    .i1(inst_dob_i28_006),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b6/B0_14 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_15  (
    .i0(inst_dob_i30_006),
    .i1(inst_dob_i30_006),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b6/B0_15 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_16  (
    .i0(inst_dob_i32_006),
    .i1(inst_dob_i32_006),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b6/B0_16 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_17  (
    .i0(inst_dob_i34_006),
    .i1(inst_dob_i34_006),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b6/B0_17 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_18  (
    .i0(inst_dob_i36_006),
    .i1(inst_dob_i36_006),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b6/B0_18 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_19  (
    .i0(inst_dob_i38_006),
    .i1(inst_dob_i38_006),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b6/B0_19 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_2  (
    .i0(inst_dob_i4_006),
    .i1(inst_dob_i4_006),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b6/B0_2 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_20  (
    .i0(inst_dob_i40_006),
    .i1(inst_dob_i40_006),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b6/B0_20 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_21  (
    .i0(inst_dob_i42_006),
    .i1(inst_dob_i42_006),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b6/B0_21 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_22  (
    .i0(inst_dob_i44_006),
    .i1(inst_dob_i44_006),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b6/B0_22 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_23  (
    .i0(inst_dob_i46_006),
    .i1(inst_dob_i46_006),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b6/B0_23 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_24  (
    .i0(inst_dob_i48_006),
    .i1(inst_dob_i48_006),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b6/B0_24 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_25  (
    .i0(inst_dob_i50_006),
    .i1(inst_dob_i50_006),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b6/B0_25 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_26  (
    .i0(inst_dob_i52_006),
    .i1(inst_dob_i52_006),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b6/B0_26 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_27  (
    .i0(inst_dob_i54_006),
    .i1(inst_dob_i54_006),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b6/B0_27 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_28  (
    .i0(inst_dob_i56_006),
    .i1(inst_dob_i56_006),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b6/B0_28 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_29  (
    .i0(inst_dob_i58_006),
    .i1(inst_dob_i58_006),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b6/B0_29 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_3  (
    .i0(inst_dob_i6_006),
    .i1(inst_dob_i6_006),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b6/B0_3 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_30  (
    .i0(inst_dob_i60_006),
    .i1(inst_dob_i60_006),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b6/B0_30 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_31  (
    .i0(inst_dob_i62_006),
    .i1(inst_dob_i62_006),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b6/B0_31 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_32  (
    .i0(inst_dob_i64_006),
    .i1(inst_dob_i64_006),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b6/B0_32 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_33  (
    .i0(inst_dob_i64_006),
    .i1(inst_dob_i64_006),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b6/B0_33 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_34  (
    .i0(inst_dob_i64_006),
    .i1(inst_dob_i64_006),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b6/B0_34 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_35  (
    .i0(inst_dob_i64_006),
    .i1(inst_dob_i64_006),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b6/B0_35 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_36  (
    .i0(inst_dob_i64_006),
    .i1(inst_dob_i64_006),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b6/B0_36 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_37  (
    .i0(inst_dob_i64_006),
    .i1(inst_dob_i64_006),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b6/B0_37 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_38  (
    .i0(inst_dob_i64_006),
    .i1(inst_dob_i64_006),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b6/B0_38 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_39  (
    .i0(inst_dob_i64_006),
    .i1(inst_dob_i64_006),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b6/B0_39 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_4  (
    .i0(inst_dob_i8_006),
    .i1(inst_dob_i8_006),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b6/B0_4 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_40  (
    .i0(inst_dob_i64_006),
    .i1(inst_dob_i64_006),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b6/B0_40 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_41  (
    .i0(inst_dob_i64_006),
    .i1(inst_dob_i64_006),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b6/B0_41 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_42  (
    .i0(inst_dob_i64_006),
    .i1(inst_dob_i64_006),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b6/B0_42 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_43  (
    .i0(inst_dob_i64_006),
    .i1(inst_dob_i64_006),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b6/B0_43 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_44  (
    .i0(inst_dob_i64_006),
    .i1(inst_dob_i64_006),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b6/B0_44 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_45  (
    .i0(inst_dob_i64_006),
    .i1(inst_dob_i64_006),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b6/B0_45 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_46  (
    .i0(inst_dob_i64_006),
    .i1(inst_dob_i64_006),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b6/B0_46 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_47  (
    .i0(inst_dob_i64_006),
    .i1(inst_dob_i64_006),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b6/B0_47 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_48  (
    .i0(inst_dob_i64_006),
    .i1(inst_dob_i64_006),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b6/B0_48 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_49  (
    .i0(inst_dob_i64_006),
    .i1(inst_dob_i64_006),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b6/B0_49 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_5  (
    .i0(inst_dob_i10_006),
    .i1(inst_dob_i10_006),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b6/B0_5 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_50  (
    .i0(inst_dob_i64_006),
    .i1(inst_dob_i64_006),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b6/B0_50 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_51  (
    .i0(inst_dob_i64_006),
    .i1(inst_dob_i64_006),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b6/B0_51 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_52  (
    .i0(inst_dob_i64_006),
    .i1(inst_dob_i64_006),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b6/B0_52 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_53  (
    .i0(inst_dob_i64_006),
    .i1(inst_dob_i64_006),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b6/B0_53 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_54  (
    .i0(inst_dob_i64_006),
    .i1(inst_dob_i64_006),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b6/B0_54 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_55  (
    .i0(inst_dob_i64_006),
    .i1(inst_dob_i64_006),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b6/B0_55 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_56  (
    .i0(inst_dob_i64_006),
    .i1(inst_dob_i64_006),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b6/B0_56 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_57  (
    .i0(inst_dob_i64_006),
    .i1(inst_dob_i64_006),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b6/B0_57 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_58  (
    .i0(inst_dob_i64_006),
    .i1(inst_dob_i64_006),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b6/B0_58 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_59  (
    .i0(inst_dob_i64_006),
    .i1(inst_dob_i64_006),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b6/B0_59 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_6  (
    .i0(inst_dob_i12_006),
    .i1(inst_dob_i12_006),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b6/B0_6 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_60  (
    .i0(inst_dob_i64_006),
    .i1(inst_dob_i64_006),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b6/B0_60 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_61  (
    .i0(inst_dob_i64_006),
    .i1(inst_dob_i64_006),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b6/B0_61 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_62  (
    .i0(inst_dob_i64_006),
    .i1(inst_dob_i64_006),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b6/B0_62 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_63  (
    .i0(inst_dob_i64_006),
    .i1(inst_dob_i64_006),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b6/B0_63 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_7  (
    .i0(inst_dob_i14_006),
    .i1(inst_dob_i14_006),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b6/B0_7 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_8  (
    .i0(inst_dob_i16_006),
    .i1(inst_dob_i16_006),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b6/B0_8 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_9  (
    .i0(inst_dob_i18_006),
    .i1(inst_dob_i18_006),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b6/B0_9 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_1_0  (
    .i0(\inst_dob_mux_b6/B0_0 ),
    .i1(\inst_dob_mux_b6/B0_1 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b6/B1_0 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_1_1  (
    .i0(\inst_dob_mux_b6/B0_2 ),
    .i1(\inst_dob_mux_b6/B0_3 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b6/B1_1 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_1_10  (
    .i0(\inst_dob_mux_b6/B0_20 ),
    .i1(\inst_dob_mux_b6/B0_21 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b6/B1_10 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_1_11  (
    .i0(\inst_dob_mux_b6/B0_22 ),
    .i1(\inst_dob_mux_b6/B0_23 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b6/B1_11 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_1_12  (
    .i0(\inst_dob_mux_b6/B0_24 ),
    .i1(\inst_dob_mux_b6/B0_25 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b6/B1_12 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_1_13  (
    .i0(\inst_dob_mux_b6/B0_26 ),
    .i1(\inst_dob_mux_b6/B0_27 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b6/B1_13 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_1_14  (
    .i0(\inst_dob_mux_b6/B0_28 ),
    .i1(\inst_dob_mux_b6/B0_29 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b6/B1_14 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_1_15  (
    .i0(\inst_dob_mux_b6/B0_30 ),
    .i1(\inst_dob_mux_b6/B0_31 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b6/B1_15 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_1_16  (
    .i0(\inst_dob_mux_b6/B0_32 ),
    .i1(\inst_dob_mux_b6/B0_33 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b6/B1_16 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_1_17  (
    .i0(\inst_dob_mux_b6/B0_34 ),
    .i1(\inst_dob_mux_b6/B0_35 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b6/B1_17 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_1_18  (
    .i0(\inst_dob_mux_b6/B0_36 ),
    .i1(\inst_dob_mux_b6/B0_37 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b6/B1_18 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_1_19  (
    .i0(\inst_dob_mux_b6/B0_38 ),
    .i1(\inst_dob_mux_b6/B0_39 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b6/B1_19 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_1_2  (
    .i0(\inst_dob_mux_b6/B0_4 ),
    .i1(\inst_dob_mux_b6/B0_5 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b6/B1_2 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_1_20  (
    .i0(\inst_dob_mux_b6/B0_40 ),
    .i1(\inst_dob_mux_b6/B0_41 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b6/B1_20 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_1_21  (
    .i0(\inst_dob_mux_b6/B0_42 ),
    .i1(\inst_dob_mux_b6/B0_43 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b6/B1_21 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_1_22  (
    .i0(\inst_dob_mux_b6/B0_44 ),
    .i1(\inst_dob_mux_b6/B0_45 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b6/B1_22 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_1_23  (
    .i0(\inst_dob_mux_b6/B0_46 ),
    .i1(\inst_dob_mux_b6/B0_47 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b6/B1_23 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_1_24  (
    .i0(\inst_dob_mux_b6/B0_48 ),
    .i1(\inst_dob_mux_b6/B0_49 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b6/B1_24 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_1_25  (
    .i0(\inst_dob_mux_b6/B0_50 ),
    .i1(\inst_dob_mux_b6/B0_51 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b6/B1_25 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_1_26  (
    .i0(\inst_dob_mux_b6/B0_52 ),
    .i1(\inst_dob_mux_b6/B0_53 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b6/B1_26 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_1_27  (
    .i0(\inst_dob_mux_b6/B0_54 ),
    .i1(\inst_dob_mux_b6/B0_55 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b6/B1_27 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_1_28  (
    .i0(\inst_dob_mux_b6/B0_56 ),
    .i1(\inst_dob_mux_b6/B0_57 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b6/B1_28 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_1_29  (
    .i0(\inst_dob_mux_b6/B0_58 ),
    .i1(\inst_dob_mux_b6/B0_59 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b6/B1_29 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_1_3  (
    .i0(\inst_dob_mux_b6/B0_6 ),
    .i1(\inst_dob_mux_b6/B0_7 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b6/B1_3 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_1_30  (
    .i0(\inst_dob_mux_b6/B0_60 ),
    .i1(\inst_dob_mux_b6/B0_61 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b6/B1_30 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_1_31  (
    .i0(\inst_dob_mux_b6/B0_62 ),
    .i1(\inst_dob_mux_b6/B0_63 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b6/B1_31 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_1_4  (
    .i0(\inst_dob_mux_b6/B0_8 ),
    .i1(\inst_dob_mux_b6/B0_9 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b6/B1_4 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_1_5  (
    .i0(\inst_dob_mux_b6/B0_10 ),
    .i1(\inst_dob_mux_b6/B0_11 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b6/B1_5 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_1_6  (
    .i0(\inst_dob_mux_b6/B0_12 ),
    .i1(\inst_dob_mux_b6/B0_13 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b6/B1_6 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_1_7  (
    .i0(\inst_dob_mux_b6/B0_14 ),
    .i1(\inst_dob_mux_b6/B0_15 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b6/B1_7 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_1_8  (
    .i0(\inst_dob_mux_b6/B0_16 ),
    .i1(\inst_dob_mux_b6/B0_17 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b6/B1_8 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_1_9  (
    .i0(\inst_dob_mux_b6/B0_18 ),
    .i1(\inst_dob_mux_b6/B0_19 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b6/B1_9 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_2_0  (
    .i0(\inst_dob_mux_b6/B1_0 ),
    .i1(\inst_dob_mux_b6/B1_1 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b6/B2_0 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_2_1  (
    .i0(\inst_dob_mux_b6/B1_2 ),
    .i1(\inst_dob_mux_b6/B1_3 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b6/B2_1 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_2_10  (
    .i0(\inst_dob_mux_b6/B1_20 ),
    .i1(\inst_dob_mux_b6/B1_21 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b6/B2_10 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_2_11  (
    .i0(\inst_dob_mux_b6/B1_22 ),
    .i1(\inst_dob_mux_b6/B1_23 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b6/B2_11 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_2_12  (
    .i0(\inst_dob_mux_b6/B1_24 ),
    .i1(\inst_dob_mux_b6/B1_25 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b6/B2_12 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_2_13  (
    .i0(\inst_dob_mux_b6/B1_26 ),
    .i1(\inst_dob_mux_b6/B1_27 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b6/B2_13 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_2_14  (
    .i0(\inst_dob_mux_b6/B1_28 ),
    .i1(\inst_dob_mux_b6/B1_29 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b6/B2_14 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_2_15  (
    .i0(\inst_dob_mux_b6/B1_30 ),
    .i1(\inst_dob_mux_b6/B1_31 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b6/B2_15 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_2_2  (
    .i0(\inst_dob_mux_b6/B1_4 ),
    .i1(\inst_dob_mux_b6/B1_5 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b6/B2_2 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_2_3  (
    .i0(\inst_dob_mux_b6/B1_6 ),
    .i1(\inst_dob_mux_b6/B1_7 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b6/B2_3 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_2_4  (
    .i0(\inst_dob_mux_b6/B1_8 ),
    .i1(\inst_dob_mux_b6/B1_9 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b6/B2_4 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_2_5  (
    .i0(\inst_dob_mux_b6/B1_10 ),
    .i1(\inst_dob_mux_b6/B1_11 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b6/B2_5 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_2_6  (
    .i0(\inst_dob_mux_b6/B1_12 ),
    .i1(\inst_dob_mux_b6/B1_13 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b6/B2_6 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_2_7  (
    .i0(\inst_dob_mux_b6/B1_14 ),
    .i1(\inst_dob_mux_b6/B1_15 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b6/B2_7 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_2_8  (
    .i0(\inst_dob_mux_b6/B1_16 ),
    .i1(\inst_dob_mux_b6/B1_17 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b6/B2_8 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_2_9  (
    .i0(\inst_dob_mux_b6/B1_18 ),
    .i1(\inst_dob_mux_b6/B1_19 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b6/B2_9 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_3_0  (
    .i0(\inst_dob_mux_b6/B2_0 ),
    .i1(\inst_dob_mux_b6/B2_1 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b6/B3_0 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_3_1  (
    .i0(\inst_dob_mux_b6/B2_2 ),
    .i1(\inst_dob_mux_b6/B2_3 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b6/B3_1 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_3_2  (
    .i0(\inst_dob_mux_b6/B2_4 ),
    .i1(\inst_dob_mux_b6/B2_5 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b6/B3_2 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_3_3  (
    .i0(\inst_dob_mux_b6/B2_6 ),
    .i1(\inst_dob_mux_b6/B2_7 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b6/B3_3 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_3_4  (
    .i0(\inst_dob_mux_b6/B2_8 ),
    .i1(\inst_dob_mux_b6/B2_9 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b6/B3_4 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_3_5  (
    .i0(\inst_dob_mux_b6/B2_10 ),
    .i1(\inst_dob_mux_b6/B2_11 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b6/B3_5 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_3_6  (
    .i0(\inst_dob_mux_b6/B2_12 ),
    .i1(\inst_dob_mux_b6/B2_13 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b6/B3_6 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_3_7  (
    .i0(\inst_dob_mux_b6/B2_14 ),
    .i1(\inst_dob_mux_b6/B2_15 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b6/B3_7 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_4_0  (
    .i0(\inst_dob_mux_b6/B3_0 ),
    .i1(\inst_dob_mux_b6/B3_1 ),
    .sel(addrb_piped_piped[4]),
    .o(\inst_dob_mux_b6/B4_0 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_4_1  (
    .i0(\inst_dob_mux_b6/B3_2 ),
    .i1(\inst_dob_mux_b6/B3_3 ),
    .sel(addrb_piped_piped[4]),
    .o(\inst_dob_mux_b6/B4_1 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_4_2  (
    .i0(\inst_dob_mux_b6/B3_4 ),
    .i1(\inst_dob_mux_b6/B3_5 ),
    .sel(addrb_piped_piped[4]),
    .o(\inst_dob_mux_b6/B4_2 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_4_3  (
    .i0(\inst_dob_mux_b6/B3_6 ),
    .i1(\inst_dob_mux_b6/B3_7 ),
    .sel(addrb_piped_piped[4]),
    .o(\inst_dob_mux_b6/B4_3 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_5_0  (
    .i0(\inst_dob_mux_b6/B4_0 ),
    .i1(\inst_dob_mux_b6/B4_1 ),
    .sel(addrb_piped_piped[5]),
    .o(\inst_dob_mux_b6/B5_0 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_5_1  (
    .i0(\inst_dob_mux_b6/B4_2 ),
    .i1(\inst_dob_mux_b6/B4_3 ),
    .sel(addrb_piped_piped[5]),
    .o(\inst_dob_mux_b6/B5_1 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_6_0  (
    .i0(\inst_dob_mux_b6/B5_0 ),
    .i1(\inst_dob_mux_b6/B5_1 ),
    .sel(addrb_piped_piped[6]),
    .o(dob[6]));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_0  (
    .i0(inst_dob_i0_007),
    .i1(inst_dob_i0_007),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b7/B0_0 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_1  (
    .i0(inst_dob_i2_007),
    .i1(inst_dob_i2_007),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b7/B0_1 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_10  (
    .i0(inst_dob_i20_007),
    .i1(inst_dob_i20_007),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b7/B0_10 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_11  (
    .i0(inst_dob_i22_007),
    .i1(inst_dob_i22_007),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b7/B0_11 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_12  (
    .i0(inst_dob_i24_007),
    .i1(inst_dob_i24_007),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b7/B0_12 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_13  (
    .i0(inst_dob_i26_007),
    .i1(inst_dob_i26_007),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b7/B0_13 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_14  (
    .i0(inst_dob_i28_007),
    .i1(inst_dob_i28_007),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b7/B0_14 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_15  (
    .i0(inst_dob_i30_007),
    .i1(inst_dob_i30_007),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b7/B0_15 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_16  (
    .i0(inst_dob_i32_007),
    .i1(inst_dob_i32_007),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b7/B0_16 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_17  (
    .i0(inst_dob_i34_007),
    .i1(inst_dob_i34_007),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b7/B0_17 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_18  (
    .i0(inst_dob_i36_007),
    .i1(inst_dob_i36_007),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b7/B0_18 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_19  (
    .i0(inst_dob_i38_007),
    .i1(inst_dob_i38_007),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b7/B0_19 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_2  (
    .i0(inst_dob_i4_007),
    .i1(inst_dob_i4_007),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b7/B0_2 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_20  (
    .i0(inst_dob_i40_007),
    .i1(inst_dob_i40_007),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b7/B0_20 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_21  (
    .i0(inst_dob_i42_007),
    .i1(inst_dob_i42_007),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b7/B0_21 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_22  (
    .i0(inst_dob_i44_007),
    .i1(inst_dob_i44_007),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b7/B0_22 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_23  (
    .i0(inst_dob_i46_007),
    .i1(inst_dob_i46_007),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b7/B0_23 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_24  (
    .i0(inst_dob_i48_007),
    .i1(inst_dob_i48_007),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b7/B0_24 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_25  (
    .i0(inst_dob_i50_007),
    .i1(inst_dob_i50_007),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b7/B0_25 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_26  (
    .i0(inst_dob_i52_007),
    .i1(inst_dob_i52_007),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b7/B0_26 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_27  (
    .i0(inst_dob_i54_007),
    .i1(inst_dob_i54_007),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b7/B0_27 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_28  (
    .i0(inst_dob_i56_007),
    .i1(inst_dob_i56_007),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b7/B0_28 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_29  (
    .i0(inst_dob_i58_007),
    .i1(inst_dob_i58_007),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b7/B0_29 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_3  (
    .i0(inst_dob_i6_007),
    .i1(inst_dob_i6_007),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b7/B0_3 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_30  (
    .i0(inst_dob_i60_007),
    .i1(inst_dob_i60_007),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b7/B0_30 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_31  (
    .i0(inst_dob_i62_007),
    .i1(inst_dob_i62_007),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b7/B0_31 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_32  (
    .i0(inst_dob_i64_007),
    .i1(inst_dob_i64_007),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b7/B0_32 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_33  (
    .i0(inst_dob_i64_007),
    .i1(inst_dob_i64_007),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b7/B0_33 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_34  (
    .i0(inst_dob_i64_007),
    .i1(inst_dob_i64_007),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b7/B0_34 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_35  (
    .i0(inst_dob_i64_007),
    .i1(inst_dob_i64_007),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b7/B0_35 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_36  (
    .i0(inst_dob_i64_007),
    .i1(inst_dob_i64_007),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b7/B0_36 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_37  (
    .i0(inst_dob_i64_007),
    .i1(inst_dob_i64_007),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b7/B0_37 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_38  (
    .i0(inst_dob_i64_007),
    .i1(inst_dob_i64_007),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b7/B0_38 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_39  (
    .i0(inst_dob_i64_007),
    .i1(inst_dob_i64_007),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b7/B0_39 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_4  (
    .i0(inst_dob_i8_007),
    .i1(inst_dob_i8_007),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b7/B0_4 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_40  (
    .i0(inst_dob_i64_007),
    .i1(inst_dob_i64_007),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b7/B0_40 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_41  (
    .i0(inst_dob_i64_007),
    .i1(inst_dob_i64_007),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b7/B0_41 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_42  (
    .i0(inst_dob_i64_007),
    .i1(inst_dob_i64_007),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b7/B0_42 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_43  (
    .i0(inst_dob_i64_007),
    .i1(inst_dob_i64_007),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b7/B0_43 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_44  (
    .i0(inst_dob_i64_007),
    .i1(inst_dob_i64_007),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b7/B0_44 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_45  (
    .i0(inst_dob_i64_007),
    .i1(inst_dob_i64_007),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b7/B0_45 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_46  (
    .i0(inst_dob_i64_007),
    .i1(inst_dob_i64_007),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b7/B0_46 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_47  (
    .i0(inst_dob_i64_007),
    .i1(inst_dob_i64_007),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b7/B0_47 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_48  (
    .i0(inst_dob_i64_007),
    .i1(inst_dob_i64_007),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b7/B0_48 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_49  (
    .i0(inst_dob_i64_007),
    .i1(inst_dob_i64_007),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b7/B0_49 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_5  (
    .i0(inst_dob_i10_007),
    .i1(inst_dob_i10_007),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b7/B0_5 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_50  (
    .i0(inst_dob_i64_007),
    .i1(inst_dob_i64_007),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b7/B0_50 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_51  (
    .i0(inst_dob_i64_007),
    .i1(inst_dob_i64_007),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b7/B0_51 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_52  (
    .i0(inst_dob_i64_007),
    .i1(inst_dob_i64_007),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b7/B0_52 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_53  (
    .i0(inst_dob_i64_007),
    .i1(inst_dob_i64_007),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b7/B0_53 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_54  (
    .i0(inst_dob_i64_007),
    .i1(inst_dob_i64_007),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b7/B0_54 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_55  (
    .i0(inst_dob_i64_007),
    .i1(inst_dob_i64_007),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b7/B0_55 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_56  (
    .i0(inst_dob_i64_007),
    .i1(inst_dob_i64_007),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b7/B0_56 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_57  (
    .i0(inst_dob_i64_007),
    .i1(inst_dob_i64_007),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b7/B0_57 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_58  (
    .i0(inst_dob_i64_007),
    .i1(inst_dob_i64_007),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b7/B0_58 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_59  (
    .i0(inst_dob_i64_007),
    .i1(inst_dob_i64_007),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b7/B0_59 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_6  (
    .i0(inst_dob_i12_007),
    .i1(inst_dob_i12_007),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b7/B0_6 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_60  (
    .i0(inst_dob_i64_007),
    .i1(inst_dob_i64_007),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b7/B0_60 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_61  (
    .i0(inst_dob_i64_007),
    .i1(inst_dob_i64_007),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b7/B0_61 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_62  (
    .i0(inst_dob_i64_007),
    .i1(inst_dob_i64_007),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b7/B0_62 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_63  (
    .i0(inst_dob_i64_007),
    .i1(inst_dob_i64_007),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b7/B0_63 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_7  (
    .i0(inst_dob_i14_007),
    .i1(inst_dob_i14_007),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b7/B0_7 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_8  (
    .i0(inst_dob_i16_007),
    .i1(inst_dob_i16_007),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b7/B0_8 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_9  (
    .i0(inst_dob_i18_007),
    .i1(inst_dob_i18_007),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b7/B0_9 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_1_0  (
    .i0(\inst_dob_mux_b7/B0_0 ),
    .i1(\inst_dob_mux_b7/B0_1 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b7/B1_0 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_1_1  (
    .i0(\inst_dob_mux_b7/B0_2 ),
    .i1(\inst_dob_mux_b7/B0_3 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b7/B1_1 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_1_10  (
    .i0(\inst_dob_mux_b7/B0_20 ),
    .i1(\inst_dob_mux_b7/B0_21 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b7/B1_10 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_1_11  (
    .i0(\inst_dob_mux_b7/B0_22 ),
    .i1(\inst_dob_mux_b7/B0_23 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b7/B1_11 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_1_12  (
    .i0(\inst_dob_mux_b7/B0_24 ),
    .i1(\inst_dob_mux_b7/B0_25 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b7/B1_12 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_1_13  (
    .i0(\inst_dob_mux_b7/B0_26 ),
    .i1(\inst_dob_mux_b7/B0_27 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b7/B1_13 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_1_14  (
    .i0(\inst_dob_mux_b7/B0_28 ),
    .i1(\inst_dob_mux_b7/B0_29 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b7/B1_14 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_1_15  (
    .i0(\inst_dob_mux_b7/B0_30 ),
    .i1(\inst_dob_mux_b7/B0_31 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b7/B1_15 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_1_16  (
    .i0(\inst_dob_mux_b7/B0_32 ),
    .i1(\inst_dob_mux_b7/B0_33 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b7/B1_16 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_1_17  (
    .i0(\inst_dob_mux_b7/B0_34 ),
    .i1(\inst_dob_mux_b7/B0_35 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b7/B1_17 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_1_18  (
    .i0(\inst_dob_mux_b7/B0_36 ),
    .i1(\inst_dob_mux_b7/B0_37 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b7/B1_18 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_1_19  (
    .i0(\inst_dob_mux_b7/B0_38 ),
    .i1(\inst_dob_mux_b7/B0_39 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b7/B1_19 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_1_2  (
    .i0(\inst_dob_mux_b7/B0_4 ),
    .i1(\inst_dob_mux_b7/B0_5 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b7/B1_2 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_1_20  (
    .i0(\inst_dob_mux_b7/B0_40 ),
    .i1(\inst_dob_mux_b7/B0_41 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b7/B1_20 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_1_21  (
    .i0(\inst_dob_mux_b7/B0_42 ),
    .i1(\inst_dob_mux_b7/B0_43 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b7/B1_21 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_1_22  (
    .i0(\inst_dob_mux_b7/B0_44 ),
    .i1(\inst_dob_mux_b7/B0_45 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b7/B1_22 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_1_23  (
    .i0(\inst_dob_mux_b7/B0_46 ),
    .i1(\inst_dob_mux_b7/B0_47 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b7/B1_23 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_1_24  (
    .i0(\inst_dob_mux_b7/B0_48 ),
    .i1(\inst_dob_mux_b7/B0_49 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b7/B1_24 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_1_25  (
    .i0(\inst_dob_mux_b7/B0_50 ),
    .i1(\inst_dob_mux_b7/B0_51 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b7/B1_25 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_1_26  (
    .i0(\inst_dob_mux_b7/B0_52 ),
    .i1(\inst_dob_mux_b7/B0_53 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b7/B1_26 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_1_27  (
    .i0(\inst_dob_mux_b7/B0_54 ),
    .i1(\inst_dob_mux_b7/B0_55 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b7/B1_27 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_1_28  (
    .i0(\inst_dob_mux_b7/B0_56 ),
    .i1(\inst_dob_mux_b7/B0_57 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b7/B1_28 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_1_29  (
    .i0(\inst_dob_mux_b7/B0_58 ),
    .i1(\inst_dob_mux_b7/B0_59 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b7/B1_29 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_1_3  (
    .i0(\inst_dob_mux_b7/B0_6 ),
    .i1(\inst_dob_mux_b7/B0_7 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b7/B1_3 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_1_30  (
    .i0(\inst_dob_mux_b7/B0_60 ),
    .i1(\inst_dob_mux_b7/B0_61 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b7/B1_30 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_1_31  (
    .i0(\inst_dob_mux_b7/B0_62 ),
    .i1(\inst_dob_mux_b7/B0_63 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b7/B1_31 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_1_4  (
    .i0(\inst_dob_mux_b7/B0_8 ),
    .i1(\inst_dob_mux_b7/B0_9 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b7/B1_4 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_1_5  (
    .i0(\inst_dob_mux_b7/B0_10 ),
    .i1(\inst_dob_mux_b7/B0_11 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b7/B1_5 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_1_6  (
    .i0(\inst_dob_mux_b7/B0_12 ),
    .i1(\inst_dob_mux_b7/B0_13 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b7/B1_6 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_1_7  (
    .i0(\inst_dob_mux_b7/B0_14 ),
    .i1(\inst_dob_mux_b7/B0_15 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b7/B1_7 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_1_8  (
    .i0(\inst_dob_mux_b7/B0_16 ),
    .i1(\inst_dob_mux_b7/B0_17 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b7/B1_8 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_1_9  (
    .i0(\inst_dob_mux_b7/B0_18 ),
    .i1(\inst_dob_mux_b7/B0_19 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b7/B1_9 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_2_0  (
    .i0(\inst_dob_mux_b7/B1_0 ),
    .i1(\inst_dob_mux_b7/B1_1 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b7/B2_0 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_2_1  (
    .i0(\inst_dob_mux_b7/B1_2 ),
    .i1(\inst_dob_mux_b7/B1_3 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b7/B2_1 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_2_10  (
    .i0(\inst_dob_mux_b7/B1_20 ),
    .i1(\inst_dob_mux_b7/B1_21 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b7/B2_10 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_2_11  (
    .i0(\inst_dob_mux_b7/B1_22 ),
    .i1(\inst_dob_mux_b7/B1_23 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b7/B2_11 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_2_12  (
    .i0(\inst_dob_mux_b7/B1_24 ),
    .i1(\inst_dob_mux_b7/B1_25 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b7/B2_12 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_2_13  (
    .i0(\inst_dob_mux_b7/B1_26 ),
    .i1(\inst_dob_mux_b7/B1_27 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b7/B2_13 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_2_14  (
    .i0(\inst_dob_mux_b7/B1_28 ),
    .i1(\inst_dob_mux_b7/B1_29 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b7/B2_14 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_2_15  (
    .i0(\inst_dob_mux_b7/B1_30 ),
    .i1(\inst_dob_mux_b7/B1_31 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b7/B2_15 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_2_2  (
    .i0(\inst_dob_mux_b7/B1_4 ),
    .i1(\inst_dob_mux_b7/B1_5 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b7/B2_2 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_2_3  (
    .i0(\inst_dob_mux_b7/B1_6 ),
    .i1(\inst_dob_mux_b7/B1_7 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b7/B2_3 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_2_4  (
    .i0(\inst_dob_mux_b7/B1_8 ),
    .i1(\inst_dob_mux_b7/B1_9 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b7/B2_4 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_2_5  (
    .i0(\inst_dob_mux_b7/B1_10 ),
    .i1(\inst_dob_mux_b7/B1_11 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b7/B2_5 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_2_6  (
    .i0(\inst_dob_mux_b7/B1_12 ),
    .i1(\inst_dob_mux_b7/B1_13 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b7/B2_6 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_2_7  (
    .i0(\inst_dob_mux_b7/B1_14 ),
    .i1(\inst_dob_mux_b7/B1_15 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b7/B2_7 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_2_8  (
    .i0(\inst_dob_mux_b7/B1_16 ),
    .i1(\inst_dob_mux_b7/B1_17 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b7/B2_8 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_2_9  (
    .i0(\inst_dob_mux_b7/B1_18 ),
    .i1(\inst_dob_mux_b7/B1_19 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b7/B2_9 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_3_0  (
    .i0(\inst_dob_mux_b7/B2_0 ),
    .i1(\inst_dob_mux_b7/B2_1 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b7/B3_0 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_3_1  (
    .i0(\inst_dob_mux_b7/B2_2 ),
    .i1(\inst_dob_mux_b7/B2_3 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b7/B3_1 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_3_2  (
    .i0(\inst_dob_mux_b7/B2_4 ),
    .i1(\inst_dob_mux_b7/B2_5 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b7/B3_2 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_3_3  (
    .i0(\inst_dob_mux_b7/B2_6 ),
    .i1(\inst_dob_mux_b7/B2_7 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b7/B3_3 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_3_4  (
    .i0(\inst_dob_mux_b7/B2_8 ),
    .i1(\inst_dob_mux_b7/B2_9 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b7/B3_4 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_3_5  (
    .i0(\inst_dob_mux_b7/B2_10 ),
    .i1(\inst_dob_mux_b7/B2_11 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b7/B3_5 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_3_6  (
    .i0(\inst_dob_mux_b7/B2_12 ),
    .i1(\inst_dob_mux_b7/B2_13 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b7/B3_6 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_3_7  (
    .i0(\inst_dob_mux_b7/B2_14 ),
    .i1(\inst_dob_mux_b7/B2_15 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b7/B3_7 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_4_0  (
    .i0(\inst_dob_mux_b7/B3_0 ),
    .i1(\inst_dob_mux_b7/B3_1 ),
    .sel(addrb_piped_piped[4]),
    .o(\inst_dob_mux_b7/B4_0 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_4_1  (
    .i0(\inst_dob_mux_b7/B3_2 ),
    .i1(\inst_dob_mux_b7/B3_3 ),
    .sel(addrb_piped_piped[4]),
    .o(\inst_dob_mux_b7/B4_1 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_4_2  (
    .i0(\inst_dob_mux_b7/B3_4 ),
    .i1(\inst_dob_mux_b7/B3_5 ),
    .sel(addrb_piped_piped[4]),
    .o(\inst_dob_mux_b7/B4_2 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_4_3  (
    .i0(\inst_dob_mux_b7/B3_6 ),
    .i1(\inst_dob_mux_b7/B3_7 ),
    .sel(addrb_piped_piped[4]),
    .o(\inst_dob_mux_b7/B4_3 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_5_0  (
    .i0(\inst_dob_mux_b7/B4_0 ),
    .i1(\inst_dob_mux_b7/B4_1 ),
    .sel(addrb_piped_piped[5]),
    .o(\inst_dob_mux_b7/B5_0 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_5_1  (
    .i0(\inst_dob_mux_b7/B4_2 ),
    .i1(\inst_dob_mux_b7/B4_3 ),
    .sel(addrb_piped_piped[5]),
    .o(\inst_dob_mux_b7/B5_1 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_6_0  (
    .i0(\inst_dob_mux_b7/B5_0 ),
    .i1(\inst_dob_mux_b7/B5_1 ),
    .sel(addrb_piped_piped[6]),
    .o(dob[7]));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_0  (
    .i0(inst_dob_i0_008),
    .i1(inst_dob_i0_008),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b8/B0_0 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_1  (
    .i0(inst_dob_i2_008),
    .i1(inst_dob_i2_008),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b8/B0_1 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_10  (
    .i0(inst_dob_i20_008),
    .i1(inst_dob_i20_008),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b8/B0_10 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_11  (
    .i0(inst_dob_i22_008),
    .i1(inst_dob_i22_008),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b8/B0_11 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_12  (
    .i0(inst_dob_i24_008),
    .i1(inst_dob_i24_008),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b8/B0_12 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_13  (
    .i0(inst_dob_i26_008),
    .i1(inst_dob_i26_008),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b8/B0_13 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_14  (
    .i0(inst_dob_i28_008),
    .i1(inst_dob_i28_008),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b8/B0_14 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_15  (
    .i0(inst_dob_i30_008),
    .i1(inst_dob_i30_008),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b8/B0_15 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_16  (
    .i0(inst_dob_i32_008),
    .i1(inst_dob_i32_008),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b8/B0_16 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_17  (
    .i0(inst_dob_i34_008),
    .i1(inst_dob_i34_008),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b8/B0_17 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_18  (
    .i0(inst_dob_i36_008),
    .i1(inst_dob_i36_008),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b8/B0_18 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_19  (
    .i0(inst_dob_i38_008),
    .i1(inst_dob_i38_008),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b8/B0_19 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_2  (
    .i0(inst_dob_i4_008),
    .i1(inst_dob_i4_008),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b8/B0_2 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_20  (
    .i0(inst_dob_i40_008),
    .i1(inst_dob_i40_008),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b8/B0_20 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_21  (
    .i0(inst_dob_i42_008),
    .i1(inst_dob_i42_008),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b8/B0_21 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_22  (
    .i0(inst_dob_i44_008),
    .i1(inst_dob_i44_008),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b8/B0_22 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_23  (
    .i0(inst_dob_i46_008),
    .i1(inst_dob_i46_008),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b8/B0_23 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_24  (
    .i0(inst_dob_i48_008),
    .i1(inst_dob_i48_008),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b8/B0_24 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_25  (
    .i0(inst_dob_i50_008),
    .i1(inst_dob_i50_008),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b8/B0_25 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_26  (
    .i0(inst_dob_i52_008),
    .i1(inst_dob_i52_008),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b8/B0_26 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_27  (
    .i0(inst_dob_i54_008),
    .i1(inst_dob_i54_008),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b8/B0_27 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_28  (
    .i0(inst_dob_i56_008),
    .i1(inst_dob_i56_008),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b8/B0_28 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_29  (
    .i0(inst_dob_i58_008),
    .i1(inst_dob_i58_008),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b8/B0_29 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_3  (
    .i0(inst_dob_i6_008),
    .i1(inst_dob_i6_008),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b8/B0_3 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_30  (
    .i0(inst_dob_i60_008),
    .i1(inst_dob_i60_008),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b8/B0_30 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_31  (
    .i0(inst_dob_i62_008),
    .i1(inst_dob_i62_008),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b8/B0_31 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_32  (
    .i0(inst_dob_i64_008),
    .i1(inst_dob_i64_008),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b8/B0_32 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_33  (
    .i0(inst_dob_i64_008),
    .i1(inst_dob_i64_008),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b8/B0_33 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_34  (
    .i0(inst_dob_i64_008),
    .i1(inst_dob_i64_008),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b8/B0_34 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_35  (
    .i0(inst_dob_i64_008),
    .i1(inst_dob_i64_008),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b8/B0_35 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_36  (
    .i0(inst_dob_i64_008),
    .i1(inst_dob_i64_008),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b8/B0_36 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_37  (
    .i0(inst_dob_i64_008),
    .i1(inst_dob_i64_008),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b8/B0_37 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_38  (
    .i0(inst_dob_i64_008),
    .i1(inst_dob_i64_008),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b8/B0_38 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_39  (
    .i0(inst_dob_i64_008),
    .i1(inst_dob_i64_008),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b8/B0_39 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_4  (
    .i0(inst_dob_i8_008),
    .i1(inst_dob_i8_008),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b8/B0_4 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_40  (
    .i0(inst_dob_i64_008),
    .i1(inst_dob_i64_008),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b8/B0_40 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_41  (
    .i0(inst_dob_i64_008),
    .i1(inst_dob_i64_008),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b8/B0_41 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_42  (
    .i0(inst_dob_i64_008),
    .i1(inst_dob_i64_008),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b8/B0_42 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_43  (
    .i0(inst_dob_i64_008),
    .i1(inst_dob_i64_008),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b8/B0_43 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_44  (
    .i0(inst_dob_i64_008),
    .i1(inst_dob_i64_008),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b8/B0_44 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_45  (
    .i0(inst_dob_i64_008),
    .i1(inst_dob_i64_008),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b8/B0_45 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_46  (
    .i0(inst_dob_i64_008),
    .i1(inst_dob_i64_008),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b8/B0_46 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_47  (
    .i0(inst_dob_i64_008),
    .i1(inst_dob_i64_008),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b8/B0_47 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_48  (
    .i0(inst_dob_i64_008),
    .i1(inst_dob_i64_008),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b8/B0_48 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_49  (
    .i0(inst_dob_i64_008),
    .i1(inst_dob_i64_008),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b8/B0_49 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_5  (
    .i0(inst_dob_i10_008),
    .i1(inst_dob_i10_008),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b8/B0_5 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_50  (
    .i0(inst_dob_i64_008),
    .i1(inst_dob_i64_008),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b8/B0_50 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_51  (
    .i0(inst_dob_i64_008),
    .i1(inst_dob_i64_008),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b8/B0_51 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_52  (
    .i0(inst_dob_i64_008),
    .i1(inst_dob_i64_008),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b8/B0_52 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_53  (
    .i0(inst_dob_i64_008),
    .i1(inst_dob_i64_008),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b8/B0_53 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_54  (
    .i0(inst_dob_i64_008),
    .i1(inst_dob_i64_008),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b8/B0_54 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_55  (
    .i0(inst_dob_i64_008),
    .i1(inst_dob_i64_008),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b8/B0_55 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_56  (
    .i0(inst_dob_i64_008),
    .i1(inst_dob_i64_008),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b8/B0_56 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_57  (
    .i0(inst_dob_i64_008),
    .i1(inst_dob_i64_008),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b8/B0_57 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_58  (
    .i0(inst_dob_i64_008),
    .i1(inst_dob_i64_008),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b8/B0_58 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_59  (
    .i0(inst_dob_i64_008),
    .i1(inst_dob_i64_008),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b8/B0_59 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_6  (
    .i0(inst_dob_i12_008),
    .i1(inst_dob_i12_008),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b8/B0_6 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_60  (
    .i0(inst_dob_i64_008),
    .i1(inst_dob_i64_008),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b8/B0_60 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_61  (
    .i0(inst_dob_i64_008),
    .i1(inst_dob_i64_008),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b8/B0_61 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_62  (
    .i0(inst_dob_i64_008),
    .i1(inst_dob_i64_008),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b8/B0_62 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_63  (
    .i0(inst_dob_i64_008),
    .i1(inst_dob_i64_008),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b8/B0_63 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_7  (
    .i0(inst_dob_i14_008),
    .i1(inst_dob_i14_008),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b8/B0_7 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_8  (
    .i0(inst_dob_i16_008),
    .i1(inst_dob_i16_008),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b8/B0_8 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_9  (
    .i0(inst_dob_i18_008),
    .i1(inst_dob_i18_008),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b8/B0_9 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_1_0  (
    .i0(\inst_dob_mux_b8/B0_0 ),
    .i1(\inst_dob_mux_b8/B0_1 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b8/B1_0 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_1_1  (
    .i0(\inst_dob_mux_b8/B0_2 ),
    .i1(\inst_dob_mux_b8/B0_3 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b8/B1_1 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_1_10  (
    .i0(\inst_dob_mux_b8/B0_20 ),
    .i1(\inst_dob_mux_b8/B0_21 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b8/B1_10 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_1_11  (
    .i0(\inst_dob_mux_b8/B0_22 ),
    .i1(\inst_dob_mux_b8/B0_23 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b8/B1_11 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_1_12  (
    .i0(\inst_dob_mux_b8/B0_24 ),
    .i1(\inst_dob_mux_b8/B0_25 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b8/B1_12 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_1_13  (
    .i0(\inst_dob_mux_b8/B0_26 ),
    .i1(\inst_dob_mux_b8/B0_27 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b8/B1_13 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_1_14  (
    .i0(\inst_dob_mux_b8/B0_28 ),
    .i1(\inst_dob_mux_b8/B0_29 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b8/B1_14 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_1_15  (
    .i0(\inst_dob_mux_b8/B0_30 ),
    .i1(\inst_dob_mux_b8/B0_31 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b8/B1_15 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_1_16  (
    .i0(\inst_dob_mux_b8/B0_32 ),
    .i1(\inst_dob_mux_b8/B0_33 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b8/B1_16 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_1_17  (
    .i0(\inst_dob_mux_b8/B0_34 ),
    .i1(\inst_dob_mux_b8/B0_35 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b8/B1_17 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_1_18  (
    .i0(\inst_dob_mux_b8/B0_36 ),
    .i1(\inst_dob_mux_b8/B0_37 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b8/B1_18 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_1_19  (
    .i0(\inst_dob_mux_b8/B0_38 ),
    .i1(\inst_dob_mux_b8/B0_39 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b8/B1_19 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_1_2  (
    .i0(\inst_dob_mux_b8/B0_4 ),
    .i1(\inst_dob_mux_b8/B0_5 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b8/B1_2 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_1_20  (
    .i0(\inst_dob_mux_b8/B0_40 ),
    .i1(\inst_dob_mux_b8/B0_41 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b8/B1_20 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_1_21  (
    .i0(\inst_dob_mux_b8/B0_42 ),
    .i1(\inst_dob_mux_b8/B0_43 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b8/B1_21 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_1_22  (
    .i0(\inst_dob_mux_b8/B0_44 ),
    .i1(\inst_dob_mux_b8/B0_45 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b8/B1_22 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_1_23  (
    .i0(\inst_dob_mux_b8/B0_46 ),
    .i1(\inst_dob_mux_b8/B0_47 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b8/B1_23 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_1_24  (
    .i0(\inst_dob_mux_b8/B0_48 ),
    .i1(\inst_dob_mux_b8/B0_49 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b8/B1_24 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_1_25  (
    .i0(\inst_dob_mux_b8/B0_50 ),
    .i1(\inst_dob_mux_b8/B0_51 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b8/B1_25 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_1_26  (
    .i0(\inst_dob_mux_b8/B0_52 ),
    .i1(\inst_dob_mux_b8/B0_53 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b8/B1_26 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_1_27  (
    .i0(\inst_dob_mux_b8/B0_54 ),
    .i1(\inst_dob_mux_b8/B0_55 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b8/B1_27 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_1_28  (
    .i0(\inst_dob_mux_b8/B0_56 ),
    .i1(\inst_dob_mux_b8/B0_57 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b8/B1_28 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_1_29  (
    .i0(\inst_dob_mux_b8/B0_58 ),
    .i1(\inst_dob_mux_b8/B0_59 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b8/B1_29 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_1_3  (
    .i0(\inst_dob_mux_b8/B0_6 ),
    .i1(\inst_dob_mux_b8/B0_7 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b8/B1_3 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_1_30  (
    .i0(\inst_dob_mux_b8/B0_60 ),
    .i1(\inst_dob_mux_b8/B0_61 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b8/B1_30 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_1_31  (
    .i0(\inst_dob_mux_b8/B0_62 ),
    .i1(\inst_dob_mux_b8/B0_63 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b8/B1_31 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_1_4  (
    .i0(\inst_dob_mux_b8/B0_8 ),
    .i1(\inst_dob_mux_b8/B0_9 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b8/B1_4 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_1_5  (
    .i0(\inst_dob_mux_b8/B0_10 ),
    .i1(\inst_dob_mux_b8/B0_11 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b8/B1_5 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_1_6  (
    .i0(\inst_dob_mux_b8/B0_12 ),
    .i1(\inst_dob_mux_b8/B0_13 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b8/B1_6 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_1_7  (
    .i0(\inst_dob_mux_b8/B0_14 ),
    .i1(\inst_dob_mux_b8/B0_15 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b8/B1_7 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_1_8  (
    .i0(\inst_dob_mux_b8/B0_16 ),
    .i1(\inst_dob_mux_b8/B0_17 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b8/B1_8 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_1_9  (
    .i0(\inst_dob_mux_b8/B0_18 ),
    .i1(\inst_dob_mux_b8/B0_19 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b8/B1_9 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_2_0  (
    .i0(\inst_dob_mux_b8/B1_0 ),
    .i1(\inst_dob_mux_b8/B1_1 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b8/B2_0 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_2_1  (
    .i0(\inst_dob_mux_b8/B1_2 ),
    .i1(\inst_dob_mux_b8/B1_3 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b8/B2_1 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_2_10  (
    .i0(\inst_dob_mux_b8/B1_20 ),
    .i1(\inst_dob_mux_b8/B1_21 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b8/B2_10 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_2_11  (
    .i0(\inst_dob_mux_b8/B1_22 ),
    .i1(\inst_dob_mux_b8/B1_23 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b8/B2_11 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_2_12  (
    .i0(\inst_dob_mux_b8/B1_24 ),
    .i1(\inst_dob_mux_b8/B1_25 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b8/B2_12 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_2_13  (
    .i0(\inst_dob_mux_b8/B1_26 ),
    .i1(\inst_dob_mux_b8/B1_27 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b8/B2_13 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_2_14  (
    .i0(\inst_dob_mux_b8/B1_28 ),
    .i1(\inst_dob_mux_b8/B1_29 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b8/B2_14 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_2_15  (
    .i0(\inst_dob_mux_b8/B1_30 ),
    .i1(\inst_dob_mux_b8/B1_31 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b8/B2_15 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_2_2  (
    .i0(\inst_dob_mux_b8/B1_4 ),
    .i1(\inst_dob_mux_b8/B1_5 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b8/B2_2 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_2_3  (
    .i0(\inst_dob_mux_b8/B1_6 ),
    .i1(\inst_dob_mux_b8/B1_7 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b8/B2_3 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_2_4  (
    .i0(\inst_dob_mux_b8/B1_8 ),
    .i1(\inst_dob_mux_b8/B1_9 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b8/B2_4 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_2_5  (
    .i0(\inst_dob_mux_b8/B1_10 ),
    .i1(\inst_dob_mux_b8/B1_11 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b8/B2_5 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_2_6  (
    .i0(\inst_dob_mux_b8/B1_12 ),
    .i1(\inst_dob_mux_b8/B1_13 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b8/B2_6 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_2_7  (
    .i0(\inst_dob_mux_b8/B1_14 ),
    .i1(\inst_dob_mux_b8/B1_15 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b8/B2_7 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_2_8  (
    .i0(\inst_dob_mux_b8/B1_16 ),
    .i1(\inst_dob_mux_b8/B1_17 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b8/B2_8 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_2_9  (
    .i0(\inst_dob_mux_b8/B1_18 ),
    .i1(\inst_dob_mux_b8/B1_19 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b8/B2_9 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_3_0  (
    .i0(\inst_dob_mux_b8/B2_0 ),
    .i1(\inst_dob_mux_b8/B2_1 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b8/B3_0 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_3_1  (
    .i0(\inst_dob_mux_b8/B2_2 ),
    .i1(\inst_dob_mux_b8/B2_3 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b8/B3_1 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_3_2  (
    .i0(\inst_dob_mux_b8/B2_4 ),
    .i1(\inst_dob_mux_b8/B2_5 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b8/B3_2 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_3_3  (
    .i0(\inst_dob_mux_b8/B2_6 ),
    .i1(\inst_dob_mux_b8/B2_7 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b8/B3_3 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_3_4  (
    .i0(\inst_dob_mux_b8/B2_8 ),
    .i1(\inst_dob_mux_b8/B2_9 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b8/B3_4 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_3_5  (
    .i0(\inst_dob_mux_b8/B2_10 ),
    .i1(\inst_dob_mux_b8/B2_11 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b8/B3_5 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_3_6  (
    .i0(\inst_dob_mux_b8/B2_12 ),
    .i1(\inst_dob_mux_b8/B2_13 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b8/B3_6 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_3_7  (
    .i0(\inst_dob_mux_b8/B2_14 ),
    .i1(\inst_dob_mux_b8/B2_15 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b8/B3_7 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_4_0  (
    .i0(\inst_dob_mux_b8/B3_0 ),
    .i1(\inst_dob_mux_b8/B3_1 ),
    .sel(addrb_piped_piped[4]),
    .o(\inst_dob_mux_b8/B4_0 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_4_1  (
    .i0(\inst_dob_mux_b8/B3_2 ),
    .i1(\inst_dob_mux_b8/B3_3 ),
    .sel(addrb_piped_piped[4]),
    .o(\inst_dob_mux_b8/B4_1 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_4_2  (
    .i0(\inst_dob_mux_b8/B3_4 ),
    .i1(\inst_dob_mux_b8/B3_5 ),
    .sel(addrb_piped_piped[4]),
    .o(\inst_dob_mux_b8/B4_2 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_4_3  (
    .i0(\inst_dob_mux_b8/B3_6 ),
    .i1(\inst_dob_mux_b8/B3_7 ),
    .sel(addrb_piped_piped[4]),
    .o(\inst_dob_mux_b8/B4_3 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_5_0  (
    .i0(\inst_dob_mux_b8/B4_0 ),
    .i1(\inst_dob_mux_b8/B4_1 ),
    .sel(addrb_piped_piped[5]),
    .o(\inst_dob_mux_b8/B5_0 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_5_1  (
    .i0(\inst_dob_mux_b8/B4_2 ),
    .i1(\inst_dob_mux_b8/B4_3 ),
    .sel(addrb_piped_piped[5]),
    .o(\inst_dob_mux_b8/B5_1 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_6_0  (
    .i0(\inst_dob_mux_b8/B5_0 ),
    .i1(\inst_dob_mux_b8/B5_1 ),
    .sel(addrb_piped_piped[6]),
    .o(dob[8]));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_0  (
    .i0(inst_dob_i0_009),
    .i1(inst_dob_i0_009),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b9/B0_0 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_1  (
    .i0(inst_dob_i0_009),
    .i1(inst_dob_i0_009),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b9/B0_1 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_10  (
    .i0(inst_dob_i16_009),
    .i1(inst_dob_i16_009),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b9/B0_10 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_11  (
    .i0(inst_dob_i16_009),
    .i1(inst_dob_i16_009),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b9/B0_11 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_12  (
    .i0(inst_dob_i16_009),
    .i1(inst_dob_i16_009),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b9/B0_12 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_13  (
    .i0(inst_dob_i16_009),
    .i1(inst_dob_i16_009),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b9/B0_13 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_14  (
    .i0(inst_dob_i16_009),
    .i1(inst_dob_i16_009),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b9/B0_14 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_15  (
    .i0(inst_dob_i16_009),
    .i1(inst_dob_i16_009),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b9/B0_15 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_16  (
    .i0(inst_dob_i32_009),
    .i1(inst_dob_i32_009),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b9/B0_16 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_17  (
    .i0(inst_dob_i32_009),
    .i1(inst_dob_i32_009),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b9/B0_17 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_18  (
    .i0(inst_dob_i32_009),
    .i1(inst_dob_i32_009),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b9/B0_18 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_19  (
    .i0(inst_dob_i32_009),
    .i1(inst_dob_i32_009),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b9/B0_19 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_2  (
    .i0(inst_dob_i0_009),
    .i1(inst_dob_i0_009),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b9/B0_2 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_20  (
    .i0(inst_dob_i32_009),
    .i1(inst_dob_i32_009),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b9/B0_20 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_21  (
    .i0(inst_dob_i32_009),
    .i1(inst_dob_i32_009),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b9/B0_21 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_22  (
    .i0(inst_dob_i32_009),
    .i1(inst_dob_i32_009),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b9/B0_22 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_23  (
    .i0(inst_dob_i32_009),
    .i1(inst_dob_i32_009),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b9/B0_23 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_24  (
    .i0(inst_dob_i48_009),
    .i1(inst_dob_i48_009),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b9/B0_24 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_25  (
    .i0(inst_dob_i48_009),
    .i1(inst_dob_i48_009),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b9/B0_25 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_26  (
    .i0(inst_dob_i48_009),
    .i1(inst_dob_i48_009),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b9/B0_26 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_27  (
    .i0(inst_dob_i48_009),
    .i1(inst_dob_i48_009),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b9/B0_27 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_28  (
    .i0(inst_dob_i48_009),
    .i1(inst_dob_i48_009),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b9/B0_28 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_29  (
    .i0(inst_dob_i48_009),
    .i1(inst_dob_i48_009),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b9/B0_29 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_3  (
    .i0(inst_dob_i0_009),
    .i1(inst_dob_i0_009),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b9/B0_3 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_30  (
    .i0(inst_dob_i48_009),
    .i1(inst_dob_i48_009),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b9/B0_30 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_31  (
    .i0(inst_dob_i48_009),
    .i1(inst_dob_i48_009),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b9/B0_31 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_32  (
    .i0(inst_dob_i64_009),
    .i1(inst_dob_i64_009),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b9/B0_32 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_33  (
    .i0(inst_dob_i64_009),
    .i1(inst_dob_i64_009),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b9/B0_33 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_34  (
    .i0(inst_dob_i64_009),
    .i1(inst_dob_i64_009),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b9/B0_34 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_35  (
    .i0(inst_dob_i64_009),
    .i1(inst_dob_i64_009),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b9/B0_35 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_36  (
    .i0(inst_dob_i64_009),
    .i1(inst_dob_i64_009),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b9/B0_36 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_37  (
    .i0(inst_dob_i64_009),
    .i1(inst_dob_i64_009),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b9/B0_37 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_38  (
    .i0(inst_dob_i64_009),
    .i1(inst_dob_i64_009),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b9/B0_38 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_39  (
    .i0(inst_dob_i64_009),
    .i1(inst_dob_i64_009),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b9/B0_39 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_4  (
    .i0(inst_dob_i0_009),
    .i1(inst_dob_i0_009),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b9/B0_4 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_40  (
    .i0(inst_dob_i64_009),
    .i1(inst_dob_i64_009),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b9/B0_40 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_41  (
    .i0(inst_dob_i64_009),
    .i1(inst_dob_i64_009),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b9/B0_41 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_42  (
    .i0(inst_dob_i64_009),
    .i1(inst_dob_i64_009),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b9/B0_42 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_43  (
    .i0(inst_dob_i64_009),
    .i1(inst_dob_i64_009),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b9/B0_43 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_44  (
    .i0(inst_dob_i64_009),
    .i1(inst_dob_i64_009),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b9/B0_44 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_45  (
    .i0(inst_dob_i64_009),
    .i1(inst_dob_i64_009),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b9/B0_45 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_46  (
    .i0(inst_dob_i64_009),
    .i1(inst_dob_i64_009),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b9/B0_46 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_47  (
    .i0(inst_dob_i64_009),
    .i1(inst_dob_i64_009),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b9/B0_47 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_48  (
    .i0(inst_dob_i64_009),
    .i1(inst_dob_i64_009),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b9/B0_48 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_49  (
    .i0(inst_dob_i64_009),
    .i1(inst_dob_i64_009),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b9/B0_49 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_5  (
    .i0(inst_dob_i0_009),
    .i1(inst_dob_i0_009),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b9/B0_5 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_50  (
    .i0(inst_dob_i64_009),
    .i1(inst_dob_i64_009),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b9/B0_50 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_51  (
    .i0(inst_dob_i64_009),
    .i1(inst_dob_i64_009),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b9/B0_51 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_52  (
    .i0(inst_dob_i64_009),
    .i1(inst_dob_i64_009),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b9/B0_52 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_53  (
    .i0(inst_dob_i64_009),
    .i1(inst_dob_i64_009),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b9/B0_53 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_54  (
    .i0(inst_dob_i64_009),
    .i1(inst_dob_i64_009),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b9/B0_54 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_55  (
    .i0(inst_dob_i64_009),
    .i1(inst_dob_i64_009),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b9/B0_55 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_56  (
    .i0(inst_dob_i64_009),
    .i1(inst_dob_i64_009),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b9/B0_56 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_57  (
    .i0(inst_dob_i64_009),
    .i1(inst_dob_i64_009),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b9/B0_57 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_58  (
    .i0(inst_dob_i64_009),
    .i1(inst_dob_i64_009),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b9/B0_58 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_59  (
    .i0(inst_dob_i64_009),
    .i1(inst_dob_i64_009),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b9/B0_59 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_6  (
    .i0(inst_dob_i0_009),
    .i1(inst_dob_i0_009),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b9/B0_6 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_60  (
    .i0(inst_dob_i64_009),
    .i1(inst_dob_i64_009),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b9/B0_60 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_61  (
    .i0(inst_dob_i64_009),
    .i1(inst_dob_i64_009),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b9/B0_61 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_62  (
    .i0(inst_dob_i64_009),
    .i1(inst_dob_i64_009),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b9/B0_62 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_63  (
    .i0(inst_dob_i64_009),
    .i1(inst_dob_i64_009),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b9/B0_63 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_7  (
    .i0(inst_dob_i0_009),
    .i1(inst_dob_i0_009),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b9/B0_7 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_8  (
    .i0(inst_dob_i16_009),
    .i1(inst_dob_i16_009),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b9/B0_8 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_9  (
    .i0(inst_dob_i16_009),
    .i1(inst_dob_i16_009),
    .sel(addrb_piped_piped[0]),
    .o(\inst_dob_mux_b9/B0_9 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_1_0  (
    .i0(\inst_dob_mux_b9/B0_0 ),
    .i1(\inst_dob_mux_b9/B0_1 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b9/B1_0 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_1_1  (
    .i0(\inst_dob_mux_b9/B0_2 ),
    .i1(\inst_dob_mux_b9/B0_3 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b9/B1_1 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_1_10  (
    .i0(\inst_dob_mux_b9/B0_20 ),
    .i1(\inst_dob_mux_b9/B0_21 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b9/B1_10 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_1_11  (
    .i0(\inst_dob_mux_b9/B0_22 ),
    .i1(\inst_dob_mux_b9/B0_23 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b9/B1_11 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_1_12  (
    .i0(\inst_dob_mux_b9/B0_24 ),
    .i1(\inst_dob_mux_b9/B0_25 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b9/B1_12 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_1_13  (
    .i0(\inst_dob_mux_b9/B0_26 ),
    .i1(\inst_dob_mux_b9/B0_27 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b9/B1_13 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_1_14  (
    .i0(\inst_dob_mux_b9/B0_28 ),
    .i1(\inst_dob_mux_b9/B0_29 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b9/B1_14 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_1_15  (
    .i0(\inst_dob_mux_b9/B0_30 ),
    .i1(\inst_dob_mux_b9/B0_31 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b9/B1_15 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_1_16  (
    .i0(\inst_dob_mux_b9/B0_32 ),
    .i1(\inst_dob_mux_b9/B0_33 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b9/B1_16 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_1_17  (
    .i0(\inst_dob_mux_b9/B0_34 ),
    .i1(\inst_dob_mux_b9/B0_35 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b9/B1_17 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_1_18  (
    .i0(\inst_dob_mux_b9/B0_36 ),
    .i1(\inst_dob_mux_b9/B0_37 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b9/B1_18 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_1_19  (
    .i0(\inst_dob_mux_b9/B0_38 ),
    .i1(\inst_dob_mux_b9/B0_39 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b9/B1_19 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_1_2  (
    .i0(\inst_dob_mux_b9/B0_4 ),
    .i1(\inst_dob_mux_b9/B0_5 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b9/B1_2 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_1_20  (
    .i0(\inst_dob_mux_b9/B0_40 ),
    .i1(\inst_dob_mux_b9/B0_41 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b9/B1_20 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_1_21  (
    .i0(\inst_dob_mux_b9/B0_42 ),
    .i1(\inst_dob_mux_b9/B0_43 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b9/B1_21 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_1_22  (
    .i0(\inst_dob_mux_b9/B0_44 ),
    .i1(\inst_dob_mux_b9/B0_45 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b9/B1_22 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_1_23  (
    .i0(\inst_dob_mux_b9/B0_46 ),
    .i1(\inst_dob_mux_b9/B0_47 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b9/B1_23 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_1_24  (
    .i0(\inst_dob_mux_b9/B0_48 ),
    .i1(\inst_dob_mux_b9/B0_49 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b9/B1_24 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_1_25  (
    .i0(\inst_dob_mux_b9/B0_50 ),
    .i1(\inst_dob_mux_b9/B0_51 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b9/B1_25 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_1_26  (
    .i0(\inst_dob_mux_b9/B0_52 ),
    .i1(\inst_dob_mux_b9/B0_53 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b9/B1_26 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_1_27  (
    .i0(\inst_dob_mux_b9/B0_54 ),
    .i1(\inst_dob_mux_b9/B0_55 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b9/B1_27 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_1_28  (
    .i0(\inst_dob_mux_b9/B0_56 ),
    .i1(\inst_dob_mux_b9/B0_57 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b9/B1_28 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_1_29  (
    .i0(\inst_dob_mux_b9/B0_58 ),
    .i1(\inst_dob_mux_b9/B0_59 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b9/B1_29 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_1_3  (
    .i0(\inst_dob_mux_b9/B0_6 ),
    .i1(\inst_dob_mux_b9/B0_7 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b9/B1_3 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_1_30  (
    .i0(\inst_dob_mux_b9/B0_60 ),
    .i1(\inst_dob_mux_b9/B0_61 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b9/B1_30 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_1_31  (
    .i0(\inst_dob_mux_b9/B0_62 ),
    .i1(\inst_dob_mux_b9/B0_63 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b9/B1_31 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_1_4  (
    .i0(\inst_dob_mux_b9/B0_8 ),
    .i1(\inst_dob_mux_b9/B0_9 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b9/B1_4 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_1_5  (
    .i0(\inst_dob_mux_b9/B0_10 ),
    .i1(\inst_dob_mux_b9/B0_11 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b9/B1_5 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_1_6  (
    .i0(\inst_dob_mux_b9/B0_12 ),
    .i1(\inst_dob_mux_b9/B0_13 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b9/B1_6 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_1_7  (
    .i0(\inst_dob_mux_b9/B0_14 ),
    .i1(\inst_dob_mux_b9/B0_15 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b9/B1_7 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_1_8  (
    .i0(\inst_dob_mux_b9/B0_16 ),
    .i1(\inst_dob_mux_b9/B0_17 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b9/B1_8 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_1_9  (
    .i0(\inst_dob_mux_b9/B0_18 ),
    .i1(\inst_dob_mux_b9/B0_19 ),
    .sel(addrb_piped_piped[1]),
    .o(\inst_dob_mux_b9/B1_9 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_2_0  (
    .i0(\inst_dob_mux_b9/B1_0 ),
    .i1(\inst_dob_mux_b9/B1_1 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b9/B2_0 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_2_1  (
    .i0(\inst_dob_mux_b9/B1_2 ),
    .i1(\inst_dob_mux_b9/B1_3 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b9/B2_1 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_2_10  (
    .i0(\inst_dob_mux_b9/B1_20 ),
    .i1(\inst_dob_mux_b9/B1_21 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b9/B2_10 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_2_11  (
    .i0(\inst_dob_mux_b9/B1_22 ),
    .i1(\inst_dob_mux_b9/B1_23 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b9/B2_11 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_2_12  (
    .i0(\inst_dob_mux_b9/B1_24 ),
    .i1(\inst_dob_mux_b9/B1_25 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b9/B2_12 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_2_13  (
    .i0(\inst_dob_mux_b9/B1_26 ),
    .i1(\inst_dob_mux_b9/B1_27 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b9/B2_13 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_2_14  (
    .i0(\inst_dob_mux_b9/B1_28 ),
    .i1(\inst_dob_mux_b9/B1_29 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b9/B2_14 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_2_15  (
    .i0(\inst_dob_mux_b9/B1_30 ),
    .i1(\inst_dob_mux_b9/B1_31 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b9/B2_15 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_2_2  (
    .i0(\inst_dob_mux_b9/B1_4 ),
    .i1(\inst_dob_mux_b9/B1_5 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b9/B2_2 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_2_3  (
    .i0(\inst_dob_mux_b9/B1_6 ),
    .i1(\inst_dob_mux_b9/B1_7 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b9/B2_3 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_2_4  (
    .i0(\inst_dob_mux_b9/B1_8 ),
    .i1(\inst_dob_mux_b9/B1_9 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b9/B2_4 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_2_5  (
    .i0(\inst_dob_mux_b9/B1_10 ),
    .i1(\inst_dob_mux_b9/B1_11 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b9/B2_5 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_2_6  (
    .i0(\inst_dob_mux_b9/B1_12 ),
    .i1(\inst_dob_mux_b9/B1_13 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b9/B2_6 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_2_7  (
    .i0(\inst_dob_mux_b9/B1_14 ),
    .i1(\inst_dob_mux_b9/B1_15 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b9/B2_7 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_2_8  (
    .i0(\inst_dob_mux_b9/B1_16 ),
    .i1(\inst_dob_mux_b9/B1_17 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b9/B2_8 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_2_9  (
    .i0(\inst_dob_mux_b9/B1_18 ),
    .i1(\inst_dob_mux_b9/B1_19 ),
    .sel(addrb_piped_piped[2]),
    .o(\inst_dob_mux_b9/B2_9 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_3_0  (
    .i0(\inst_dob_mux_b9/B2_0 ),
    .i1(\inst_dob_mux_b9/B2_1 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b9/B3_0 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_3_1  (
    .i0(\inst_dob_mux_b9/B2_2 ),
    .i1(\inst_dob_mux_b9/B2_3 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b9/B3_1 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_3_2  (
    .i0(\inst_dob_mux_b9/B2_4 ),
    .i1(\inst_dob_mux_b9/B2_5 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b9/B3_2 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_3_3  (
    .i0(\inst_dob_mux_b9/B2_6 ),
    .i1(\inst_dob_mux_b9/B2_7 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b9/B3_3 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_3_4  (
    .i0(\inst_dob_mux_b9/B2_8 ),
    .i1(\inst_dob_mux_b9/B2_9 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b9/B3_4 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_3_5  (
    .i0(\inst_dob_mux_b9/B2_10 ),
    .i1(\inst_dob_mux_b9/B2_11 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b9/B3_5 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_3_6  (
    .i0(\inst_dob_mux_b9/B2_12 ),
    .i1(\inst_dob_mux_b9/B2_13 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b9/B3_6 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_3_7  (
    .i0(\inst_dob_mux_b9/B2_14 ),
    .i1(\inst_dob_mux_b9/B2_15 ),
    .sel(addrb_piped_piped[3]),
    .o(\inst_dob_mux_b9/B3_7 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_4_0  (
    .i0(\inst_dob_mux_b9/B3_0 ),
    .i1(\inst_dob_mux_b9/B3_1 ),
    .sel(addrb_piped_piped[4]),
    .o(\inst_dob_mux_b9/B4_0 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_4_1  (
    .i0(\inst_dob_mux_b9/B3_2 ),
    .i1(\inst_dob_mux_b9/B3_3 ),
    .sel(addrb_piped_piped[4]),
    .o(\inst_dob_mux_b9/B4_1 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_4_2  (
    .i0(\inst_dob_mux_b9/B3_4 ),
    .i1(\inst_dob_mux_b9/B3_5 ),
    .sel(addrb_piped_piped[4]),
    .o(\inst_dob_mux_b9/B4_2 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_4_3  (
    .i0(\inst_dob_mux_b9/B3_6 ),
    .i1(\inst_dob_mux_b9/B3_7 ),
    .sel(addrb_piped_piped[4]),
    .o(\inst_dob_mux_b9/B4_3 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_5_0  (
    .i0(\inst_dob_mux_b9/B4_0 ),
    .i1(\inst_dob_mux_b9/B4_1 ),
    .sel(addrb_piped_piped[5]),
    .o(\inst_dob_mux_b9/B5_0 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_5_1  (
    .i0(\inst_dob_mux_b9/B4_2 ),
    .i1(\inst_dob_mux_b9/B4_3 ),
    .sel(addrb_piped_piped[5]),
    .o(\inst_dob_mux_b9/B5_1 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_6_0  (
    .i0(\inst_dob_mux_b9/B5_0 ),
    .i1(\inst_dob_mux_b9/B5_1 ),
    .sel(addrb_piped_piped[6]),
    .o(dob[9]));

endmodule 

module reg_sr_as_w1
  (
  clk,
  d,
  en,
  reset,
  set,
  q
  );

  input clk;
  input d;
  input en;
  input reset;
  input set;
  output q;

  parameter REGSET = "RESET";
  wire enout;
  wire resetout;

  AL_MUX u_en0 (
    .i0(q),
    .i1(d),
    .sel(en),
    .o(enout));
  AL_MUX u_reset0 (
    .i0(enout),
    .i1(1'b0),
    .sel(reset),
    .o(resetout));
  AL_DFF #(
    .INI((REGSET == "SET") ? 1'b1 : 1'b0))
    u_seq0 (
    .clk(clk),
    .d(resetout),
    .reset(1'b0),
    .set(set),
    .q(q));

endmodule 

module AL_MUX
  (
  input i0,
  input i1,
  input sel,
  output o
  );

  wire not_sel, sel_i0, sel_i1;
  not u0 (not_sel, sel);
  and u1 (sel_i1, sel, i1);
  and u2 (sel_i0, not_sel, i0);
  or u3 (o, sel_i1, sel_i0);

endmodule

module AL_DFF
  (
  input reset,
  input set,
  input clk,
  input d,
  output reg q
  );

  parameter INI = 1'b0;

  tri0 gsrn = glbl.gsrn;

  always @(gsrn)
  begin
    if(!gsrn)
      assign q = INI;
    else
      deassign q;
  end

  always @(posedge reset or posedge set or posedge clk)
  begin
    if (reset)
      q <= 1'b0;
    else if (set)
      q <= 1'b1;
    else
      q <= d;
  end

endmodule

