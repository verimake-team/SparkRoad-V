// Verilog netlist created by TD v4.6.12906
// Tue Jul 30 09:10:06 2019

`timescale 1ns / 1ps
module test_camera  // sources/rtl/test_camera.v(14)
  (
  cam_data,
  cam_href,
  cam_pclk,
  cam_vsync,
  clk_24m,
  rst_n,
  cam_pwdn,
  cam_rst,
  cam_soic,
  cam_xclk,
  vga_b,
  vga_clk,
  vga_g,
  vga_hsync,
  vga_r,
  vga_vsync,
  cam_soid
  );

  input [7:0] cam_data;  // sources/rtl/test_camera.v(27)
  input cam_href;  // sources/rtl/test_camera.v(21)
  input cam_pclk;  // sources/rtl/test_camera.v(19)
  input cam_vsync;  // sources/rtl/test_camera.v(22)
  input clk_24m;  // sources/rtl/test_camera.v(16)
  input rst_n;  // sources/rtl/test_camera.v(17)
  output cam_pwdn;  // sources/rtl/test_camera.v(23)
  output cam_rst;  // sources/rtl/test_camera.v(24)
  output cam_soic;  // sources/rtl/test_camera.v(25)
  output cam_xclk;  // sources/rtl/test_camera.v(20)
  output [7:0] vga_b;  // sources/rtl/test_camera.v(31)
  output vga_clk;  // sources/rtl/test_camera.v(32)
  output [7:0] vga_g;  // sources/rtl/test_camera.v(30)
  output vga_hsync;  // sources/rtl/test_camera.v(33)
  output [7:0] vga_r;  // sources/rtl/test_camera.v(29)
  output vga_vsync;  // sources/rtl/test_camera.v(34)
  inout cam_soid;  // sources/rtl/test_camera.v(26)

  wire [7:0] cam_data_pad;  // sources/rtl/test_camera.v(27)
  wire [19:0] camera_addr;  // sources/rtl/test_camera.v(45)
  wire [15:0] camera_wrdat;  // sources/rtl/test_camera.v(44)
  wire [15:0] \u_camera_reader/current_pixel ;  // sources/rtl/camera_reader.v(37)
  wire [19:0] \u_camera_reader/n19 ;
  wire [19:0] \u_camera_reader/n21 ;
  wire [19:0] \u_camera_reader/n8 ;
  wire [19:0] \u_camera_reader/n9 ;
  wire [19:0] \u_camera_reader/pixel_counter ;  // sources/rtl/camera_reader.v(32)
  wire [7:0] \u_camera_reader/subpixel ;  // sources/rtl/camera_reader.v(36)
  wire [7:0] vga_b_pad;  // sources/rtl/test_camera.v(31)
  wire [7:0] vga_g_pad;  // sources/rtl/test_camera.v(30)
  wire [7:0] vga_r_pad;  // sources/rtl/test_camera.v(29)
  wire [15:0] vga_rdaddr;  // sources/rtl/test_camera.v(59)
  wire [0:6] vga_rdaddr_piped;
  wire [0:6] vga_rdaddr_piped_piped;
  wire _al_u430_o;
  wire _al_u440_o;
  wire _al_u487_o;
  wire _al_u488_o;
  wire _al_u489_o;
  wire _al_u491_o;
  wire _al_u492_o;
  wire _al_u493_o;
  wire _al_u494_o;
  wire _al_u495_o;
  wire _al_u496_o;
  wire _al_u497_o;
  wire _al_u498_o;
  wire _al_u499_o;
  wire _al_u500_o;
  wire _al_u501_o;
  wire _al_u502_o;
  wire _al_u503_o;
  wire _al_u504_o;
  wire _al_u505_o;
  wire _al_u506_o;
  wire _al_u507_o;
  wire _al_u508_o;
  wire _al_u509_o;
  wire _al_u510_o;
  wire _al_u511_o;
  wire _al_u512_o;
  wire _al_u513_o;
  wire _al_u514_o;
  wire _al_u515_o;
  wire _al_u516_o;
  wire _al_u517_o;
  wire _al_u519_o;
  wire _al_u520_o;
  wire _al_u521_o;
  wire _al_u522_o;
  wire _al_u523_o;
  wire _al_u524_o;
  wire _al_u525_o;
  wire _al_u526_o;
  wire _al_u527_o;
  wire _al_u528_o;
  wire _al_u529_o;
  wire _al_u530_o;
  wire _al_u531_o;
  wire _al_u532_o;
  wire _al_u533_o;
  wire _al_u534_o;
  wire _al_u535_o;
  wire _al_u536_o;
  wire _al_u537_o;
  wire _al_u538_o;
  wire _al_u539_o;
  wire _al_u540_o;
  wire _al_u541_o;
  wire _al_u542_o;
  wire _al_u543_o;
  wire _al_u544_o;
  wire _al_u545_o;
  wire _al_u547_o;
  wire _al_u548_o;
  wire _al_u549_o;
  wire _al_u550_o;
  wire _al_u551_o;
  wire _al_u552_o;
  wire _al_u553_o;
  wire _al_u554_o;
  wire _al_u555_o;
  wire _al_u556_o;
  wire _al_u557_o;
  wire _al_u558_o;
  wire _al_u559_o;
  wire _al_u560_o;
  wire _al_u561_o;
  wire _al_u562_o;
  wire _al_u563_o;
  wire _al_u564_o;
  wire _al_u565_o;
  wire _al_u566_o;
  wire _al_u567_o;
  wire _al_u568_o;
  wire _al_u569_o;
  wire _al_u570_o;
  wire _al_u571_o;
  wire _al_u572_o;
  wire _al_u573_o;
  wire _al_u575_o;
  wire _al_u576_o;
  wire _al_u577_o;
  wire _al_u578_o;
  wire _al_u579_o;
  wire _al_u580_o;
  wire _al_u581_o;
  wire _al_u582_o;
  wire _al_u583_o;
  wire _al_u584_o;
  wire _al_u585_o;
  wire _al_u586_o;
  wire _al_u587_o;
  wire _al_u588_o;
  wire _al_u589_o;
  wire _al_u590_o;
  wire _al_u591_o;
  wire _al_u592_o;
  wire _al_u593_o;
  wire _al_u594_o;
  wire _al_u595_o;
  wire _al_u596_o;
  wire _al_u597_o;
  wire _al_u598_o;
  wire _al_u599_o;
  wire _al_u600_o;
  wire _al_u601_o;
  wire _al_u603_o;
  wire _al_u604_o;
  wire _al_u605_o;
  wire _al_u606_o;
  wire _al_u607_o;
  wire _al_u608_o;
  wire _al_u609_o;
  wire _al_u610_o;
  wire _al_u611_o;
  wire _al_u612_o;
  wire _al_u613_o;
  wire _al_u614_o;
  wire _al_u615_o;
  wire _al_u616_o;
  wire _al_u617_o;
  wire _al_u618_o;
  wire _al_u619_o;
  wire _al_u620_o;
  wire _al_u621_o;
  wire _al_u622_o;
  wire _al_u623_o;
  wire _al_u624_o;
  wire _al_u625_o;
  wire _al_u626_o;
  wire _al_u627_o;
  wire _al_u628_o;
  wire _al_u629_o;
  wire _al_u631_o;
  wire _al_u632_o;
  wire _al_u633_o;
  wire _al_u634_o;
  wire _al_u635_o;
  wire _al_u636_o;
  wire _al_u637_o;
  wire _al_u638_o;
  wire _al_u639_o;
  wire _al_u640_o;
  wire _al_u641_o;
  wire _al_u642_o;
  wire _al_u643_o;
  wire _al_u644_o;
  wire _al_u645_o;
  wire _al_u646_o;
  wire _al_u647_o;
  wire _al_u648_o;
  wire _al_u649_o;
  wire _al_u650_o;
  wire _al_u651_o;
  wire _al_u652_o;
  wire _al_u653_o;
  wire _al_u654_o;
  wire _al_u655_o;
  wire _al_u656_o;
  wire _al_u657_o;
  wire _al_u659_o;
  wire _al_u660_o;
  wire _al_u661_o;
  wire _al_u662_o;
  wire _al_u663_o;
  wire _al_u664_o;
  wire _al_u665_o;
  wire _al_u666_o;
  wire _al_u667_o;
  wire _al_u668_o;
  wire _al_u669_o;
  wire _al_u670_o;
  wire _al_u671_o;
  wire _al_u672_o;
  wire _al_u673_o;
  wire _al_u674_o;
  wire _al_u675_o;
  wire _al_u676_o;
  wire _al_u677_o;
  wire _al_u678_o;
  wire _al_u679_o;
  wire _al_u680_o;
  wire _al_u681_o;
  wire _al_u682_o;
  wire _al_u683_o;
  wire _al_u684_o;
  wire _al_u685_o;
  wire _al_u687_o;
  wire _al_u688_o;
  wire _al_u689_o;
  wire _al_u691_o;
  wire _al_u692_o;
  wire _al_u693_o;
  wire _al_u695_o;
  wire _al_u696_o;
  wire _al_u697_o;
  wire _al_u699_o;
  wire _al_u700_o;
  wire _al_u701_o;
  wire _al_u703_o;
  wire _al_u704_o;
  wire _al_u705_o;
  wire _al_u707_o;
  wire _al_u708_o;
  wire _al_u709_o;
  wire _al_u711_o;
  wire _al_u712_o;
  wire _al_u713_o;
  wire _al_u714_o;
  wire _al_u715_o;
  wire _al_u716_o;
  wire _al_u717_o;
  wire _al_u718_o;
  wire _al_u719_o;
  wire _al_u720_o;
  wire _al_u721_o;
  wire _al_u722_o;
  wire _al_u723_o;
  wire _al_u724_o;
  wire _al_u725_o;
  wire _al_u726_o;
  wire _al_u727_o;
  wire _al_u728_o;
  wire _al_u729_o;
  wire _al_u730_o;
  wire _al_u731_o;
  wire _al_u732_o;
  wire _al_u733_o;
  wire _al_u734_o;
  wire _al_u735_o;
  wire _al_u736_o;
  wire _al_u737_o;
  wire _al_u739_o;
  wire _al_u740_o;
  wire _al_u741_o;
  wire _al_u742_o;
  wire _al_u743_o;
  wire _al_u744_o;
  wire _al_u745_o;
  wire _al_u746_o;
  wire _al_u747_o;
  wire _al_u748_o;
  wire _al_u749_o;
  wire _al_u750_o;
  wire _al_u751_o;
  wire _al_u752_o;
  wire _al_u753_o;
  wire _al_u754_o;
  wire _al_u755_o;
  wire _al_u756_o;
  wire _al_u757_o;
  wire _al_u758_o;
  wire _al_u759_o;
  wire _al_u760_o;
  wire _al_u761_o;
  wire _al_u762_o;
  wire _al_u763_o;
  wire _al_u764_o;
  wire _al_u765_o;
  wire \and_Ncamera_addr[11]_o_and_camera_wrreq ;
  wire \and_Ncamera_addr[12]_o ;
  wire \and_Ncamera_addr[12]_o_al_n177 ;
  wire \and_Ncamera_addr[12]_o_al_n208 ;
  wire \and_Ncamera_addr[12]_o_al_n240 ;
  wire \and_Nvga_rdaddr[11]__o_and_vga_rden ;
  wire \and_Nvga_rdaddr[12]__o ;
  wire \and_Nvga_rdaddr[12]__o_al_n180 ;
  wire \and_Nvga_rdaddr[12]__o_al_n211 ;
  wire \and_Nvga_rdaddr[12]__o_al_n243 ;
  wire \and_camera_addr[12]__o ;
  wire \and_camera_addr[12]__o_al_n193 ;
  wire \and_camera_addr[12]__o_al_n224 ;
  wire \and_camera_addr[12]__o_al_n256 ;
  wire \and_vga_rdaddr[12]_N_o ;
  wire \and_vga_rdaddr[12]_N_o_al_n227 ;
  wire \and_vga_rdaddr[12]_v_o ;
  wire \and_vga_rdaddr[12]_v_o_al_n259 ;
  wire cam_pclk_pad;  // sources/rtl/test_camera.v(19)
  wire cam_rst_pad;  // sources/rtl/test_camera.v(24)
  wire cam_rst_pad_neg;
  wire cam_soid_pad;  // sources/rtl/test_camera.v(26)
  wire cam_vsync_pad;  // sources/rtl/test_camera.v(22)
  wire cam_xclk_pad;  // sources/rtl/test_camera.v(20)
  wire camera_wrreq;  // sources/rtl/test_camera.v(42)
  wire clk_24m_pad;  // sources/rtl/test_camera.v(16)
  wire clk_cam;  // sources/rtl/test_camera.v(39)
  wire clk_lcd;  // sources/rtl/test_camera.v(38)
  wire clk_sccb;  // sources/rtl/test_camera.v(40)
  wire sda;  // sources/rtl/test_camera.v(50)
  wire sda_oe;  // sources/rtl/test_camera.v(49)
  wire \u_camera_reader/add0/c0 ;
  wire \u_camera_reader/add0/c1 ;
  wire \u_camera_reader/add0/c10 ;
  wire \u_camera_reader/add0/c11 ;
  wire \u_camera_reader/add0/c12 ;
  wire \u_camera_reader/add0/c13 ;
  wire \u_camera_reader/add0/c14 ;
  wire \u_camera_reader/add0/c15 ;
  wire \u_camera_reader/add0/c16 ;
  wire \u_camera_reader/add0/c17 ;
  wire \u_camera_reader/add0/c18 ;
  wire \u_camera_reader/add0/c19 ;
  wire \u_camera_reader/add0/c2 ;
  wire \u_camera_reader/add0/c3 ;
  wire \u_camera_reader/add0/c4 ;
  wire \u_camera_reader/add0/c5 ;
  wire \u_camera_reader/add0/c6 ;
  wire \u_camera_reader/add0/c7 ;
  wire \u_camera_reader/add0/c8 ;
  wire \u_camera_reader/add0/c9 ;
  wire \u_camera_reader/add1/c0 ;
  wire \u_camera_reader/add1/c1 ;
  wire \u_camera_reader/add1/c10 ;
  wire \u_camera_reader/add1/c11 ;
  wire \u_camera_reader/add1/c12 ;
  wire \u_camera_reader/add1/c13 ;
  wire \u_camera_reader/add1/c14 ;
  wire \u_camera_reader/add1/c15 ;
  wire \u_camera_reader/add1/c2 ;
  wire \u_camera_reader/add1/c3 ;
  wire \u_camera_reader/add1/c4 ;
  wire \u_camera_reader/add1/c5 ;
  wire \u_camera_reader/add1/c6 ;
  wire \u_camera_reader/add1/c7 ;
  wire \u_camera_reader/add1/c8 ;
  wire \u_camera_reader/add1/c9 ;
  wire \u_camera_reader/lt0_c0 ;
  wire \u_camera_reader/lt0_c1 ;
  wire \u_camera_reader/lt0_c10 ;
  wire \u_camera_reader/lt0_c11 ;
  wire \u_camera_reader/lt0_c12 ;
  wire \u_camera_reader/lt0_c13 ;
  wire \u_camera_reader/lt0_c14 ;
  wire \u_camera_reader/lt0_c15 ;
  wire \u_camera_reader/lt0_c16 ;
  wire \u_camera_reader/lt0_c17 ;
  wire \u_camera_reader/lt0_c18 ;
  wire \u_camera_reader/lt0_c19 ;
  wire \u_camera_reader/lt0_c2 ;
  wire \u_camera_reader/lt0_c20 ;
  wire \u_camera_reader/lt0_c3 ;
  wire \u_camera_reader/lt0_c4 ;
  wire \u_camera_reader/lt0_c5 ;
  wire \u_camera_reader/lt0_c6 ;
  wire \u_camera_reader/lt0_c7 ;
  wire \u_camera_reader/lt0_c8 ;
  wire \u_camera_reader/lt0_c9 ;
  wire \u_camera_reader/mux13_b0_sel_is_2_o ;
  wire \u_camera_reader/mux14_b0_sel_is_2_o ;
  wire \u_camera_reader/mux5_b0_sel_is_3_o ;
  wire \u_camera_reader/mux6_b0_sel_is_1_o ;
  wire \u_camera_reader/mux8_b0_sel_is_0_o ;
  wire \u_camera_reader/n1 ;
  wire \u_camera_reader/n2 ;
  wire \u_camera_reader/n27 ;
  wire \u_camera_reader/vsync_passed ;  // sources/rtl/camera_reader.v(34)
  wire \u_camera_reader/vsync_passed_d ;
  wire \u_camera_reader/wrclk1 ;  // sources/rtl/camera_reader.v(38)
  wire \u_camera_reader/write_pixel ;  // sources/rtl/camera_reader.v(35)
  wire \u_img/inst_dob_i0_000 ;
  wire \u_img/inst_dob_i0_001 ;
  wire \u_img/inst_dob_i0_002 ;
  wire \u_img/inst_dob_i0_003 ;
  wire \u_img/inst_dob_i0_004 ;
  wire \u_img/inst_dob_i0_005 ;
  wire \u_img/inst_dob_i0_006 ;
  wire \u_img/inst_dob_i0_007 ;
  wire \u_img/inst_dob_i0_008 ;
  wire \u_img/inst_dob_i0_009 ;
  wire \u_img/inst_dob_i0_010 ;
  wire \u_img/inst_dob_i0_011 ;
  wire \u_img/inst_dob_i0_012 ;
  wire \u_img/inst_dob_i0_013 ;
  wire \u_img/inst_dob_i0_014 ;
  wire \u_img/inst_dob_i0_015 ;
  wire \u_img/inst_dob_i10_000 ;
  wire \u_img/inst_dob_i10_001 ;
  wire \u_img/inst_dob_i10_002 ;
  wire \u_img/inst_dob_i10_003 ;
  wire \u_img/inst_dob_i10_004 ;
  wire \u_img/inst_dob_i10_005 ;
  wire \u_img/inst_dob_i10_006 ;
  wire \u_img/inst_dob_i10_007 ;
  wire \u_img/inst_dob_i10_008 ;
  wire \u_img/inst_dob_i12_000 ;
  wire \u_img/inst_dob_i12_001 ;
  wire \u_img/inst_dob_i12_002 ;
  wire \u_img/inst_dob_i12_003 ;
  wire \u_img/inst_dob_i12_004 ;
  wire \u_img/inst_dob_i12_005 ;
  wire \u_img/inst_dob_i12_006 ;
  wire \u_img/inst_dob_i12_007 ;
  wire \u_img/inst_dob_i12_008 ;
  wire \u_img/inst_dob_i14_000 ;
  wire \u_img/inst_dob_i14_001 ;
  wire \u_img/inst_dob_i14_002 ;
  wire \u_img/inst_dob_i14_003 ;
  wire \u_img/inst_dob_i14_004 ;
  wire \u_img/inst_dob_i14_005 ;
  wire \u_img/inst_dob_i14_006 ;
  wire \u_img/inst_dob_i14_007 ;
  wire \u_img/inst_dob_i14_008 ;
  wire \u_img/inst_dob_i16_000 ;
  wire \u_img/inst_dob_i16_001 ;
  wire \u_img/inst_dob_i16_002 ;
  wire \u_img/inst_dob_i16_003 ;
  wire \u_img/inst_dob_i16_004 ;
  wire \u_img/inst_dob_i16_005 ;
  wire \u_img/inst_dob_i16_006 ;
  wire \u_img/inst_dob_i16_007 ;
  wire \u_img/inst_dob_i16_008 ;
  wire \u_img/inst_dob_i16_009 ;
  wire \u_img/inst_dob_i16_010 ;
  wire \u_img/inst_dob_i16_011 ;
  wire \u_img/inst_dob_i16_012 ;
  wire \u_img/inst_dob_i16_013 ;
  wire \u_img/inst_dob_i16_014 ;
  wire \u_img/inst_dob_i16_015 ;
  wire \u_img/inst_dob_i18_000 ;
  wire \u_img/inst_dob_i18_001 ;
  wire \u_img/inst_dob_i18_002 ;
  wire \u_img/inst_dob_i18_003 ;
  wire \u_img/inst_dob_i18_004 ;
  wire \u_img/inst_dob_i18_005 ;
  wire \u_img/inst_dob_i18_006 ;
  wire \u_img/inst_dob_i18_007 ;
  wire \u_img/inst_dob_i18_008 ;
  wire \u_img/inst_dob_i20_000 ;
  wire \u_img/inst_dob_i20_001 ;
  wire \u_img/inst_dob_i20_002 ;
  wire \u_img/inst_dob_i20_003 ;
  wire \u_img/inst_dob_i20_004 ;
  wire \u_img/inst_dob_i20_005 ;
  wire \u_img/inst_dob_i20_006 ;
  wire \u_img/inst_dob_i20_007 ;
  wire \u_img/inst_dob_i20_008 ;
  wire \u_img/inst_dob_i22_000 ;
  wire \u_img/inst_dob_i22_001 ;
  wire \u_img/inst_dob_i22_002 ;
  wire \u_img/inst_dob_i22_003 ;
  wire \u_img/inst_dob_i22_004 ;
  wire \u_img/inst_dob_i22_005 ;
  wire \u_img/inst_dob_i22_006 ;
  wire \u_img/inst_dob_i22_007 ;
  wire \u_img/inst_dob_i22_008 ;
  wire \u_img/inst_dob_i24_000 ;
  wire \u_img/inst_dob_i24_001 ;
  wire \u_img/inst_dob_i24_002 ;
  wire \u_img/inst_dob_i24_003 ;
  wire \u_img/inst_dob_i24_004 ;
  wire \u_img/inst_dob_i24_005 ;
  wire \u_img/inst_dob_i24_006 ;
  wire \u_img/inst_dob_i24_007 ;
  wire \u_img/inst_dob_i24_008 ;
  wire \u_img/inst_dob_i26_000 ;
  wire \u_img/inst_dob_i26_001 ;
  wire \u_img/inst_dob_i26_002 ;
  wire \u_img/inst_dob_i26_003 ;
  wire \u_img/inst_dob_i26_004 ;
  wire \u_img/inst_dob_i26_005 ;
  wire \u_img/inst_dob_i26_006 ;
  wire \u_img/inst_dob_i26_007 ;
  wire \u_img/inst_dob_i26_008 ;
  wire \u_img/inst_dob_i28_000 ;
  wire \u_img/inst_dob_i28_001 ;
  wire \u_img/inst_dob_i28_002 ;
  wire \u_img/inst_dob_i28_003 ;
  wire \u_img/inst_dob_i28_004 ;
  wire \u_img/inst_dob_i28_005 ;
  wire \u_img/inst_dob_i28_006 ;
  wire \u_img/inst_dob_i28_007 ;
  wire \u_img/inst_dob_i28_008 ;
  wire \u_img/inst_dob_i2_000 ;
  wire \u_img/inst_dob_i2_001 ;
  wire \u_img/inst_dob_i2_002 ;
  wire \u_img/inst_dob_i2_003 ;
  wire \u_img/inst_dob_i2_004 ;
  wire \u_img/inst_dob_i2_005 ;
  wire \u_img/inst_dob_i2_006 ;
  wire \u_img/inst_dob_i2_007 ;
  wire \u_img/inst_dob_i2_008 ;
  wire \u_img/inst_dob_i30_000 ;
  wire \u_img/inst_dob_i30_001 ;
  wire \u_img/inst_dob_i30_002 ;
  wire \u_img/inst_dob_i30_003 ;
  wire \u_img/inst_dob_i30_004 ;
  wire \u_img/inst_dob_i30_005 ;
  wire \u_img/inst_dob_i30_006 ;
  wire \u_img/inst_dob_i30_007 ;
  wire \u_img/inst_dob_i30_008 ;
  wire \u_img/inst_dob_i32_000 ;
  wire \u_img/inst_dob_i32_001 ;
  wire \u_img/inst_dob_i32_002 ;
  wire \u_img/inst_dob_i32_003 ;
  wire \u_img/inst_dob_i32_004 ;
  wire \u_img/inst_dob_i32_005 ;
  wire \u_img/inst_dob_i32_006 ;
  wire \u_img/inst_dob_i32_007 ;
  wire \u_img/inst_dob_i32_008 ;
  wire \u_img/inst_dob_i32_009 ;
  wire \u_img/inst_dob_i32_010 ;
  wire \u_img/inst_dob_i32_011 ;
  wire \u_img/inst_dob_i32_012 ;
  wire \u_img/inst_dob_i32_013 ;
  wire \u_img/inst_dob_i32_014 ;
  wire \u_img/inst_dob_i32_015 ;
  wire \u_img/inst_dob_i34_000 ;
  wire \u_img/inst_dob_i34_001 ;
  wire \u_img/inst_dob_i34_002 ;
  wire \u_img/inst_dob_i34_003 ;
  wire \u_img/inst_dob_i34_004 ;
  wire \u_img/inst_dob_i34_005 ;
  wire \u_img/inst_dob_i34_006 ;
  wire \u_img/inst_dob_i34_007 ;
  wire \u_img/inst_dob_i34_008 ;
  wire \u_img/inst_dob_i36_000 ;
  wire \u_img/inst_dob_i36_001 ;
  wire \u_img/inst_dob_i36_002 ;
  wire \u_img/inst_dob_i36_003 ;
  wire \u_img/inst_dob_i36_004 ;
  wire \u_img/inst_dob_i36_005 ;
  wire \u_img/inst_dob_i36_006 ;
  wire \u_img/inst_dob_i36_007 ;
  wire \u_img/inst_dob_i36_008 ;
  wire \u_img/inst_dob_i38_000 ;
  wire \u_img/inst_dob_i38_001 ;
  wire \u_img/inst_dob_i38_002 ;
  wire \u_img/inst_dob_i38_003 ;
  wire \u_img/inst_dob_i38_004 ;
  wire \u_img/inst_dob_i38_005 ;
  wire \u_img/inst_dob_i38_006 ;
  wire \u_img/inst_dob_i38_007 ;
  wire \u_img/inst_dob_i38_008 ;
  wire \u_img/inst_dob_i40_000 ;
  wire \u_img/inst_dob_i40_001 ;
  wire \u_img/inst_dob_i40_002 ;
  wire \u_img/inst_dob_i40_003 ;
  wire \u_img/inst_dob_i40_004 ;
  wire \u_img/inst_dob_i40_005 ;
  wire \u_img/inst_dob_i40_006 ;
  wire \u_img/inst_dob_i40_007 ;
  wire \u_img/inst_dob_i40_008 ;
  wire \u_img/inst_dob_i42_000 ;
  wire \u_img/inst_dob_i42_001 ;
  wire \u_img/inst_dob_i42_002 ;
  wire \u_img/inst_dob_i42_003 ;
  wire \u_img/inst_dob_i42_004 ;
  wire \u_img/inst_dob_i42_005 ;
  wire \u_img/inst_dob_i42_006 ;
  wire \u_img/inst_dob_i42_007 ;
  wire \u_img/inst_dob_i42_008 ;
  wire \u_img/inst_dob_i44_000 ;
  wire \u_img/inst_dob_i44_001 ;
  wire \u_img/inst_dob_i44_002 ;
  wire \u_img/inst_dob_i44_003 ;
  wire \u_img/inst_dob_i44_004 ;
  wire \u_img/inst_dob_i44_005 ;
  wire \u_img/inst_dob_i44_006 ;
  wire \u_img/inst_dob_i44_007 ;
  wire \u_img/inst_dob_i44_008 ;
  wire \u_img/inst_dob_i46_000 ;
  wire \u_img/inst_dob_i46_001 ;
  wire \u_img/inst_dob_i46_002 ;
  wire \u_img/inst_dob_i46_003 ;
  wire \u_img/inst_dob_i46_004 ;
  wire \u_img/inst_dob_i46_005 ;
  wire \u_img/inst_dob_i46_006 ;
  wire \u_img/inst_dob_i46_007 ;
  wire \u_img/inst_dob_i46_008 ;
  wire \u_img/inst_dob_i48_000 ;
  wire \u_img/inst_dob_i48_001 ;
  wire \u_img/inst_dob_i48_002 ;
  wire \u_img/inst_dob_i48_003 ;
  wire \u_img/inst_dob_i48_004 ;
  wire \u_img/inst_dob_i48_005 ;
  wire \u_img/inst_dob_i48_006 ;
  wire \u_img/inst_dob_i48_007 ;
  wire \u_img/inst_dob_i48_008 ;
  wire \u_img/inst_dob_i48_009 ;
  wire \u_img/inst_dob_i48_010 ;
  wire \u_img/inst_dob_i48_011 ;
  wire \u_img/inst_dob_i48_012 ;
  wire \u_img/inst_dob_i48_013 ;
  wire \u_img/inst_dob_i48_014 ;
  wire \u_img/inst_dob_i48_015 ;
  wire \u_img/inst_dob_i4_000 ;
  wire \u_img/inst_dob_i4_001 ;
  wire \u_img/inst_dob_i4_002 ;
  wire \u_img/inst_dob_i4_003 ;
  wire \u_img/inst_dob_i4_004 ;
  wire \u_img/inst_dob_i4_005 ;
  wire \u_img/inst_dob_i4_006 ;
  wire \u_img/inst_dob_i4_007 ;
  wire \u_img/inst_dob_i4_008 ;
  wire \u_img/inst_dob_i50_000 ;
  wire \u_img/inst_dob_i50_001 ;
  wire \u_img/inst_dob_i50_002 ;
  wire \u_img/inst_dob_i50_003 ;
  wire \u_img/inst_dob_i50_004 ;
  wire \u_img/inst_dob_i50_005 ;
  wire \u_img/inst_dob_i50_006 ;
  wire \u_img/inst_dob_i50_007 ;
  wire \u_img/inst_dob_i50_008 ;
  wire \u_img/inst_dob_i52_000 ;
  wire \u_img/inst_dob_i52_001 ;
  wire \u_img/inst_dob_i52_002 ;
  wire \u_img/inst_dob_i52_003 ;
  wire \u_img/inst_dob_i52_004 ;
  wire \u_img/inst_dob_i52_005 ;
  wire \u_img/inst_dob_i52_006 ;
  wire \u_img/inst_dob_i52_007 ;
  wire \u_img/inst_dob_i52_008 ;
  wire \u_img/inst_dob_i54_000 ;
  wire \u_img/inst_dob_i54_001 ;
  wire \u_img/inst_dob_i54_002 ;
  wire \u_img/inst_dob_i54_003 ;
  wire \u_img/inst_dob_i54_004 ;
  wire \u_img/inst_dob_i54_005 ;
  wire \u_img/inst_dob_i54_006 ;
  wire \u_img/inst_dob_i54_007 ;
  wire \u_img/inst_dob_i54_008 ;
  wire \u_img/inst_dob_i56_000 ;
  wire \u_img/inst_dob_i56_001 ;
  wire \u_img/inst_dob_i56_002 ;
  wire \u_img/inst_dob_i56_003 ;
  wire \u_img/inst_dob_i56_004 ;
  wire \u_img/inst_dob_i56_005 ;
  wire \u_img/inst_dob_i56_006 ;
  wire \u_img/inst_dob_i56_007 ;
  wire \u_img/inst_dob_i56_008 ;
  wire \u_img/inst_dob_i58_000 ;
  wire \u_img/inst_dob_i58_001 ;
  wire \u_img/inst_dob_i58_002 ;
  wire \u_img/inst_dob_i58_003 ;
  wire \u_img/inst_dob_i58_004 ;
  wire \u_img/inst_dob_i58_005 ;
  wire \u_img/inst_dob_i58_006 ;
  wire \u_img/inst_dob_i58_007 ;
  wire \u_img/inst_dob_i58_008 ;
  wire \u_img/inst_dob_i60_000 ;
  wire \u_img/inst_dob_i60_001 ;
  wire \u_img/inst_dob_i60_002 ;
  wire \u_img/inst_dob_i60_003 ;
  wire \u_img/inst_dob_i60_004 ;
  wire \u_img/inst_dob_i60_005 ;
  wire \u_img/inst_dob_i60_006 ;
  wire \u_img/inst_dob_i60_007 ;
  wire \u_img/inst_dob_i60_008 ;
  wire \u_img/inst_dob_i62_000 ;
  wire \u_img/inst_dob_i62_001 ;
  wire \u_img/inst_dob_i62_002 ;
  wire \u_img/inst_dob_i62_003 ;
  wire \u_img/inst_dob_i62_004 ;
  wire \u_img/inst_dob_i62_005 ;
  wire \u_img/inst_dob_i62_006 ;
  wire \u_img/inst_dob_i62_007 ;
  wire \u_img/inst_dob_i62_008 ;
  wire \u_img/inst_dob_i64_000 ;
  wire \u_img/inst_dob_i64_001 ;
  wire \u_img/inst_dob_i64_002 ;
  wire \u_img/inst_dob_i64_003 ;
  wire \u_img/inst_dob_i64_004 ;
  wire \u_img/inst_dob_i64_005 ;
  wire \u_img/inst_dob_i64_006 ;
  wire \u_img/inst_dob_i64_007 ;
  wire \u_img/inst_dob_i64_008 ;
  wire \u_img/inst_dob_i64_009 ;
  wire \u_img/inst_dob_i64_010 ;
  wire \u_img/inst_dob_i64_011 ;
  wire \u_img/inst_dob_i64_012 ;
  wire \u_img/inst_dob_i64_013 ;
  wire \u_img/inst_dob_i64_014 ;
  wire \u_img/inst_dob_i64_015 ;
  wire \u_img/inst_dob_i6_000 ;
  wire \u_img/inst_dob_i6_001 ;
  wire \u_img/inst_dob_i6_002 ;
  wire \u_img/inst_dob_i6_003 ;
  wire \u_img/inst_dob_i6_004 ;
  wire \u_img/inst_dob_i6_005 ;
  wire \u_img/inst_dob_i6_006 ;
  wire \u_img/inst_dob_i6_007 ;
  wire \u_img/inst_dob_i6_008 ;
  wire \u_img/inst_dob_i8_000 ;
  wire \u_img/inst_dob_i8_001 ;
  wire \u_img/inst_dob_i8_002 ;
  wire \u_img/inst_dob_i8_003 ;
  wire \u_img/inst_dob_i8_004 ;
  wire \u_img/inst_dob_i8_005 ;
  wire \u_img/inst_dob_i8_006 ;
  wire \u_img/inst_dob_i8_007 ;
  wire \u_img/inst_dob_i8_008 ;
  wire \u_pll/clk0_buf ;  // al_ip/ip_pll.v(34)
  wire vga_clk_pad;  // sources/rtl/test_camera.v(32)
  wire vga_hsync_pad;  // sources/rtl/test_camera.v(33)
  wire vga_rden;  // sources/rtl/test_camera.v(57)
  wire vga_vsync_pad;  // sources/rtl/test_camera.v(34)

  EG_PHY_PAD #(
    //.LOCATION("H13"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS33"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u151 (
    .ipad(cam_data[7]),
    .di(cam_data_pad[7]));  // sources/rtl/test_camera.v(27)
  EG_PHY_PAD #(
    //.LOCATION("G16"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS33"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u152 (
    .ipad(cam_data[6]),
    .di(cam_data_pad[6]));  // sources/rtl/test_camera.v(27)
  EG_PHY_PAD #(
    //.LOCATION("H16"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS33"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u153 (
    .ipad(cam_data[5]),
    .di(cam_data_pad[5]));  // sources/rtl/test_camera.v(27)
  EG_PHY_PAD #(
    //.LOCATION("G14"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS33"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u154 (
    .ipad(cam_data[4]),
    .di(cam_data_pad[4]));  // sources/rtl/test_camera.v(27)
  EG_PHY_PAD #(
    //.LOCATION("K15"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS33"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u155 (
    .ipad(cam_data[3]),
    .di(cam_data_pad[3]));  // sources/rtl/test_camera.v(27)
  EG_PHY_PAD #(
    //.LOCATION("K16"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS33"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u156 (
    .ipad(cam_data[2]),
    .di(cam_data_pad[2]));  // sources/rtl/test_camera.v(27)
  EG_PHY_PAD #(
    //.LOCATION("J16"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS33"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u157 (
    .ipad(cam_data[1]),
    .di(cam_data_pad[1]));  // sources/rtl/test_camera.v(27)
  EG_PHY_PAD #(
    //.LOCATION("H15"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS33"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u158 (
    .ipad(cam_data[0]),
    .di(cam_data_pad[0]));  // sources/rtl/test_camera.v(27)
  EG_PHY_PAD #(
    //.LOCATION("F15"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u159 (
    .ipad(cam_href),
    .di(\u_camera_reader/n2 ));  // sources/rtl/test_camera.v(21)
  EG_PHY_PAD #(
    //.LOCATION("K12"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u160 (
    .ipad(cam_pclk),
    .di(cam_pclk_pad));  // sources/rtl/test_camera.v(19)
  EG_PHY_PAD #(
    //.LOCATION("F14"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u161 (
    .do({open_n171,open_n172,open_n173,1'b0}),
    .opad(cam_pwdn));  // sources/rtl/test_camera.v(23)
  EG_PHY_PAD #(
    //.LOCATION("F13"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u162 (
    .do({open_n188,open_n189,open_n190,cam_rst_pad}),
    .opad(cam_rst));  // sources/rtl/test_camera.v(24)
  EG_PHY_PAD #(
    //.LOCATION("D14"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("BI"),
    .TSMUX("INV"))
    _al_u163 (
    .do({open_n205,open_n206,open_n207,sda}),
    .ts(sda_oe),
    .di(cam_soid_pad),
    .bpad(cam_soid));  // sources/rtl/test_camera.v(61)
  EG_PHY_PAD #(
    //.LOCATION("E15"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u164 (
    .ipad(cam_vsync),
    .di(cam_vsync_pad));  // sources/rtl/test_camera.v(22)
  EG_PHY_PAD #(
    //.LOCATION("J12"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u165 (
    .do({open_n237,open_n238,open_n239,cam_xclk_pad}),
    .opad(cam_xclk));  // sources/rtl/test_camera.v(20)
  EG_PHY_PAD #(
    //.LOCATION("K14"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u166 (
    .ipad(clk_24m),
    .di(clk_24m_pad));  // sources/rtl/test_camera.v(16)
  EG_PHY_PAD #(
    //.LOCATION("G11"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u167 (
    .ipad(rst_n),
    .di(cam_rst_pad));  // sources/rtl/test_camera.v(17)
  EG_PHY_PAD #(
    //.LOCATION("C1"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("FAST"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u168 (
    .do({open_n288,open_n289,open_n290,vga_b_pad[7]}),
    .opad(vga_b[7]));  // sources/rtl/test_camera.v(31)
  EG_PHY_PAD #(
    //.LOCATION("D1"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("FAST"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u169 (
    .do({open_n305,open_n306,open_n307,vga_b_pad[6]}),
    .opad(vga_b[6]));  // sources/rtl/test_camera.v(31)
  EG_PHY_PAD #(
    //.LOCATION("E2"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("FAST"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u170 (
    .do({open_n322,open_n323,open_n324,vga_b_pad[5]}),
    .opad(vga_b[5]));  // sources/rtl/test_camera.v(31)
  EG_PHY_PAD #(
    //.LOCATION("G3"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("FAST"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u171 (
    .do({open_n339,open_n340,open_n341,vga_b_pad[4]}),
    .opad(vga_b[4]));  // sources/rtl/test_camera.v(31)
  EG_PHY_PAD #(
    //.LOCATION("E1"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("FAST"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u172 (
    .do({open_n356,open_n357,open_n358,vga_b_pad[3]}),
    .opad(vga_b[3]));  // sources/rtl/test_camera.v(31)
  EG_PHY_PAD #(
    //.LOCATION("F2"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("FAST"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u173 (
    .do({open_n373,open_n374,open_n375,1'b0}),
    .opad(vga_b[2]));  // sources/rtl/test_camera.v(31)
  EG_PHY_PAD #(
    //.LOCATION("F1"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("FAST"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u174 (
    .do({open_n390,open_n391,open_n392,1'b0}),
    .opad(vga_b[1]));  // sources/rtl/test_camera.v(31)
  EG_PHY_PAD #(
    //.LOCATION("G1"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("FAST"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u175 (
    .do({open_n407,open_n408,open_n409,1'b0}),
    .opad(vga_b[0]));  // sources/rtl/test_camera.v(31)
  EG_PHY_PAD #(
    //.LOCATION("H2"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u176 (
    .do({open_n424,open_n425,open_n426,vga_clk_pad}),
    .opad(vga_clk));  // sources/rtl/test_camera.v(32)
  EG_PHY_PAD #(
    //.LOCATION("H5"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u177 (
    .do({open_n441,open_n442,open_n443,vga_g_pad[7]}),
    .opad(vga_g[7]));  // sources/rtl/test_camera.v(30)
  EG_PHY_PAD #(
    //.LOCATION("H1"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u178 (
    .do({open_n458,open_n459,open_n460,vga_g_pad[6]}),
    .opad(vga_g[6]));  // sources/rtl/test_camera.v(30)
  EG_PHY_PAD #(
    //.LOCATION("J6"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u179 (
    .do({open_n475,open_n476,open_n477,vga_g_pad[5]}),
    .opad(vga_g[5]));  // sources/rtl/test_camera.v(30)
  EG_PHY_PAD #(
    //.LOCATION("H3"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u180 (
    .do({open_n492,open_n493,open_n494,vga_g_pad[4]}),
    .opad(vga_g[4]));  // sources/rtl/test_camera.v(30)
  EG_PHY_PAD #(
    //.LOCATION("J1"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u181 (
    .do({open_n509,open_n510,open_n511,vga_g_pad[3]}),
    .opad(vga_g[3]));  // sources/rtl/test_camera.v(30)
  EG_PHY_PAD #(
    //.LOCATION("K1"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u182 (
    .do({open_n526,open_n527,open_n528,vga_g_pad[2]}),
    .opad(vga_g[2]));  // sources/rtl/test_camera.v(30)
  EG_PHY_PAD #(
    //.LOCATION("K2"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u183 (
    .do({open_n543,open_n544,open_n545,1'b0}),
    .opad(vga_g[1]));  // sources/rtl/test_camera.v(30)
  EG_PHY_PAD #(
    //.LOCATION("L1"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u184 (
    .do({open_n560,open_n561,open_n562,1'b0}),
    .opad(vga_g[0]));  // sources/rtl/test_camera.v(30)
  EG_PHY_PAD #(
    //.LOCATION("J3"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u185 (
    .do({open_n577,open_n578,open_n579,vga_hsync_pad}),
    .opad(vga_hsync));  // sources/rtl/test_camera.v(33)
  EG_PHY_PAD #(
    //.LOCATION("L5"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u186 (
    .do({open_n594,open_n595,open_n596,vga_r_pad[7]}),
    .opad(vga_r[7]));  // sources/rtl/test_camera.v(29)
  EG_PHY_PAD #(
    //.LOCATION("L3"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u187 (
    .do({open_n611,open_n612,open_n613,vga_r_pad[6]}),
    .opad(vga_r[6]));  // sources/rtl/test_camera.v(29)
  EG_PHY_PAD #(
    //.LOCATION("M2"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u188 (
    .do({open_n628,open_n629,open_n630,vga_r_pad[5]}),
    .opad(vga_r[5]));  // sources/rtl/test_camera.v(29)
  EG_PHY_PAD #(
    //.LOCATION("M1"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u189 (
    .do({open_n645,open_n646,open_n647,vga_r_pad[4]}),
    .opad(vga_r[4]));  // sources/rtl/test_camera.v(29)
  EG_PHY_PAD #(
    //.LOCATION("L4"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u190 (
    .do({open_n662,open_n663,open_n664,vga_r_pad[3]}),
    .opad(vga_r[3]));  // sources/rtl/test_camera.v(29)
  EG_PHY_PAD #(
    //.LOCATION("K5"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u191 (
    .do({open_n679,open_n680,open_n681,1'b0}),
    .opad(vga_r[2]));  // sources/rtl/test_camera.v(29)
  EG_PHY_PAD #(
    //.LOCATION("K3"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u192 (
    .do({open_n696,open_n697,open_n698,1'b0}),
    .opad(vga_r[1]));  // sources/rtl/test_camera.v(29)
  EG_PHY_PAD #(
    //.LOCATION("K6"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u193 (
    .do({open_n713,open_n714,open_n715,1'b0}),
    .opad(vga_r[0]));  // sources/rtl/test_camera.v(29)
  EG_PHY_PAD #(
    //.LOCATION("J4"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u194 (
    .do({open_n730,open_n731,open_n732,vga_vsync_pad}),
    .opad(vga_vsync));  // sources/rtl/test_camera.v(34)
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*A)"),
    .INIT(16'h0080))
    _al_u423 (
    .a(camera_addr[12]),
    .b(camera_addr[13]),
    .c(camera_addr[14]),
    .d(camera_addr[15]),
    .o(\and_camera_addr[12]__o_al_n256 ));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*~B*A)"),
    .INIT(16'h0020))
    _al_u424 (
    .a(camera_addr[12]),
    .b(camera_addr[13]),
    .c(camera_addr[14]),
    .d(camera_addr[15]),
    .o(\and_camera_addr[12]__o_al_n224 ));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    _al_u425 (
    .a(camera_addr[12]),
    .b(camera_addr[13]),
    .c(camera_addr[14]),
    .d(camera_addr[15]),
    .o(\and_camera_addr[12]__o_al_n193 ));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*A)"),
    .INIT(16'h0002))
    _al_u426 (
    .a(camera_addr[12]),
    .b(camera_addr[13]),
    .c(camera_addr[14]),
    .d(camera_addr[15]),
    .o(\and_camera_addr[12]__o ));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*~A)"),
    .INIT(16'h0040))
    _al_u427 (
    .a(camera_addr[12]),
    .b(camera_addr[13]),
    .c(camera_addr[14]),
    .d(camera_addr[15]),
    .o(\and_Ncamera_addr[12]_o_al_n240 ));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*~B*~A)"),
    .INIT(16'h0010))
    _al_u428 (
    .a(camera_addr[12]),
    .b(camera_addr[13]),
    .c(camera_addr[14]),
    .d(camera_addr[15]),
    .o(\and_Ncamera_addr[12]_o_al_n208 ));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*~A)"),
    .INIT(16'h0004))
    _al_u429 (
    .a(camera_addr[12]),
    .b(camera_addr[13]),
    .c(camera_addr[14]),
    .d(camera_addr[15]),
    .o(\and_Ncamera_addr[12]_o_al_n177 ));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u430 (
    .a(camera_addr[12]),
    .b(camera_addr[13]),
    .c(camera_addr[14]),
    .o(_al_u430_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u431 (
    .a(_al_u430_o),
    .b(camera_addr[15]),
    .o(\and_Ncamera_addr[12]_o ));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*~A)"),
    .INIT(16'h4000))
    _al_u432 (
    .a(vga_rdaddr[15]),
    .b(vga_rdaddr[14]),
    .c(vga_rdaddr[13]),
    .d(vga_rdaddr[12]),
    .o(\and_vga_rdaddr[12]_v_o_al_n259 ));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*~A)"),
    .INIT(16'h1000))
    _al_u433 (
    .a(vga_rdaddr[15]),
    .b(vga_rdaddr[14]),
    .c(vga_rdaddr[13]),
    .d(vga_rdaddr[12]),
    .o(\and_vga_rdaddr[12]_v_o ));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*B*~A)"),
    .INIT(16'h0400))
    _al_u434 (
    .a(vga_rdaddr[15]),
    .b(vga_rdaddr[14]),
    .c(vga_rdaddr[13]),
    .d(vga_rdaddr[12]),
    .o(\and_vga_rdaddr[12]_N_o_al_n227 ));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*~A)"),
    .INIT(16'h0100))
    _al_u435 (
    .a(vga_rdaddr[15]),
    .b(vga_rdaddr[14]),
    .c(vga_rdaddr[13]),
    .d(vga_rdaddr[12]),
    .o(\and_vga_rdaddr[12]_N_o ));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*~A)"),
    .INIT(16'h0040))
    _al_u436 (
    .a(vga_rdaddr[15]),
    .b(vga_rdaddr[14]),
    .c(vga_rdaddr[13]),
    .d(vga_rdaddr[12]),
    .o(\and_Nvga_rdaddr[12]__o_al_n243 ));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*~A)"),
    .INIT(16'h0004))
    _al_u437 (
    .a(vga_rdaddr[15]),
    .b(vga_rdaddr[14]),
    .c(vga_rdaddr[13]),
    .d(vga_rdaddr[12]),
    .o(\and_Nvga_rdaddr[12]__o_al_n211 ));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*~B*~A)"),
    .INIT(16'h0010))
    _al_u438 (
    .a(vga_rdaddr[15]),
    .b(vga_rdaddr[14]),
    .c(vga_rdaddr[13]),
    .d(vga_rdaddr[12]),
    .o(\and_Nvga_rdaddr[12]__o_al_n180 ));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u439 (
    .a(vga_rdaddr[15]),
    .b(vga_rdaddr[14]),
    .c(vga_rdaddr[13]),
    .d(vga_rdaddr[12]),
    .o(\and_Nvga_rdaddr[12]__o ));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*A)"),
    .INIT(16'h0200))
    _al_u440 (
    .a(vga_rdaddr[15]),
    .b(vga_rdaddr[14]),
    .c(vga_rdaddr[11]),
    .d(vga_rden),
    .o(_al_u440_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u441 (
    .a(_al_u440_o),
    .b(vga_rdaddr[13]),
    .c(vga_rdaddr[12]),
    .o(\and_Nvga_rdaddr[11]__o_and_vga_rden ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u442 (
    .a(cam_rst_pad),
    .b(clk_cam),
    .o(cam_xclk_pad));
  AL_MAP_LUT2 #(
    .EQN("~(~B*A)"),
    .INIT(4'hd))
    _al_u443 (
    .a(cam_vsync_pad),
    .b(\u_camera_reader/vsync_passed ),
    .o(\u_camera_reader/vsync_passed_d ));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u444 (
    .a(\u_camera_reader/n27 ),
    .b(\u_camera_reader/wrclk1 ),
    .c(\u_camera_reader/write_pixel ),
    .o(camera_wrreq));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*B*A)"),
    .INIT(16'h0800))
    _al_u445 (
    .a(_al_u430_o),
    .b(camera_wrreq),
    .c(camera_addr[11]),
    .d(camera_addr[15]),
    .o(\and_Ncamera_addr[11]_o_and_camera_wrreq ));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u446 (
    .a(\u_camera_reader/n2 ),
    .b(\u_camera_reader/pixel_counter [0]),
    .c(\u_camera_reader/vsync_passed ),
    .o(\u_camera_reader/mux6_b0_sel_is_1_o ));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u447 (
    .a(\u_camera_reader/mux6_b0_sel_is_1_o ),
    .b(cam_vsync_pad),
    .c(\u_camera_reader/n9 [9]),
    .d(camera_addr[9]),
    .o(\u_camera_reader/n21 [9]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u448 (
    .a(\u_camera_reader/mux6_b0_sel_is_1_o ),
    .b(cam_vsync_pad),
    .c(\u_camera_reader/n9 [8]),
    .d(camera_addr[8]),
    .o(\u_camera_reader/n21 [8]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u449 (
    .a(\u_camera_reader/mux6_b0_sel_is_1_o ),
    .b(cam_vsync_pad),
    .c(\u_camera_reader/n9 [7]),
    .d(camera_addr[7]),
    .o(\u_camera_reader/n21 [7]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u450 (
    .a(\u_camera_reader/mux6_b0_sel_is_1_o ),
    .b(cam_vsync_pad),
    .c(\u_camera_reader/n9 [6]),
    .d(camera_addr[6]),
    .o(\u_camera_reader/n21 [6]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u451 (
    .a(\u_camera_reader/mux6_b0_sel_is_1_o ),
    .b(cam_vsync_pad),
    .c(\u_camera_reader/n9 [5]),
    .d(camera_addr[5]),
    .o(\u_camera_reader/n21 [5]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u452 (
    .a(\u_camera_reader/mux6_b0_sel_is_1_o ),
    .b(cam_vsync_pad),
    .c(\u_camera_reader/n9 [4]),
    .d(camera_addr[4]),
    .o(\u_camera_reader/n21 [4]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u453 (
    .a(\u_camera_reader/mux6_b0_sel_is_1_o ),
    .b(cam_vsync_pad),
    .c(\u_camera_reader/n9 [3]),
    .d(camera_addr[3]),
    .o(\u_camera_reader/n21 [3]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u454 (
    .a(\u_camera_reader/mux6_b0_sel_is_1_o ),
    .b(cam_vsync_pad),
    .c(\u_camera_reader/n9 [2]),
    .d(camera_addr[2]),
    .o(\u_camera_reader/n21 [2]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u455 (
    .a(\u_camera_reader/mux6_b0_sel_is_1_o ),
    .b(cam_vsync_pad),
    .c(\u_camera_reader/n9 [1]),
    .d(camera_addr[1]),
    .o(\u_camera_reader/n21 [1]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u456 (
    .a(\u_camera_reader/mux6_b0_sel_is_1_o ),
    .b(cam_vsync_pad),
    .c(\u_camera_reader/n9 [15]),
    .d(camera_addr[15]),
    .o(\u_camera_reader/n21 [15]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u457 (
    .a(\u_camera_reader/mux6_b0_sel_is_1_o ),
    .b(cam_vsync_pad),
    .c(\u_camera_reader/n9 [14]),
    .d(camera_addr[14]),
    .o(\u_camera_reader/n21 [14]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u458 (
    .a(\u_camera_reader/mux6_b0_sel_is_1_o ),
    .b(cam_vsync_pad),
    .c(\u_camera_reader/n9 [13]),
    .d(camera_addr[13]),
    .o(\u_camera_reader/n21 [13]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u459 (
    .a(\u_camera_reader/mux6_b0_sel_is_1_o ),
    .b(cam_vsync_pad),
    .c(\u_camera_reader/n9 [12]),
    .d(camera_addr[12]),
    .o(\u_camera_reader/n21 [12]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u460 (
    .a(\u_camera_reader/mux6_b0_sel_is_1_o ),
    .b(cam_vsync_pad),
    .c(\u_camera_reader/n9 [11]),
    .d(camera_addr[11]),
    .o(\u_camera_reader/n21 [11]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u461 (
    .a(\u_camera_reader/mux6_b0_sel_is_1_o ),
    .b(cam_vsync_pad),
    .c(\u_camera_reader/n9 [10]),
    .d(camera_addr[10]),
    .o(\u_camera_reader/n21 [10]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u462 (
    .a(\u_camera_reader/mux6_b0_sel_is_1_o ),
    .b(cam_vsync_pad),
    .c(\u_camera_reader/n9 [0]),
    .d(camera_addr[0]),
    .o(\u_camera_reader/n21 [0]));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u463 (
    .a(\u_camera_reader/mux6_b0_sel_is_1_o ),
    .b(cam_vsync_pad),
    .c(cam_rst_pad),
    .o(\u_camera_reader/mux14_b0_sel_is_2_o ));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u464 (
    .a(\u_camera_reader/n2 ),
    .b(\u_camera_reader/pixel_counter [0]),
    .c(\u_camera_reader/vsync_passed ),
    .o(\u_camera_reader/mux5_b0_sel_is_3_o ));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u465 (
    .a(\u_camera_reader/mux5_b0_sel_is_3_o ),
    .b(cam_vsync_pad),
    .c(cam_rst_pad),
    .o(\u_camera_reader/mux13_b0_sel_is_2_o ));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~D*~(C*A)))"),
    .INIT(16'hcc80))
    _al_u466 (
    .a(\u_camera_reader/n2 ),
    .b(cam_vsync_pad),
    .c(\u_camera_reader/vsync_passed ),
    .d(\u_camera_reader/write_pixel ),
    .o(\u_camera_reader/mux8_b0_sel_is_0_o ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u467 (
    .a(\u_camera_reader/mux8_b0_sel_is_0_o ),
    .b(\u_camera_reader/n8 [9]),
    .o(\u_camera_reader/n19 [9]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u468 (
    .a(\u_camera_reader/mux8_b0_sel_is_0_o ),
    .b(\u_camera_reader/n8 [8]),
    .o(\u_camera_reader/n19 [8]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u469 (
    .a(\u_camera_reader/mux8_b0_sel_is_0_o ),
    .b(\u_camera_reader/n8 [7]),
    .o(\u_camera_reader/n19 [7]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u470 (
    .a(\u_camera_reader/mux8_b0_sel_is_0_o ),
    .b(\u_camera_reader/n8 [6]),
    .o(\u_camera_reader/n19 [6]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u471 (
    .a(\u_camera_reader/mux8_b0_sel_is_0_o ),
    .b(\u_camera_reader/n8 [5]),
    .o(\u_camera_reader/n19 [5]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u472 (
    .a(\u_camera_reader/mux8_b0_sel_is_0_o ),
    .b(\u_camera_reader/n8 [4]),
    .o(\u_camera_reader/n19 [4]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u473 (
    .a(\u_camera_reader/mux8_b0_sel_is_0_o ),
    .b(\u_camera_reader/n8 [3]),
    .o(\u_camera_reader/n19 [3]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u474 (
    .a(\u_camera_reader/mux8_b0_sel_is_0_o ),
    .b(\u_camera_reader/n8 [2]),
    .o(\u_camera_reader/n19 [2]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u475 (
    .a(\u_camera_reader/mux8_b0_sel_is_0_o ),
    .b(\u_camera_reader/n8 [1]),
    .o(\u_camera_reader/n19 [1]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u476 (
    .a(\u_camera_reader/mux8_b0_sel_is_0_o ),
    .b(\u_camera_reader/n8 [19]),
    .o(\u_camera_reader/n19 [19]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u477 (
    .a(\u_camera_reader/mux8_b0_sel_is_0_o ),
    .b(\u_camera_reader/n8 [18]),
    .o(\u_camera_reader/n19 [18]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u478 (
    .a(\u_camera_reader/mux8_b0_sel_is_0_o ),
    .b(\u_camera_reader/n8 [17]),
    .o(\u_camera_reader/n19 [17]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u479 (
    .a(\u_camera_reader/mux8_b0_sel_is_0_o ),
    .b(\u_camera_reader/n8 [16]),
    .o(\u_camera_reader/n19 [16]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u480 (
    .a(\u_camera_reader/mux8_b0_sel_is_0_o ),
    .b(\u_camera_reader/n8 [15]),
    .o(\u_camera_reader/n19 [15]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u481 (
    .a(\u_camera_reader/mux8_b0_sel_is_0_o ),
    .b(\u_camera_reader/n8 [14]),
    .o(\u_camera_reader/n19 [14]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u482 (
    .a(\u_camera_reader/mux8_b0_sel_is_0_o ),
    .b(\u_camera_reader/n8 [13]),
    .o(\u_camera_reader/n19 [13]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u483 (
    .a(\u_camera_reader/mux8_b0_sel_is_0_o ),
    .b(\u_camera_reader/n8 [12]),
    .o(\u_camera_reader/n19 [12]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u484 (
    .a(\u_camera_reader/mux8_b0_sel_is_0_o ),
    .b(\u_camera_reader/n8 [11]),
    .o(\u_camera_reader/n19 [11]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u485 (
    .a(\u_camera_reader/mux8_b0_sel_is_0_o ),
    .b(\u_camera_reader/n8 [10]),
    .o(\u_camera_reader/n19 [10]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u486 (
    .a(\u_camera_reader/mux8_b0_sel_is_0_o ),
    .b(\u_camera_reader/n8 [0]),
    .o(\u_camera_reader/n19 [0]));
  AL_MAP_LUT4 #(
    .EQN("(~D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h00ca))
    _al_u487 (
    .a(\u_img/inst_dob_i0_009 ),
    .b(\u_img/inst_dob_i16_009 ),
    .c(vga_rdaddr_piped_piped[4]),
    .d(vga_rdaddr_piped_piped[5]),
    .o(_al_u487_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'hca00))
    _al_u488 (
    .a(\u_img/inst_dob_i32_009 ),
    .b(\u_img/inst_dob_i48_009 ),
    .c(vga_rdaddr_piped_piped[4]),
    .d(vga_rdaddr_piped_piped[5]),
    .o(_al_u488_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*~A))"),
    .INIT(8'h8c))
    _al_u489 (
    .a(\u_img/inst_dob_i64_009 ),
    .b(vga_rden),
    .c(vga_rdaddr_piped_piped[6]),
    .o(_al_u489_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(~D*~B*~A))"),
    .INIT(16'hf0e0))
    _al_u490 (
    .a(_al_u487_o),
    .b(_al_u488_o),
    .c(_al_u489_o),
    .d(vga_rdaddr_piped_piped[6]),
    .o(vga_g_pad[6]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h0035))
    _al_u491 (
    .a(\u_img/inst_dob_i24_008 ),
    .b(\u_img/inst_dob_i26_008 ),
    .c(vga_rdaddr_piped_piped[1]),
    .d(vga_rdaddr_piped_piped[2]),
    .o(_al_u491_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h3500))
    _al_u492 (
    .a(\u_img/inst_dob_i28_008 ),
    .b(\u_img/inst_dob_i30_008 ),
    .c(vga_rdaddr_piped_piped[1]),
    .d(vga_rdaddr_piped_piped[2]),
    .o(_al_u492_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h0035))
    _al_u493 (
    .a(\u_img/inst_dob_i16_008 ),
    .b(\u_img/inst_dob_i18_008 ),
    .c(vga_rdaddr_piped_piped[1]),
    .d(vga_rdaddr_piped_piped[2]),
    .o(_al_u493_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h3500))
    _al_u494 (
    .a(\u_img/inst_dob_i20_008 ),
    .b(\u_img/inst_dob_i22_008 ),
    .c(vga_rdaddr_piped_piped[1]),
    .d(vga_rdaddr_piped_piped[2]),
    .o(_al_u494_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u495 (
    .a(_al_u493_o),
    .b(_al_u494_o),
    .c(vga_rdaddr_piped_piped[3]),
    .o(_al_u495_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(D*~C*~B))"),
    .INIT(16'h5455))
    _al_u496 (
    .a(_al_u495_o),
    .b(_al_u491_o),
    .c(_al_u492_o),
    .d(vga_rdaddr_piped_piped[3]),
    .o(_al_u496_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h0035))
    _al_u497 (
    .a(\u_img/inst_dob_i8_008 ),
    .b(\u_img/inst_dob_i10_008 ),
    .c(vga_rdaddr_piped_piped[1]),
    .d(vga_rdaddr_piped_piped[2]),
    .o(_al_u497_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h3500))
    _al_u498 (
    .a(\u_img/inst_dob_i12_008 ),
    .b(\u_img/inst_dob_i14_008 ),
    .c(vga_rdaddr_piped_piped[1]),
    .d(vga_rdaddr_piped_piped[2]),
    .o(_al_u498_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h0035))
    _al_u499 (
    .a(\u_img/inst_dob_i0_008 ),
    .b(\u_img/inst_dob_i2_008 ),
    .c(vga_rdaddr_piped_piped[1]),
    .d(vga_rdaddr_piped_piped[2]),
    .o(_al_u499_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h3500))
    _al_u500 (
    .a(\u_img/inst_dob_i4_008 ),
    .b(\u_img/inst_dob_i6_008 ),
    .c(vga_rdaddr_piped_piped[1]),
    .d(vga_rdaddr_piped_piped[2]),
    .o(_al_u500_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u501 (
    .a(_al_u499_o),
    .b(_al_u500_o),
    .c(vga_rdaddr_piped_piped[3]),
    .o(_al_u501_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(D*~C*~B))"),
    .INIT(16'h5455))
    _al_u502 (
    .a(_al_u501_o),
    .b(_al_u497_o),
    .c(_al_u498_o),
    .d(vga_rdaddr_piped_piped[3]),
    .o(_al_u502_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'h00ac))
    _al_u503 (
    .a(_al_u496_o),
    .b(_al_u502_o),
    .c(vga_rdaddr_piped_piped[4]),
    .d(vga_rdaddr_piped_piped[5]),
    .o(_al_u503_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h0035))
    _al_u504 (
    .a(\u_img/inst_dob_i40_008 ),
    .b(\u_img/inst_dob_i42_008 ),
    .c(vga_rdaddr_piped_piped[1]),
    .d(vga_rdaddr_piped_piped[2]),
    .o(_al_u504_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h3500))
    _al_u505 (
    .a(\u_img/inst_dob_i44_008 ),
    .b(\u_img/inst_dob_i46_008 ),
    .c(vga_rdaddr_piped_piped[1]),
    .d(vga_rdaddr_piped_piped[2]),
    .o(_al_u505_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h0035))
    _al_u506 (
    .a(\u_img/inst_dob_i32_008 ),
    .b(\u_img/inst_dob_i34_008 ),
    .c(vga_rdaddr_piped_piped[1]),
    .d(vga_rdaddr_piped_piped[2]),
    .o(_al_u506_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h3500))
    _al_u507 (
    .a(\u_img/inst_dob_i36_008 ),
    .b(\u_img/inst_dob_i38_008 ),
    .c(vga_rdaddr_piped_piped[1]),
    .d(vga_rdaddr_piped_piped[2]),
    .o(_al_u507_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u508 (
    .a(_al_u506_o),
    .b(_al_u507_o),
    .c(vga_rdaddr_piped_piped[3]),
    .o(_al_u508_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(D*~C*~B))"),
    .INIT(16'h5455))
    _al_u509 (
    .a(_al_u508_o),
    .b(_al_u504_o),
    .c(_al_u505_o),
    .d(vga_rdaddr_piped_piped[3]),
    .o(_al_u509_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h0035))
    _al_u510 (
    .a(\u_img/inst_dob_i56_008 ),
    .b(\u_img/inst_dob_i58_008 ),
    .c(vga_rdaddr_piped_piped[1]),
    .d(vga_rdaddr_piped_piped[2]),
    .o(_al_u510_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h3500))
    _al_u511 (
    .a(\u_img/inst_dob_i60_008 ),
    .b(\u_img/inst_dob_i62_008 ),
    .c(vga_rdaddr_piped_piped[1]),
    .d(vga_rdaddr_piped_piped[2]),
    .o(_al_u511_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h0035))
    _al_u512 (
    .a(\u_img/inst_dob_i48_008 ),
    .b(\u_img/inst_dob_i50_008 ),
    .c(vga_rdaddr_piped_piped[1]),
    .d(vga_rdaddr_piped_piped[2]),
    .o(_al_u512_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h3500))
    _al_u513 (
    .a(\u_img/inst_dob_i52_008 ),
    .b(\u_img/inst_dob_i54_008 ),
    .c(vga_rdaddr_piped_piped[1]),
    .d(vga_rdaddr_piped_piped[2]),
    .o(_al_u513_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u514 (
    .a(_al_u512_o),
    .b(_al_u513_o),
    .c(vga_rdaddr_piped_piped[3]),
    .o(_al_u514_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(D*~C*~B))"),
    .INIT(16'h5455))
    _al_u515 (
    .a(_al_u514_o),
    .b(_al_u510_o),
    .c(_al_u511_o),
    .d(vga_rdaddr_piped_piped[3]),
    .o(_al_u515_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'hca00))
    _al_u516 (
    .a(_al_u509_o),
    .b(_al_u515_o),
    .c(vga_rdaddr_piped_piped[4]),
    .d(vga_rdaddr_piped_piped[5]),
    .o(_al_u516_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*~A))"),
    .INIT(8'h8c))
    _al_u517 (
    .a(\u_img/inst_dob_i64_008 ),
    .b(vga_rden),
    .c(vga_rdaddr_piped_piped[6]),
    .o(_al_u517_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(~D*~(~B*~A)))"),
    .INIT(16'hf010))
    _al_u518 (
    .a(_al_u503_o),
    .b(_al_u516_o),
    .c(_al_u517_o),
    .d(vga_rdaddr_piped_piped[6]),
    .o(vga_g_pad[5]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h0035))
    _al_u519 (
    .a(\u_img/inst_dob_i56_007 ),
    .b(\u_img/inst_dob_i58_007 ),
    .c(vga_rdaddr_piped_piped[1]),
    .d(vga_rdaddr_piped_piped[2]),
    .o(_al_u519_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h3500))
    _al_u520 (
    .a(\u_img/inst_dob_i60_007 ),
    .b(\u_img/inst_dob_i62_007 ),
    .c(vga_rdaddr_piped_piped[1]),
    .d(vga_rdaddr_piped_piped[2]),
    .o(_al_u520_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h0035))
    _al_u521 (
    .a(\u_img/inst_dob_i48_007 ),
    .b(\u_img/inst_dob_i50_007 ),
    .c(vga_rdaddr_piped_piped[1]),
    .d(vga_rdaddr_piped_piped[2]),
    .o(_al_u521_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h3500))
    _al_u522 (
    .a(\u_img/inst_dob_i52_007 ),
    .b(\u_img/inst_dob_i54_007 ),
    .c(vga_rdaddr_piped_piped[1]),
    .d(vga_rdaddr_piped_piped[2]),
    .o(_al_u522_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u523 (
    .a(_al_u521_o),
    .b(_al_u522_o),
    .c(vga_rdaddr_piped_piped[3]),
    .o(_al_u523_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(D*~C*~B))"),
    .INIT(16'h5455))
    _al_u524 (
    .a(_al_u523_o),
    .b(_al_u519_o),
    .c(_al_u520_o),
    .d(vga_rdaddr_piped_piped[3]),
    .o(_al_u524_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h0035))
    _al_u525 (
    .a(\u_img/inst_dob_i40_007 ),
    .b(\u_img/inst_dob_i42_007 ),
    .c(vga_rdaddr_piped_piped[1]),
    .d(vga_rdaddr_piped_piped[2]),
    .o(_al_u525_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h3500))
    _al_u526 (
    .a(\u_img/inst_dob_i44_007 ),
    .b(\u_img/inst_dob_i46_007 ),
    .c(vga_rdaddr_piped_piped[1]),
    .d(vga_rdaddr_piped_piped[2]),
    .o(_al_u526_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h0035))
    _al_u527 (
    .a(\u_img/inst_dob_i32_007 ),
    .b(\u_img/inst_dob_i34_007 ),
    .c(vga_rdaddr_piped_piped[1]),
    .d(vga_rdaddr_piped_piped[2]),
    .o(_al_u527_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h3500))
    _al_u528 (
    .a(\u_img/inst_dob_i36_007 ),
    .b(\u_img/inst_dob_i38_007 ),
    .c(vga_rdaddr_piped_piped[1]),
    .d(vga_rdaddr_piped_piped[2]),
    .o(_al_u528_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u529 (
    .a(_al_u527_o),
    .b(_al_u528_o),
    .c(vga_rdaddr_piped_piped[3]),
    .o(_al_u529_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(D*~C*~B))"),
    .INIT(16'h5455))
    _al_u530 (
    .a(_al_u529_o),
    .b(_al_u525_o),
    .c(_al_u526_o),
    .d(vga_rdaddr_piped_piped[3]),
    .o(_al_u530_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'hac00))
    _al_u531 (
    .a(_al_u524_o),
    .b(_al_u530_o),
    .c(vga_rdaddr_piped_piped[4]),
    .d(vga_rdaddr_piped_piped[5]),
    .o(_al_u531_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h0035))
    _al_u532 (
    .a(\u_img/inst_dob_i24_007 ),
    .b(\u_img/inst_dob_i26_007 ),
    .c(vga_rdaddr_piped_piped[1]),
    .d(vga_rdaddr_piped_piped[2]),
    .o(_al_u532_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h3500))
    _al_u533 (
    .a(\u_img/inst_dob_i28_007 ),
    .b(\u_img/inst_dob_i30_007 ),
    .c(vga_rdaddr_piped_piped[1]),
    .d(vga_rdaddr_piped_piped[2]),
    .o(_al_u533_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h0035))
    _al_u534 (
    .a(\u_img/inst_dob_i16_007 ),
    .b(\u_img/inst_dob_i18_007 ),
    .c(vga_rdaddr_piped_piped[1]),
    .d(vga_rdaddr_piped_piped[2]),
    .o(_al_u534_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h3500))
    _al_u535 (
    .a(\u_img/inst_dob_i20_007 ),
    .b(\u_img/inst_dob_i22_007 ),
    .c(vga_rdaddr_piped_piped[1]),
    .d(vga_rdaddr_piped_piped[2]),
    .o(_al_u535_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u536 (
    .a(_al_u534_o),
    .b(_al_u535_o),
    .c(vga_rdaddr_piped_piped[3]),
    .o(_al_u536_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(D*~C*~B))"),
    .INIT(16'h5455))
    _al_u537 (
    .a(_al_u536_o),
    .b(_al_u532_o),
    .c(_al_u533_o),
    .d(vga_rdaddr_piped_piped[3]),
    .o(_al_u537_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h0035))
    _al_u538 (
    .a(\u_img/inst_dob_i8_007 ),
    .b(\u_img/inst_dob_i10_007 ),
    .c(vga_rdaddr_piped_piped[1]),
    .d(vga_rdaddr_piped_piped[2]),
    .o(_al_u538_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h3500))
    _al_u539 (
    .a(\u_img/inst_dob_i12_007 ),
    .b(\u_img/inst_dob_i14_007 ),
    .c(vga_rdaddr_piped_piped[1]),
    .d(vga_rdaddr_piped_piped[2]),
    .o(_al_u539_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h0035))
    _al_u540 (
    .a(\u_img/inst_dob_i0_007 ),
    .b(\u_img/inst_dob_i2_007 ),
    .c(vga_rdaddr_piped_piped[1]),
    .d(vga_rdaddr_piped_piped[2]),
    .o(_al_u540_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h3500))
    _al_u541 (
    .a(\u_img/inst_dob_i4_007 ),
    .b(\u_img/inst_dob_i6_007 ),
    .c(vga_rdaddr_piped_piped[1]),
    .d(vga_rdaddr_piped_piped[2]),
    .o(_al_u541_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u542 (
    .a(_al_u540_o),
    .b(_al_u541_o),
    .c(vga_rdaddr_piped_piped[3]),
    .o(_al_u542_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(D*~C*~B))"),
    .INIT(16'h5455))
    _al_u543 (
    .a(_al_u542_o),
    .b(_al_u538_o),
    .c(_al_u539_o),
    .d(vga_rdaddr_piped_piped[3]),
    .o(_al_u543_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'h00ac))
    _al_u544 (
    .a(_al_u537_o),
    .b(_al_u543_o),
    .c(vga_rdaddr_piped_piped[4]),
    .d(vga_rdaddr_piped_piped[5]),
    .o(_al_u544_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*~A))"),
    .INIT(8'h8c))
    _al_u545 (
    .a(\u_img/inst_dob_i64_007 ),
    .b(vga_rden),
    .c(vga_rdaddr_piped_piped[6]),
    .o(_al_u545_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(~D*~(~B*~A)))"),
    .INIT(16'hf010))
    _al_u546 (
    .a(_al_u531_o),
    .b(_al_u544_o),
    .c(_al_u545_o),
    .d(vga_rdaddr_piped_piped[6]),
    .o(vga_g_pad[4]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u547 (
    .a(\u_img/inst_dob_i4_006 ),
    .b(\u_img/inst_dob_i6_006 ),
    .c(vga_rdaddr_piped_piped[1]),
    .o(_al_u547_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u548 (
    .a(\u_img/inst_dob_i0_006 ),
    .b(\u_img/inst_dob_i2_006 ),
    .c(vga_rdaddr_piped_piped[1]),
    .o(_al_u548_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'h00ac))
    _al_u549 (
    .a(_al_u547_o),
    .b(_al_u548_o),
    .c(vga_rdaddr_piped_piped[2]),
    .d(vga_rdaddr_piped_piped[3]),
    .o(_al_u549_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'hca00))
    _al_u550 (
    .a(\u_img/inst_dob_i12_006 ),
    .b(\u_img/inst_dob_i14_006 ),
    .c(vga_rdaddr_piped_piped[1]),
    .d(vga_rdaddr_piped_piped[2]),
    .o(_al_u550_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h00ca))
    _al_u551 (
    .a(\u_img/inst_dob_i8_006 ),
    .b(\u_img/inst_dob_i10_006 ),
    .c(vga_rdaddr_piped_piped[1]),
    .d(vga_rdaddr_piped_piped[2]),
    .o(_al_u551_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(C*~B*~A))"),
    .INIT(16'h00ef))
    _al_u552 (
    .a(_al_u550_o),
    .b(_al_u551_o),
    .c(vga_rdaddr_piped_piped[3]),
    .d(vga_rdaddr_piped_piped[4]),
    .o(_al_u552_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u553 (
    .a(\u_img/inst_dob_i28_006 ),
    .b(\u_img/inst_dob_i30_006 ),
    .c(vga_rdaddr_piped_piped[1]),
    .o(_al_u553_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u554 (
    .a(\u_img/inst_dob_i24_006 ),
    .b(\u_img/inst_dob_i26_006 ),
    .c(vga_rdaddr_piped_piped[1]),
    .o(_al_u554_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'hac00))
    _al_u555 (
    .a(_al_u553_o),
    .b(_al_u554_o),
    .c(vga_rdaddr_piped_piped[2]),
    .d(vga_rdaddr_piped_piped[3]),
    .o(_al_u555_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'hca00))
    _al_u556 (
    .a(\u_img/inst_dob_i20_006 ),
    .b(\u_img/inst_dob_i22_006 ),
    .c(vga_rdaddr_piped_piped[1]),
    .d(vga_rdaddr_piped_piped[2]),
    .o(_al_u556_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h00ca))
    _al_u557 (
    .a(\u_img/inst_dob_i16_006 ),
    .b(\u_img/inst_dob_i18_006 ),
    .c(vga_rdaddr_piped_piped[1]),
    .d(vga_rdaddr_piped_piped[2]),
    .o(_al_u557_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(~C*~B*~A))"),
    .INIT(16'hfe00))
    _al_u558 (
    .a(_al_u556_o),
    .b(_al_u557_o),
    .c(vga_rdaddr_piped_piped[3]),
    .d(vga_rdaddr_piped_piped[4]),
    .o(_al_u558_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~C)*~(B*~A))"),
    .INIT(16'hb0bb))
    _al_u559 (
    .a(_al_u549_o),
    .b(_al_u552_o),
    .c(_al_u555_o),
    .d(_al_u558_o),
    .o(_al_u559_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u560 (
    .a(\u_img/inst_dob_i36_006 ),
    .b(\u_img/inst_dob_i38_006 ),
    .c(vga_rdaddr_piped_piped[1]),
    .o(_al_u560_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u561 (
    .a(\u_img/inst_dob_i32_006 ),
    .b(\u_img/inst_dob_i34_006 ),
    .c(vga_rdaddr_piped_piped[1]),
    .o(_al_u561_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'h00ac))
    _al_u562 (
    .a(_al_u560_o),
    .b(_al_u561_o),
    .c(vga_rdaddr_piped_piped[2]),
    .d(vga_rdaddr_piped_piped[3]),
    .o(_al_u562_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'hca00))
    _al_u563 (
    .a(\u_img/inst_dob_i44_006 ),
    .b(\u_img/inst_dob_i46_006 ),
    .c(vga_rdaddr_piped_piped[1]),
    .d(vga_rdaddr_piped_piped[2]),
    .o(_al_u563_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h00ca))
    _al_u564 (
    .a(\u_img/inst_dob_i40_006 ),
    .b(\u_img/inst_dob_i42_006 ),
    .c(vga_rdaddr_piped_piped[1]),
    .d(vga_rdaddr_piped_piped[2]),
    .o(_al_u564_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(C*~B*~A))"),
    .INIT(16'h00ef))
    _al_u565 (
    .a(_al_u563_o),
    .b(_al_u564_o),
    .c(vga_rdaddr_piped_piped[3]),
    .d(vga_rdaddr_piped_piped[4]),
    .o(_al_u565_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u566 (
    .a(\u_img/inst_dob_i52_006 ),
    .b(\u_img/inst_dob_i54_006 ),
    .c(vga_rdaddr_piped_piped[1]),
    .o(_al_u566_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u567 (
    .a(\u_img/inst_dob_i48_006 ),
    .b(\u_img/inst_dob_i50_006 ),
    .c(vga_rdaddr_piped_piped[1]),
    .o(_al_u567_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'h00ac))
    _al_u568 (
    .a(_al_u566_o),
    .b(_al_u567_o),
    .c(vga_rdaddr_piped_piped[2]),
    .d(vga_rdaddr_piped_piped[3]),
    .o(_al_u568_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'hca00))
    _al_u569 (
    .a(\u_img/inst_dob_i60_006 ),
    .b(\u_img/inst_dob_i62_006 ),
    .c(vga_rdaddr_piped_piped[1]),
    .d(vga_rdaddr_piped_piped[2]),
    .o(_al_u569_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h00ca))
    _al_u570 (
    .a(\u_img/inst_dob_i56_006 ),
    .b(\u_img/inst_dob_i58_006 ),
    .c(vga_rdaddr_piped_piped[1]),
    .d(vga_rdaddr_piped_piped[2]),
    .o(_al_u570_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C*~B*~A))"),
    .INIT(16'hef00))
    _al_u571 (
    .a(_al_u569_o),
    .b(_al_u570_o),
    .c(vga_rdaddr_piped_piped[3]),
    .d(vga_rdaddr_piped_piped[4]),
    .o(_al_u571_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~C)*~(B*~A))"),
    .INIT(16'hb0bb))
    _al_u572 (
    .a(_al_u562_o),
    .b(_al_u565_o),
    .c(_al_u568_o),
    .d(_al_u571_o),
    .o(_al_u572_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h00ca))
    _al_u573 (
    .a(_al_u559_o),
    .b(_al_u572_o),
    .c(vga_rdaddr_piped_piped[5]),
    .d(vga_rdaddr_piped_piped[6]),
    .o(_al_u573_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*~(D*~B))"),
    .INIT(16'h4050))
    _al_u574 (
    .a(_al_u573_o),
    .b(\u_img/inst_dob_i64_006 ),
    .c(vga_rden),
    .d(vga_rdaddr_piped_piped[6]),
    .o(vga_g_pad[3]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h0035))
    _al_u575 (
    .a(\u_img/inst_dob_i56_005 ),
    .b(\u_img/inst_dob_i58_005 ),
    .c(vga_rdaddr_piped_piped[1]),
    .d(vga_rdaddr_piped_piped[2]),
    .o(_al_u575_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h3500))
    _al_u576 (
    .a(\u_img/inst_dob_i60_005 ),
    .b(\u_img/inst_dob_i62_005 ),
    .c(vga_rdaddr_piped_piped[1]),
    .d(vga_rdaddr_piped_piped[2]),
    .o(_al_u576_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h0035))
    _al_u577 (
    .a(\u_img/inst_dob_i48_005 ),
    .b(\u_img/inst_dob_i50_005 ),
    .c(vga_rdaddr_piped_piped[1]),
    .d(vga_rdaddr_piped_piped[2]),
    .o(_al_u577_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h3500))
    _al_u578 (
    .a(\u_img/inst_dob_i52_005 ),
    .b(\u_img/inst_dob_i54_005 ),
    .c(vga_rdaddr_piped_piped[1]),
    .d(vga_rdaddr_piped_piped[2]),
    .o(_al_u578_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u579 (
    .a(_al_u577_o),
    .b(_al_u578_o),
    .c(vga_rdaddr_piped_piped[3]),
    .o(_al_u579_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(D*~C*~B))"),
    .INIT(16'h5455))
    _al_u580 (
    .a(_al_u579_o),
    .b(_al_u575_o),
    .c(_al_u576_o),
    .d(vga_rdaddr_piped_piped[3]),
    .o(_al_u580_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h0035))
    _al_u581 (
    .a(\u_img/inst_dob_i40_005 ),
    .b(\u_img/inst_dob_i42_005 ),
    .c(vga_rdaddr_piped_piped[1]),
    .d(vga_rdaddr_piped_piped[2]),
    .o(_al_u581_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h3500))
    _al_u582 (
    .a(\u_img/inst_dob_i44_005 ),
    .b(\u_img/inst_dob_i46_005 ),
    .c(vga_rdaddr_piped_piped[1]),
    .d(vga_rdaddr_piped_piped[2]),
    .o(_al_u582_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h0035))
    _al_u583 (
    .a(\u_img/inst_dob_i32_005 ),
    .b(\u_img/inst_dob_i34_005 ),
    .c(vga_rdaddr_piped_piped[1]),
    .d(vga_rdaddr_piped_piped[2]),
    .o(_al_u583_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h3500))
    _al_u584 (
    .a(\u_img/inst_dob_i36_005 ),
    .b(\u_img/inst_dob_i38_005 ),
    .c(vga_rdaddr_piped_piped[1]),
    .d(vga_rdaddr_piped_piped[2]),
    .o(_al_u584_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u585 (
    .a(_al_u583_o),
    .b(_al_u584_o),
    .c(vga_rdaddr_piped_piped[3]),
    .o(_al_u585_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(D*~C*~B))"),
    .INIT(16'h5455))
    _al_u586 (
    .a(_al_u585_o),
    .b(_al_u581_o),
    .c(_al_u582_o),
    .d(vga_rdaddr_piped_piped[3]),
    .o(_al_u586_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'hac00))
    _al_u587 (
    .a(_al_u580_o),
    .b(_al_u586_o),
    .c(vga_rdaddr_piped_piped[4]),
    .d(vga_rdaddr_piped_piped[5]),
    .o(_al_u587_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h0035))
    _al_u588 (
    .a(\u_img/inst_dob_i24_005 ),
    .b(\u_img/inst_dob_i26_005 ),
    .c(vga_rdaddr_piped_piped[1]),
    .d(vga_rdaddr_piped_piped[2]),
    .o(_al_u588_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h3500))
    _al_u589 (
    .a(\u_img/inst_dob_i28_005 ),
    .b(\u_img/inst_dob_i30_005 ),
    .c(vga_rdaddr_piped_piped[1]),
    .d(vga_rdaddr_piped_piped[2]),
    .o(_al_u589_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h0035))
    _al_u590 (
    .a(\u_img/inst_dob_i16_005 ),
    .b(\u_img/inst_dob_i18_005 ),
    .c(vga_rdaddr_piped_piped[1]),
    .d(vga_rdaddr_piped_piped[2]),
    .o(_al_u590_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h3500))
    _al_u591 (
    .a(\u_img/inst_dob_i20_005 ),
    .b(\u_img/inst_dob_i22_005 ),
    .c(vga_rdaddr_piped_piped[1]),
    .d(vga_rdaddr_piped_piped[2]),
    .o(_al_u591_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u592 (
    .a(_al_u590_o),
    .b(_al_u591_o),
    .c(vga_rdaddr_piped_piped[3]),
    .o(_al_u592_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(D*~C*~B))"),
    .INIT(16'h5455))
    _al_u593 (
    .a(_al_u592_o),
    .b(_al_u588_o),
    .c(_al_u589_o),
    .d(vga_rdaddr_piped_piped[3]),
    .o(_al_u593_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h0035))
    _al_u594 (
    .a(\u_img/inst_dob_i8_005 ),
    .b(\u_img/inst_dob_i10_005 ),
    .c(vga_rdaddr_piped_piped[1]),
    .d(vga_rdaddr_piped_piped[2]),
    .o(_al_u594_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h3500))
    _al_u595 (
    .a(\u_img/inst_dob_i12_005 ),
    .b(\u_img/inst_dob_i14_005 ),
    .c(vga_rdaddr_piped_piped[1]),
    .d(vga_rdaddr_piped_piped[2]),
    .o(_al_u595_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h0035))
    _al_u596 (
    .a(\u_img/inst_dob_i0_005 ),
    .b(\u_img/inst_dob_i2_005 ),
    .c(vga_rdaddr_piped_piped[1]),
    .d(vga_rdaddr_piped_piped[2]),
    .o(_al_u596_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h3500))
    _al_u597 (
    .a(\u_img/inst_dob_i4_005 ),
    .b(\u_img/inst_dob_i6_005 ),
    .c(vga_rdaddr_piped_piped[1]),
    .d(vga_rdaddr_piped_piped[2]),
    .o(_al_u597_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u598 (
    .a(_al_u596_o),
    .b(_al_u597_o),
    .c(vga_rdaddr_piped_piped[3]),
    .o(_al_u598_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(D*~C*~B))"),
    .INIT(16'h5455))
    _al_u599 (
    .a(_al_u598_o),
    .b(_al_u594_o),
    .c(_al_u595_o),
    .d(vga_rdaddr_piped_piped[3]),
    .o(_al_u599_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'h00ac))
    _al_u600 (
    .a(_al_u593_o),
    .b(_al_u599_o),
    .c(vga_rdaddr_piped_piped[4]),
    .d(vga_rdaddr_piped_piped[5]),
    .o(_al_u600_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*~A))"),
    .INIT(8'h8c))
    _al_u601 (
    .a(\u_img/inst_dob_i64_005 ),
    .b(vga_rden),
    .c(vga_rdaddr_piped_piped[6]),
    .o(_al_u601_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(~D*~(~B*~A)))"),
    .INIT(16'hf010))
    _al_u602 (
    .a(_al_u587_o),
    .b(_al_u600_o),
    .c(_al_u601_o),
    .d(vga_rdaddr_piped_piped[6]),
    .o(vga_g_pad[2]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h0035))
    _al_u603 (
    .a(\u_img/inst_dob_i56_004 ),
    .b(\u_img/inst_dob_i58_004 ),
    .c(vga_rdaddr_piped_piped[1]),
    .d(vga_rdaddr_piped_piped[2]),
    .o(_al_u603_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h3500))
    _al_u604 (
    .a(\u_img/inst_dob_i60_004 ),
    .b(\u_img/inst_dob_i62_004 ),
    .c(vga_rdaddr_piped_piped[1]),
    .d(vga_rdaddr_piped_piped[2]),
    .o(_al_u604_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h0035))
    _al_u605 (
    .a(\u_img/inst_dob_i48_004 ),
    .b(\u_img/inst_dob_i50_004 ),
    .c(vga_rdaddr_piped_piped[1]),
    .d(vga_rdaddr_piped_piped[2]),
    .o(_al_u605_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h3500))
    _al_u606 (
    .a(\u_img/inst_dob_i52_004 ),
    .b(\u_img/inst_dob_i54_004 ),
    .c(vga_rdaddr_piped_piped[1]),
    .d(vga_rdaddr_piped_piped[2]),
    .o(_al_u606_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u607 (
    .a(_al_u605_o),
    .b(_al_u606_o),
    .c(vga_rdaddr_piped_piped[3]),
    .o(_al_u607_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(D*~C*~B))"),
    .INIT(16'h5455))
    _al_u608 (
    .a(_al_u607_o),
    .b(_al_u603_o),
    .c(_al_u604_o),
    .d(vga_rdaddr_piped_piped[3]),
    .o(_al_u608_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h0035))
    _al_u609 (
    .a(\u_img/inst_dob_i40_004 ),
    .b(\u_img/inst_dob_i42_004 ),
    .c(vga_rdaddr_piped_piped[1]),
    .d(vga_rdaddr_piped_piped[2]),
    .o(_al_u609_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h3500))
    _al_u610 (
    .a(\u_img/inst_dob_i44_004 ),
    .b(\u_img/inst_dob_i46_004 ),
    .c(vga_rdaddr_piped_piped[1]),
    .d(vga_rdaddr_piped_piped[2]),
    .o(_al_u610_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h0035))
    _al_u611 (
    .a(\u_img/inst_dob_i32_004 ),
    .b(\u_img/inst_dob_i34_004 ),
    .c(vga_rdaddr_piped_piped[1]),
    .d(vga_rdaddr_piped_piped[2]),
    .o(_al_u611_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h3500))
    _al_u612 (
    .a(\u_img/inst_dob_i36_004 ),
    .b(\u_img/inst_dob_i38_004 ),
    .c(vga_rdaddr_piped_piped[1]),
    .d(vga_rdaddr_piped_piped[2]),
    .o(_al_u612_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u613 (
    .a(_al_u611_o),
    .b(_al_u612_o),
    .c(vga_rdaddr_piped_piped[3]),
    .o(_al_u613_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(D*~C*~B))"),
    .INIT(16'h5455))
    _al_u614 (
    .a(_al_u613_o),
    .b(_al_u609_o),
    .c(_al_u610_o),
    .d(vga_rdaddr_piped_piped[3]),
    .o(_al_u614_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'hac00))
    _al_u615 (
    .a(_al_u608_o),
    .b(_al_u614_o),
    .c(vga_rdaddr_piped_piped[4]),
    .d(vga_rdaddr_piped_piped[5]),
    .o(_al_u615_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h0035))
    _al_u616 (
    .a(\u_img/inst_dob_i24_004 ),
    .b(\u_img/inst_dob_i26_004 ),
    .c(vga_rdaddr_piped_piped[1]),
    .d(vga_rdaddr_piped_piped[2]),
    .o(_al_u616_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h3500))
    _al_u617 (
    .a(\u_img/inst_dob_i28_004 ),
    .b(\u_img/inst_dob_i30_004 ),
    .c(vga_rdaddr_piped_piped[1]),
    .d(vga_rdaddr_piped_piped[2]),
    .o(_al_u617_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h0035))
    _al_u618 (
    .a(\u_img/inst_dob_i16_004 ),
    .b(\u_img/inst_dob_i18_004 ),
    .c(vga_rdaddr_piped_piped[1]),
    .d(vga_rdaddr_piped_piped[2]),
    .o(_al_u618_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h3500))
    _al_u619 (
    .a(\u_img/inst_dob_i20_004 ),
    .b(\u_img/inst_dob_i22_004 ),
    .c(vga_rdaddr_piped_piped[1]),
    .d(vga_rdaddr_piped_piped[2]),
    .o(_al_u619_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u620 (
    .a(_al_u618_o),
    .b(_al_u619_o),
    .c(vga_rdaddr_piped_piped[3]),
    .o(_al_u620_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(D*~C*~B))"),
    .INIT(16'h5455))
    _al_u621 (
    .a(_al_u620_o),
    .b(_al_u616_o),
    .c(_al_u617_o),
    .d(vga_rdaddr_piped_piped[3]),
    .o(_al_u621_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h0035))
    _al_u622 (
    .a(\u_img/inst_dob_i8_004 ),
    .b(\u_img/inst_dob_i10_004 ),
    .c(vga_rdaddr_piped_piped[1]),
    .d(vga_rdaddr_piped_piped[2]),
    .o(_al_u622_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h3500))
    _al_u623 (
    .a(\u_img/inst_dob_i12_004 ),
    .b(\u_img/inst_dob_i14_004 ),
    .c(vga_rdaddr_piped_piped[1]),
    .d(vga_rdaddr_piped_piped[2]),
    .o(_al_u623_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h0035))
    _al_u624 (
    .a(\u_img/inst_dob_i0_004 ),
    .b(\u_img/inst_dob_i2_004 ),
    .c(vga_rdaddr_piped_piped[1]),
    .d(vga_rdaddr_piped_piped[2]),
    .o(_al_u624_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h3500))
    _al_u625 (
    .a(\u_img/inst_dob_i4_004 ),
    .b(\u_img/inst_dob_i6_004 ),
    .c(vga_rdaddr_piped_piped[1]),
    .d(vga_rdaddr_piped_piped[2]),
    .o(_al_u625_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u626 (
    .a(_al_u624_o),
    .b(_al_u625_o),
    .c(vga_rdaddr_piped_piped[3]),
    .o(_al_u626_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(D*~C*~B))"),
    .INIT(16'h5455))
    _al_u627 (
    .a(_al_u626_o),
    .b(_al_u622_o),
    .c(_al_u623_o),
    .d(vga_rdaddr_piped_piped[3]),
    .o(_al_u627_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'h00ac))
    _al_u628 (
    .a(_al_u621_o),
    .b(_al_u627_o),
    .c(vga_rdaddr_piped_piped[4]),
    .d(vga_rdaddr_piped_piped[5]),
    .o(_al_u628_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*~A))"),
    .INIT(8'h8c))
    _al_u629 (
    .a(\u_img/inst_dob_i64_004 ),
    .b(vga_rden),
    .c(vga_rdaddr_piped_piped[6]),
    .o(_al_u629_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(~D*~(~B*~A)))"),
    .INIT(16'hf010))
    _al_u630 (
    .a(_al_u615_o),
    .b(_al_u628_o),
    .c(_al_u629_o),
    .d(vga_rdaddr_piped_piped[6]),
    .o(vga_b_pad[7]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u631 (
    .a(\u_img/inst_dob_i8_003 ),
    .b(\u_img/inst_dob_i10_003 ),
    .c(vga_rdaddr_piped_piped[1]),
    .o(_al_u631_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u632 (
    .a(\u_img/inst_dob_i12_003 ),
    .b(\u_img/inst_dob_i14_003 ),
    .c(vga_rdaddr_piped_piped[1]),
    .o(_al_u632_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'hca00))
    _al_u633 (
    .a(_al_u631_o),
    .b(_al_u632_o),
    .c(vga_rdaddr_piped_piped[2]),
    .d(vga_rdaddr_piped_piped[3]),
    .o(_al_u633_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'hca00))
    _al_u634 (
    .a(\u_img/inst_dob_i4_003 ),
    .b(\u_img/inst_dob_i6_003 ),
    .c(vga_rdaddr_piped_piped[1]),
    .d(vga_rdaddr_piped_piped[2]),
    .o(_al_u634_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h00ca))
    _al_u635 (
    .a(\u_img/inst_dob_i0_003 ),
    .b(\u_img/inst_dob_i2_003 ),
    .c(vga_rdaddr_piped_piped[1]),
    .d(vga_rdaddr_piped_piped[2]),
    .o(_al_u635_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(~C*~B*~A))"),
    .INIT(16'h00fe))
    _al_u636 (
    .a(_al_u634_o),
    .b(_al_u635_o),
    .c(vga_rdaddr_piped_piped[3]),
    .d(vga_rdaddr_piped_piped[4]),
    .o(_al_u636_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u637 (
    .a(\u_img/inst_dob_i20_003 ),
    .b(\u_img/inst_dob_i22_003 ),
    .c(vga_rdaddr_piped_piped[1]),
    .o(_al_u637_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u638 (
    .a(\u_img/inst_dob_i16_003 ),
    .b(\u_img/inst_dob_i18_003 ),
    .c(vga_rdaddr_piped_piped[1]),
    .o(_al_u638_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'h00ac))
    _al_u639 (
    .a(_al_u637_o),
    .b(_al_u638_o),
    .c(vga_rdaddr_piped_piped[2]),
    .d(vga_rdaddr_piped_piped[3]),
    .o(_al_u639_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h00ca))
    _al_u640 (
    .a(\u_img/inst_dob_i24_003 ),
    .b(\u_img/inst_dob_i26_003 ),
    .c(vga_rdaddr_piped_piped[1]),
    .d(vga_rdaddr_piped_piped[2]),
    .o(_al_u640_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'hca00))
    _al_u641 (
    .a(\u_img/inst_dob_i28_003 ),
    .b(\u_img/inst_dob_i30_003 ),
    .c(vga_rdaddr_piped_piped[1]),
    .d(vga_rdaddr_piped_piped[2]),
    .o(_al_u641_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C*~B*~A))"),
    .INIT(16'hef00))
    _al_u642 (
    .a(_al_u640_o),
    .b(_al_u641_o),
    .c(vga_rdaddr_piped_piped[3]),
    .d(vga_rdaddr_piped_piped[4]),
    .o(_al_u642_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~C)*~(B*~A))"),
    .INIT(16'hb0bb))
    _al_u643 (
    .a(_al_u633_o),
    .b(_al_u636_o),
    .c(_al_u639_o),
    .d(_al_u642_o),
    .o(_al_u643_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u644 (
    .a(\u_img/inst_dob_i36_003 ),
    .b(\u_img/inst_dob_i38_003 ),
    .c(vga_rdaddr_piped_piped[1]),
    .o(_al_u644_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u645 (
    .a(\u_img/inst_dob_i32_003 ),
    .b(\u_img/inst_dob_i34_003 ),
    .c(vga_rdaddr_piped_piped[1]),
    .o(_al_u645_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'h00ac))
    _al_u646 (
    .a(_al_u644_o),
    .b(_al_u645_o),
    .c(vga_rdaddr_piped_piped[2]),
    .d(vga_rdaddr_piped_piped[3]),
    .o(_al_u646_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'hca00))
    _al_u647 (
    .a(\u_img/inst_dob_i44_003 ),
    .b(\u_img/inst_dob_i46_003 ),
    .c(vga_rdaddr_piped_piped[1]),
    .d(vga_rdaddr_piped_piped[2]),
    .o(_al_u647_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h00ca))
    _al_u648 (
    .a(\u_img/inst_dob_i40_003 ),
    .b(\u_img/inst_dob_i42_003 ),
    .c(vga_rdaddr_piped_piped[1]),
    .d(vga_rdaddr_piped_piped[2]),
    .o(_al_u648_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(C*~B*~A))"),
    .INIT(16'h00ef))
    _al_u649 (
    .a(_al_u647_o),
    .b(_al_u648_o),
    .c(vga_rdaddr_piped_piped[3]),
    .d(vga_rdaddr_piped_piped[4]),
    .o(_al_u649_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u650 (
    .a(\u_img/inst_dob_i52_003 ),
    .b(\u_img/inst_dob_i54_003 ),
    .c(vga_rdaddr_piped_piped[1]),
    .o(_al_u650_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u651 (
    .a(\u_img/inst_dob_i48_003 ),
    .b(\u_img/inst_dob_i50_003 ),
    .c(vga_rdaddr_piped_piped[1]),
    .o(_al_u651_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'h00ac))
    _al_u652 (
    .a(_al_u650_o),
    .b(_al_u651_o),
    .c(vga_rdaddr_piped_piped[2]),
    .d(vga_rdaddr_piped_piped[3]),
    .o(_al_u652_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h00ca))
    _al_u653 (
    .a(\u_img/inst_dob_i56_003 ),
    .b(\u_img/inst_dob_i58_003 ),
    .c(vga_rdaddr_piped_piped[1]),
    .d(vga_rdaddr_piped_piped[2]),
    .o(_al_u653_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'hca00))
    _al_u654 (
    .a(\u_img/inst_dob_i60_003 ),
    .b(\u_img/inst_dob_i62_003 ),
    .c(vga_rdaddr_piped_piped[1]),
    .d(vga_rdaddr_piped_piped[2]),
    .o(_al_u654_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C*~B*~A))"),
    .INIT(16'hef00))
    _al_u655 (
    .a(_al_u653_o),
    .b(_al_u654_o),
    .c(vga_rdaddr_piped_piped[3]),
    .d(vga_rdaddr_piped_piped[4]),
    .o(_al_u655_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~C)*~(B*~A))"),
    .INIT(16'hb0bb))
    _al_u656 (
    .a(_al_u646_o),
    .b(_al_u649_o),
    .c(_al_u652_o),
    .d(_al_u655_o),
    .o(_al_u656_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h00ca))
    _al_u657 (
    .a(_al_u643_o),
    .b(_al_u656_o),
    .c(vga_rdaddr_piped_piped[5]),
    .d(vga_rdaddr_piped_piped[6]),
    .o(_al_u657_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*~(D*~B))"),
    .INIT(16'h4050))
    _al_u658 (
    .a(_al_u657_o),
    .b(\u_img/inst_dob_i64_003 ),
    .c(vga_rden),
    .d(vga_rdaddr_piped_piped[6]),
    .o(vga_b_pad[6]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u659 (
    .a(\u_img/inst_dob_i4_002 ),
    .b(\u_img/inst_dob_i6_002 ),
    .c(vga_rdaddr_piped_piped[1]),
    .o(_al_u659_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u660 (
    .a(\u_img/inst_dob_i0_002 ),
    .b(\u_img/inst_dob_i2_002 ),
    .c(vga_rdaddr_piped_piped[1]),
    .o(_al_u660_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'h00ac))
    _al_u661 (
    .a(_al_u659_o),
    .b(_al_u660_o),
    .c(vga_rdaddr_piped_piped[2]),
    .d(vga_rdaddr_piped_piped[3]),
    .o(_al_u661_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'hca00))
    _al_u662 (
    .a(\u_img/inst_dob_i12_002 ),
    .b(\u_img/inst_dob_i14_002 ),
    .c(vga_rdaddr_piped_piped[1]),
    .d(vga_rdaddr_piped_piped[2]),
    .o(_al_u662_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h00ca))
    _al_u663 (
    .a(\u_img/inst_dob_i8_002 ),
    .b(\u_img/inst_dob_i10_002 ),
    .c(vga_rdaddr_piped_piped[1]),
    .d(vga_rdaddr_piped_piped[2]),
    .o(_al_u663_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(C*~B*~A))"),
    .INIT(16'h00ef))
    _al_u664 (
    .a(_al_u662_o),
    .b(_al_u663_o),
    .c(vga_rdaddr_piped_piped[3]),
    .d(vga_rdaddr_piped_piped[4]),
    .o(_al_u664_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u665 (
    .a(\u_img/inst_dob_i20_002 ),
    .b(\u_img/inst_dob_i22_002 ),
    .c(vga_rdaddr_piped_piped[1]),
    .o(_al_u665_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u666 (
    .a(\u_img/inst_dob_i16_002 ),
    .b(\u_img/inst_dob_i18_002 ),
    .c(vga_rdaddr_piped_piped[1]),
    .o(_al_u666_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'h00ac))
    _al_u667 (
    .a(_al_u665_o),
    .b(_al_u666_o),
    .c(vga_rdaddr_piped_piped[2]),
    .d(vga_rdaddr_piped_piped[3]),
    .o(_al_u667_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h00ca))
    _al_u668 (
    .a(\u_img/inst_dob_i24_002 ),
    .b(\u_img/inst_dob_i26_002 ),
    .c(vga_rdaddr_piped_piped[1]),
    .d(vga_rdaddr_piped_piped[2]),
    .o(_al_u668_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'hca00))
    _al_u669 (
    .a(\u_img/inst_dob_i28_002 ),
    .b(\u_img/inst_dob_i30_002 ),
    .c(vga_rdaddr_piped_piped[1]),
    .d(vga_rdaddr_piped_piped[2]),
    .o(_al_u669_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C*~B*~A))"),
    .INIT(16'hef00))
    _al_u670 (
    .a(_al_u668_o),
    .b(_al_u669_o),
    .c(vga_rdaddr_piped_piped[3]),
    .d(vga_rdaddr_piped_piped[4]),
    .o(_al_u670_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~C)*~(B*~A))"),
    .INIT(16'hb0bb))
    _al_u671 (
    .a(_al_u661_o),
    .b(_al_u664_o),
    .c(_al_u667_o),
    .d(_al_u670_o),
    .o(_al_u671_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u672 (
    .a(\u_img/inst_dob_i36_002 ),
    .b(\u_img/inst_dob_i38_002 ),
    .c(vga_rdaddr_piped_piped[1]),
    .o(_al_u672_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u673 (
    .a(\u_img/inst_dob_i32_002 ),
    .b(\u_img/inst_dob_i34_002 ),
    .c(vga_rdaddr_piped_piped[1]),
    .o(_al_u673_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'h00ac))
    _al_u674 (
    .a(_al_u672_o),
    .b(_al_u673_o),
    .c(vga_rdaddr_piped_piped[2]),
    .d(vga_rdaddr_piped_piped[3]),
    .o(_al_u674_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'hca00))
    _al_u675 (
    .a(\u_img/inst_dob_i44_002 ),
    .b(\u_img/inst_dob_i46_002 ),
    .c(vga_rdaddr_piped_piped[1]),
    .d(vga_rdaddr_piped_piped[2]),
    .o(_al_u675_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h00ca))
    _al_u676 (
    .a(\u_img/inst_dob_i40_002 ),
    .b(\u_img/inst_dob_i42_002 ),
    .c(vga_rdaddr_piped_piped[1]),
    .d(vga_rdaddr_piped_piped[2]),
    .o(_al_u676_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(C*~B*~A))"),
    .INIT(16'h00ef))
    _al_u677 (
    .a(_al_u675_o),
    .b(_al_u676_o),
    .c(vga_rdaddr_piped_piped[3]),
    .d(vga_rdaddr_piped_piped[4]),
    .o(_al_u677_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u678 (
    .a(\u_img/inst_dob_i60_002 ),
    .b(\u_img/inst_dob_i62_002 ),
    .c(vga_rdaddr_piped_piped[1]),
    .o(_al_u678_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u679 (
    .a(\u_img/inst_dob_i56_002 ),
    .b(\u_img/inst_dob_i58_002 ),
    .c(vga_rdaddr_piped_piped[1]),
    .o(_al_u679_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'hac00))
    _al_u680 (
    .a(_al_u678_o),
    .b(_al_u679_o),
    .c(vga_rdaddr_piped_piped[2]),
    .d(vga_rdaddr_piped_piped[3]),
    .o(_al_u680_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'hca00))
    _al_u681 (
    .a(\u_img/inst_dob_i52_002 ),
    .b(\u_img/inst_dob_i54_002 ),
    .c(vga_rdaddr_piped_piped[1]),
    .d(vga_rdaddr_piped_piped[2]),
    .o(_al_u681_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h00ca))
    _al_u682 (
    .a(\u_img/inst_dob_i48_002 ),
    .b(\u_img/inst_dob_i50_002 ),
    .c(vga_rdaddr_piped_piped[1]),
    .d(vga_rdaddr_piped_piped[2]),
    .o(_al_u682_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(~C*~B*~A))"),
    .INIT(16'hfe00))
    _al_u683 (
    .a(_al_u681_o),
    .b(_al_u682_o),
    .c(vga_rdaddr_piped_piped[3]),
    .d(vga_rdaddr_piped_piped[4]),
    .o(_al_u683_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~C)*~(B*~A))"),
    .INIT(16'hb0bb))
    _al_u684 (
    .a(_al_u674_o),
    .b(_al_u677_o),
    .c(_al_u680_o),
    .d(_al_u683_o),
    .o(_al_u684_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h00ca))
    _al_u685 (
    .a(_al_u671_o),
    .b(_al_u684_o),
    .c(vga_rdaddr_piped_piped[5]),
    .d(vga_rdaddr_piped_piped[6]),
    .o(_al_u685_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*~(D*~B))"),
    .INIT(16'h4050))
    _al_u686 (
    .a(_al_u685_o),
    .b(\u_img/inst_dob_i64_002 ),
    .c(vga_rden),
    .d(vga_rdaddr_piped_piped[6]),
    .o(vga_b_pad[5]));
  AL_MAP_LUT4 #(
    .EQN("(~D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h00ca))
    _al_u687 (
    .a(\u_img/inst_dob_i0_015 ),
    .b(\u_img/inst_dob_i16_015 ),
    .c(vga_rdaddr_piped_piped[4]),
    .d(vga_rdaddr_piped_piped[5]),
    .o(_al_u687_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'hca00))
    _al_u688 (
    .a(\u_img/inst_dob_i32_015 ),
    .b(\u_img/inst_dob_i48_015 ),
    .c(vga_rdaddr_piped_piped[4]),
    .d(vga_rdaddr_piped_piped[5]),
    .o(_al_u688_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*~A))"),
    .INIT(8'h8c))
    _al_u689 (
    .a(\u_img/inst_dob_i64_015 ),
    .b(vga_rden),
    .c(vga_rdaddr_piped_piped[6]),
    .o(_al_u689_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(~D*~B*~A))"),
    .INIT(16'hf0e0))
    _al_u690 (
    .a(_al_u687_o),
    .b(_al_u688_o),
    .c(_al_u689_o),
    .d(vga_rdaddr_piped_piped[6]),
    .o(vga_r_pad[7]));
  AL_MAP_LUT4 #(
    .EQN("(~D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h00ca))
    _al_u691 (
    .a(\u_img/inst_dob_i0_014 ),
    .b(\u_img/inst_dob_i16_014 ),
    .c(vga_rdaddr_piped_piped[4]),
    .d(vga_rdaddr_piped_piped[5]),
    .o(_al_u691_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'hca00))
    _al_u692 (
    .a(\u_img/inst_dob_i32_014 ),
    .b(\u_img/inst_dob_i48_014 ),
    .c(vga_rdaddr_piped_piped[4]),
    .d(vga_rdaddr_piped_piped[5]),
    .o(_al_u692_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*~A))"),
    .INIT(8'h8c))
    _al_u693 (
    .a(\u_img/inst_dob_i64_014 ),
    .b(vga_rden),
    .c(vga_rdaddr_piped_piped[6]),
    .o(_al_u693_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(~D*~B*~A))"),
    .INIT(16'hf0e0))
    _al_u694 (
    .a(_al_u691_o),
    .b(_al_u692_o),
    .c(_al_u693_o),
    .d(vga_rdaddr_piped_piped[6]),
    .o(vga_r_pad[6]));
  AL_MAP_LUT4 #(
    .EQN("(~D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h00ca))
    _al_u695 (
    .a(\u_img/inst_dob_i0_013 ),
    .b(\u_img/inst_dob_i16_013 ),
    .c(vga_rdaddr_piped_piped[4]),
    .d(vga_rdaddr_piped_piped[5]),
    .o(_al_u695_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'hca00))
    _al_u696 (
    .a(\u_img/inst_dob_i32_013 ),
    .b(\u_img/inst_dob_i48_013 ),
    .c(vga_rdaddr_piped_piped[4]),
    .d(vga_rdaddr_piped_piped[5]),
    .o(_al_u696_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*~A))"),
    .INIT(8'h8c))
    _al_u697 (
    .a(\u_img/inst_dob_i64_013 ),
    .b(vga_rden),
    .c(vga_rdaddr_piped_piped[6]),
    .o(_al_u697_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(~D*~B*~A))"),
    .INIT(16'hf0e0))
    _al_u698 (
    .a(_al_u695_o),
    .b(_al_u696_o),
    .c(_al_u697_o),
    .d(vga_rdaddr_piped_piped[6]),
    .o(vga_r_pad[5]));
  AL_MAP_LUT4 #(
    .EQN("(~D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h00ca))
    _al_u699 (
    .a(\u_img/inst_dob_i0_012 ),
    .b(\u_img/inst_dob_i16_012 ),
    .c(vga_rdaddr_piped_piped[4]),
    .d(vga_rdaddr_piped_piped[5]),
    .o(_al_u699_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'hca00))
    _al_u700 (
    .a(\u_img/inst_dob_i32_012 ),
    .b(\u_img/inst_dob_i48_012 ),
    .c(vga_rdaddr_piped_piped[4]),
    .d(vga_rdaddr_piped_piped[5]),
    .o(_al_u700_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*~A))"),
    .INIT(8'h8c))
    _al_u701 (
    .a(\u_img/inst_dob_i64_012 ),
    .b(vga_rden),
    .c(vga_rdaddr_piped_piped[6]),
    .o(_al_u701_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(~D*~B*~A))"),
    .INIT(16'hf0e0))
    _al_u702 (
    .a(_al_u699_o),
    .b(_al_u700_o),
    .c(_al_u701_o),
    .d(vga_rdaddr_piped_piped[6]),
    .o(vga_r_pad[4]));
  AL_MAP_LUT4 #(
    .EQN("(~D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h00ca))
    _al_u703 (
    .a(\u_img/inst_dob_i0_011 ),
    .b(\u_img/inst_dob_i16_011 ),
    .c(vga_rdaddr_piped_piped[4]),
    .d(vga_rdaddr_piped_piped[5]),
    .o(_al_u703_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'hca00))
    _al_u704 (
    .a(\u_img/inst_dob_i32_011 ),
    .b(\u_img/inst_dob_i48_011 ),
    .c(vga_rdaddr_piped_piped[4]),
    .d(vga_rdaddr_piped_piped[5]),
    .o(_al_u704_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*~A))"),
    .INIT(8'h8c))
    _al_u705 (
    .a(\u_img/inst_dob_i64_011 ),
    .b(vga_rden),
    .c(vga_rdaddr_piped_piped[6]),
    .o(_al_u705_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(~D*~B*~A))"),
    .INIT(16'hf0e0))
    _al_u706 (
    .a(_al_u703_o),
    .b(_al_u704_o),
    .c(_al_u705_o),
    .d(vga_rdaddr_piped_piped[6]),
    .o(vga_r_pad[3]));
  AL_MAP_LUT4 #(
    .EQN("(~D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h00ca))
    _al_u707 (
    .a(\u_img/inst_dob_i0_010 ),
    .b(\u_img/inst_dob_i16_010 ),
    .c(vga_rdaddr_piped_piped[4]),
    .d(vga_rdaddr_piped_piped[5]),
    .o(_al_u707_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'hca00))
    _al_u708 (
    .a(\u_img/inst_dob_i32_010 ),
    .b(\u_img/inst_dob_i48_010 ),
    .c(vga_rdaddr_piped_piped[4]),
    .d(vga_rdaddr_piped_piped[5]),
    .o(_al_u708_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*~A))"),
    .INIT(8'h8c))
    _al_u709 (
    .a(\u_img/inst_dob_i64_010 ),
    .b(vga_rden),
    .c(vga_rdaddr_piped_piped[6]),
    .o(_al_u709_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(~D*~B*~A))"),
    .INIT(16'hf0e0))
    _al_u710 (
    .a(_al_u707_o),
    .b(_al_u708_o),
    .c(_al_u709_o),
    .d(vga_rdaddr_piped_piped[6]),
    .o(vga_g_pad[7]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u711 (
    .a(\u_img/inst_dob_i36_001 ),
    .b(\u_img/inst_dob_i38_001 ),
    .c(vga_rdaddr_piped_piped[1]),
    .o(_al_u711_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u712 (
    .a(\u_img/inst_dob_i32_001 ),
    .b(\u_img/inst_dob_i34_001 ),
    .c(vga_rdaddr_piped_piped[1]),
    .o(_al_u712_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'h00ac))
    _al_u713 (
    .a(_al_u711_o),
    .b(_al_u712_o),
    .c(vga_rdaddr_piped_piped[2]),
    .d(vga_rdaddr_piped_piped[3]),
    .o(_al_u713_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'hca00))
    _al_u714 (
    .a(\u_img/inst_dob_i44_001 ),
    .b(\u_img/inst_dob_i46_001 ),
    .c(vga_rdaddr_piped_piped[1]),
    .d(vga_rdaddr_piped_piped[2]),
    .o(_al_u714_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h00ca))
    _al_u715 (
    .a(\u_img/inst_dob_i40_001 ),
    .b(\u_img/inst_dob_i42_001 ),
    .c(vga_rdaddr_piped_piped[1]),
    .d(vga_rdaddr_piped_piped[2]),
    .o(_al_u715_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(C*~B*~A))"),
    .INIT(16'h00ef))
    _al_u716 (
    .a(_al_u714_o),
    .b(_al_u715_o),
    .c(vga_rdaddr_piped_piped[3]),
    .d(vga_rdaddr_piped_piped[4]),
    .o(_al_u716_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u717 (
    .a(\u_img/inst_dob_i52_001 ),
    .b(\u_img/inst_dob_i54_001 ),
    .c(vga_rdaddr_piped_piped[1]),
    .o(_al_u717_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u718 (
    .a(\u_img/inst_dob_i48_001 ),
    .b(\u_img/inst_dob_i50_001 ),
    .c(vga_rdaddr_piped_piped[1]),
    .o(_al_u718_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'h00ac))
    _al_u719 (
    .a(_al_u717_o),
    .b(_al_u718_o),
    .c(vga_rdaddr_piped_piped[2]),
    .d(vga_rdaddr_piped_piped[3]),
    .o(_al_u719_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h00ca))
    _al_u720 (
    .a(\u_img/inst_dob_i56_001 ),
    .b(\u_img/inst_dob_i58_001 ),
    .c(vga_rdaddr_piped_piped[1]),
    .d(vga_rdaddr_piped_piped[2]),
    .o(_al_u720_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'hca00))
    _al_u721 (
    .a(\u_img/inst_dob_i60_001 ),
    .b(\u_img/inst_dob_i62_001 ),
    .c(vga_rdaddr_piped_piped[1]),
    .d(vga_rdaddr_piped_piped[2]),
    .o(_al_u721_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C*~B*~A))"),
    .INIT(16'hef00))
    _al_u722 (
    .a(_al_u720_o),
    .b(_al_u721_o),
    .c(vga_rdaddr_piped_piped[3]),
    .d(vga_rdaddr_piped_piped[4]),
    .o(_al_u722_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~C)*~(B*~A))"),
    .INIT(16'hb0bb))
    _al_u723 (
    .a(_al_u713_o),
    .b(_al_u716_o),
    .c(_al_u719_o),
    .d(_al_u722_o),
    .o(_al_u723_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u724 (
    .a(\u_img/inst_dob_i4_001 ),
    .b(\u_img/inst_dob_i6_001 ),
    .c(vga_rdaddr_piped_piped[1]),
    .o(_al_u724_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u725 (
    .a(\u_img/inst_dob_i0_001 ),
    .b(\u_img/inst_dob_i2_001 ),
    .c(vga_rdaddr_piped_piped[1]),
    .o(_al_u725_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'h00ac))
    _al_u726 (
    .a(_al_u724_o),
    .b(_al_u725_o),
    .c(vga_rdaddr_piped_piped[2]),
    .d(vga_rdaddr_piped_piped[3]),
    .o(_al_u726_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'hca00))
    _al_u727 (
    .a(\u_img/inst_dob_i12_001 ),
    .b(\u_img/inst_dob_i14_001 ),
    .c(vga_rdaddr_piped_piped[1]),
    .d(vga_rdaddr_piped_piped[2]),
    .o(_al_u727_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h00ca))
    _al_u728 (
    .a(\u_img/inst_dob_i8_001 ),
    .b(\u_img/inst_dob_i10_001 ),
    .c(vga_rdaddr_piped_piped[1]),
    .d(vga_rdaddr_piped_piped[2]),
    .o(_al_u728_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(C*~B*~A))"),
    .INIT(16'h00ef))
    _al_u729 (
    .a(_al_u727_o),
    .b(_al_u728_o),
    .c(vga_rdaddr_piped_piped[3]),
    .d(vga_rdaddr_piped_piped[4]),
    .o(_al_u729_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u730 (
    .a(\u_img/inst_dob_i20_001 ),
    .b(\u_img/inst_dob_i22_001 ),
    .c(vga_rdaddr_piped_piped[1]),
    .o(_al_u730_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u731 (
    .a(\u_img/inst_dob_i16_001 ),
    .b(\u_img/inst_dob_i18_001 ),
    .c(vga_rdaddr_piped_piped[1]),
    .o(_al_u731_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'h00ac))
    _al_u732 (
    .a(_al_u730_o),
    .b(_al_u731_o),
    .c(vga_rdaddr_piped_piped[2]),
    .d(vga_rdaddr_piped_piped[3]),
    .o(_al_u732_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h00ca))
    _al_u733 (
    .a(\u_img/inst_dob_i24_001 ),
    .b(\u_img/inst_dob_i26_001 ),
    .c(vga_rdaddr_piped_piped[1]),
    .d(vga_rdaddr_piped_piped[2]),
    .o(_al_u733_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'hca00))
    _al_u734 (
    .a(\u_img/inst_dob_i28_001 ),
    .b(\u_img/inst_dob_i30_001 ),
    .c(vga_rdaddr_piped_piped[1]),
    .d(vga_rdaddr_piped_piped[2]),
    .o(_al_u734_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C*~B*~A))"),
    .INIT(16'hef00))
    _al_u735 (
    .a(_al_u733_o),
    .b(_al_u734_o),
    .c(vga_rdaddr_piped_piped[3]),
    .d(vga_rdaddr_piped_piped[4]),
    .o(_al_u735_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~C)*~(B*~A))"),
    .INIT(16'hb0bb))
    _al_u736 (
    .a(_al_u726_o),
    .b(_al_u729_o),
    .c(_al_u732_o),
    .d(_al_u735_o),
    .o(_al_u736_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'h00ac))
    _al_u737 (
    .a(_al_u723_o),
    .b(_al_u736_o),
    .c(vga_rdaddr_piped_piped[5]),
    .d(vga_rdaddr_piped_piped[6]),
    .o(_al_u737_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*~(D*~B))"),
    .INIT(16'h4050))
    _al_u738 (
    .a(_al_u737_o),
    .b(\u_img/inst_dob_i64_001 ),
    .c(vga_rden),
    .d(vga_rdaddr_piped_piped[6]),
    .o(vga_b_pad[4]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u739 (
    .a(\u_img/inst_dob_i36_000 ),
    .b(\u_img/inst_dob_i38_000 ),
    .c(vga_rdaddr_piped_piped[1]),
    .o(_al_u739_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u740 (
    .a(\u_img/inst_dob_i32_000 ),
    .b(\u_img/inst_dob_i34_000 ),
    .c(vga_rdaddr_piped_piped[1]),
    .o(_al_u740_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'h00ac))
    _al_u741 (
    .a(_al_u739_o),
    .b(_al_u740_o),
    .c(vga_rdaddr_piped_piped[2]),
    .d(vga_rdaddr_piped_piped[3]),
    .o(_al_u741_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'hca00))
    _al_u742 (
    .a(\u_img/inst_dob_i44_000 ),
    .b(\u_img/inst_dob_i46_000 ),
    .c(vga_rdaddr_piped_piped[1]),
    .d(vga_rdaddr_piped_piped[2]),
    .o(_al_u742_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h00ca))
    _al_u743 (
    .a(\u_img/inst_dob_i40_000 ),
    .b(\u_img/inst_dob_i42_000 ),
    .c(vga_rdaddr_piped_piped[1]),
    .d(vga_rdaddr_piped_piped[2]),
    .o(_al_u743_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(C*~B*~A))"),
    .INIT(16'h00ef))
    _al_u744 (
    .a(_al_u742_o),
    .b(_al_u743_o),
    .c(vga_rdaddr_piped_piped[3]),
    .d(vga_rdaddr_piped_piped[4]),
    .o(_al_u744_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u745 (
    .a(\u_img/inst_dob_i52_000 ),
    .b(\u_img/inst_dob_i54_000 ),
    .c(vga_rdaddr_piped_piped[1]),
    .o(_al_u745_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u746 (
    .a(\u_img/inst_dob_i48_000 ),
    .b(\u_img/inst_dob_i50_000 ),
    .c(vga_rdaddr_piped_piped[1]),
    .o(_al_u746_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'h00ac))
    _al_u747 (
    .a(_al_u745_o),
    .b(_al_u746_o),
    .c(vga_rdaddr_piped_piped[2]),
    .d(vga_rdaddr_piped_piped[3]),
    .o(_al_u747_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'hca00))
    _al_u748 (
    .a(\u_img/inst_dob_i60_000 ),
    .b(\u_img/inst_dob_i62_000 ),
    .c(vga_rdaddr_piped_piped[1]),
    .d(vga_rdaddr_piped_piped[2]),
    .o(_al_u748_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h00ca))
    _al_u749 (
    .a(\u_img/inst_dob_i56_000 ),
    .b(\u_img/inst_dob_i58_000 ),
    .c(vga_rdaddr_piped_piped[1]),
    .d(vga_rdaddr_piped_piped[2]),
    .o(_al_u749_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C*~B*~A))"),
    .INIT(16'hef00))
    _al_u750 (
    .a(_al_u748_o),
    .b(_al_u749_o),
    .c(vga_rdaddr_piped_piped[3]),
    .d(vga_rdaddr_piped_piped[4]),
    .o(_al_u750_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~C)*~(B*~A))"),
    .INIT(16'hb0bb))
    _al_u751 (
    .a(_al_u741_o),
    .b(_al_u744_o),
    .c(_al_u747_o),
    .d(_al_u750_o),
    .o(_al_u751_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u752 (
    .a(\u_img/inst_dob_i4_000 ),
    .b(\u_img/inst_dob_i6_000 ),
    .c(vga_rdaddr_piped_piped[1]),
    .o(_al_u752_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u753 (
    .a(\u_img/inst_dob_i0_000 ),
    .b(\u_img/inst_dob_i2_000 ),
    .c(vga_rdaddr_piped_piped[1]),
    .o(_al_u753_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'h00ac))
    _al_u754 (
    .a(_al_u752_o),
    .b(_al_u753_o),
    .c(vga_rdaddr_piped_piped[2]),
    .d(vga_rdaddr_piped_piped[3]),
    .o(_al_u754_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'hca00))
    _al_u755 (
    .a(\u_img/inst_dob_i12_000 ),
    .b(\u_img/inst_dob_i14_000 ),
    .c(vga_rdaddr_piped_piped[1]),
    .d(vga_rdaddr_piped_piped[2]),
    .o(_al_u755_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h00ca))
    _al_u756 (
    .a(\u_img/inst_dob_i8_000 ),
    .b(\u_img/inst_dob_i10_000 ),
    .c(vga_rdaddr_piped_piped[1]),
    .d(vga_rdaddr_piped_piped[2]),
    .o(_al_u756_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(C*~B*~A))"),
    .INIT(16'h00ef))
    _al_u757 (
    .a(_al_u755_o),
    .b(_al_u756_o),
    .c(vga_rdaddr_piped_piped[3]),
    .d(vga_rdaddr_piped_piped[4]),
    .o(_al_u757_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u758 (
    .a(\u_img/inst_dob_i28_000 ),
    .b(\u_img/inst_dob_i30_000 ),
    .c(vga_rdaddr_piped_piped[1]),
    .o(_al_u758_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u759 (
    .a(\u_img/inst_dob_i24_000 ),
    .b(\u_img/inst_dob_i26_000 ),
    .c(vga_rdaddr_piped_piped[1]),
    .o(_al_u759_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'hac00))
    _al_u760 (
    .a(_al_u758_o),
    .b(_al_u759_o),
    .c(vga_rdaddr_piped_piped[2]),
    .d(vga_rdaddr_piped_piped[3]),
    .o(_al_u760_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'hca00))
    _al_u761 (
    .a(\u_img/inst_dob_i20_000 ),
    .b(\u_img/inst_dob_i22_000 ),
    .c(vga_rdaddr_piped_piped[1]),
    .d(vga_rdaddr_piped_piped[2]),
    .o(_al_u761_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h00ca))
    _al_u762 (
    .a(\u_img/inst_dob_i16_000 ),
    .b(\u_img/inst_dob_i18_000 ),
    .c(vga_rdaddr_piped_piped[1]),
    .d(vga_rdaddr_piped_piped[2]),
    .o(_al_u762_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(~C*~B*~A))"),
    .INIT(16'hfe00))
    _al_u763 (
    .a(_al_u761_o),
    .b(_al_u762_o),
    .c(vga_rdaddr_piped_piped[3]),
    .d(vga_rdaddr_piped_piped[4]),
    .o(_al_u763_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~C)*~(B*~A))"),
    .INIT(16'hb0bb))
    _al_u764 (
    .a(_al_u754_o),
    .b(_al_u757_o),
    .c(_al_u760_o),
    .d(_al_u763_o),
    .o(_al_u764_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'h00ac))
    _al_u765 (
    .a(_al_u751_o),
    .b(_al_u764_o),
    .c(vga_rdaddr_piped_piped[5]),
    .d(vga_rdaddr_piped_piped[6]),
    .o(_al_u765_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*~(D*~B))"),
    .INIT(16'h4050))
    _al_u766 (
    .a(_al_u765_o),
    .b(\u_img/inst_dob_i64_000 ),
    .c(vga_rden),
    .d(vga_rdaddr_piped_piped[6]),
    .o(vga_b_pad[3]));
  AL_MAP_LUT1 #(
    .EQN("(~A)"),
    .INIT(2'h1))
    _al_u767 (
    .a(cam_rst_pad),
    .o(cam_rst_pad_neg));
  AL_MAP_LUT1 #(
    .EQN("(~A)"),
    .INIT(2'h1))
    _al_u768 (
    .a(\u_camera_reader/wrclk1 ),
    .o(\u_camera_reader/n1 ));
  EG_PHY_CONFIG #(
    .DONE_PERSISTN("ENABLE"),
    .INIT_PERSISTN("ENABLE"),
    .JTAG_PERSISTN("DISABLE"),
    .PROGRAMN_PERSISTN("DISABLE"))
    config_inst ();
  camera_init u_camera_init (
    .clk(clk_sccb),
    .reset_n(cam_rst_pad),
    .sda_in(cam_soid_pad),
    .scl(cam_soic),
    .sda(sda),
    .sda_oe(sda_oe));  // sources/rtl/test_camera.v(84)
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_camera_reader/add0/u0  (
    .a(\u_camera_reader/pixel_counter [0]),
    .b(1'b1),
    .c(\u_camera_reader/add0/c0 ),
    .o({\u_camera_reader/add0/c1 ,\u_camera_reader/n8 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_camera_reader/add0/u1  (
    .a(\u_camera_reader/pixel_counter [1]),
    .b(1'b0),
    .c(\u_camera_reader/add0/c1 ),
    .o({\u_camera_reader/add0/c2 ,\u_camera_reader/n8 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_camera_reader/add0/u10  (
    .a(\u_camera_reader/pixel_counter [10]),
    .b(1'b0),
    .c(\u_camera_reader/add0/c10 ),
    .o({\u_camera_reader/add0/c11 ,\u_camera_reader/n8 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_camera_reader/add0/u11  (
    .a(\u_camera_reader/pixel_counter [11]),
    .b(1'b0),
    .c(\u_camera_reader/add0/c11 ),
    .o({\u_camera_reader/add0/c12 ,\u_camera_reader/n8 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_camera_reader/add0/u12  (
    .a(\u_camera_reader/pixel_counter [12]),
    .b(1'b0),
    .c(\u_camera_reader/add0/c12 ),
    .o({\u_camera_reader/add0/c13 ,\u_camera_reader/n8 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_camera_reader/add0/u13  (
    .a(\u_camera_reader/pixel_counter [13]),
    .b(1'b0),
    .c(\u_camera_reader/add0/c13 ),
    .o({\u_camera_reader/add0/c14 ,\u_camera_reader/n8 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_camera_reader/add0/u14  (
    .a(\u_camera_reader/pixel_counter [14]),
    .b(1'b0),
    .c(\u_camera_reader/add0/c14 ),
    .o({\u_camera_reader/add0/c15 ,\u_camera_reader/n8 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_camera_reader/add0/u15  (
    .a(\u_camera_reader/pixel_counter [15]),
    .b(1'b0),
    .c(\u_camera_reader/add0/c15 ),
    .o({\u_camera_reader/add0/c16 ,\u_camera_reader/n8 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_camera_reader/add0/u16  (
    .a(\u_camera_reader/pixel_counter [16]),
    .b(1'b0),
    .c(\u_camera_reader/add0/c16 ),
    .o({\u_camera_reader/add0/c17 ,\u_camera_reader/n8 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_camera_reader/add0/u17  (
    .a(\u_camera_reader/pixel_counter [17]),
    .b(1'b0),
    .c(\u_camera_reader/add0/c17 ),
    .o({\u_camera_reader/add0/c18 ,\u_camera_reader/n8 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_camera_reader/add0/u18  (
    .a(\u_camera_reader/pixel_counter [18]),
    .b(1'b0),
    .c(\u_camera_reader/add0/c18 ),
    .o({\u_camera_reader/add0/c19 ,\u_camera_reader/n8 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_camera_reader/add0/u19  (
    .a(\u_camera_reader/pixel_counter [19]),
    .b(1'b0),
    .c(\u_camera_reader/add0/c19 ),
    .o({open_n794,\u_camera_reader/n8 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_camera_reader/add0/u2  (
    .a(\u_camera_reader/pixel_counter [2]),
    .b(1'b0),
    .c(\u_camera_reader/add0/c2 ),
    .o({\u_camera_reader/add0/c3 ,\u_camera_reader/n8 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_camera_reader/add0/u3  (
    .a(\u_camera_reader/pixel_counter [3]),
    .b(1'b0),
    .c(\u_camera_reader/add0/c3 ),
    .o({\u_camera_reader/add0/c4 ,\u_camera_reader/n8 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_camera_reader/add0/u4  (
    .a(\u_camera_reader/pixel_counter [4]),
    .b(1'b0),
    .c(\u_camera_reader/add0/c4 ),
    .o({\u_camera_reader/add0/c5 ,\u_camera_reader/n8 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_camera_reader/add0/u5  (
    .a(\u_camera_reader/pixel_counter [5]),
    .b(1'b0),
    .c(\u_camera_reader/add0/c5 ),
    .o({\u_camera_reader/add0/c6 ,\u_camera_reader/n8 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_camera_reader/add0/u6  (
    .a(\u_camera_reader/pixel_counter [6]),
    .b(1'b0),
    .c(\u_camera_reader/add0/c6 ),
    .o({\u_camera_reader/add0/c7 ,\u_camera_reader/n8 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_camera_reader/add0/u7  (
    .a(\u_camera_reader/pixel_counter [7]),
    .b(1'b0),
    .c(\u_camera_reader/add0/c7 ),
    .o({\u_camera_reader/add0/c8 ,\u_camera_reader/n8 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_camera_reader/add0/u8  (
    .a(\u_camera_reader/pixel_counter [8]),
    .b(1'b0),
    .c(\u_camera_reader/add0/c8 ),
    .o({\u_camera_reader/add0/c9 ,\u_camera_reader/n8 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_camera_reader/add0/u9  (
    .a(\u_camera_reader/pixel_counter [9]),
    .b(1'b0),
    .c(\u_camera_reader/add0/c9 ),
    .o({\u_camera_reader/add0/c10 ,\u_camera_reader/n8 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u_camera_reader/add0/ucin  (
    .a(1'b0),
    .o({\u_camera_reader/add0/c0 ,open_n797}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_camera_reader/add1/u0  (
    .a(camera_addr[0]),
    .b(1'b1),
    .c(\u_camera_reader/add1/c0 ),
    .o({\u_camera_reader/add1/c1 ,\u_camera_reader/n9 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_camera_reader/add1/u1  (
    .a(camera_addr[1]),
    .b(1'b0),
    .c(\u_camera_reader/add1/c1 ),
    .o({\u_camera_reader/add1/c2 ,\u_camera_reader/n9 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_camera_reader/add1/u10  (
    .a(camera_addr[10]),
    .b(1'b0),
    .c(\u_camera_reader/add1/c10 ),
    .o({\u_camera_reader/add1/c11 ,\u_camera_reader/n9 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_camera_reader/add1/u11  (
    .a(camera_addr[11]),
    .b(1'b0),
    .c(\u_camera_reader/add1/c11 ),
    .o({\u_camera_reader/add1/c12 ,\u_camera_reader/n9 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_camera_reader/add1/u12  (
    .a(camera_addr[12]),
    .b(1'b0),
    .c(\u_camera_reader/add1/c12 ),
    .o({\u_camera_reader/add1/c13 ,\u_camera_reader/n9 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_camera_reader/add1/u13  (
    .a(camera_addr[13]),
    .b(1'b0),
    .c(\u_camera_reader/add1/c13 ),
    .o({\u_camera_reader/add1/c14 ,\u_camera_reader/n9 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_camera_reader/add1/u14  (
    .a(camera_addr[14]),
    .b(1'b0),
    .c(\u_camera_reader/add1/c14 ),
    .o({\u_camera_reader/add1/c15 ,\u_camera_reader/n9 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_camera_reader/add1/u15  (
    .a(camera_addr[15]),
    .b(1'b0),
    .c(\u_camera_reader/add1/c15 ),
    .o({open_n798,\u_camera_reader/n9 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_camera_reader/add1/u2  (
    .a(camera_addr[2]),
    .b(1'b0),
    .c(\u_camera_reader/add1/c2 ),
    .o({\u_camera_reader/add1/c3 ,\u_camera_reader/n9 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_camera_reader/add1/u3  (
    .a(camera_addr[3]),
    .b(1'b0),
    .c(\u_camera_reader/add1/c3 ),
    .o({\u_camera_reader/add1/c4 ,\u_camera_reader/n9 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_camera_reader/add1/u4  (
    .a(camera_addr[4]),
    .b(1'b0),
    .c(\u_camera_reader/add1/c4 ),
    .o({\u_camera_reader/add1/c5 ,\u_camera_reader/n9 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_camera_reader/add1/u5  (
    .a(camera_addr[5]),
    .b(1'b0),
    .c(\u_camera_reader/add1/c5 ),
    .o({\u_camera_reader/add1/c6 ,\u_camera_reader/n9 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_camera_reader/add1/u6  (
    .a(camera_addr[6]),
    .b(1'b0),
    .c(\u_camera_reader/add1/c6 ),
    .o({\u_camera_reader/add1/c7 ,\u_camera_reader/n9 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_camera_reader/add1/u7  (
    .a(camera_addr[7]),
    .b(1'b0),
    .c(\u_camera_reader/add1/c7 ),
    .o({\u_camera_reader/add1/c8 ,\u_camera_reader/n9 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_camera_reader/add1/u8  (
    .a(camera_addr[8]),
    .b(1'b0),
    .c(\u_camera_reader/add1/c8 ),
    .o({\u_camera_reader/add1/c9 ,\u_camera_reader/n9 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_camera_reader/add1/u9  (
    .a(camera_addr[9]),
    .b(1'b0),
    .c(\u_camera_reader/add1/c9 ),
    .o({\u_camera_reader/add1/c10 ,\u_camera_reader/n9 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u_camera_reader/add1/ucin  (
    .a(1'b0),
    .o({\u_camera_reader/add1/c0 ,open_n801}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_camera_reader/lt0_0  (
    .a(1'b0),
    .b(\u_camera_reader/pixel_counter [0]),
    .c(\u_camera_reader/lt0_c0 ),
    .o({\u_camera_reader/lt0_c1 ,open_n802}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_camera_reader/lt0_1  (
    .a(1'b1),
    .b(\u_camera_reader/pixel_counter [1]),
    .c(\u_camera_reader/lt0_c1 ),
    .o({\u_camera_reader/lt0_c2 ,open_n803}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_camera_reader/lt0_10  (
    .a(1'b0),
    .b(\u_camera_reader/pixel_counter [10]),
    .c(\u_camera_reader/lt0_c10 ),
    .o({\u_camera_reader/lt0_c11 ,open_n804}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_camera_reader/lt0_11  (
    .a(1'b0),
    .b(\u_camera_reader/pixel_counter [11]),
    .c(\u_camera_reader/lt0_c11 ),
    .o({\u_camera_reader/lt0_c12 ,open_n805}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_camera_reader/lt0_12  (
    .a(1'b0),
    .b(\u_camera_reader/pixel_counter [12]),
    .c(\u_camera_reader/lt0_c12 ),
    .o({\u_camera_reader/lt0_c13 ,open_n806}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_camera_reader/lt0_13  (
    .a(1'b0),
    .b(\u_camera_reader/pixel_counter [13]),
    .c(\u_camera_reader/lt0_c13 ),
    .o({\u_camera_reader/lt0_c14 ,open_n807}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_camera_reader/lt0_14  (
    .a(1'b0),
    .b(\u_camera_reader/pixel_counter [14]),
    .c(\u_camera_reader/lt0_c14 ),
    .o({\u_camera_reader/lt0_c15 ,open_n808}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_camera_reader/lt0_15  (
    .a(1'b0),
    .b(\u_camera_reader/pixel_counter [15]),
    .c(\u_camera_reader/lt0_c15 ),
    .o({\u_camera_reader/lt0_c16 ,open_n809}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_camera_reader/lt0_16  (
    .a(1'b0),
    .b(\u_camera_reader/pixel_counter [16]),
    .c(\u_camera_reader/lt0_c16 ),
    .o({\u_camera_reader/lt0_c17 ,open_n810}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_camera_reader/lt0_17  (
    .a(1'b0),
    .b(\u_camera_reader/pixel_counter [17]),
    .c(\u_camera_reader/lt0_c17 ),
    .o({\u_camera_reader/lt0_c18 ,open_n811}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_camera_reader/lt0_18  (
    .a(1'b0),
    .b(\u_camera_reader/pixel_counter [18]),
    .c(\u_camera_reader/lt0_c18 ),
    .o({\u_camera_reader/lt0_c19 ,open_n812}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_camera_reader/lt0_19  (
    .a(1'b0),
    .b(\u_camera_reader/pixel_counter [19]),
    .c(\u_camera_reader/lt0_c19 ),
    .o({\u_camera_reader/lt0_c20 ,open_n813}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_camera_reader/lt0_2  (
    .a(1'b0),
    .b(\u_camera_reader/pixel_counter [2]),
    .c(\u_camera_reader/lt0_c2 ),
    .o({\u_camera_reader/lt0_c3 ,open_n814}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_camera_reader/lt0_3  (
    .a(1'b0),
    .b(\u_camera_reader/pixel_counter [3]),
    .c(\u_camera_reader/lt0_c3 ),
    .o({\u_camera_reader/lt0_c4 ,open_n815}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_camera_reader/lt0_4  (
    .a(1'b0),
    .b(\u_camera_reader/pixel_counter [4]),
    .c(\u_camera_reader/lt0_c4 ),
    .o({\u_camera_reader/lt0_c5 ,open_n816}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_camera_reader/lt0_5  (
    .a(1'b0),
    .b(\u_camera_reader/pixel_counter [5]),
    .c(\u_camera_reader/lt0_c5 ),
    .o({\u_camera_reader/lt0_c6 ,open_n817}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_camera_reader/lt0_6  (
    .a(1'b0),
    .b(\u_camera_reader/pixel_counter [6]),
    .c(\u_camera_reader/lt0_c6 ),
    .o({\u_camera_reader/lt0_c7 ,open_n818}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_camera_reader/lt0_7  (
    .a(1'b0),
    .b(\u_camera_reader/pixel_counter [7]),
    .c(\u_camera_reader/lt0_c7 ),
    .o({\u_camera_reader/lt0_c8 ,open_n819}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_camera_reader/lt0_8  (
    .a(1'b0),
    .b(\u_camera_reader/pixel_counter [8]),
    .c(\u_camera_reader/lt0_c8 ),
    .o({\u_camera_reader/lt0_c9 ,open_n820}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_camera_reader/lt0_9  (
    .a(1'b0),
    .b(\u_camera_reader/pixel_counter [9]),
    .c(\u_camera_reader/lt0_c9 ),
    .o({\u_camera_reader/lt0_c10 ,open_n821}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u_camera_reader/lt0_cin  (
    .a(1'b0),
    .o({\u_camera_reader/lt0_c0 ,open_n824}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_camera_reader/lt0_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u_camera_reader/lt0_c20 ),
    .o({open_n825,\u_camera_reader/n27 }));
  reg_ar_as_w1 \u_camera_reader/reg0_b0  (
    .clk(camera_wrreq),
    .d(\u_camera_reader/current_pixel [0]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(camera_wrdat[0]));  // sources/rtl/camera_reader.v(56)
  reg_ar_as_w1 \u_camera_reader/reg0_b1  (
    .clk(camera_wrreq),
    .d(\u_camera_reader/current_pixel [1]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(camera_wrdat[1]));  // sources/rtl/camera_reader.v(56)
  reg_ar_as_w1 \u_camera_reader/reg0_b10  (
    .clk(camera_wrreq),
    .d(\u_camera_reader/current_pixel [10]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(camera_wrdat[10]));  // sources/rtl/camera_reader.v(56)
  reg_ar_as_w1 \u_camera_reader/reg0_b11  (
    .clk(camera_wrreq),
    .d(\u_camera_reader/current_pixel [11]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(camera_wrdat[11]));  // sources/rtl/camera_reader.v(56)
  reg_ar_as_w1 \u_camera_reader/reg0_b12  (
    .clk(camera_wrreq),
    .d(\u_camera_reader/current_pixel [12]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(camera_wrdat[12]));  // sources/rtl/camera_reader.v(56)
  reg_ar_as_w1 \u_camera_reader/reg0_b13  (
    .clk(camera_wrreq),
    .d(\u_camera_reader/current_pixel [13]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(camera_wrdat[13]));  // sources/rtl/camera_reader.v(56)
  reg_ar_as_w1 \u_camera_reader/reg0_b14  (
    .clk(camera_wrreq),
    .d(\u_camera_reader/current_pixel [14]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(camera_wrdat[14]));  // sources/rtl/camera_reader.v(56)
  reg_ar_as_w1 \u_camera_reader/reg0_b15  (
    .clk(camera_wrreq),
    .d(\u_camera_reader/current_pixel [15]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(camera_wrdat[15]));  // sources/rtl/camera_reader.v(56)
  reg_ar_as_w1 \u_camera_reader/reg0_b2  (
    .clk(camera_wrreq),
    .d(\u_camera_reader/current_pixel [2]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(camera_wrdat[2]));  // sources/rtl/camera_reader.v(56)
  reg_ar_as_w1 \u_camera_reader/reg0_b3  (
    .clk(camera_wrreq),
    .d(\u_camera_reader/current_pixel [3]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(camera_wrdat[3]));  // sources/rtl/camera_reader.v(56)
  reg_ar_as_w1 \u_camera_reader/reg0_b4  (
    .clk(camera_wrreq),
    .d(\u_camera_reader/current_pixel [4]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(camera_wrdat[4]));  // sources/rtl/camera_reader.v(56)
  reg_ar_as_w1 \u_camera_reader/reg0_b5  (
    .clk(camera_wrreq),
    .d(\u_camera_reader/current_pixel [5]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(camera_wrdat[5]));  // sources/rtl/camera_reader.v(56)
  reg_ar_as_w1 \u_camera_reader/reg0_b6  (
    .clk(camera_wrreq),
    .d(\u_camera_reader/current_pixel [6]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(camera_wrdat[6]));  // sources/rtl/camera_reader.v(56)
  reg_ar_as_w1 \u_camera_reader/reg0_b7  (
    .clk(camera_wrreq),
    .d(\u_camera_reader/current_pixel [7]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(camera_wrdat[7]));  // sources/rtl/camera_reader.v(56)
  reg_ar_as_w1 \u_camera_reader/reg0_b8  (
    .clk(camera_wrreq),
    .d(\u_camera_reader/current_pixel [8]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(camera_wrdat[8]));  // sources/rtl/camera_reader.v(56)
  reg_ar_as_w1 \u_camera_reader/reg0_b9  (
    .clk(camera_wrreq),
    .d(\u_camera_reader/current_pixel [9]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(camera_wrdat[9]));  // sources/rtl/camera_reader.v(56)
  reg_ar_as_w1 \u_camera_reader/reg1_b0  (
    .clk(cam_pclk_pad),
    .d(\u_camera_reader/n19 [0]),
    .en(1'b1),
    .reset(cam_rst_pad_neg),
    .set(1'b0),
    .q(\u_camera_reader/pixel_counter [0]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg1_b1  (
    .clk(cam_pclk_pad),
    .d(\u_camera_reader/n19 [1]),
    .en(1'b1),
    .reset(cam_rst_pad_neg),
    .set(1'b0),
    .q(\u_camera_reader/pixel_counter [1]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg1_b10  (
    .clk(cam_pclk_pad),
    .d(\u_camera_reader/n19 [10]),
    .en(1'b1),
    .reset(cam_rst_pad_neg),
    .set(1'b0),
    .q(\u_camera_reader/pixel_counter [10]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg1_b11  (
    .clk(cam_pclk_pad),
    .d(\u_camera_reader/n19 [11]),
    .en(1'b1),
    .reset(cam_rst_pad_neg),
    .set(1'b0),
    .q(\u_camera_reader/pixel_counter [11]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg1_b12  (
    .clk(cam_pclk_pad),
    .d(\u_camera_reader/n19 [12]),
    .en(1'b1),
    .reset(cam_rst_pad_neg),
    .set(1'b0),
    .q(\u_camera_reader/pixel_counter [12]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg1_b13  (
    .clk(cam_pclk_pad),
    .d(\u_camera_reader/n19 [13]),
    .en(1'b1),
    .reset(cam_rst_pad_neg),
    .set(1'b0),
    .q(\u_camera_reader/pixel_counter [13]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg1_b14  (
    .clk(cam_pclk_pad),
    .d(\u_camera_reader/n19 [14]),
    .en(1'b1),
    .reset(cam_rst_pad_neg),
    .set(1'b0),
    .q(\u_camera_reader/pixel_counter [14]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg1_b15  (
    .clk(cam_pclk_pad),
    .d(\u_camera_reader/n19 [15]),
    .en(1'b1),
    .reset(cam_rst_pad_neg),
    .set(1'b0),
    .q(\u_camera_reader/pixel_counter [15]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg1_b16  (
    .clk(cam_pclk_pad),
    .d(\u_camera_reader/n19 [16]),
    .en(1'b1),
    .reset(cam_rst_pad_neg),
    .set(1'b0),
    .q(\u_camera_reader/pixel_counter [16]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg1_b17  (
    .clk(cam_pclk_pad),
    .d(\u_camera_reader/n19 [17]),
    .en(1'b1),
    .reset(cam_rst_pad_neg),
    .set(1'b0),
    .q(\u_camera_reader/pixel_counter [17]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg1_b18  (
    .clk(cam_pclk_pad),
    .d(\u_camera_reader/n19 [18]),
    .en(1'b1),
    .reset(cam_rst_pad_neg),
    .set(1'b0),
    .q(\u_camera_reader/pixel_counter [18]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg1_b19  (
    .clk(cam_pclk_pad),
    .d(\u_camera_reader/n19 [19]),
    .en(1'b1),
    .reset(cam_rst_pad_neg),
    .set(1'b0),
    .q(\u_camera_reader/pixel_counter [19]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg1_b2  (
    .clk(cam_pclk_pad),
    .d(\u_camera_reader/n19 [2]),
    .en(1'b1),
    .reset(cam_rst_pad_neg),
    .set(1'b0),
    .q(\u_camera_reader/pixel_counter [2]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg1_b3  (
    .clk(cam_pclk_pad),
    .d(\u_camera_reader/n19 [3]),
    .en(1'b1),
    .reset(cam_rst_pad_neg),
    .set(1'b0),
    .q(\u_camera_reader/pixel_counter [3]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg1_b4  (
    .clk(cam_pclk_pad),
    .d(\u_camera_reader/n19 [4]),
    .en(1'b1),
    .reset(cam_rst_pad_neg),
    .set(1'b0),
    .q(\u_camera_reader/pixel_counter [4]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg1_b5  (
    .clk(cam_pclk_pad),
    .d(\u_camera_reader/n19 [5]),
    .en(1'b1),
    .reset(cam_rst_pad_neg),
    .set(1'b0),
    .q(\u_camera_reader/pixel_counter [5]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg1_b6  (
    .clk(cam_pclk_pad),
    .d(\u_camera_reader/n19 [6]),
    .en(1'b1),
    .reset(cam_rst_pad_neg),
    .set(1'b0),
    .q(\u_camera_reader/pixel_counter [6]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg1_b7  (
    .clk(cam_pclk_pad),
    .d(\u_camera_reader/n19 [7]),
    .en(1'b1),
    .reset(cam_rst_pad_neg),
    .set(1'b0),
    .q(\u_camera_reader/pixel_counter [7]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg1_b8  (
    .clk(cam_pclk_pad),
    .d(\u_camera_reader/n19 [8]),
    .en(1'b1),
    .reset(cam_rst_pad_neg),
    .set(1'b0),
    .q(\u_camera_reader/pixel_counter [8]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg1_b9  (
    .clk(cam_pclk_pad),
    .d(\u_camera_reader/n19 [9]),
    .en(1'b1),
    .reset(cam_rst_pad_neg),
    .set(1'b0),
    .q(\u_camera_reader/pixel_counter [9]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg2_b0  (
    .clk(cam_pclk_pad),
    .d(\u_camera_reader/n21 [0]),
    .en(~cam_rst_pad_neg),
    .reset(1'b0),
    .set(1'b0),
    .q(camera_addr[0]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg2_b1  (
    .clk(cam_pclk_pad),
    .d(\u_camera_reader/n21 [1]),
    .en(~cam_rst_pad_neg),
    .reset(1'b0),
    .set(1'b0),
    .q(camera_addr[1]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg2_b10  (
    .clk(cam_pclk_pad),
    .d(\u_camera_reader/n21 [10]),
    .en(~cam_rst_pad_neg),
    .reset(1'b0),
    .set(1'b0),
    .q(camera_addr[10]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg2_b11  (
    .clk(cam_pclk_pad),
    .d(\u_camera_reader/n21 [11]),
    .en(~cam_rst_pad_neg),
    .reset(1'b0),
    .set(1'b0),
    .q(camera_addr[11]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg2_b12  (
    .clk(cam_pclk_pad),
    .d(\u_camera_reader/n21 [12]),
    .en(~cam_rst_pad_neg),
    .reset(1'b0),
    .set(1'b0),
    .q(camera_addr[12]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg2_b13  (
    .clk(cam_pclk_pad),
    .d(\u_camera_reader/n21 [13]),
    .en(~cam_rst_pad_neg),
    .reset(1'b0),
    .set(1'b0),
    .q(camera_addr[13]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg2_b14  (
    .clk(cam_pclk_pad),
    .d(\u_camera_reader/n21 [14]),
    .en(~cam_rst_pad_neg),
    .reset(1'b0),
    .set(1'b0),
    .q(camera_addr[14]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg2_b15  (
    .clk(cam_pclk_pad),
    .d(\u_camera_reader/n21 [15]),
    .en(~cam_rst_pad_neg),
    .reset(1'b0),
    .set(1'b0),
    .q(camera_addr[15]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg2_b2  (
    .clk(cam_pclk_pad),
    .d(\u_camera_reader/n21 [2]),
    .en(~cam_rst_pad_neg),
    .reset(1'b0),
    .set(1'b0),
    .q(camera_addr[2]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg2_b3  (
    .clk(cam_pclk_pad),
    .d(\u_camera_reader/n21 [3]),
    .en(~cam_rst_pad_neg),
    .reset(1'b0),
    .set(1'b0),
    .q(camera_addr[3]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg2_b4  (
    .clk(cam_pclk_pad),
    .d(\u_camera_reader/n21 [4]),
    .en(~cam_rst_pad_neg),
    .reset(1'b0),
    .set(1'b0),
    .q(camera_addr[4]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg2_b5  (
    .clk(cam_pclk_pad),
    .d(\u_camera_reader/n21 [5]),
    .en(~cam_rst_pad_neg),
    .reset(1'b0),
    .set(1'b0),
    .q(camera_addr[5]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg2_b6  (
    .clk(cam_pclk_pad),
    .d(\u_camera_reader/n21 [6]),
    .en(~cam_rst_pad_neg),
    .reset(1'b0),
    .set(1'b0),
    .q(camera_addr[6]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg2_b7  (
    .clk(cam_pclk_pad),
    .d(\u_camera_reader/n21 [7]),
    .en(~cam_rst_pad_neg),
    .reset(1'b0),
    .set(1'b0),
    .q(camera_addr[7]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg2_b8  (
    .clk(cam_pclk_pad),
    .d(\u_camera_reader/n21 [8]),
    .en(~cam_rst_pad_neg),
    .reset(1'b0),
    .set(1'b0),
    .q(camera_addr[8]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg2_b9  (
    .clk(cam_pclk_pad),
    .d(\u_camera_reader/n21 [9]),
    .en(~cam_rst_pad_neg),
    .reset(1'b0),
    .set(1'b0),
    .q(camera_addr[9]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg3_b0  (
    .clk(cam_pclk_pad),
    .d(cam_data_pad[0]),
    .en(\u_camera_reader/mux13_b0_sel_is_2_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_camera_reader/subpixel [0]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg3_b1  (
    .clk(cam_pclk_pad),
    .d(cam_data_pad[1]),
    .en(\u_camera_reader/mux13_b0_sel_is_2_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_camera_reader/subpixel [1]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg3_b2  (
    .clk(cam_pclk_pad),
    .d(cam_data_pad[2]),
    .en(\u_camera_reader/mux13_b0_sel_is_2_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_camera_reader/subpixel [2]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg3_b3  (
    .clk(cam_pclk_pad),
    .d(cam_data_pad[3]),
    .en(\u_camera_reader/mux13_b0_sel_is_2_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_camera_reader/subpixel [3]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg3_b4  (
    .clk(cam_pclk_pad),
    .d(cam_data_pad[4]),
    .en(\u_camera_reader/mux13_b0_sel_is_2_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_camera_reader/subpixel [4]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg3_b5  (
    .clk(cam_pclk_pad),
    .d(cam_data_pad[5]),
    .en(\u_camera_reader/mux13_b0_sel_is_2_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_camera_reader/subpixel [5]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg3_b6  (
    .clk(cam_pclk_pad),
    .d(cam_data_pad[6]),
    .en(\u_camera_reader/mux13_b0_sel_is_2_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_camera_reader/subpixel [6]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg3_b7  (
    .clk(cam_pclk_pad),
    .d(cam_data_pad[7]),
    .en(\u_camera_reader/mux13_b0_sel_is_2_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_camera_reader/subpixel [7]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg4_b0  (
    .clk(cam_pclk_pad),
    .d(cam_data_pad[0]),
    .en(\u_camera_reader/mux14_b0_sel_is_2_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_camera_reader/current_pixel [0]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg4_b1  (
    .clk(cam_pclk_pad),
    .d(cam_data_pad[1]),
    .en(\u_camera_reader/mux14_b0_sel_is_2_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_camera_reader/current_pixel [1]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg4_b10  (
    .clk(cam_pclk_pad),
    .d(\u_camera_reader/subpixel [2]),
    .en(\u_camera_reader/mux14_b0_sel_is_2_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_camera_reader/current_pixel [10]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg4_b11  (
    .clk(cam_pclk_pad),
    .d(\u_camera_reader/subpixel [3]),
    .en(\u_camera_reader/mux14_b0_sel_is_2_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_camera_reader/current_pixel [11]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg4_b12  (
    .clk(cam_pclk_pad),
    .d(\u_camera_reader/subpixel [4]),
    .en(\u_camera_reader/mux14_b0_sel_is_2_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_camera_reader/current_pixel [12]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg4_b13  (
    .clk(cam_pclk_pad),
    .d(\u_camera_reader/subpixel [5]),
    .en(\u_camera_reader/mux14_b0_sel_is_2_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_camera_reader/current_pixel [13]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg4_b14  (
    .clk(cam_pclk_pad),
    .d(\u_camera_reader/subpixel [6]),
    .en(\u_camera_reader/mux14_b0_sel_is_2_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_camera_reader/current_pixel [14]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg4_b15  (
    .clk(cam_pclk_pad),
    .d(\u_camera_reader/subpixel [7]),
    .en(\u_camera_reader/mux14_b0_sel_is_2_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_camera_reader/current_pixel [15]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg4_b2  (
    .clk(cam_pclk_pad),
    .d(cam_data_pad[2]),
    .en(\u_camera_reader/mux14_b0_sel_is_2_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_camera_reader/current_pixel [2]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg4_b3  (
    .clk(cam_pclk_pad),
    .d(cam_data_pad[3]),
    .en(\u_camera_reader/mux14_b0_sel_is_2_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_camera_reader/current_pixel [3]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg4_b4  (
    .clk(cam_pclk_pad),
    .d(cam_data_pad[4]),
    .en(\u_camera_reader/mux14_b0_sel_is_2_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_camera_reader/current_pixel [4]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg4_b5  (
    .clk(cam_pclk_pad),
    .d(cam_data_pad[5]),
    .en(\u_camera_reader/mux14_b0_sel_is_2_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_camera_reader/current_pixel [5]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg4_b6  (
    .clk(cam_pclk_pad),
    .d(cam_data_pad[6]),
    .en(\u_camera_reader/mux14_b0_sel_is_2_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_camera_reader/current_pixel [6]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg4_b7  (
    .clk(cam_pclk_pad),
    .d(cam_data_pad[7]),
    .en(\u_camera_reader/mux14_b0_sel_is_2_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_camera_reader/current_pixel [7]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg4_b8  (
    .clk(cam_pclk_pad),
    .d(\u_camera_reader/subpixel [0]),
    .en(\u_camera_reader/mux14_b0_sel_is_2_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_camera_reader/current_pixel [8]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg4_b9  (
    .clk(cam_pclk_pad),
    .d(\u_camera_reader/subpixel [1]),
    .en(\u_camera_reader/mux14_b0_sel_is_2_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_camera_reader/current_pixel [9]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/vsync_passed_reg  (
    .clk(cam_pclk_pad),
    .d(\u_camera_reader/vsync_passed_d ),
    .en(1'b1),
    .reset(cam_rst_pad_neg),
    .set(1'b0),
    .q(\u_camera_reader/vsync_passed ));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/wrclk1_reg  (
    .clk(cam_pclk_pad),
    .d(\u_camera_reader/n1 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_camera_reader/wrclk1 ));  // sources/rtl/camera_reader.v(43)
  reg_ar_as_w1 \u_camera_reader/write_pixel_reg  (
    .clk(~\u_camera_reader/wrclk1 ),
    .d(\u_camera_reader/n2 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_camera_reader/write_pixel ));  // sources/rtl/camera_reader.v(51)
  // address_offset=0;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("INV"),
    .CSB1("INV"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_img/inst_32800x16_sub_000000_000  (
    .addra({camera_addr[9:0],3'b111}),
    .addrb({vga_rdaddr[9:0],3'b111}),
    .cea(camera_wrreq),
    .ceb(vga_rden),
    .clka(cam_pclk_pad),
    .clkb(clk_lcd),
    .csa({\and_Ncamera_addr[12]_o ,camera_addr[11:10]}),
    .csb({\and_Nvga_rdaddr[12]__o ,vga_rdaddr[11:10]}),
    .dia(camera_wrdat[8:0]),
    .rsta(cam_rst_pad),
    .rstb(cam_rst_pad),
    .dob({\u_img/inst_dob_i0_008 ,\u_img/inst_dob_i0_007 ,\u_img/inst_dob_i0_006 ,\u_img/inst_dob_i0_005 ,\u_img/inst_dob_i0_004 ,\u_img/inst_dob_i0_003 ,\u_img/inst_dob_i0_002 ,\u_img/inst_dob_i0_001 ,\u_img/inst_dob_i0_000 }));
  // address_offset=0;data_offset=9;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("INV"),
    .CSB1("INV"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_img/inst_32800x16_sub_000000_009  (
    .addra(camera_addr[12:0]),
    .addrb(vga_rdaddr[12:0]),
    .cea(camera_wrreq),
    .ceb(vga_rden),
    .clka(cam_pclk_pad),
    .clkb(clk_lcd),
    .csa(camera_addr[15:13]),
    .csb(vga_rdaddr[15:13]),
    .dia({open_n848,open_n849,open_n850,open_n851,open_n852,open_n853,open_n854,camera_wrdat[9],open_n855}),
    .rsta(cam_rst_pad),
    .rstb(cam_rst_pad),
    .dob({open_n878,open_n879,open_n880,open_n881,open_n882,open_n883,open_n884,open_n885,\u_img/inst_dob_i0_009 }));
  // address_offset=0;data_offset=10;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("INV"),
    .CSB1("INV"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_img/inst_32800x16_sub_000000_010  (
    .addra(camera_addr[12:0]),
    .addrb(vga_rdaddr[12:0]),
    .cea(camera_wrreq),
    .ceb(vga_rden),
    .clka(cam_pclk_pad),
    .clkb(clk_lcd),
    .csa(camera_addr[15:13]),
    .csb(vga_rdaddr[15:13]),
    .dia({open_n886,open_n887,open_n888,open_n889,open_n890,open_n891,open_n892,camera_wrdat[10],open_n893}),
    .rsta(cam_rst_pad),
    .rstb(cam_rst_pad),
    .dob({open_n916,open_n917,open_n918,open_n919,open_n920,open_n921,open_n922,open_n923,\u_img/inst_dob_i0_010 }));
  // address_offset=0;data_offset=11;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("INV"),
    .CSB1("INV"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_img/inst_32800x16_sub_000000_011  (
    .addra(camera_addr[12:0]),
    .addrb(vga_rdaddr[12:0]),
    .cea(camera_wrreq),
    .ceb(vga_rden),
    .clka(cam_pclk_pad),
    .clkb(clk_lcd),
    .csa(camera_addr[15:13]),
    .csb(vga_rdaddr[15:13]),
    .dia({open_n924,open_n925,open_n926,open_n927,open_n928,open_n929,open_n930,camera_wrdat[11],open_n931}),
    .rsta(cam_rst_pad),
    .rstb(cam_rst_pad),
    .dob({open_n954,open_n955,open_n956,open_n957,open_n958,open_n959,open_n960,open_n961,\u_img/inst_dob_i0_011 }));
  // address_offset=0;data_offset=12;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("INV"),
    .CSB1("INV"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_img/inst_32800x16_sub_000000_012  (
    .addra(camera_addr[12:0]),
    .addrb(vga_rdaddr[12:0]),
    .cea(camera_wrreq),
    .ceb(vga_rden),
    .clka(cam_pclk_pad),
    .clkb(clk_lcd),
    .csa(camera_addr[15:13]),
    .csb(vga_rdaddr[15:13]),
    .dia({open_n962,open_n963,open_n964,open_n965,open_n966,open_n967,open_n968,camera_wrdat[12],open_n969}),
    .rsta(cam_rst_pad),
    .rstb(cam_rst_pad),
    .dob({open_n992,open_n993,open_n994,open_n995,open_n996,open_n997,open_n998,open_n999,\u_img/inst_dob_i0_012 }));
  // address_offset=0;data_offset=13;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("INV"),
    .CSB1("INV"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_img/inst_32800x16_sub_000000_013  (
    .addra(camera_addr[12:0]),
    .addrb(vga_rdaddr[12:0]),
    .cea(camera_wrreq),
    .ceb(vga_rden),
    .clka(cam_pclk_pad),
    .clkb(clk_lcd),
    .csa(camera_addr[15:13]),
    .csb(vga_rdaddr[15:13]),
    .dia({open_n1000,open_n1001,open_n1002,open_n1003,open_n1004,open_n1005,open_n1006,camera_wrdat[13],open_n1007}),
    .rsta(cam_rst_pad),
    .rstb(cam_rst_pad),
    .dob({open_n1030,open_n1031,open_n1032,open_n1033,open_n1034,open_n1035,open_n1036,open_n1037,\u_img/inst_dob_i0_013 }));
  // address_offset=0;data_offset=14;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("INV"),
    .CSB1("INV"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_img/inst_32800x16_sub_000000_014  (
    .addra(camera_addr[12:0]),
    .addrb(vga_rdaddr[12:0]),
    .cea(camera_wrreq),
    .ceb(vga_rden),
    .clka(cam_pclk_pad),
    .clkb(clk_lcd),
    .csa(camera_addr[15:13]),
    .csb(vga_rdaddr[15:13]),
    .dia({open_n1038,open_n1039,open_n1040,open_n1041,open_n1042,open_n1043,open_n1044,camera_wrdat[14],open_n1045}),
    .rsta(cam_rst_pad),
    .rstb(cam_rst_pad),
    .dob({open_n1068,open_n1069,open_n1070,open_n1071,open_n1072,open_n1073,open_n1074,open_n1075,\u_img/inst_dob_i0_014 }));
  // address_offset=0;data_offset=15;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("INV"),
    .CSB1("INV"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_img/inst_32800x16_sub_000000_015  (
    .addra(camera_addr[12:0]),
    .addrb(vga_rdaddr[12:0]),
    .cea(camera_wrreq),
    .ceb(vga_rden),
    .clka(cam_pclk_pad),
    .clkb(clk_lcd),
    .csa(camera_addr[15:13]),
    .csb(vga_rdaddr[15:13]),
    .dia({open_n1076,open_n1077,open_n1078,open_n1079,open_n1080,open_n1081,open_n1082,camera_wrdat[15],open_n1083}),
    .rsta(cam_rst_pad),
    .rstb(cam_rst_pad),
    .dob({open_n1106,open_n1107,open_n1108,open_n1109,open_n1110,open_n1111,open_n1112,open_n1113,\u_img/inst_dob_i0_015 }));
  // address_offset=1024;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("SIG"),
    .CSB1("INV"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_img/inst_32800x16_sub_001024_000  (
    .addra({camera_addr[9:0],3'b111}),
    .addrb({vga_rdaddr[9:0],3'b111}),
    .cea(camera_wrreq),
    .ceb(vga_rden),
    .clka(cam_pclk_pad),
    .clkb(clk_lcd),
    .csa({\and_Ncamera_addr[12]_o ,camera_addr[11:10]}),
    .csb({\and_Nvga_rdaddr[12]__o ,vga_rdaddr[11:10]}),
    .dia(camera_wrdat[8:0]),
    .rsta(cam_rst_pad),
    .rstb(cam_rst_pad),
    .dob({\u_img/inst_dob_i2_008 ,\u_img/inst_dob_i2_007 ,\u_img/inst_dob_i2_006 ,\u_img/inst_dob_i2_005 ,\u_img/inst_dob_i2_004 ,\u_img/inst_dob_i2_003 ,\u_img/inst_dob_i2_002 ,\u_img/inst_dob_i2_001 ,\u_img/inst_dob_i2_000 }));
  // address_offset=2048;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("INV"),
    .CSB1("SIG"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_img/inst_32800x16_sub_002048_000  (
    .addra({camera_addr[9:0],3'b111}),
    .addrb({vga_rdaddr[9:0],3'b111}),
    .cea(camera_wrreq),
    .ceb(vga_rden),
    .clka(cam_pclk_pad),
    .clkb(clk_lcd),
    .csa({\and_Ncamera_addr[12]_o ,camera_addr[11:10]}),
    .csb({\and_Nvga_rdaddr[12]__o ,vga_rdaddr[11:10]}),
    .dia(camera_wrdat[8:0]),
    .rsta(cam_rst_pad),
    .rstb(cam_rst_pad),
    .dob({\u_img/inst_dob_i4_008 ,\u_img/inst_dob_i4_007 ,\u_img/inst_dob_i4_006 ,\u_img/inst_dob_i4_005 ,\u_img/inst_dob_i4_004 ,\u_img/inst_dob_i4_003 ,\u_img/inst_dob_i4_002 ,\u_img/inst_dob_i4_001 ,\u_img/inst_dob_i4_000 }));
  // address_offset=3072;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("SIG"),
    .CSB1("SIG"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_img/inst_32800x16_sub_003072_000  (
    .addra({camera_addr[9:0],3'b111}),
    .addrb({vga_rdaddr[9:0],3'b111}),
    .cea(camera_wrreq),
    .ceb(vga_rden),
    .clka(cam_pclk_pad),
    .clkb(clk_lcd),
    .csa({\and_Ncamera_addr[12]_o ,camera_addr[11:10]}),
    .csb({\and_Nvga_rdaddr[12]__o ,vga_rdaddr[11:10]}),
    .dia(camera_wrdat[8:0]),
    .rsta(cam_rst_pad),
    .rstb(cam_rst_pad),
    .dob({\u_img/inst_dob_i6_008 ,\u_img/inst_dob_i6_007 ,\u_img/inst_dob_i6_006 ,\u_img/inst_dob_i6_005 ,\u_img/inst_dob_i6_004 ,\u_img/inst_dob_i6_003 ,\u_img/inst_dob_i6_002 ,\u_img/inst_dob_i6_001 ,\u_img/inst_dob_i6_000 }));
  // address_offset=4096;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("INV"),
    .CSB1("INV"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_img/inst_32800x16_sub_004096_000  (
    .addra({camera_addr[9:0],3'b111}),
    .addrb({vga_rdaddr[9:0],3'b111}),
    .cea(camera_wrreq),
    .ceb(vga_rden),
    .clka(cam_pclk_pad),
    .clkb(clk_lcd),
    .csa({\and_camera_addr[12]__o ,camera_addr[11:10]}),
    .csb({\and_vga_rdaddr[12]_N_o ,vga_rdaddr[11:10]}),
    .dia(camera_wrdat[8:0]),
    .rsta(cam_rst_pad),
    .rstb(cam_rst_pad),
    .dob({\u_img/inst_dob_i8_008 ,\u_img/inst_dob_i8_007 ,\u_img/inst_dob_i8_006 ,\u_img/inst_dob_i8_005 ,\u_img/inst_dob_i8_004 ,\u_img/inst_dob_i8_003 ,\u_img/inst_dob_i8_002 ,\u_img/inst_dob_i8_001 ,\u_img/inst_dob_i8_000 }));
  // address_offset=5120;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("SIG"),
    .CSB1("INV"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_img/inst_32800x16_sub_005120_000  (
    .addra({camera_addr[9:0],3'b111}),
    .addrb({vga_rdaddr[9:0],3'b111}),
    .cea(camera_wrreq),
    .ceb(vga_rden),
    .clka(cam_pclk_pad),
    .clkb(clk_lcd),
    .csa({\and_camera_addr[12]__o ,camera_addr[11:10]}),
    .csb({\and_vga_rdaddr[12]_N_o ,vga_rdaddr[11:10]}),
    .dia(camera_wrdat[8:0]),
    .rsta(cam_rst_pad),
    .rstb(cam_rst_pad),
    .dob({\u_img/inst_dob_i10_008 ,\u_img/inst_dob_i10_007 ,\u_img/inst_dob_i10_006 ,\u_img/inst_dob_i10_005 ,\u_img/inst_dob_i10_004 ,\u_img/inst_dob_i10_003 ,\u_img/inst_dob_i10_002 ,\u_img/inst_dob_i10_001 ,\u_img/inst_dob_i10_000 }));
  // address_offset=6144;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("INV"),
    .CSB1("SIG"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_img/inst_32800x16_sub_006144_000  (
    .addra({camera_addr[9:0],3'b111}),
    .addrb({vga_rdaddr[9:0],3'b111}),
    .cea(camera_wrreq),
    .ceb(vga_rden),
    .clka(cam_pclk_pad),
    .clkb(clk_lcd),
    .csa({\and_camera_addr[12]__o ,camera_addr[11:10]}),
    .csb({\and_vga_rdaddr[12]_N_o ,vga_rdaddr[11:10]}),
    .dia(camera_wrdat[8:0]),
    .rsta(cam_rst_pad),
    .rstb(cam_rst_pad),
    .dob({\u_img/inst_dob_i12_008 ,\u_img/inst_dob_i12_007 ,\u_img/inst_dob_i12_006 ,\u_img/inst_dob_i12_005 ,\u_img/inst_dob_i12_004 ,\u_img/inst_dob_i12_003 ,\u_img/inst_dob_i12_002 ,\u_img/inst_dob_i12_001 ,\u_img/inst_dob_i12_000 }));
  // address_offset=7168;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("SIG"),
    .CSB1("SIG"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_img/inst_32800x16_sub_007168_000  (
    .addra({camera_addr[9:0],3'b111}),
    .addrb({vga_rdaddr[9:0],3'b111}),
    .cea(camera_wrreq),
    .ceb(vga_rden),
    .clka(cam_pclk_pad),
    .clkb(clk_lcd),
    .csa({\and_camera_addr[12]__o ,camera_addr[11:10]}),
    .csb({\and_vga_rdaddr[12]_N_o ,vga_rdaddr[11:10]}),
    .dia(camera_wrdat[8:0]),
    .rsta(cam_rst_pad),
    .rstb(cam_rst_pad),
    .dob({\u_img/inst_dob_i14_008 ,\u_img/inst_dob_i14_007 ,\u_img/inst_dob_i14_006 ,\u_img/inst_dob_i14_005 ,\u_img/inst_dob_i14_004 ,\u_img/inst_dob_i14_003 ,\u_img/inst_dob_i14_002 ,\u_img/inst_dob_i14_001 ,\u_img/inst_dob_i14_000 }));
  // address_offset=8192;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("INV"),
    .CSB1("INV"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_img/inst_32800x16_sub_008192_000  (
    .addra({camera_addr[9:0],3'b111}),
    .addrb({vga_rdaddr[9:0],3'b111}),
    .cea(camera_wrreq),
    .ceb(vga_rden),
    .clka(cam_pclk_pad),
    .clkb(clk_lcd),
    .csa({\and_Ncamera_addr[12]_o_al_n177 ,camera_addr[11:10]}),
    .csb({\and_Nvga_rdaddr[12]__o_al_n180 ,vga_rdaddr[11:10]}),
    .dia(camera_wrdat[8:0]),
    .rsta(cam_rst_pad),
    .rstb(cam_rst_pad),
    .dob({\u_img/inst_dob_i16_008 ,\u_img/inst_dob_i16_007 ,\u_img/inst_dob_i16_006 ,\u_img/inst_dob_i16_005 ,\u_img/inst_dob_i16_004 ,\u_img/inst_dob_i16_003 ,\u_img/inst_dob_i16_002 ,\u_img/inst_dob_i16_001 ,\u_img/inst_dob_i16_000 }));
  // address_offset=8192;data_offset=9;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("SIG"),
    .CSB1("INV"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_img/inst_32800x16_sub_008192_009  (
    .addra(camera_addr[12:0]),
    .addrb(vga_rdaddr[12:0]),
    .cea(camera_wrreq),
    .ceb(vga_rden),
    .clka(cam_pclk_pad),
    .clkb(clk_lcd),
    .csa(camera_addr[15:13]),
    .csb(vga_rdaddr[15:13]),
    .dia({open_n1290,open_n1291,open_n1292,open_n1293,open_n1294,open_n1295,open_n1296,camera_wrdat[9],open_n1297}),
    .rsta(cam_rst_pad),
    .rstb(cam_rst_pad),
    .dob({open_n1320,open_n1321,open_n1322,open_n1323,open_n1324,open_n1325,open_n1326,open_n1327,\u_img/inst_dob_i16_009 }));
  // address_offset=8192;data_offset=10;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("SIG"),
    .CSB1("INV"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_img/inst_32800x16_sub_008192_010  (
    .addra(camera_addr[12:0]),
    .addrb(vga_rdaddr[12:0]),
    .cea(camera_wrreq),
    .ceb(vga_rden),
    .clka(cam_pclk_pad),
    .clkb(clk_lcd),
    .csa(camera_addr[15:13]),
    .csb(vga_rdaddr[15:13]),
    .dia({open_n1328,open_n1329,open_n1330,open_n1331,open_n1332,open_n1333,open_n1334,camera_wrdat[10],open_n1335}),
    .rsta(cam_rst_pad),
    .rstb(cam_rst_pad),
    .dob({open_n1358,open_n1359,open_n1360,open_n1361,open_n1362,open_n1363,open_n1364,open_n1365,\u_img/inst_dob_i16_010 }));
  // address_offset=8192;data_offset=11;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("SIG"),
    .CSB1("INV"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_img/inst_32800x16_sub_008192_011  (
    .addra(camera_addr[12:0]),
    .addrb(vga_rdaddr[12:0]),
    .cea(camera_wrreq),
    .ceb(vga_rden),
    .clka(cam_pclk_pad),
    .clkb(clk_lcd),
    .csa(camera_addr[15:13]),
    .csb(vga_rdaddr[15:13]),
    .dia({open_n1366,open_n1367,open_n1368,open_n1369,open_n1370,open_n1371,open_n1372,camera_wrdat[11],open_n1373}),
    .rsta(cam_rst_pad),
    .rstb(cam_rst_pad),
    .dob({open_n1396,open_n1397,open_n1398,open_n1399,open_n1400,open_n1401,open_n1402,open_n1403,\u_img/inst_dob_i16_011 }));
  // address_offset=8192;data_offset=12;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("SIG"),
    .CSB1("INV"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_img/inst_32800x16_sub_008192_012  (
    .addra(camera_addr[12:0]),
    .addrb(vga_rdaddr[12:0]),
    .cea(camera_wrreq),
    .ceb(vga_rden),
    .clka(cam_pclk_pad),
    .clkb(clk_lcd),
    .csa(camera_addr[15:13]),
    .csb(vga_rdaddr[15:13]),
    .dia({open_n1404,open_n1405,open_n1406,open_n1407,open_n1408,open_n1409,open_n1410,camera_wrdat[12],open_n1411}),
    .rsta(cam_rst_pad),
    .rstb(cam_rst_pad),
    .dob({open_n1434,open_n1435,open_n1436,open_n1437,open_n1438,open_n1439,open_n1440,open_n1441,\u_img/inst_dob_i16_012 }));
  // address_offset=8192;data_offset=13;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("SIG"),
    .CSB1("INV"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_img/inst_32800x16_sub_008192_013  (
    .addra(camera_addr[12:0]),
    .addrb(vga_rdaddr[12:0]),
    .cea(camera_wrreq),
    .ceb(vga_rden),
    .clka(cam_pclk_pad),
    .clkb(clk_lcd),
    .csa(camera_addr[15:13]),
    .csb(vga_rdaddr[15:13]),
    .dia({open_n1442,open_n1443,open_n1444,open_n1445,open_n1446,open_n1447,open_n1448,camera_wrdat[13],open_n1449}),
    .rsta(cam_rst_pad),
    .rstb(cam_rst_pad),
    .dob({open_n1472,open_n1473,open_n1474,open_n1475,open_n1476,open_n1477,open_n1478,open_n1479,\u_img/inst_dob_i16_013 }));
  // address_offset=8192;data_offset=14;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("SIG"),
    .CSB1("INV"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_img/inst_32800x16_sub_008192_014  (
    .addra(camera_addr[12:0]),
    .addrb(vga_rdaddr[12:0]),
    .cea(camera_wrreq),
    .ceb(vga_rden),
    .clka(cam_pclk_pad),
    .clkb(clk_lcd),
    .csa(camera_addr[15:13]),
    .csb(vga_rdaddr[15:13]),
    .dia({open_n1480,open_n1481,open_n1482,open_n1483,open_n1484,open_n1485,open_n1486,camera_wrdat[14],open_n1487}),
    .rsta(cam_rst_pad),
    .rstb(cam_rst_pad),
    .dob({open_n1510,open_n1511,open_n1512,open_n1513,open_n1514,open_n1515,open_n1516,open_n1517,\u_img/inst_dob_i16_014 }));
  // address_offset=8192;data_offset=15;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("SIG"),
    .CSB1("INV"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_img/inst_32800x16_sub_008192_015  (
    .addra(camera_addr[12:0]),
    .addrb(vga_rdaddr[12:0]),
    .cea(camera_wrreq),
    .ceb(vga_rden),
    .clka(cam_pclk_pad),
    .clkb(clk_lcd),
    .csa(camera_addr[15:13]),
    .csb(vga_rdaddr[15:13]),
    .dia({open_n1518,open_n1519,open_n1520,open_n1521,open_n1522,open_n1523,open_n1524,camera_wrdat[15],open_n1525}),
    .rsta(cam_rst_pad),
    .rstb(cam_rst_pad),
    .dob({open_n1548,open_n1549,open_n1550,open_n1551,open_n1552,open_n1553,open_n1554,open_n1555,\u_img/inst_dob_i16_015 }));
  // address_offset=9216;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("SIG"),
    .CSB1("INV"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_img/inst_32800x16_sub_009216_000  (
    .addra({camera_addr[9:0],3'b111}),
    .addrb({vga_rdaddr[9:0],3'b111}),
    .cea(camera_wrreq),
    .ceb(vga_rden),
    .clka(cam_pclk_pad),
    .clkb(clk_lcd),
    .csa({\and_Ncamera_addr[12]_o_al_n177 ,camera_addr[11:10]}),
    .csb({\and_Nvga_rdaddr[12]__o_al_n180 ,vga_rdaddr[11:10]}),
    .dia(camera_wrdat[8:0]),
    .rsta(cam_rst_pad),
    .rstb(cam_rst_pad),
    .dob({\u_img/inst_dob_i18_008 ,\u_img/inst_dob_i18_007 ,\u_img/inst_dob_i18_006 ,\u_img/inst_dob_i18_005 ,\u_img/inst_dob_i18_004 ,\u_img/inst_dob_i18_003 ,\u_img/inst_dob_i18_002 ,\u_img/inst_dob_i18_001 ,\u_img/inst_dob_i18_000 }));
  // address_offset=10240;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("INV"),
    .CSB1("SIG"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_img/inst_32800x16_sub_010240_000  (
    .addra({camera_addr[9:0],3'b111}),
    .addrb({vga_rdaddr[9:0],3'b111}),
    .cea(camera_wrreq),
    .ceb(vga_rden),
    .clka(cam_pclk_pad),
    .clkb(clk_lcd),
    .csa({\and_Ncamera_addr[12]_o_al_n177 ,camera_addr[11:10]}),
    .csb({\and_Nvga_rdaddr[12]__o_al_n180 ,vga_rdaddr[11:10]}),
    .dia(camera_wrdat[8:0]),
    .rsta(cam_rst_pad),
    .rstb(cam_rst_pad),
    .dob({\u_img/inst_dob_i20_008 ,\u_img/inst_dob_i20_007 ,\u_img/inst_dob_i20_006 ,\u_img/inst_dob_i20_005 ,\u_img/inst_dob_i20_004 ,\u_img/inst_dob_i20_003 ,\u_img/inst_dob_i20_002 ,\u_img/inst_dob_i20_001 ,\u_img/inst_dob_i20_000 }));
  // address_offset=11264;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("SIG"),
    .CSB1("SIG"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_img/inst_32800x16_sub_011264_000  (
    .addra({camera_addr[9:0],3'b111}),
    .addrb({vga_rdaddr[9:0],3'b111}),
    .cea(camera_wrreq),
    .ceb(vga_rden),
    .clka(cam_pclk_pad),
    .clkb(clk_lcd),
    .csa({\and_Ncamera_addr[12]_o_al_n177 ,camera_addr[11:10]}),
    .csb({\and_Nvga_rdaddr[12]__o_al_n180 ,vga_rdaddr[11:10]}),
    .dia(camera_wrdat[8:0]),
    .rsta(cam_rst_pad),
    .rstb(cam_rst_pad),
    .dob({\u_img/inst_dob_i22_008 ,\u_img/inst_dob_i22_007 ,\u_img/inst_dob_i22_006 ,\u_img/inst_dob_i22_005 ,\u_img/inst_dob_i22_004 ,\u_img/inst_dob_i22_003 ,\u_img/inst_dob_i22_002 ,\u_img/inst_dob_i22_001 ,\u_img/inst_dob_i22_000 }));
  // address_offset=12288;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("INV"),
    .CSB1("INV"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_img/inst_32800x16_sub_012288_000  (
    .addra({camera_addr[9:0],3'b111}),
    .addrb({vga_rdaddr[9:0],3'b111}),
    .cea(camera_wrreq),
    .ceb(vga_rden),
    .clka(cam_pclk_pad),
    .clkb(clk_lcd),
    .csa({\and_camera_addr[12]__o_al_n193 ,camera_addr[11:10]}),
    .csb({\and_vga_rdaddr[12]_v_o ,vga_rdaddr[11:10]}),
    .dia(camera_wrdat[8:0]),
    .rsta(cam_rst_pad),
    .rstb(cam_rst_pad),
    .dob({\u_img/inst_dob_i24_008 ,\u_img/inst_dob_i24_007 ,\u_img/inst_dob_i24_006 ,\u_img/inst_dob_i24_005 ,\u_img/inst_dob_i24_004 ,\u_img/inst_dob_i24_003 ,\u_img/inst_dob_i24_002 ,\u_img/inst_dob_i24_001 ,\u_img/inst_dob_i24_000 }));
  // address_offset=13312;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("SIG"),
    .CSB1("INV"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_img/inst_32800x16_sub_013312_000  (
    .addra({camera_addr[9:0],3'b111}),
    .addrb({vga_rdaddr[9:0],3'b111}),
    .cea(camera_wrreq),
    .ceb(vga_rden),
    .clka(cam_pclk_pad),
    .clkb(clk_lcd),
    .csa({\and_camera_addr[12]__o_al_n193 ,camera_addr[11:10]}),
    .csb({\and_vga_rdaddr[12]_v_o ,vga_rdaddr[11:10]}),
    .dia(camera_wrdat[8:0]),
    .rsta(cam_rst_pad),
    .rstb(cam_rst_pad),
    .dob({\u_img/inst_dob_i26_008 ,\u_img/inst_dob_i26_007 ,\u_img/inst_dob_i26_006 ,\u_img/inst_dob_i26_005 ,\u_img/inst_dob_i26_004 ,\u_img/inst_dob_i26_003 ,\u_img/inst_dob_i26_002 ,\u_img/inst_dob_i26_001 ,\u_img/inst_dob_i26_000 }));
  // address_offset=14336;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("INV"),
    .CSB1("SIG"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_img/inst_32800x16_sub_014336_000  (
    .addra({camera_addr[9:0],3'b111}),
    .addrb({vga_rdaddr[9:0],3'b111}),
    .cea(camera_wrreq),
    .ceb(vga_rden),
    .clka(cam_pclk_pad),
    .clkb(clk_lcd),
    .csa({\and_camera_addr[12]__o_al_n193 ,camera_addr[11:10]}),
    .csb({\and_vga_rdaddr[12]_v_o ,vga_rdaddr[11:10]}),
    .dia(camera_wrdat[8:0]),
    .rsta(cam_rst_pad),
    .rstb(cam_rst_pad),
    .dob({\u_img/inst_dob_i28_008 ,\u_img/inst_dob_i28_007 ,\u_img/inst_dob_i28_006 ,\u_img/inst_dob_i28_005 ,\u_img/inst_dob_i28_004 ,\u_img/inst_dob_i28_003 ,\u_img/inst_dob_i28_002 ,\u_img/inst_dob_i28_001 ,\u_img/inst_dob_i28_000 }));
  // address_offset=15360;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("SIG"),
    .CSB1("SIG"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_img/inst_32800x16_sub_015360_000  (
    .addra({camera_addr[9:0],3'b111}),
    .addrb({vga_rdaddr[9:0],3'b111}),
    .cea(camera_wrreq),
    .ceb(vga_rden),
    .clka(cam_pclk_pad),
    .clkb(clk_lcd),
    .csa({\and_camera_addr[12]__o_al_n193 ,camera_addr[11:10]}),
    .csb({\and_vga_rdaddr[12]_v_o ,vga_rdaddr[11:10]}),
    .dia(camera_wrdat[8:0]),
    .rsta(cam_rst_pad),
    .rstb(cam_rst_pad),
    .dob({\u_img/inst_dob_i30_008 ,\u_img/inst_dob_i30_007 ,\u_img/inst_dob_i30_006 ,\u_img/inst_dob_i30_005 ,\u_img/inst_dob_i30_004 ,\u_img/inst_dob_i30_003 ,\u_img/inst_dob_i30_002 ,\u_img/inst_dob_i30_001 ,\u_img/inst_dob_i30_000 }));
  // address_offset=16384;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("INV"),
    .CSB1("INV"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_img/inst_32800x16_sub_016384_000  (
    .addra({camera_addr[9:0],3'b111}),
    .addrb({vga_rdaddr[9:0],3'b111}),
    .cea(camera_wrreq),
    .ceb(vga_rden),
    .clka(cam_pclk_pad),
    .clkb(clk_lcd),
    .csa({\and_Ncamera_addr[12]_o_al_n208 ,camera_addr[11:10]}),
    .csb({\and_Nvga_rdaddr[12]__o_al_n211 ,vga_rdaddr[11:10]}),
    .dia(camera_wrdat[8:0]),
    .rsta(cam_rst_pad),
    .rstb(cam_rst_pad),
    .dob({\u_img/inst_dob_i32_008 ,\u_img/inst_dob_i32_007 ,\u_img/inst_dob_i32_006 ,\u_img/inst_dob_i32_005 ,\u_img/inst_dob_i32_004 ,\u_img/inst_dob_i32_003 ,\u_img/inst_dob_i32_002 ,\u_img/inst_dob_i32_001 ,\u_img/inst_dob_i32_000 }));
  // address_offset=16384;data_offset=9;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("INV"),
    .CSB1("SIG"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_img/inst_32800x16_sub_016384_009  (
    .addra(camera_addr[12:0]),
    .addrb(vga_rdaddr[12:0]),
    .cea(camera_wrreq),
    .ceb(vga_rden),
    .clka(cam_pclk_pad),
    .clkb(clk_lcd),
    .csa(camera_addr[15:13]),
    .csb(vga_rdaddr[15:13]),
    .dia({open_n1732,open_n1733,open_n1734,open_n1735,open_n1736,open_n1737,open_n1738,camera_wrdat[9],open_n1739}),
    .rsta(cam_rst_pad),
    .rstb(cam_rst_pad),
    .dob({open_n1762,open_n1763,open_n1764,open_n1765,open_n1766,open_n1767,open_n1768,open_n1769,\u_img/inst_dob_i32_009 }));
  // address_offset=16384;data_offset=10;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("INV"),
    .CSB1("SIG"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_img/inst_32800x16_sub_016384_010  (
    .addra(camera_addr[12:0]),
    .addrb(vga_rdaddr[12:0]),
    .cea(camera_wrreq),
    .ceb(vga_rden),
    .clka(cam_pclk_pad),
    .clkb(clk_lcd),
    .csa(camera_addr[15:13]),
    .csb(vga_rdaddr[15:13]),
    .dia({open_n1770,open_n1771,open_n1772,open_n1773,open_n1774,open_n1775,open_n1776,camera_wrdat[10],open_n1777}),
    .rsta(cam_rst_pad),
    .rstb(cam_rst_pad),
    .dob({open_n1800,open_n1801,open_n1802,open_n1803,open_n1804,open_n1805,open_n1806,open_n1807,\u_img/inst_dob_i32_010 }));
  // address_offset=16384;data_offset=11;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("INV"),
    .CSB1("SIG"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_img/inst_32800x16_sub_016384_011  (
    .addra(camera_addr[12:0]),
    .addrb(vga_rdaddr[12:0]),
    .cea(camera_wrreq),
    .ceb(vga_rden),
    .clka(cam_pclk_pad),
    .clkb(clk_lcd),
    .csa(camera_addr[15:13]),
    .csb(vga_rdaddr[15:13]),
    .dia({open_n1808,open_n1809,open_n1810,open_n1811,open_n1812,open_n1813,open_n1814,camera_wrdat[11],open_n1815}),
    .rsta(cam_rst_pad),
    .rstb(cam_rst_pad),
    .dob({open_n1838,open_n1839,open_n1840,open_n1841,open_n1842,open_n1843,open_n1844,open_n1845,\u_img/inst_dob_i32_011 }));
  // address_offset=16384;data_offset=12;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("INV"),
    .CSB1("SIG"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_img/inst_32800x16_sub_016384_012  (
    .addra(camera_addr[12:0]),
    .addrb(vga_rdaddr[12:0]),
    .cea(camera_wrreq),
    .ceb(vga_rden),
    .clka(cam_pclk_pad),
    .clkb(clk_lcd),
    .csa(camera_addr[15:13]),
    .csb(vga_rdaddr[15:13]),
    .dia({open_n1846,open_n1847,open_n1848,open_n1849,open_n1850,open_n1851,open_n1852,camera_wrdat[12],open_n1853}),
    .rsta(cam_rst_pad),
    .rstb(cam_rst_pad),
    .dob({open_n1876,open_n1877,open_n1878,open_n1879,open_n1880,open_n1881,open_n1882,open_n1883,\u_img/inst_dob_i32_012 }));
  // address_offset=16384;data_offset=13;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("INV"),
    .CSB1("SIG"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_img/inst_32800x16_sub_016384_013  (
    .addra(camera_addr[12:0]),
    .addrb(vga_rdaddr[12:0]),
    .cea(camera_wrreq),
    .ceb(vga_rden),
    .clka(cam_pclk_pad),
    .clkb(clk_lcd),
    .csa(camera_addr[15:13]),
    .csb(vga_rdaddr[15:13]),
    .dia({open_n1884,open_n1885,open_n1886,open_n1887,open_n1888,open_n1889,open_n1890,camera_wrdat[13],open_n1891}),
    .rsta(cam_rst_pad),
    .rstb(cam_rst_pad),
    .dob({open_n1914,open_n1915,open_n1916,open_n1917,open_n1918,open_n1919,open_n1920,open_n1921,\u_img/inst_dob_i32_013 }));
  // address_offset=16384;data_offset=14;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("INV"),
    .CSB1("SIG"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_img/inst_32800x16_sub_016384_014  (
    .addra(camera_addr[12:0]),
    .addrb(vga_rdaddr[12:0]),
    .cea(camera_wrreq),
    .ceb(vga_rden),
    .clka(cam_pclk_pad),
    .clkb(clk_lcd),
    .csa(camera_addr[15:13]),
    .csb(vga_rdaddr[15:13]),
    .dia({open_n1922,open_n1923,open_n1924,open_n1925,open_n1926,open_n1927,open_n1928,camera_wrdat[14],open_n1929}),
    .rsta(cam_rst_pad),
    .rstb(cam_rst_pad),
    .dob({open_n1952,open_n1953,open_n1954,open_n1955,open_n1956,open_n1957,open_n1958,open_n1959,\u_img/inst_dob_i32_014 }));
  // address_offset=16384;data_offset=15;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("INV"),
    .CSB1("SIG"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_img/inst_32800x16_sub_016384_015  (
    .addra(camera_addr[12:0]),
    .addrb(vga_rdaddr[12:0]),
    .cea(camera_wrreq),
    .ceb(vga_rden),
    .clka(cam_pclk_pad),
    .clkb(clk_lcd),
    .csa(camera_addr[15:13]),
    .csb(vga_rdaddr[15:13]),
    .dia({open_n1960,open_n1961,open_n1962,open_n1963,open_n1964,open_n1965,open_n1966,camera_wrdat[15],open_n1967}),
    .rsta(cam_rst_pad),
    .rstb(cam_rst_pad),
    .dob({open_n1990,open_n1991,open_n1992,open_n1993,open_n1994,open_n1995,open_n1996,open_n1997,\u_img/inst_dob_i32_015 }));
  // address_offset=17408;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("SIG"),
    .CSB1("INV"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_img/inst_32800x16_sub_017408_000  (
    .addra({camera_addr[9:0],3'b111}),
    .addrb({vga_rdaddr[9:0],3'b111}),
    .cea(camera_wrreq),
    .ceb(vga_rden),
    .clka(cam_pclk_pad),
    .clkb(clk_lcd),
    .csa({\and_Ncamera_addr[12]_o_al_n208 ,camera_addr[11:10]}),
    .csb({\and_Nvga_rdaddr[12]__o_al_n211 ,vga_rdaddr[11:10]}),
    .dia(camera_wrdat[8:0]),
    .rsta(cam_rst_pad),
    .rstb(cam_rst_pad),
    .dob({\u_img/inst_dob_i34_008 ,\u_img/inst_dob_i34_007 ,\u_img/inst_dob_i34_006 ,\u_img/inst_dob_i34_005 ,\u_img/inst_dob_i34_004 ,\u_img/inst_dob_i34_003 ,\u_img/inst_dob_i34_002 ,\u_img/inst_dob_i34_001 ,\u_img/inst_dob_i34_000 }));
  // address_offset=18432;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("INV"),
    .CSB1("SIG"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_img/inst_32800x16_sub_018432_000  (
    .addra({camera_addr[9:0],3'b111}),
    .addrb({vga_rdaddr[9:0],3'b111}),
    .cea(camera_wrreq),
    .ceb(vga_rden),
    .clka(cam_pclk_pad),
    .clkb(clk_lcd),
    .csa({\and_Ncamera_addr[12]_o_al_n208 ,camera_addr[11:10]}),
    .csb({\and_Nvga_rdaddr[12]__o_al_n211 ,vga_rdaddr[11:10]}),
    .dia(camera_wrdat[8:0]),
    .rsta(cam_rst_pad),
    .rstb(cam_rst_pad),
    .dob({\u_img/inst_dob_i36_008 ,\u_img/inst_dob_i36_007 ,\u_img/inst_dob_i36_006 ,\u_img/inst_dob_i36_005 ,\u_img/inst_dob_i36_004 ,\u_img/inst_dob_i36_003 ,\u_img/inst_dob_i36_002 ,\u_img/inst_dob_i36_001 ,\u_img/inst_dob_i36_000 }));
  // address_offset=19456;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("SIG"),
    .CSB1("SIG"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_img/inst_32800x16_sub_019456_000  (
    .addra({camera_addr[9:0],3'b111}),
    .addrb({vga_rdaddr[9:0],3'b111}),
    .cea(camera_wrreq),
    .ceb(vga_rden),
    .clka(cam_pclk_pad),
    .clkb(clk_lcd),
    .csa({\and_Ncamera_addr[12]_o_al_n208 ,camera_addr[11:10]}),
    .csb({\and_Nvga_rdaddr[12]__o_al_n211 ,vga_rdaddr[11:10]}),
    .dia(camera_wrdat[8:0]),
    .rsta(cam_rst_pad),
    .rstb(cam_rst_pad),
    .dob({\u_img/inst_dob_i38_008 ,\u_img/inst_dob_i38_007 ,\u_img/inst_dob_i38_006 ,\u_img/inst_dob_i38_005 ,\u_img/inst_dob_i38_004 ,\u_img/inst_dob_i38_003 ,\u_img/inst_dob_i38_002 ,\u_img/inst_dob_i38_001 ,\u_img/inst_dob_i38_000 }));
  // address_offset=20480;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("INV"),
    .CSB1("INV"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_img/inst_32800x16_sub_020480_000  (
    .addra({camera_addr[9:0],3'b111}),
    .addrb({vga_rdaddr[9:0],3'b111}),
    .cea(camera_wrreq),
    .ceb(vga_rden),
    .clka(cam_pclk_pad),
    .clkb(clk_lcd),
    .csa({\and_camera_addr[12]__o_al_n224 ,camera_addr[11:10]}),
    .csb({\and_vga_rdaddr[12]_N_o_al_n227 ,vga_rdaddr[11:10]}),
    .dia(camera_wrdat[8:0]),
    .rsta(cam_rst_pad),
    .rstb(cam_rst_pad),
    .dob({\u_img/inst_dob_i40_008 ,\u_img/inst_dob_i40_007 ,\u_img/inst_dob_i40_006 ,\u_img/inst_dob_i40_005 ,\u_img/inst_dob_i40_004 ,\u_img/inst_dob_i40_003 ,\u_img/inst_dob_i40_002 ,\u_img/inst_dob_i40_001 ,\u_img/inst_dob_i40_000 }));
  // address_offset=21504;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("SIG"),
    .CSB1("INV"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_img/inst_32800x16_sub_021504_000  (
    .addra({camera_addr[9:0],3'b111}),
    .addrb({vga_rdaddr[9:0],3'b111}),
    .cea(camera_wrreq),
    .ceb(vga_rden),
    .clka(cam_pclk_pad),
    .clkb(clk_lcd),
    .csa({\and_camera_addr[12]__o_al_n224 ,camera_addr[11:10]}),
    .csb({\and_vga_rdaddr[12]_N_o_al_n227 ,vga_rdaddr[11:10]}),
    .dia(camera_wrdat[8:0]),
    .rsta(cam_rst_pad),
    .rstb(cam_rst_pad),
    .dob({\u_img/inst_dob_i42_008 ,\u_img/inst_dob_i42_007 ,\u_img/inst_dob_i42_006 ,\u_img/inst_dob_i42_005 ,\u_img/inst_dob_i42_004 ,\u_img/inst_dob_i42_003 ,\u_img/inst_dob_i42_002 ,\u_img/inst_dob_i42_001 ,\u_img/inst_dob_i42_000 }));
  // address_offset=22528;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("INV"),
    .CSB1("SIG"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_img/inst_32800x16_sub_022528_000  (
    .addra({camera_addr[9:0],3'b111}),
    .addrb({vga_rdaddr[9:0],3'b111}),
    .cea(camera_wrreq),
    .ceb(vga_rden),
    .clka(cam_pclk_pad),
    .clkb(clk_lcd),
    .csa({\and_camera_addr[12]__o_al_n224 ,camera_addr[11:10]}),
    .csb({\and_vga_rdaddr[12]_N_o_al_n227 ,vga_rdaddr[11:10]}),
    .dia(camera_wrdat[8:0]),
    .rsta(cam_rst_pad),
    .rstb(cam_rst_pad),
    .dob({\u_img/inst_dob_i44_008 ,\u_img/inst_dob_i44_007 ,\u_img/inst_dob_i44_006 ,\u_img/inst_dob_i44_005 ,\u_img/inst_dob_i44_004 ,\u_img/inst_dob_i44_003 ,\u_img/inst_dob_i44_002 ,\u_img/inst_dob_i44_001 ,\u_img/inst_dob_i44_000 }));
  // address_offset=23552;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("SIG"),
    .CSB1("SIG"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_img/inst_32800x16_sub_023552_000  (
    .addra({camera_addr[9:0],3'b111}),
    .addrb({vga_rdaddr[9:0],3'b111}),
    .cea(camera_wrreq),
    .ceb(vga_rden),
    .clka(cam_pclk_pad),
    .clkb(clk_lcd),
    .csa({\and_camera_addr[12]__o_al_n224 ,camera_addr[11:10]}),
    .csb({\and_vga_rdaddr[12]_N_o_al_n227 ,vga_rdaddr[11:10]}),
    .dia(camera_wrdat[8:0]),
    .rsta(cam_rst_pad),
    .rstb(cam_rst_pad),
    .dob({\u_img/inst_dob_i46_008 ,\u_img/inst_dob_i46_007 ,\u_img/inst_dob_i46_006 ,\u_img/inst_dob_i46_005 ,\u_img/inst_dob_i46_004 ,\u_img/inst_dob_i46_003 ,\u_img/inst_dob_i46_002 ,\u_img/inst_dob_i46_001 ,\u_img/inst_dob_i46_000 }));
  // address_offset=24576;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("INV"),
    .CSB1("INV"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_img/inst_32800x16_sub_024576_000  (
    .addra({camera_addr[9:0],3'b111}),
    .addrb({vga_rdaddr[9:0],3'b111}),
    .cea(camera_wrreq),
    .ceb(vga_rden),
    .clka(cam_pclk_pad),
    .clkb(clk_lcd),
    .csa({\and_Ncamera_addr[12]_o_al_n240 ,camera_addr[11:10]}),
    .csb({\and_Nvga_rdaddr[12]__o_al_n243 ,vga_rdaddr[11:10]}),
    .dia(camera_wrdat[8:0]),
    .rsta(cam_rst_pad),
    .rstb(cam_rst_pad),
    .dob({\u_img/inst_dob_i48_008 ,\u_img/inst_dob_i48_007 ,\u_img/inst_dob_i48_006 ,\u_img/inst_dob_i48_005 ,\u_img/inst_dob_i48_004 ,\u_img/inst_dob_i48_003 ,\u_img/inst_dob_i48_002 ,\u_img/inst_dob_i48_001 ,\u_img/inst_dob_i48_000 }));
  // address_offset=24576;data_offset=9;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("SIG"),
    .CSB1("SIG"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_img/inst_32800x16_sub_024576_009  (
    .addra(camera_addr[12:0]),
    .addrb(vga_rdaddr[12:0]),
    .cea(camera_wrreq),
    .ceb(vga_rden),
    .clka(cam_pclk_pad),
    .clkb(clk_lcd),
    .csa(camera_addr[15:13]),
    .csb(vga_rdaddr[15:13]),
    .dia({open_n2174,open_n2175,open_n2176,open_n2177,open_n2178,open_n2179,open_n2180,camera_wrdat[9],open_n2181}),
    .rsta(cam_rst_pad),
    .rstb(cam_rst_pad),
    .dob({open_n2204,open_n2205,open_n2206,open_n2207,open_n2208,open_n2209,open_n2210,open_n2211,\u_img/inst_dob_i48_009 }));
  // address_offset=24576;data_offset=10;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("SIG"),
    .CSB1("SIG"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_img/inst_32800x16_sub_024576_010  (
    .addra(camera_addr[12:0]),
    .addrb(vga_rdaddr[12:0]),
    .cea(camera_wrreq),
    .ceb(vga_rden),
    .clka(cam_pclk_pad),
    .clkb(clk_lcd),
    .csa(camera_addr[15:13]),
    .csb(vga_rdaddr[15:13]),
    .dia({open_n2212,open_n2213,open_n2214,open_n2215,open_n2216,open_n2217,open_n2218,camera_wrdat[10],open_n2219}),
    .rsta(cam_rst_pad),
    .rstb(cam_rst_pad),
    .dob({open_n2242,open_n2243,open_n2244,open_n2245,open_n2246,open_n2247,open_n2248,open_n2249,\u_img/inst_dob_i48_010 }));
  // address_offset=24576;data_offset=11;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("SIG"),
    .CSB1("SIG"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_img/inst_32800x16_sub_024576_011  (
    .addra(camera_addr[12:0]),
    .addrb(vga_rdaddr[12:0]),
    .cea(camera_wrreq),
    .ceb(vga_rden),
    .clka(cam_pclk_pad),
    .clkb(clk_lcd),
    .csa(camera_addr[15:13]),
    .csb(vga_rdaddr[15:13]),
    .dia({open_n2250,open_n2251,open_n2252,open_n2253,open_n2254,open_n2255,open_n2256,camera_wrdat[11],open_n2257}),
    .rsta(cam_rst_pad),
    .rstb(cam_rst_pad),
    .dob({open_n2280,open_n2281,open_n2282,open_n2283,open_n2284,open_n2285,open_n2286,open_n2287,\u_img/inst_dob_i48_011 }));
  // address_offset=24576;data_offset=12;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("SIG"),
    .CSB1("SIG"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_img/inst_32800x16_sub_024576_012  (
    .addra(camera_addr[12:0]),
    .addrb(vga_rdaddr[12:0]),
    .cea(camera_wrreq),
    .ceb(vga_rden),
    .clka(cam_pclk_pad),
    .clkb(clk_lcd),
    .csa(camera_addr[15:13]),
    .csb(vga_rdaddr[15:13]),
    .dia({open_n2288,open_n2289,open_n2290,open_n2291,open_n2292,open_n2293,open_n2294,camera_wrdat[12],open_n2295}),
    .rsta(cam_rst_pad),
    .rstb(cam_rst_pad),
    .dob({open_n2318,open_n2319,open_n2320,open_n2321,open_n2322,open_n2323,open_n2324,open_n2325,\u_img/inst_dob_i48_012 }));
  // address_offset=24576;data_offset=13;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("SIG"),
    .CSB1("SIG"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_img/inst_32800x16_sub_024576_013  (
    .addra(camera_addr[12:0]),
    .addrb(vga_rdaddr[12:0]),
    .cea(camera_wrreq),
    .ceb(vga_rden),
    .clka(cam_pclk_pad),
    .clkb(clk_lcd),
    .csa(camera_addr[15:13]),
    .csb(vga_rdaddr[15:13]),
    .dia({open_n2326,open_n2327,open_n2328,open_n2329,open_n2330,open_n2331,open_n2332,camera_wrdat[13],open_n2333}),
    .rsta(cam_rst_pad),
    .rstb(cam_rst_pad),
    .dob({open_n2356,open_n2357,open_n2358,open_n2359,open_n2360,open_n2361,open_n2362,open_n2363,\u_img/inst_dob_i48_013 }));
  // address_offset=24576;data_offset=14;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("SIG"),
    .CSB1("SIG"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_img/inst_32800x16_sub_024576_014  (
    .addra(camera_addr[12:0]),
    .addrb(vga_rdaddr[12:0]),
    .cea(camera_wrreq),
    .ceb(vga_rden),
    .clka(cam_pclk_pad),
    .clkb(clk_lcd),
    .csa(camera_addr[15:13]),
    .csb(vga_rdaddr[15:13]),
    .dia({open_n2364,open_n2365,open_n2366,open_n2367,open_n2368,open_n2369,open_n2370,camera_wrdat[14],open_n2371}),
    .rsta(cam_rst_pad),
    .rstb(cam_rst_pad),
    .dob({open_n2394,open_n2395,open_n2396,open_n2397,open_n2398,open_n2399,open_n2400,open_n2401,\u_img/inst_dob_i48_014 }));
  // address_offset=24576;data_offset=15;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("SIG"),
    .CSB1("SIG"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_img/inst_32800x16_sub_024576_015  (
    .addra(camera_addr[12:0]),
    .addrb(vga_rdaddr[12:0]),
    .cea(camera_wrreq),
    .ceb(vga_rden),
    .clka(cam_pclk_pad),
    .clkb(clk_lcd),
    .csa(camera_addr[15:13]),
    .csb(vga_rdaddr[15:13]),
    .dia({open_n2402,open_n2403,open_n2404,open_n2405,open_n2406,open_n2407,open_n2408,camera_wrdat[15],open_n2409}),
    .rsta(cam_rst_pad),
    .rstb(cam_rst_pad),
    .dob({open_n2432,open_n2433,open_n2434,open_n2435,open_n2436,open_n2437,open_n2438,open_n2439,\u_img/inst_dob_i48_015 }));
  // address_offset=25600;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("SIG"),
    .CSB1("INV"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_img/inst_32800x16_sub_025600_000  (
    .addra({camera_addr[9:0],3'b111}),
    .addrb({vga_rdaddr[9:0],3'b111}),
    .cea(camera_wrreq),
    .ceb(vga_rden),
    .clka(cam_pclk_pad),
    .clkb(clk_lcd),
    .csa({\and_Ncamera_addr[12]_o_al_n240 ,camera_addr[11:10]}),
    .csb({\and_Nvga_rdaddr[12]__o_al_n243 ,vga_rdaddr[11:10]}),
    .dia(camera_wrdat[8:0]),
    .rsta(cam_rst_pad),
    .rstb(cam_rst_pad),
    .dob({\u_img/inst_dob_i50_008 ,\u_img/inst_dob_i50_007 ,\u_img/inst_dob_i50_006 ,\u_img/inst_dob_i50_005 ,\u_img/inst_dob_i50_004 ,\u_img/inst_dob_i50_003 ,\u_img/inst_dob_i50_002 ,\u_img/inst_dob_i50_001 ,\u_img/inst_dob_i50_000 }));
  // address_offset=26624;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("INV"),
    .CSB1("SIG"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_img/inst_32800x16_sub_026624_000  (
    .addra({camera_addr[9:0],3'b111}),
    .addrb({vga_rdaddr[9:0],3'b111}),
    .cea(camera_wrreq),
    .ceb(vga_rden),
    .clka(cam_pclk_pad),
    .clkb(clk_lcd),
    .csa({\and_Ncamera_addr[12]_o_al_n240 ,camera_addr[11:10]}),
    .csb({\and_Nvga_rdaddr[12]__o_al_n243 ,vga_rdaddr[11:10]}),
    .dia(camera_wrdat[8:0]),
    .rsta(cam_rst_pad),
    .rstb(cam_rst_pad),
    .dob({\u_img/inst_dob_i52_008 ,\u_img/inst_dob_i52_007 ,\u_img/inst_dob_i52_006 ,\u_img/inst_dob_i52_005 ,\u_img/inst_dob_i52_004 ,\u_img/inst_dob_i52_003 ,\u_img/inst_dob_i52_002 ,\u_img/inst_dob_i52_001 ,\u_img/inst_dob_i52_000 }));
  // address_offset=27648;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("SIG"),
    .CSB1("SIG"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_img/inst_32800x16_sub_027648_000  (
    .addra({camera_addr[9:0],3'b111}),
    .addrb({vga_rdaddr[9:0],3'b111}),
    .cea(camera_wrreq),
    .ceb(vga_rden),
    .clka(cam_pclk_pad),
    .clkb(clk_lcd),
    .csa({\and_Ncamera_addr[12]_o_al_n240 ,camera_addr[11:10]}),
    .csb({\and_Nvga_rdaddr[12]__o_al_n243 ,vga_rdaddr[11:10]}),
    .dia(camera_wrdat[8:0]),
    .rsta(cam_rst_pad),
    .rstb(cam_rst_pad),
    .dob({\u_img/inst_dob_i54_008 ,\u_img/inst_dob_i54_007 ,\u_img/inst_dob_i54_006 ,\u_img/inst_dob_i54_005 ,\u_img/inst_dob_i54_004 ,\u_img/inst_dob_i54_003 ,\u_img/inst_dob_i54_002 ,\u_img/inst_dob_i54_001 ,\u_img/inst_dob_i54_000 }));
  // address_offset=28672;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("INV"),
    .CSB1("INV"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_img/inst_32800x16_sub_028672_000  (
    .addra({camera_addr[9:0],3'b111}),
    .addrb({vga_rdaddr[9:0],3'b111}),
    .cea(camera_wrreq),
    .ceb(vga_rden),
    .clka(cam_pclk_pad),
    .clkb(clk_lcd),
    .csa({\and_camera_addr[12]__o_al_n256 ,camera_addr[11:10]}),
    .csb({\and_vga_rdaddr[12]_v_o_al_n259 ,vga_rdaddr[11:10]}),
    .dia(camera_wrdat[8:0]),
    .rsta(cam_rst_pad),
    .rstb(cam_rst_pad),
    .dob({\u_img/inst_dob_i56_008 ,\u_img/inst_dob_i56_007 ,\u_img/inst_dob_i56_006 ,\u_img/inst_dob_i56_005 ,\u_img/inst_dob_i56_004 ,\u_img/inst_dob_i56_003 ,\u_img/inst_dob_i56_002 ,\u_img/inst_dob_i56_001 ,\u_img/inst_dob_i56_000 }));
  // address_offset=29696;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("SIG"),
    .CSB1("INV"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_img/inst_32800x16_sub_029696_000  (
    .addra({camera_addr[9:0],3'b111}),
    .addrb({vga_rdaddr[9:0],3'b111}),
    .cea(camera_wrreq),
    .ceb(vga_rden),
    .clka(cam_pclk_pad),
    .clkb(clk_lcd),
    .csa({\and_camera_addr[12]__o_al_n256 ,camera_addr[11:10]}),
    .csb({\and_vga_rdaddr[12]_v_o_al_n259 ,vga_rdaddr[11:10]}),
    .dia(camera_wrdat[8:0]),
    .rsta(cam_rst_pad),
    .rstb(cam_rst_pad),
    .dob({\u_img/inst_dob_i58_008 ,\u_img/inst_dob_i58_007 ,\u_img/inst_dob_i58_006 ,\u_img/inst_dob_i58_005 ,\u_img/inst_dob_i58_004 ,\u_img/inst_dob_i58_003 ,\u_img/inst_dob_i58_002 ,\u_img/inst_dob_i58_001 ,\u_img/inst_dob_i58_000 }));
  // address_offset=30720;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("INV"),
    .CSB1("SIG"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_img/inst_32800x16_sub_030720_000  (
    .addra({camera_addr[9:0],3'b111}),
    .addrb({vga_rdaddr[9:0],3'b111}),
    .cea(camera_wrreq),
    .ceb(vga_rden),
    .clka(cam_pclk_pad),
    .clkb(clk_lcd),
    .csa({\and_camera_addr[12]__o_al_n256 ,camera_addr[11:10]}),
    .csb({\and_vga_rdaddr[12]_v_o_al_n259 ,vga_rdaddr[11:10]}),
    .dia(camera_wrdat[8:0]),
    .rsta(cam_rst_pad),
    .rstb(cam_rst_pad),
    .dob({\u_img/inst_dob_i60_008 ,\u_img/inst_dob_i60_007 ,\u_img/inst_dob_i60_006 ,\u_img/inst_dob_i60_005 ,\u_img/inst_dob_i60_004 ,\u_img/inst_dob_i60_003 ,\u_img/inst_dob_i60_002 ,\u_img/inst_dob_i60_001 ,\u_img/inst_dob_i60_000 }));
  // address_offset=31744;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("SIG"),
    .CSB1("SIG"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_img/inst_32800x16_sub_031744_000  (
    .addra({camera_addr[9:0],3'b111}),
    .addrb({vga_rdaddr[9:0],3'b111}),
    .cea(camera_wrreq),
    .ceb(vga_rden),
    .clka(cam_pclk_pad),
    .clkb(clk_lcd),
    .csa({\and_camera_addr[12]__o_al_n256 ,camera_addr[11:10]}),
    .csb({\and_vga_rdaddr[12]_v_o_al_n259 ,vga_rdaddr[11:10]}),
    .dia(camera_wrdat[8:0]),
    .rsta(cam_rst_pad),
    .rstb(cam_rst_pad),
    .dob({\u_img/inst_dob_i62_008 ,\u_img/inst_dob_i62_007 ,\u_img/inst_dob_i62_006 ,\u_img/inst_dob_i62_005 ,\u_img/inst_dob_i62_004 ,\u_img/inst_dob_i62_003 ,\u_img/inst_dob_i62_002 ,\u_img/inst_dob_i62_001 ,\u_img/inst_dob_i62_000 }));
  // address_offset=32768;data_offset=0;depth=32;width=16;num_section=1;width_per_section=16;section_size=16;working_depth=512;working_width=18;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("1"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("INV"),
    .CSB1("INV"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("18"),
    .DATA_WIDTH_B("18"),
    .MODE("PDPW8K"),
    .OCEAMUX("1"),
    .OCEBMUX("1"),
    .REGMODE_A("OUTREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_img/inst_32800x16_sub_032768_000  (
    .addra({camera_addr[8:0],4'b1111}),
    .addrb({vga_rdaddr[8:0],4'b1111}),
    .clka(cam_pclk_pad),
    .clkb(clk_lcd),
    .csa({\and_Ncamera_addr[11]_o_and_camera_wrreq ,camera_addr[10:9]}),
    .csb({\and_Nvga_rdaddr[11]__o_and_vga_rden ,vga_rdaddr[10:9]}),
    .dia(camera_wrdat[8:0]),
    .dib({open_n2596,open_n2597,camera_wrdat[15:9]}),
    .rsta(cam_rst_pad),
    .rstb(cam_rst_pad),
    .doa({\u_img/inst_dob_i64_008 ,\u_img/inst_dob_i64_007 ,\u_img/inst_dob_i64_006 ,\u_img/inst_dob_i64_005 ,\u_img/inst_dob_i64_004 ,\u_img/inst_dob_i64_003 ,\u_img/inst_dob_i64_002 ,\u_img/inst_dob_i64_001 ,\u_img/inst_dob_i64_000 }),
    .dob({open_n2602,open_n2603,\u_img/inst_dob_i64_015 ,\u_img/inst_dob_i64_014 ,\u_img/inst_dob_i64_013 ,\u_img/inst_dob_i64_012 ,\u_img/inst_dob_i64_011 ,\u_img/inst_dob_i64_010 ,\u_img/inst_dob_i64_009 }));
  EG_PHY_GCLK \u_pll/bufg_feedback  (
    .clki(\u_pll/clk0_buf ),
    .clko(clk_lcd));  // al_ip/ip_pll.v(36)
  EG_PHY_PLL #(
    .CLKC0_CPHASE(19),
    .CLKC0_DIV(20),
    .CLKC0_DIV2_ENABLE("DISABLE"),
    .CLKC0_ENABLE("ENABLE"),
    .CLKC0_FPHASE(0),
    .CLKC1_CPHASE(41),
    .CLKC1_DIV(42),
    .CLKC1_DIV2_ENABLE("DISABLE"),
    .CLKC1_ENABLE("ENABLE"),
    .CLKC1_FPHASE(0),
    .CLKC2_CPHASE(125),
    .CLKC2_DIV(126),
    .CLKC2_DIV2_ENABLE("DISABLE"),
    .CLKC2_ENABLE("ENABLE"),
    .CLKC2_FPHASE(0),
    .CLKC3_CPHASE(1),
    .CLKC3_DIV(1),
    .CLKC3_DIV2_ENABLE("DISABLE"),
    .CLKC3_ENABLE("DISABLE"),
    .CLKC3_FPHASE(0),
    .CLKC4_CPHASE(1),
    .CLKC4_DIV(1),
    .CLKC4_DIV2_ENABLE("DISABLE"),
    .CLKC4_ENABLE("DISABLE"),
    .CLKC4_FPHASE(0),
    .DERIVE_PLL_CLOCKS("DISABLE"),
    .DPHASE_SOURCE("DISABLE"),
    .DYNCFG("DISABLE"),
    .FBCLK_DIV(17),
    .FEEDBK_MODE("NORMAL"),
    .FEEDBK_PATH("CLKC0_EXT"),
    .FIN("24.000"),
    .FREQ_LOCK_ACCURACY(2),
    .GEN_BASIC_CLOCK("DISABLE"),
    .GMC_GAIN(6),
    .GMC_TEST(14),
    .ICP_CURRENT(3),
    .IF_ESCLKSTSW("DISABLE"),
    .INTFB_WAKE("DISABLE"),
    .KVCO(6),
    .LPF_CAPACITOR(3),
    .LPF_RESISTOR(2),
    .NORESET("DISABLE"),
    .ODIV_MUXC0("DIV"),
    .ODIV_MUXC1("DIV"),
    .ODIV_MUXC2("DIV"),
    .ODIV_MUXC3("DIV"),
    .ODIV_MUXC4("DIV"),
    .PLLC2RST_ENA("DISABLE"),
    .PLLC34RST_ENA("DISABLE"),
    .PLLMRST_ENA("DISABLE"),
    .PLLRST_ENA("DISABLE"),
    .PLL_LOCK_MODE(0),
    .PREDIV_MUXC0("VCO"),
    .PREDIV_MUXC1("VCO"),
    .PREDIV_MUXC2("VCO"),
    .PREDIV_MUXC3("VCO"),
    .PREDIV_MUXC4("VCO"),
    .REFCLK_DIV(16),
    .REFCLK_SEL("INTERNAL"),
    .STDBY_ENABLE("DISABLE"),
    .STDBY_VCO_ENA("DISABLE"),
    .SYNC_ENABLE("DISABLE"),
    .VCO_NORESET("DISABLE"))
    \u_pll/pll_inst  (
    .daddr(6'b000000),
    .dclk(1'b0),
    .dcs(1'b0),
    .di(8'b00000000),
    .dwe(1'b0),
    .fbclk(clk_lcd),
    .psclk(1'b0),
    .psclksel(3'b000),
    .psdown(1'b0),
    .psstep(1'b0),
    .refclk(clk_24m_pad),
    .reset(1'b0),
    .stdby(1'b0),
    .clkc({open_n2604,open_n2605,clk_sccb,clk_cam,\u_pll/clk0_buf }));  // al_ip/ip_pll.v(67)
  \lcd_sync(IMG_Y=1)  u_vga_sync (
    .clk(clk_lcd),
    .rest_n(cam_rst_pad),
    .addr(vga_rdaddr),
    .img_ack(vga_rden),
    .lcd_clk(vga_clk_pad),
    .lcd_hsync(vga_hsync_pad),
    .lcd_vsync(vga_vsync_pad));  // sources/rtl/test_camera.v(102)
  reg_sr_as_w1 vga_rdaddr_pipe_b0 (
    .clk(clk_lcd),
    .d(vga_rdaddr[9]),
    .en(vga_rden),
    .reset(cam_rst_pad_neg),
    .set(1'b0),
    .q(vga_rdaddr_piped[0]));
  reg_sr_as_w1 vga_rdaddr_pipe_b1 (
    .clk(clk_lcd),
    .d(vga_rdaddr[10]),
    .en(vga_rden),
    .reset(cam_rst_pad_neg),
    .set(1'b0),
    .q(vga_rdaddr_piped[1]));
  reg_sr_as_w1 vga_rdaddr_pipe_b2 (
    .clk(clk_lcd),
    .d(vga_rdaddr[11]),
    .en(vga_rden),
    .reset(cam_rst_pad_neg),
    .set(1'b0),
    .q(vga_rdaddr_piped[2]));
  reg_sr_as_w1 vga_rdaddr_pipe_b3 (
    .clk(clk_lcd),
    .d(vga_rdaddr[12]),
    .en(vga_rden),
    .reset(cam_rst_pad_neg),
    .set(1'b0),
    .q(vga_rdaddr_piped[3]));
  reg_sr_as_w1 vga_rdaddr_pipe_b4 (
    .clk(clk_lcd),
    .d(vga_rdaddr[13]),
    .en(vga_rden),
    .reset(cam_rst_pad_neg),
    .set(1'b0),
    .q(vga_rdaddr_piped[4]));
  reg_sr_as_w1 vga_rdaddr_pipe_b5 (
    .clk(clk_lcd),
    .d(vga_rdaddr[14]),
    .en(vga_rden),
    .reset(cam_rst_pad_neg),
    .set(1'b0),
    .q(vga_rdaddr_piped[5]));
  reg_sr_as_w1 vga_rdaddr_pipe_b6 (
    .clk(clk_lcd),
    .d(vga_rdaddr[15]),
    .en(vga_rden),
    .reset(cam_rst_pad_neg),
    .set(1'b0),
    .q(vga_rdaddr_piped[6]));
  reg_sr_as_w1 vga_rdaddr_piped_pipe_b0 (
    .clk(clk_lcd),
    .d(vga_rdaddr_piped[0]),
    .en(vga_rden),
    .reset(cam_rst_pad_neg),
    .set(1'b0));
  reg_sr_as_w1 vga_rdaddr_piped_pipe_b1 (
    .clk(clk_lcd),
    .d(vga_rdaddr_piped[1]),
    .en(vga_rden),
    .reset(cam_rst_pad_neg),
    .set(1'b0),
    .q(vga_rdaddr_piped_piped[1]));
  reg_sr_as_w1 vga_rdaddr_piped_pipe_b2 (
    .clk(clk_lcd),
    .d(vga_rdaddr_piped[2]),
    .en(vga_rden),
    .reset(cam_rst_pad_neg),
    .set(1'b0),
    .q(vga_rdaddr_piped_piped[2]));
  reg_sr_as_w1 vga_rdaddr_piped_pipe_b3 (
    .clk(clk_lcd),
    .d(vga_rdaddr_piped[3]),
    .en(vga_rden),
    .reset(cam_rst_pad_neg),
    .set(1'b0),
    .q(vga_rdaddr_piped_piped[3]));
  reg_sr_as_w1 vga_rdaddr_piped_pipe_b4 (
    .clk(clk_lcd),
    .d(vga_rdaddr_piped[4]),
    .en(vga_rden),
    .reset(cam_rst_pad_neg),
    .set(1'b0),
    .q(vga_rdaddr_piped_piped[4]));
  reg_sr_as_w1 vga_rdaddr_piped_pipe_b5 (
    .clk(clk_lcd),
    .d(vga_rdaddr_piped[5]),
    .en(vga_rden),
    .reset(cam_rst_pad_neg),
    .set(1'b0),
    .q(vga_rdaddr_piped_piped[5]));
  reg_sr_as_w1 vga_rdaddr_piped_pipe_b6 (
    .clk(clk_lcd),
    .d(vga_rdaddr_piped[6]),
    .en(vga_rden),
    .reset(cam_rst_pad_neg),
    .set(1'b0),
    .q(vga_rdaddr_piped_piped[6]));

endmodule 

module camera_init  // sources/rtl/camera_init.v(14)
  (
  clk,
  reset_n,
  sda_in,
  ready,
  scl,
  sda,
  sda_oe
  );

  input clk;  // sources/rtl/camera_init.v(15)
  input reset_n;  // sources/rtl/camera_init.v(16)
  input sda_in;  // sources/rtl/camera_init.v(20)
  output ready;  // sources/rtl/camera_init.v(17)
  output scl;  // sources/rtl/camera_init.v(21)
  output sda;  // sources/rtl/camera_init.v(19)
  output sda_oe;  // sources/rtl/camera_init.v(18)

  parameter REGS_TO_INIT = 178;
  // localparam CAMERA_IDLE = 18;
  // localparam CAMERA_INIT_1 = 11;
  // localparam CAMERA_INIT_2 = 12;
  // localparam CAMERA_INIT_3 = 13;
  // localparam CAMERA_INIT_4 = 14;
  // localparam CAMERA_INIT_5 = 15;
  // localparam CAMERA_INIT_6 = 16;
  // localparam CAMERA_INIT_7 = 17;
  // localparam CONTROL_REG = 3'b000;
  // localparam SLAVE_ADDRESS = 3'b001;
  // localparam SLAVE_DATA_1 = 3'b011;
  // localparam SLAVE_DATA_2 = 3'b100;
  // localparam SLAVE_REG_ADDRESS = 3'b010;
  wire [7:0] cnt;  // sources/rtl/camera_init.v(64)
  wire [7:0] counter;  // sources/rtl/camera_init.v(63)
  wire [7:0] data_in_bus;  // sources/rtl/camera_init.v(42)
  wire [8:0] divider2;  // sources/rtl/camera_init.v(67)
  wire [8:0] n0;
  wire [15:0] n184;
  wire [15:0] n185;
  wire [15:0] n187;
  wire [15:0] n196;
  wire [15:0] n198;
  wire [15:0] n200;
  wire [15:0] n201;
  wire [15:0] n203;
  wire [15:0] n204;
  wire [15:0] n206;
  wire [15:0] n207;
  wire [15:0] n209;
  wire [15:0] n212;
  wire [15:0] n213;
  wire [15:0] n214;
  wire [15:0] n215;
  wire [15:0] n219;
  wire [15:0] n223;
  wire [15:0] n225;
  wire [15:0] n240;
  wire [15:0] n244;
  wire [15:0] n256;
  wire [7:0] n369;
  wire [7:0] n371;
  wire [7:0] n372;
  wire [7:0] n374;
  wire [2:0] n384;
  wire [2:0] reg_address;  // sources/rtl/camera_init.v(43)
  wire [7:0] state_next;  // sources/rtl/camera_init.v(66)
  wire _al_u2836_o;
  wire _al_u2837_o;
  wire _al_u2840_o;
  wire _al_u2841_o;
  wire _al_u2842_o;
  wire _al_u2843_o;
  wire _al_u2852_o;
  wire _al_u2853_o;
  wire _al_u2861_o;
  wire _al_u2862_o;
  wire _al_u2864_o;
  wire _al_u2865_o;
  wire _al_u2866_o;
  wire _al_u2867_o;
  wire _al_u2869_o;
  wire _al_u2870_o;
  wire _al_u2871_o;
  wire _al_u2872_o;
  wire _al_u2873_o;
  wire _al_u2874_o;
  wire _al_u2876_o;
  wire _al_u2877_o;
  wire _al_u2878_o;
  wire _al_u2881_o;
  wire _al_u2883_o;
  wire _al_u2884_o;
  wire _al_u2885_o;
  wire _al_u2886_o;
  wire _al_u2887_o;
  wire _al_u2888_o;
  wire _al_u2889_o;
  wire _al_u2890_o;
  wire _al_u2892_o;
  wire _al_u2893_o;
  wire _al_u2894_o;
  wire _al_u2896_o;
  wire _al_u2897_o;
  wire _al_u2898_o;
  wire _al_u2900_o;
  wire _al_u2901_o;
  wire _al_u2902_o;
  wire _al_u2903_o;
  wire _al_u2905_o;
  wire _al_u2907_o;
  wire _al_u2908_o;
  wire _al_u2909_o;
  wire _al_u2910_o;
  wire _al_u2911_o;
  wire _al_u2912_o;
  wire _al_u2913_o;
  wire _al_u2914_o;
  wire _al_u2917_o;
  wire _al_u2918_o;
  wire _al_u2919_o;
  wire _al_u2921_o;
  wire _al_u2922_o;
  wire _al_u2923_o;
  wire _al_u2924_o;
  wire _al_u2925_o;
  wire _al_u2926_o;
  wire _al_u2927_o;
  wire _al_u2928_o;
  wire _al_u2929_o;
  wire _al_u2930_o;
  wire _al_u2931_o;
  wire _al_u2932_o;
  wire _al_u2934_o;
  wire _al_u2935_o;
  wire _al_u2938_o;
  wire _al_u2939_o;
  wire _al_u2940_o;
  wire _al_u2942_o;
  wire _al_u2944_o;
  wire _al_u2945_o;
  wire _al_u2946_o;
  wire _al_u2949_o;
  wire _al_u2950_o;
  wire _al_u2952_o;
  wire _al_u2955_o;
  wire _al_u2956_o;
  wire _al_u2957_o;
  wire _al_u2958_o;
  wire _al_u2959_o;
  wire _al_u2960_o;
  wire _al_u2961_o;
  wire _al_u2962_o;
  wire _al_u2965_o;
  wire _al_u2967_o;
  wire _al_u2968_o;
  wire _al_u2969_o;
  wire _al_u2970_o;
  wire _al_u2971_o;
  wire _al_u2972_o;
  wire _al_u2973_o;
  wire _al_u2974_o;
  wire _al_u2975_o;
  wire _al_u2976_o;
  wire _al_u2977_o;
  wire _al_u2978_o;
  wire _al_u2979_o;
  wire _al_u2980_o;
  wire _al_u2981_o;
  wire _al_u2982_o;
  wire _al_u2983_o;
  wire _al_u2984_o;
  wire _al_u2986_o;
  wire _al_u2987_o;
  wire _al_u2988_o;
  wire _al_u2989_o;
  wire _al_u2990_o;
  wire _al_u2992_o;
  wire _al_u2993_o;
  wire _al_u2994_o;
  wire _al_u2995_o;
  wire _al_u2996_o;
  wire _al_u2997_o;
  wire _al_u2998_o;
  wire _al_u2999_o;
  wire _al_u3001_o;
  wire _al_u3002_o;
  wire _al_u3003_o;
  wire _al_u3004_o;
  wire _al_u3005_o;
  wire _al_u3006_o;
  wire _al_u3007_o;
  wire _al_u3009_o;
  wire _al_u3010_o;
  wire _al_u3011_o;
  wire _al_u3012_o;
  wire _al_u3013_o;
  wire _al_u3014_o;
  wire _al_u3015_o;
  wire _al_u3017_o;
  wire _al_u3018_o;
  wire _al_u3019_o;
  wire _al_u3020_o;
  wire _al_u3021_o;
  wire _al_u3022_o;
  wire _al_u3024_o;
  wire _al_u3027_o;
  wire _al_u3028_o;
  wire _al_u3029_o;
  wire _al_u3030_o;
  wire _al_u3031_o;
  wire _al_u3032_o;
  wire _al_u3033_o;
  wire _al_u3034_o;
  wire _al_u3036_o;
  wire _al_u3038_o;
  wire _al_u3040_o;
  wire _al_u3041_o;
  wire _al_u3042_o;
  wire _al_u3043_o;
  wire _al_u3044_o;
  wire _al_u3045_o;
  wire _al_u3046_o;
  wire _al_u3048_o;
  wire _al_u3050_o;
  wire _al_u3051_o;
  wire _al_u3052_o;
  wire _al_u3053_o;
  wire _al_u3055_o;
  wire _al_u3057_o;
  wire _al_u3058_o;
  wire _al_u3059_o;
  wire _al_u3060_o;
  wire _al_u3061_o;
  wire _al_u3062_o;
  wire _al_u3063_o;
  wire _al_u3064_o;
  wire _al_u3065_o;
  wire _al_u3066_o;
  wire _al_u3067_o;
  wire _al_u3068_o;
  wire _al_u3069_o;
  wire _al_u3072_o;
  wire _al_u3073_o;
  wire _al_u3074_o;
  wire _al_u3075_o;
  wire _al_u3076_o;
  wire _al_u3077_o;
  wire _al_u3078_o;
  wire _al_u3079_o;
  wire _al_u3080_o;
  wire _al_u3081_o;
  wire _al_u3082_o;
  wire _al_u3083_o;
  wire _al_u3084_o;
  wire _al_u3085_o;
  wire _al_u3086_o;
  wire _al_u3088_o;
  wire _al_u3089_o;
  wire _al_u3090_o;
  wire _al_u3091_o;
  wire _al_u3092_o;
  wire _al_u3094_o;
  wire _al_u3095_o;
  wire _al_u3096_o;
  wire _al_u3097_o;
  wire _al_u3098_o;
  wire _al_u3099_o;
  wire _al_u3100_o;
  wire _al_u3102_o;
  wire _al_u3103_o;
  wire _al_u3104_o;
  wire _al_u3106_o;
  wire _al_u3107_o;
  wire _al_u3109_o;
  wire _al_u3110_o;
  wire _al_u3111_o;
  wire _al_u3112_o;
  wire _al_u3115_o;
  wire _al_u3121_o;
  wire _al_u3122_o;
  wire _al_u3123_o;
  wire _al_u3125_o;
  wire _al_u3127_o;
  wire _al_u3128_o;
  wire _al_u3129_o;
  wire _al_u3131_o;
  wire _al_u3132_o;
  wire _al_u3133_o;
  wire _al_u3134_o;
  wire _al_u3135_o;
  wire _al_u3136_o;
  wire _al_u3137_o;
  wire _al_u3139_o;
  wire _al_u3140_o;
  wire _al_u3142_o;
  wire _al_u3143_o;
  wire _al_u3144_o;
  wire _al_u3145_o;
  wire _al_u3147_o;
  wire _al_u3150_o;
  wire _al_u3151_o;
  wire _al_u3152_o;
  wire _al_u3153_o;
  wire _al_u3154_o;
  wire _al_u3155_o;
  wire _al_u3157_o;
  wire _al_u3160_o;
  wire _al_u3161_o;
  wire _al_u3163_o;
  wire _al_u3164_o;
  wire _al_u3165_o;
  wire _al_u3166_o;
  wire _al_u3167_o;
  wire _al_u3168_o;
  wire _al_u3169_o;
  wire _al_u3170_o;
  wire _al_u3171_o;
  wire _al_u3172_o;
  wire _al_u3173_o;
  wire _al_u3174_o;
  wire _al_u3175_o;
  wire _al_u3176_o;
  wire _al_u3177_o;
  wire _al_u3179_o;
  wire _al_u3180_o;
  wire _al_u3181_o;
  wire _al_u3182_o;
  wire _al_u3184_o;
  wire _al_u3185_o;
  wire _al_u3186_o;
  wire _al_u3188_o;
  wire _al_u3189_o;
  wire _al_u3190_o;
  wire _al_u3191_o;
  wire _al_u3192_o;
  wire _al_u3193_o;
  wire _al_u3194_o;
  wire _al_u3195_o;
  wire _al_u3196_o;
  wire _al_u3197_o;
  wire _al_u3198_o;
  wire _al_u3199_o;
  wire _al_u3200_o;
  wire _al_u3201_o;
  wire _al_u3202_o;
  wire _al_u3203_o;
  wire _al_u3204_o;
  wire _al_u3205_o;
  wire _al_u3206_o;
  wire _al_u3207_o;
  wire _al_u3208_o;
  wire _al_u3209_o;
  wire _al_u3210_o;
  wire _al_u3211_o;
  wire _al_u3212_o;
  wire _al_u3213_o;
  wire _al_u3214_o;
  wire _al_u3215_o;
  wire _al_u3216_o;
  wire _al_u3217_o;
  wire _al_u3219_o;
  wire _al_u3220_o;
  wire _al_u3221_o;
  wire _al_u3222_o;
  wire _al_u3223_o;
  wire _al_u3224_o;
  wire _al_u3225_o;
  wire _al_u3226_o;
  wire _al_u3227_o;
  wire _al_u3231_o;
  wire _al_u3235_o;
  wire _al_u3236_o;
  wire _al_u3237_o;
  wire _al_u3238_o;
  wire _al_u3240_o;
  wire _al_u3241_o;
  wire _al_u3242_o;
  wire _al_u3243_o;
  wire _al_u3244_o;
  wire _al_u3245_o;
  wire _al_u3246_o;
  wire _al_u3247_o;
  wire _al_u3248_o;
  wire _al_u3249_o;
  wire _al_u3250_o;
  wire _al_u3251_o;
  wire _al_u3252_o;
  wire _al_u3253_o;
  wire _al_u3254_o;
  wire _al_u3255_o;
  wire _al_u3256_o;
  wire _al_u3257_o;
  wire _al_u3258_o;
  wire _al_u3259_o;
  wire _al_u3260_o;
  wire _al_u3261_o;
  wire _al_u3262_o;
  wire _al_u3263_o;
  wire _al_u3264_o;
  wire _al_u3265_o;
  wire _al_u3266_o;
  wire _al_u3268_o;
  wire _al_u3269_o;
  wire _al_u3270_o;
  wire _al_u3271_o;
  wire _al_u3272_o;
  wire _al_u3273_o;
  wire _al_u3274_o;
  wire _al_u3275_o;
  wire _al_u3276_o;
  wire _al_u3277_o;
  wire _al_u3278_o;
  wire _al_u3279_o;
  wire _al_u3280_o;
  wire _al_u3281_o;
  wire _al_u3282_o;
  wire _al_u3283_o;
  wire _al_u3288_o;
  wire _al_u3290_o;
  wire _al_u3291_o;
  wire _al_u3292_o;
  wire _al_u3293_o;
  wire _al_u3296_o;
  wire _al_u3299_o;
  wire _al_u3300_o;
  wire _al_u3301_o;
  wire _al_u3302_o;
  wire _al_u3303_o;
  wire _al_u3306_o;
  wire _al_u3307_o;
  wire _al_u3308_o;
  wire _al_u3309_o;
  wire _al_u3310_o;
  wire _al_u3311_o;
  wire _al_u3312_o;
  wire _al_u3313_o;
  wire _al_u3314_o;
  wire _al_u3315_o;
  wire _al_u3317_o;
  wire _al_u3319_o;
  wire _al_u3320_o;
  wire _al_u3321_o;
  wire _al_u3322_o;
  wire _al_u3324_o;
  wire _al_u3327_o;
  wire _al_u3328_o;
  wire _al_u3329_o;
  wire _al_u3330_o;
  wire _al_u3332_o;
  wire _al_u3333_o;
  wire _al_u3334_o;
  wire _al_u3335_o;
  wire _al_u3336_o;
  wire _al_u3337_o;
  wire _al_u3338_o;
  wire _al_u3339_o;
  wire _al_u3340_o;
  wire _al_u3341_o;
  wire _al_u3342_o;
  wire _al_u3343_o;
  wire _al_u3344_o;
  wire _al_u3345_o;
  wire _al_u3346_o;
  wire _al_u3347_o;
  wire _al_u3348_o;
  wire _al_u3349_o;
  wire _al_u3350_o;
  wire _al_u3351_o;
  wire _al_u3352_o;
  wire _al_u3353_o;
  wire _al_u3355_o;
  wire _al_u3356_o;
  wire _al_u3358_o;
  wire _al_u3359_o;
  wire _al_u3360_o;
  wire _al_u3361_o;
  wire _al_u3362_o;
  wire _al_u3363_o;
  wire _al_u3364_o;
  wire _al_u3365_o;
  wire _al_u3366_o;
  wire _al_u3368_o;
  wire _al_u3369_o;
  wire _al_u3371_o;
  wire _al_u3372_o;
  wire _al_u3376_o;
  wire _al_u3377_o;
  wire _al_u3378_o;
  wire _al_u3379_o;
  wire _al_u3380_o;
  wire _al_u3381_o;
  wire _al_u3382_o;
  wire _al_u3383_o;
  wire _al_u3384_o;
  wire _al_u3385_o;
  wire _al_u3386_o;
  wire _al_u3388_o;
  wire _al_u3390_o;
  wire _al_u3391_o;
  wire _al_u3392_o;
  wire _al_u3393_o;
  wire _al_u3395_o;
  wire _al_u3396_o;
  wire _al_u3397_o;
  wire _al_u3398_o;
  wire _al_u3399_o;
  wire _al_u3400_o;
  wire _al_u3402_o;
  wire _al_u3403_o;
  wire _al_u3404_o;
  wire _al_u3405_o;
  wire _al_u3406_o;
  wire _al_u3407_o;
  wire _al_u3408_o;
  wire _al_u3409_o;
  wire _al_u3410_o;
  wire _al_u3411_o;
  wire _al_u3412_o;
  wire _al_u3413_o;
  wire _al_u3414_o;
  wire _al_u3415_o;
  wire _al_u3416_o;
  wire _al_u3417_o;
  wire _al_u3418_o;
  wire _al_u3419_o;
  wire _al_u3420_o;
  wire _al_u3421_o;
  wire _al_u3422_o;
  wire _al_u3424_o;
  wire _al_u3425_o;
  wire _al_u3426_o;
  wire _al_u3427_o;
  wire _al_u3428_o;
  wire _al_u3429_o;
  wire _al_u3430_o;
  wire _al_u3431_o;
  wire _al_u3432_o;
  wire _al_u3433_o;
  wire _al_u3434_o;
  wire _al_u3435_o;
  wire _al_u3436_o;
  wire _al_u3437_o;
  wire _al_u3438_o;
  wire _al_u3439_o;
  wire _al_u3440_o;
  wire _al_u3441_o;
  wire _al_u3442_o;
  wire _al_u3443_o;
  wire _al_u3444_o;
  wire _al_u3445_o;
  wire _al_u3446_o;
  wire _al_u3447_o;
  wire _al_u3448_o;
  wire _al_u3449_o;
  wire _al_u3450_o;
  wire _al_u3451_o;
  wire _al_u3452_o;
  wire _al_u3453_o;
  wire _al_u3454_o;
  wire _al_u3455_o;
  wire _al_u3456_o;
  wire _al_u3457_o;
  wire _al_u3458_o;
  wire _al_u3459_o;
  wire _al_u3462_o;
  wire _al_u3464_o;
  wire _al_u3465_o;
  wire _al_u3466_o;
  wire _al_u3467_o;
  wire _al_u3468_o;
  wire _al_u3469_o;
  wire _al_u3470_o;
  wire _al_u3471_o;
  wire _al_u3472_o;
  wire _al_u3473_o;
  wire _al_u3474_o;
  wire _al_u3475_o;
  wire _al_u3476_o;
  wire _al_u3477_o;
  wire _al_u3480_o;
  wire _al_u3481_o;
  wire _al_u3482_o;
  wire _al_u3484_o;
  wire _al_u3485_o;
  wire _al_u3486_o;
  wire _al_u3487_o;
  wire _al_u3488_o;
  wire _al_u3492_o;
  wire _al_u3495_o;
  wire _al_u3496_o;
  wire _al_u3497_o;
  wire _al_u3498_o;
  wire _al_u3499_o;
  wire _al_u3500_o;
  wire _al_u3501_o;
  wire _al_u3502_o;
  wire _al_u3503_o;
  wire _al_u3504_o;
  wire _al_u3505_o;
  wire _al_u3506_o;
  wire _al_u3507_o;
  wire _al_u3508_o;
  wire _al_u3510_o;
  wire _al_u3511_o;
  wire _al_u3513_o;
  wire _al_u3514_o;
  wire _al_u3515_o;
  wire _al_u3516_o;
  wire _al_u3517_o;
  wire _al_u3518_o;
  wire _al_u3519_o;
  wire _al_u3520_o;
  wire _al_u3521_o;
  wire _al_u3522_o;
  wire _al_u3523_o;
  wire _al_u3524_o;
  wire _al_u3525_o;
  wire _al_u3526_o;
  wire _al_u3527_o;
  wire _al_u3528_o;
  wire _al_u3529_o;
  wire _al_u3531_o;
  wire _al_u3532_o;
  wire _al_u3533_o;
  wire _al_u3534_o;
  wire _al_u3536_o;
  wire _al_u3537_o;
  wire _al_u3538_o;
  wire _al_u3539_o;
  wire _al_u3540_o;
  wire _al_u3541_o;
  wire _al_u3542_o;
  wire _al_u3543_o;
  wire _al_u3544_o;
  wire _al_u3545_o;
  wire _al_u3546_o;
  wire _al_u3547_o;
  wire _al_u3548_o;
  wire _al_u3549_o;
  wire _al_u3550_o;
  wire _al_u3551_o;
  wire _al_u3553_o;
  wire _al_u3554_o;
  wire _al_u3555_o;
  wire _al_u3556_o;
  wire _al_u3557_o;
  wire _al_u3559_o;
  wire _al_u3560_o;
  wire _al_u3563_o;
  wire _al_u3564_o;
  wire _al_u3565_o;
  wire _al_u3566_o;
  wire _al_u3567_o;
  wire _al_u3568_o;
  wire _al_u3569_o;
  wire _al_u3571_o;
  wire _al_u3572_o;
  wire _al_u3573_o;
  wire _al_u3574_o;
  wire _al_u3575_o;
  wire _al_u3576_o;
  wire _al_u3577_o;
  wire _al_u3578_o;
  wire _al_u3579_o;
  wire _al_u3580_o;
  wire _al_u3581_o;
  wire _al_u3582_o;
  wire _al_u3583_o;
  wire _al_u3584_o;
  wire _al_u3585_o;
  wire \add0/c0 ;
  wire \add0/c1 ;
  wire \add0/c2 ;
  wire \add0/c3 ;
  wire \add0/c4 ;
  wire \add0/c5 ;
  wire \add0/c6 ;
  wire \add0/c7 ;
  wire \add0/c8 ;
  wire \add1/c0 ;
  wire \add1/c1 ;
  wire \add1/c2 ;
  wire \add1/c3 ;
  wire \add1/c4 ;
  wire \add1/c5 ;
  wire \add1/c6 ;
  wire \add1/c7 ;
  wire \add2/c0 ;
  wire \add2/c1 ;
  wire \add2/c2 ;
  wire \add2/c3 ;
  wire \add2/c4 ;
  wire \add2/c5 ;
  wire \add2/c6 ;
  wire \add2/c7 ;
  wire bus_write;  // sources/rtl/camera_init.v(44)
  wire mux103_b0_sel_is_2_o;
  wire mux103_b3_sel_is_0_o;
  wire mux104_b11_sel_is_2_o;
  wire mux107_b0_sel_is_2_o;
  wire mux111_b0_sel_is_2_o;
  wire mux115_b2_sel_is_2_o;
  wire mux119_b10_sel_is_2_o;
  wire mux119_b3_sel_is_0_o;
  wire mux119_b4_sel_is_2_o;
  wire mux121_b7_sel_is_2_o;
  wire mux122_b11_sel_is_2_o;
  wire mux123_b10_sel_is_2_o;
  wire mux124_b11_sel_is_2_o;
  wire mux12_b9_sel_is_2_o_neg_lutinv;
  wire mux130_b1_sel_is_2_o;
  wire mux130_b6_sel_is_2_o;
  wire mux132_b0_sel_is_0_o;
  wire mux132_b3_sel_is_2_o;
  wire mux135_b0_sel_is_2_o;
  wire mux135_b11_sel_is_0_o;
  wire mux137_b2_sel_is_2_o;
  wire mux137_b5_sel_is_2_o;
  wire mux139_b0_sel_is_2_o;
  wire mux140_b11_sel_is_2_o;
  wire mux140_b1_sel_is_2_o;
  wire mux140_b5_sel_is_0_o;
  wire mux141_b1_sel_is_2_o;
  wire mux144_b10_sel_is_2_o;
  wire mux144_b7_sel_is_2_o;
  wire mux145_b6_sel_is_2_o;
  wire mux147_b12_sel_is_2_o;
  wire mux148_b3_sel_is_2_o;
  wire mux149_b4_sel_is_2_o;
  wire mux14_b11_sel_is_2_o;
  wire mux153_b3_sel_is_2_o;
  wire mux156_b0_sel_is_2_o;
  wire mux158_b11_sel_is_0_o;
  wire mux159_b1_sel_is_2_o;
  wire mux159_b3_sel_is_2_o;
  wire mux159_b5_sel_is_2_o;
  wire mux15_b15_sel_is_2_o;
  wire mux166_b1_sel_is_2_o;
  wire mux169_b0_sel_is_2_o;
  wire mux16_b0_sel_is_2_o;
  wire mux16_b11_sel_is_2_o;
  wire mux16_b15_sel_is_2_o;
  wire mux16_b1_sel_is_0_o;
  wire mux16_b9_sel_is_2_o_neg_lutinv;
  wire mux170_b2_sel_is_2_o;
  wire mux174_b0_sel_is_0_o;
  wire mux181_b0_sel_is_2_o;
  wire mux19_b2_sel_is_0_o;
  wire mux21_b0_sel_is_0_o;
  wire mux21_b12_sel_is_2_o;
  wire mux24_b10_sel_is_2_o;
  wire mux31_b3_sel_is_2_o;
  wire mux33_b0_sel_is_2_o;
  wire mux37_b6_sel_is_2_o;
  wire mux38_b12_sel_is_2_o;
  wire mux38_b1_sel_is_2_o;
  wire mux42_b0_sel_is_2_o;
  wire mux47_b0_sel_is_2_o;
  wire mux47_b1_sel_is_2_o;
  wire mux49_b0_sel_is_2_o;
  wire mux49_b5_sel_is_0_o;
  wire mux52_b1_sel_is_2_o;
  wire mux5_b5_sel_is_2_o;
  wire mux60_b1_sel_is_2_o;
  wire mux61_b0_sel_is_2_o;
  wire mux63_b12_sel_is_2_o;
  wire mux63_b1_sel_is_2_o;
  wire mux63_b7_sel_is_2_o;
  wire mux67_b0_sel_is_2_o;
  wire mux68_b0_sel_is_2_o;
  wire mux68_b1_sel_is_2_o;
  wire mux68_b4_sel_is_2_o;
  wire mux75_b5_sel_is_2_o;
  wire mux75_b6_sel_is_2_o;
  wire mux83_b0_sel_is_2_o;
  wire mux83_b12_sel_is_2_o;
  wire mux83_b7_sel_is_2_o;
  wire mux84_b4_sel_is_2_o;
  wire mux85_b0_sel_is_2_o;
  wire mux87_b0_sel_is_2_o;
  wire mux94_b0_sel_is_2_o;
  wire mux94_b10_sel_is_0_o;
  wire mux97_b15_sel_is_2_o;
  wire mux97_b2_sel_is_2_o;
  wire n366;
  wire n375_lutinv;
  wire n376_lutinv;
  wire n377_lutinv;
  wire n378_lutinv;
  wire n379_lutinv;
  wire n380;
  wire n382;
  wire ready_out;  // sources/rtl/camera_init.v(45)
  wire sel1_b0_sel_o;  // sources/rtl/camera_init.v(388)
  wire sel1_b1_sel_o;  // sources/rtl/camera_init.v(388)
  wire \sel2_b0/or_or_B4_B5_o_or_B6__o ;
  wire \sel2_b1/or_B6_or_B7_B8_o_o ;
  wire \sel2_b2/or_B6_or_B7_B8_o_o ;
  wire \sel2_b3/or_B6_or_B7_B8_o_o ;
  wire \sel2_b4/or_B6_or_B7_B8_o_o ;
  wire \sel2_b5/or_B6_or_B7_B8_o_o ;
  wire \sel2_b6/or_B6_or_B7_B8_o_o ;
  wire \sel2_b7/or_B6_or_B7_B8_o_o ;
  wire success_out;  // sources/rtl/camera_init.v(46)

  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u2836 (
    .a(state_next[2]),
    .b(n369[6]),
    .c(n369[7]),
    .o(_al_u2836_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*~B*A)"),
    .INIT(16'h0020))
    _al_u2837 (
    .a(_al_u2836_o),
    .b(state_next[3]),
    .c(state_next[4]),
    .d(n369[5]),
    .o(_al_u2837_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u2838 (
    .a(_al_u2837_o),
    .b(state_next[0]),
    .c(state_next[1]),
    .o(n380));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u2839 (
    .a(_al_u2837_o),
    .b(state_next[0]),
    .c(state_next[1]),
    .o(n382));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u2840 (
    .a(counter[2]),
    .b(counter[3]),
    .o(_al_u2840_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*B*A)"),
    .INIT(16'h0800))
    _al_u2841 (
    .a(counter[4]),
    .b(counter[5]),
    .c(counter[6]),
    .d(counter[7]),
    .o(_al_u2841_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u2842 (
    .a(_al_u2840_o),
    .b(_al_u2841_o),
    .c(counter[1]),
    .o(_al_u2842_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2843 (
    .a(_al_u2842_o),
    .b(counter[0]),
    .o(_al_u2843_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2844 (
    .a(_al_u2843_o),
    .b(n372[7]),
    .o(n374[7]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2845 (
    .a(_al_u2843_o),
    .b(n372[6]),
    .o(n374[6]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2846 (
    .a(_al_u2843_o),
    .b(n372[5]),
    .o(n374[5]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2847 (
    .a(_al_u2843_o),
    .b(n372[4]),
    .o(n374[4]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2848 (
    .a(_al_u2843_o),
    .b(n372[3]),
    .o(n374[3]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2849 (
    .a(_al_u2843_o),
    .b(n372[2]),
    .o(n374[2]));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    _al_u2850 (
    .a(_al_u2843_o),
    .b(n372[1]),
    .o(n374[1]));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    _al_u2851 (
    .a(_al_u2843_o),
    .b(n372[0]),
    .o(n374[0]));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u2852 (
    .a(state_next[3]),
    .b(state_next[4]),
    .c(n369[5]),
    .o(_al_u2852_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    _al_u2853 (
    .a(_al_u2852_o),
    .b(state_next[2]),
    .c(n369[6]),
    .d(n369[7]),
    .o(_al_u2853_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u2854 (
    .a(_al_u2853_o),
    .b(state_next[1]),
    .o(sel1_b1_sel_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2855 (
    .a(sel1_b1_sel_o),
    .b(state_next[0]),
    .o(n377_lutinv));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u2856 (
    .a(_al_u2836_o),
    .b(_al_u2852_o),
    .c(state_next[0]),
    .d(state_next[1]),
    .o(n375_lutinv));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    _al_u2857 (
    .a(n377_lutinv),
    .b(n375_lutinv),
    .o(sel1_b0_sel_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u2858 (
    .a(_al_u2853_o),
    .b(state_next[0]),
    .c(state_next[1]),
    .o(n378_lutinv));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~B*~A)"),
    .INIT(8'hfe))
    _al_u2859 (
    .a(sel1_b1_sel_o),
    .b(n378_lutinv),
    .c(n375_lutinv),
    .o(n366));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u2860 (
    .a(n380),
    .b(_al_u2843_o),
    .c(reset_n),
    .o(mux181_b0_sel_is_2_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u2861 (
    .a(_al_u2837_o),
    .b(state_next[1]),
    .o(_al_u2861_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u2862 (
    .a(_al_u2861_o),
    .b(_al_u2853_o),
    .c(n375_lutinv),
    .o(_al_u2862_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u2863 (
    .a(_al_u2853_o),
    .b(state_next[0]),
    .c(state_next[1]),
    .o(n379_lutinv));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u2864 (
    .a(_al_u2862_o),
    .b(n379_lutinv),
    .c(ready_out),
    .o(_al_u2864_o));
  AL_MAP_LUT3 #(
    .EQN("(~(A)*~(B)*~(C)+A*B*~(C)+~(A)*~(B)*C+A*~(B)*C+A*B*C)"),
    .INIT(8'hb9))
    _al_u2865 (
    .a(_al_u2864_o),
    .b(state_next[2]),
    .c(ready_out),
    .o(_al_u2865_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u2866 (
    .a(n380),
    .b(sel1_b1_sel_o),
    .c(n375_lutinv),
    .o(_al_u2866_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*B))"),
    .INIT(8'ha2))
    _al_u2867 (
    .a(_al_u2866_o),
    .b(n379_lutinv),
    .c(success_out),
    .o(_al_u2867_o));
  AL_MAP_LUT2 #(
    .EQN("~(B*A)"),
    .INIT(4'h7))
    _al_u2868 (
    .a(_al_u2865_o),
    .b(_al_u2867_o),
    .o(n369[2]));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u2869 (
    .a(_al_u2843_o),
    .b(n379_lutinv),
    .c(success_out),
    .o(_al_u2869_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u2870 (
    .a(cnt[4]),
    .b(cnt[5]),
    .c(cnt[6]),
    .d(cnt[7]),
    .o(_al_u2870_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*~B*~A)"),
    .INIT(16'h0010))
    _al_u2871 (
    .a(cnt[0]),
    .b(cnt[1]),
    .c(cnt[2]),
    .d(cnt[3]),
    .o(_al_u2871_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2872 (
    .a(_al_u2870_o),
    .b(_al_u2871_o),
    .o(_al_u2872_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(~C*A))"),
    .INIT(16'hf531))
    _al_u2873 (
    .a(_al_u2869_o),
    .b(_al_u2853_o),
    .c(_al_u2872_o),
    .d(state_next[0]),
    .o(_al_u2873_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2874 (
    .a(_al_u2837_o),
    .b(state_next[0]),
    .o(_al_u2874_o));
  AL_MAP_LUT4 #(
    .EQN("~(B*~(D*~(~C*A)))"),
    .INIT(16'hf733))
    _al_u2875 (
    .a(_al_u2864_o),
    .b(_al_u2873_o),
    .c(_al_u2874_o),
    .d(state_next[0]),
    .o(n369[0]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~(~B*A))"),
    .INIT(16'hd000))
    _al_u2876 (
    .a(_al_u2843_o),
    .b(_al_u2872_o),
    .c(ready_out),
    .d(success_out),
    .o(_al_u2876_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u2877 (
    .a(_al_u2876_o),
    .b(n378_lutinv),
    .c(n379_lutinv),
    .o(_al_u2877_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u2878 (
    .a(_al_u2864_o),
    .b(_al_u2874_o),
    .c(ready_out),
    .o(_al_u2878_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    _al_u2879 (
    .a(state_next[3]),
    .b(_al_u2877_o),
    .c(_al_u2878_o),
    .o(n369[3]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C*~A))"),
    .INIT(8'h73))
    _al_u2880 (
    .a(_al_u2878_o),
    .b(_al_u2877_o),
    .c(state_next[4]),
    .o(n369[4]));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u2881 (
    .a(n377_lutinv),
    .b(_al_u2874_o),
    .c(ready_out),
    .o(_al_u2881_o));
  AL_MAP_LUT4 #(
    .EQN("~(~C*B*~(D*~A))"),
    .INIT(16'hf7f3))
    _al_u2882 (
    .a(_al_u2864_o),
    .b(_al_u2881_o),
    .c(_al_u2869_o),
    .d(state_next[1]),
    .o(n369[1]));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u2883 (
    .a(counter[0]),
    .b(counter[1]),
    .o(_al_u2883_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2884 (
    .a(counter[2]),
    .b(counter[3]),
    .o(_al_u2884_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2885 (
    .a(_al_u2883_o),
    .b(_al_u2884_o),
    .o(_al_u2885_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u2886 (
    .a(_al_u2884_o),
    .b(counter[0]),
    .c(counter[1]),
    .o(_al_u2886_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*~B*A)"),
    .INIT(16'h0020))
    _al_u2887 (
    .a(counter[4]),
    .b(counter[5]),
    .c(counter[6]),
    .d(counter[7]),
    .o(_al_u2887_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(~B*~A))"),
    .INIT(8'he0))
    _al_u2888 (
    .a(_al_u2885_o),
    .b(_al_u2886_o),
    .c(_al_u2887_o),
    .o(_al_u2888_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*B*A)"),
    .INIT(16'h0800))
    _al_u2889 (
    .a(counter[0]),
    .b(counter[1]),
    .c(counter[2]),
    .d(counter[3]),
    .o(_al_u2889_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2890 (
    .a(_al_u2889_o),
    .b(_al_u2887_o),
    .o(_al_u2890_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u2891 (
    .a(_al_u2888_o),
    .b(_al_u2890_o),
    .o(mux84_b4_sel_is_2_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2892 (
    .a(counter[2]),
    .b(counter[3]),
    .o(_al_u2892_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u2893 (
    .a(_al_u2892_o),
    .b(counter[0]),
    .c(counter[1]),
    .o(_al_u2893_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u2894 (
    .a(_al_u2884_o),
    .b(counter[0]),
    .c(counter[1]),
    .o(_al_u2894_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D*~(~C*~B)))"),
    .INIT(16'h02aa))
    _al_u2895 (
    .a(mux84_b4_sel_is_2_o),
    .b(_al_u2893_o),
    .c(_al_u2894_o),
    .d(_al_u2887_o),
    .o(mux85_b0_sel_is_2_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2896 (
    .a(_al_u2883_o),
    .b(_al_u2892_o),
    .o(_al_u2896_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u2897 (
    .a(_al_u2892_o),
    .b(counter[0]),
    .c(counter[1]),
    .o(_al_u2897_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(~B*~A))"),
    .INIT(8'he0))
    _al_u2898 (
    .a(_al_u2896_o),
    .b(_al_u2897_o),
    .c(_al_u2887_o),
    .o(_al_u2898_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u2899 (
    .a(mux85_b0_sel_is_2_o),
    .b(_al_u2898_o),
    .o(mux87_b0_sel_is_2_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2900 (
    .a(counter[0]),
    .b(counter[1]),
    .o(_al_u2900_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2901 (
    .a(_al_u2900_o),
    .b(_al_u2884_o),
    .o(_al_u2901_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2902 (
    .a(_al_u2901_o),
    .b(_al_u2887_o),
    .o(_al_u2902_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*B*~A)"),
    .INIT(16'h0400))
    _al_u2903 (
    .a(counter[4]),
    .b(counter[5]),
    .c(counter[6]),
    .d(counter[7]),
    .o(_al_u2903_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u2904 (
    .a(_al_u2843_o),
    .b(_al_u2901_o),
    .c(_al_u2903_o),
    .o(n184[0]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(~B*~A))"),
    .INIT(8'he0))
    _al_u2905 (
    .a(_al_u2893_o),
    .b(_al_u2889_o),
    .c(_al_u2903_o),
    .o(_al_u2905_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u2906 (
    .a(_al_u2905_o),
    .b(_al_u2886_o),
    .c(_al_u2903_o),
    .o(mux5_b5_sel_is_2_o));
  AL_MAP_LUT4 #(
    .EQN("(~((~B*~A))*~(C)*~(D)+(~B*~A)*~(C)*~(D)+(~B*~A)*C*~(D)+~((~B*~A))*~(C)*D+~((~B*~A))*C*D+(~B*~A)*C*D)"),
    .INIT(16'hfe1f))
    _al_u2907 (
    .a(counter[0]),
    .b(counter[1]),
    .c(counter[2]),
    .d(counter[3]),
    .o(_al_u2907_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u2908 (
    .a(_al_u2903_o),
    .b(_al_u2907_o),
    .o(_al_u2908_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u2909 (
    .a(n184[0]),
    .b(mux5_b5_sel_is_2_o),
    .c(_al_u2908_o),
    .o(_al_u2909_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2910 (
    .a(_al_u2840_o),
    .b(_al_u2900_o),
    .o(_al_u2910_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u2911 (
    .a(counter[2]),
    .b(counter[3]),
    .o(_al_u2911_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2912 (
    .a(_al_u2911_o),
    .b(_al_u2883_o),
    .o(_al_u2912_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u2913 (
    .a(_al_u2910_o),
    .b(_al_u2912_o),
    .o(_al_u2913_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*(D@C))"),
    .INIT(16'h0880))
    _al_u2914 (
    .a(_al_u2840_o),
    .b(_al_u2903_o),
    .c(counter[0]),
    .d(counter[1]),
    .o(_al_u2914_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*~A))"),
    .INIT(8'h23))
    _al_u2915 (
    .a(_al_u2913_o),
    .b(_al_u2914_o),
    .c(_al_u2903_o),
    .o(mux14_b11_sel_is_2_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2916 (
    .a(_al_u2909_o),
    .b(mux14_b11_sel_is_2_o),
    .o(n196[6]));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*A)"),
    .INIT(16'h0200))
    _al_u2917 (
    .a(counter[4]),
    .b(counter[5]),
    .c(counter[6]),
    .d(counter[7]),
    .o(_al_u2917_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2918 (
    .a(_al_u2893_o),
    .b(_al_u2917_o),
    .o(_al_u2918_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2919 (
    .a(_al_u2889_o),
    .b(_al_u2917_o),
    .o(_al_u2919_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u2920 (
    .a(_al_u2918_o),
    .b(_al_u2919_o),
    .o(mux21_b0_sel_is_0_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2921 (
    .a(_al_u2885_o),
    .b(_al_u2917_o),
    .o(_al_u2921_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u2922 (
    .a(mux21_b0_sel_is_0_o),
    .b(_al_u2921_o),
    .o(_al_u2922_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*A))"),
    .INIT(8'hc4))
    _al_u2923 (
    .a(n196[6]),
    .b(_al_u2922_o),
    .c(_al_u2917_o),
    .o(_al_u2923_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2924 (
    .a(_al_u2911_o),
    .b(_al_u2917_o),
    .o(_al_u2924_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u2925 (
    .a(_al_u2840_o),
    .b(_al_u2917_o),
    .c(counter[1]),
    .o(_al_u2925_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*A*~(D*B))"),
    .INIT(16'h020a))
    _al_u2926 (
    .a(_al_u2923_o),
    .b(_al_u2924_o),
    .c(_al_u2925_o),
    .d(counter[1]),
    .o(_al_u2926_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*~A)"),
    .INIT(16'h0100))
    _al_u2927 (
    .a(counter[4]),
    .b(counter[5]),
    .c(counter[6]),
    .d(counter[7]),
    .o(_al_u2927_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2928 (
    .a(_al_u2894_o),
    .b(_al_u2927_o),
    .o(_al_u2928_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2929 (
    .a(_al_u2901_o),
    .b(_al_u2927_o),
    .o(_al_u2929_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u2930 (
    .a(_al_u2928_o),
    .b(_al_u2929_o),
    .o(_al_u2930_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u2931 (
    .a(_al_u2840_o),
    .b(counter[1]),
    .o(_al_u2931_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2932 (
    .a(_al_u2931_o),
    .b(_al_u2917_o),
    .o(_al_u2932_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(A*~(D)*~(C)+A*D*~(C)+~(A)*D*C+A*D*C))"),
    .INIT(16'h04c4))
    _al_u2933 (
    .a(_al_u2926_o),
    .b(_al_u2930_o),
    .c(_al_u2932_o),
    .d(counter[0]),
    .o(n215[6]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(~B*~A))"),
    .INIT(8'he0))
    _al_u2934 (
    .a(_al_u2893_o),
    .b(_al_u2889_o),
    .c(_al_u2927_o),
    .o(_al_u2934_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2935 (
    .a(_al_u2885_o),
    .b(_al_u2927_o),
    .o(_al_u2935_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u2936 (
    .a(_al_u2934_o),
    .b(_al_u2935_o),
    .o(mux37_b6_sel_is_2_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2937 (
    .a(n215[6]),
    .b(mux37_b6_sel_is_2_o),
    .o(n219[6]));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u2938 (
    .a(_al_u2840_o),
    .b(counter[0]),
    .c(counter[1]),
    .o(_al_u2938_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2939 (
    .a(_al_u2938_o),
    .b(_al_u2927_o),
    .o(_al_u2939_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2940 (
    .a(_al_u2931_o),
    .b(_al_u2927_o),
    .o(_al_u2940_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u2941 (
    .a(_al_u2939_o),
    .b(_al_u2940_o),
    .o(mux47_b1_sel_is_2_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(~B*~A))"),
    .INIT(8'he0))
    _al_u2942 (
    .a(_al_u2896_o),
    .b(_al_u2911_o),
    .c(_al_u2927_o),
    .o(_al_u2942_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*A*~(D*C))"),
    .INIT(16'h0222))
    _al_u2943 (
    .a(mux47_b1_sel_is_2_o),
    .b(_al_u2942_o),
    .c(_al_u2910_o),
    .d(_al_u2927_o),
    .o(mux47_b0_sel_is_2_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*A)"),
    .INIT(16'h0080))
    _al_u2944 (
    .a(counter[4]),
    .b(counter[5]),
    .c(counter[6]),
    .d(counter[7]),
    .o(_al_u2944_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2945 (
    .a(_al_u2894_o),
    .b(_al_u2944_o),
    .o(_al_u2945_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2946 (
    .a(_al_u2901_o),
    .b(_al_u2944_o),
    .o(_al_u2946_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u2947 (
    .a(_al_u2945_o),
    .b(_al_u2946_o),
    .o(mux49_b5_sel_is_0_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2948 (
    .a(mux47_b0_sel_is_2_o),
    .b(mux49_b5_sel_is_0_o),
    .o(mux49_b0_sel_is_2_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(~B*~A))"),
    .INIT(8'he0))
    _al_u2949 (
    .a(_al_u2885_o),
    .b(_al_u2886_o),
    .c(_al_u2944_o),
    .o(_al_u2949_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2950 (
    .a(_al_u2889_o),
    .b(_al_u2944_o),
    .o(_al_u2950_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u2951 (
    .a(_al_u2949_o),
    .b(_al_u2950_o),
    .o(mux52_b1_sel_is_2_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2952 (
    .a(mux49_b0_sel_is_2_o),
    .b(mux52_b1_sel_is_2_o),
    .o(_al_u2952_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u2953 (
    .a(_al_u2952_o),
    .b(_al_u2944_o),
    .o(mux63_b12_sel_is_2_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2954 (
    .a(n219[6]),
    .b(mux63_b12_sel_is_2_o),
    .o(n244[6]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2955 (
    .a(_al_u2911_o),
    .b(counter[1]),
    .o(_al_u2955_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2956 (
    .a(_al_u2955_o),
    .b(counter[0]),
    .o(_al_u2956_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u2957 (
    .a(_al_u2956_o),
    .b(_al_u2896_o),
    .o(_al_u2957_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*~A)"),
    .INIT(16'h0040))
    _al_u2958 (
    .a(counter[4]),
    .b(counter[5]),
    .c(counter[6]),
    .d(counter[7]),
    .o(_al_u2958_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2959 (
    .a(_al_u2957_o),
    .b(_al_u2958_o),
    .o(_al_u2959_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u2960 (
    .a(_al_u2955_o),
    .b(_al_u2958_o),
    .c(counter[0]),
    .o(_al_u2960_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u2961 (
    .a(_al_u2911_o),
    .b(counter[1]),
    .o(_al_u2961_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2962 (
    .a(_al_u2961_o),
    .b(_al_u2958_o),
    .o(_al_u2962_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u2963 (
    .a(_al_u2960_o),
    .b(_al_u2962_o),
    .o(mux75_b5_sel_is_2_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2964 (
    .a(_al_u2959_o),
    .b(mux75_b5_sel_is_2_o),
    .o(mux75_b6_sel_is_2_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(~B*~A))"),
    .INIT(8'he0))
    _al_u2965 (
    .a(_al_u2886_o),
    .b(_al_u2894_o),
    .c(_al_u2958_o),
    .o(_al_u2965_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u2966 (
    .a(_al_u2965_o),
    .b(_al_u2885_o),
    .c(_al_u2958_o),
    .o(mux67_b0_sel_is_2_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u2967 (
    .a(n244[6]),
    .b(mux75_b6_sel_is_2_o),
    .c(mux67_b0_sel_is_2_o),
    .o(_al_u2967_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u2968 (
    .a(mux87_b0_sel_is_2_o),
    .b(_al_u2902_o),
    .c(_al_u2967_o),
    .o(_al_u2968_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*~B*~A)"),
    .INIT(16'h0010))
    _al_u2969 (
    .a(counter[4]),
    .b(counter[5]),
    .c(counter[6]),
    .d(counter[7]),
    .o(_al_u2969_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2970 (
    .a(_al_u2894_o),
    .b(_al_u2969_o),
    .o(_al_u2970_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2971 (
    .a(_al_u2901_o),
    .b(_al_u2969_o),
    .o(_al_u2971_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u2972 (
    .a(_al_u2931_o),
    .b(_al_u2887_o),
    .c(counter[0]),
    .o(_al_u2972_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u2973 (
    .a(_al_u2970_o),
    .b(_al_u2971_o),
    .c(_al_u2972_o),
    .o(_al_u2973_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u2974 (
    .a(_al_u2911_o),
    .b(counter[0]),
    .c(counter[1]),
    .o(_al_u2974_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(~C*~B*A))"),
    .INIT(16'hfd00))
    _al_u2975 (
    .a(_al_u2913_o),
    .b(_al_u2974_o),
    .c(_al_u2938_o),
    .d(_al_u2887_o),
    .o(_al_u2975_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2976 (
    .a(_al_u2885_o),
    .b(_al_u2969_o),
    .o(_al_u2976_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2977 (
    .a(_al_u2886_o),
    .b(_al_u2969_o),
    .o(_al_u2977_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u2978 (
    .a(_al_u2976_o),
    .b(_al_u2977_o),
    .o(_al_u2978_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u2979 (
    .a(_al_u2931_o),
    .b(_al_u2887_o),
    .c(counter[0]),
    .o(_al_u2979_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*~B*A)"),
    .INIT(16'h0020))
    _al_u2980 (
    .a(_al_u2973_o),
    .b(_al_u2975_o),
    .c(_al_u2978_o),
    .d(_al_u2979_o),
    .o(_al_u2980_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(B*A))"),
    .INIT(8'h07))
    _al_u2981 (
    .a(_al_u2968_o),
    .b(_al_u2980_o),
    .c(_al_u2976_o),
    .o(_al_u2981_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u2982 (
    .a(_al_u2897_o),
    .b(_al_u2893_o),
    .o(_al_u2982_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(~B*A))"),
    .INIT(8'hd0))
    _al_u2983 (
    .a(_al_u2982_o),
    .b(_al_u2889_o),
    .c(_al_u2969_o),
    .o(_al_u2983_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2984 (
    .a(_al_u2896_o),
    .b(_al_u2969_o),
    .o(_al_u2984_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u2985 (
    .a(_al_u2983_o),
    .b(_al_u2984_o),
    .o(mux103_b0_sel_is_2_o));
  AL_MAP_LUT3 #(
    .EQN("(A*(C@B))"),
    .INIT(8'h28))
    _al_u2986 (
    .a(_al_u2911_o),
    .b(counter[0]),
    .c(counter[1]),
    .o(_al_u2986_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2987 (
    .a(_al_u2986_o),
    .b(_al_u2969_o),
    .o(_al_u2987_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*~A)"),
    .INIT(8'h04))
    _al_u2988 (
    .a(_al_u2981_o),
    .b(mux103_b0_sel_is_2_o),
    .c(_al_u2987_o),
    .o(_al_u2988_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2989 (
    .a(_al_u2931_o),
    .b(_al_u2969_o),
    .o(_al_u2989_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2990 (
    .a(_al_u2938_o),
    .b(_al_u2969_o),
    .o(_al_u2990_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u2991 (
    .a(_al_u2989_o),
    .b(_al_u2990_o),
    .o(mux111_b0_sel_is_2_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    _al_u2992 (
    .a(counter[4]),
    .b(counter[5]),
    .c(counter[6]),
    .d(counter[7]),
    .o(_al_u2992_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2993 (
    .a(_al_u2901_o),
    .b(_al_u2992_o),
    .o(_al_u2993_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u2994 (
    .a(mux111_b0_sel_is_2_o),
    .b(_al_u2993_o),
    .o(_al_u2994_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2995 (
    .a(_al_u2886_o),
    .b(_al_u2992_o),
    .o(_al_u2995_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2996 (
    .a(_al_u2894_o),
    .b(_al_u2992_o),
    .o(_al_u2996_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u2997 (
    .a(_al_u2995_o),
    .b(_al_u2996_o),
    .o(_al_u2997_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2998 (
    .a(_al_u2885_o),
    .b(_al_u2992_o),
    .o(_al_u2998_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u2999 (
    .a(_al_u2997_o),
    .b(_al_u2998_o),
    .o(_al_u2999_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3000 (
    .a(_al_u2994_o),
    .b(_al_u2999_o),
    .o(mux115_b2_sel_is_2_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3001 (
    .a(_al_u2998_o),
    .b(_al_u2995_o),
    .o(_al_u3001_o));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    _al_u3002 (
    .a(_al_u2988_o),
    .b(mux115_b2_sel_is_2_o),
    .c(_al_u3001_o),
    .o(_al_u3002_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u3003 (
    .a(_al_u3002_o),
    .b(_al_u2889_o),
    .c(_al_u2992_o),
    .o(_al_u3003_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3004 (
    .a(_al_u2897_o),
    .b(_al_u2992_o),
    .o(_al_u3004_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3005 (
    .a(_al_u3003_o),
    .b(_al_u3004_o),
    .o(_al_u3005_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3006 (
    .a(_al_u2955_o),
    .b(_al_u2992_o),
    .o(_al_u3006_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3007 (
    .a(_al_u2974_o),
    .b(_al_u2992_o),
    .o(_al_u3007_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3008 (
    .a(_al_u3006_o),
    .b(_al_u3007_o),
    .o(mux122_b11_sel_is_2_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*~B))"),
    .INIT(8'ha8))
    _al_u3009 (
    .a(_al_u3005_o),
    .b(mux122_b11_sel_is_2_o),
    .c(_al_u2986_o),
    .o(_al_u3009_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*~A)"),
    .INIT(16'h0004))
    _al_u3010 (
    .a(counter[4]),
    .b(counter[5]),
    .c(counter[6]),
    .d(counter[7]),
    .o(_al_u3010_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3011 (
    .a(_al_u2886_o),
    .b(_al_u3010_o),
    .o(_al_u3011_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(~B*~A))"),
    .INIT(8'he0))
    _al_u3012 (
    .a(_al_u2894_o),
    .b(_al_u2901_o),
    .c(_al_u3010_o),
    .o(_al_u3012_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3013 (
    .a(_al_u3011_o),
    .b(_al_u3012_o),
    .o(_al_u3013_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3014 (
    .a(_al_u2912_o),
    .b(_al_u2992_o),
    .o(_al_u3014_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3015 (
    .a(_al_u2840_o),
    .b(_al_u2992_o),
    .o(_al_u3015_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u3016 (
    .a(_al_u3013_o),
    .b(_al_u3014_o),
    .c(_al_u3015_o),
    .o(mux130_b6_sel_is_2_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3017 (
    .a(_al_u2885_o),
    .b(_al_u3010_o),
    .o(_al_u3017_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3018 (
    .a(_al_u3009_o),
    .b(mux130_b6_sel_is_2_o),
    .c(_al_u3017_o),
    .o(_al_u3018_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u3019 (
    .a(_al_u2982_o),
    .b(_al_u2955_o),
    .c(_al_u2896_o),
    .o(_al_u3019_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D*~(~C*B)))"),
    .INIT(16'h08aa))
    _al_u3020 (
    .a(_al_u3018_o),
    .b(_al_u3019_o),
    .c(_al_u2961_o),
    .d(_al_u3010_o),
    .o(_al_u3020_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3021 (
    .a(_al_u2931_o),
    .b(_al_u3010_o),
    .o(_al_u3021_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*A)"),
    .INIT(16'h0002))
    _al_u3022 (
    .a(counter[4]),
    .b(counter[5]),
    .c(counter[6]),
    .d(counter[7]),
    .o(_al_u3022_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u3023 (
    .a(_al_u3021_o),
    .b(_al_u2901_o),
    .c(_al_u3022_o),
    .o(mux144_b7_sel_is_2_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3024 (
    .a(_al_u2840_o),
    .b(_al_u3010_o),
    .c(counter[1]),
    .o(_al_u3024_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3025 (
    .a(mux144_b7_sel_is_2_o),
    .b(_al_u3024_o),
    .o(mux144_b10_sel_is_2_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u3026 (
    .a(mux144_b10_sel_is_2_o),
    .b(_al_u2894_o),
    .c(_al_u3022_o),
    .o(mux145_b6_sel_is_2_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3027 (
    .a(_al_u2912_o),
    .b(_al_u3010_o),
    .o(_al_u3027_o));
  AL_MAP_LUT3 #(
    .EQN("(~(A)*~(B)*~(C)+A*B*~(C)+~(A)*~(B)*C+~(A)*B*C+A*B*C)"),
    .INIT(8'hd9))
    _al_u3028 (
    .a(_al_u3020_o),
    .b(mux145_b6_sel_is_2_o),
    .c(_al_u3027_o),
    .o(_al_u3028_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u3029 (
    .a(_al_u3028_o),
    .b(_al_u2885_o),
    .c(_al_u3022_o),
    .o(_al_u3029_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*~B))"),
    .INIT(8'h8a))
    _al_u3030 (
    .a(_al_u3029_o),
    .b(_al_u2982_o),
    .c(_al_u3022_o),
    .o(_al_u3030_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3031 (
    .a(_al_u2955_o),
    .b(_al_u3022_o),
    .o(_al_u3031_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    _al_u3032 (
    .a(_al_u3030_o),
    .b(_al_u3031_o),
    .c(counter[0]),
    .o(_al_u3032_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3033 (
    .a(_al_u2931_o),
    .b(_al_u3022_o),
    .c(counter[0]),
    .o(_al_u3033_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3034 (
    .a(_al_u2938_o),
    .b(_al_u3022_o),
    .o(_al_u3034_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3035 (
    .a(_al_u3033_o),
    .b(_al_u3034_o),
    .o(mux158_b11_sel_is_0_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3036 (
    .a(_al_u2931_o),
    .b(_al_u3022_o),
    .c(counter[0]),
    .o(_al_u3036_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3037 (
    .a(mux158_b11_sel_is_0_o),
    .b(_al_u3036_o),
    .o(mux159_b1_sel_is_2_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3038 (
    .a(_al_u2910_o),
    .b(_al_u3022_o),
    .o(_al_u3038_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3039 (
    .a(mux159_b1_sel_is_2_o),
    .b(_al_u3038_o),
    .o(mux159_b3_sel_is_2_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3040 (
    .a(_al_u2974_o),
    .b(_al_u3022_o),
    .o(_al_u3040_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*~A)"),
    .INIT(8'h04))
    _al_u3041 (
    .a(_al_u3032_o),
    .b(mux159_b3_sel_is_2_o),
    .c(_al_u3040_o),
    .o(_al_u3041_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u3042 (
    .a(counter[4]),
    .b(counter[5]),
    .c(counter[6]),
    .d(counter[7]),
    .o(_al_u3042_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3043 (
    .a(_al_u2894_o),
    .b(_al_u3042_o),
    .o(_al_u3043_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3044 (
    .a(_al_u3041_o),
    .b(_al_u3043_o),
    .o(_al_u3044_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3045 (
    .a(_al_u2955_o),
    .b(_al_u3042_o),
    .o(_al_u3045_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(~B*~A))"),
    .INIT(8'he0))
    _al_u3046 (
    .a(_al_u2896_o),
    .b(_al_u2897_o),
    .c(_al_u3042_o),
    .o(_al_u3046_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3047 (
    .a(_al_u3045_o),
    .b(_al_u3046_o),
    .o(mux169_b0_sel_is_2_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3048 (
    .a(_al_u2974_o),
    .b(_al_u3042_o),
    .o(_al_u3048_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3049 (
    .a(mux169_b0_sel_is_2_o),
    .b(_al_u3048_o),
    .o(mux170_b2_sel_is_2_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3050 (
    .a(_al_u2885_o),
    .b(_al_u3042_o),
    .o(_al_u3050_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3051 (
    .a(_al_u3044_o),
    .b(mux170_b2_sel_is_2_o),
    .c(_al_u3050_o),
    .o(_al_u3051_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(~B*~A))"),
    .INIT(8'he0))
    _al_u3052 (
    .a(_al_u2956_o),
    .b(_al_u2986_o),
    .c(_al_u2903_o),
    .o(_al_u3052_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3053 (
    .a(_al_u2931_o),
    .b(_al_u2903_o),
    .o(_al_u3053_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u3054 (
    .a(mux14_b11_sel_is_2_o),
    .b(_al_u3052_o),
    .c(_al_u3053_o),
    .o(mux15_b15_sel_is_2_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3055 (
    .a(_al_u2901_o),
    .b(_al_u2917_o),
    .o(_al_u3055_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3056 (
    .a(mux15_b15_sel_is_2_o),
    .b(_al_u3055_o),
    .o(mux16_b15_sel_is_2_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3057 (
    .a(_al_u2892_o),
    .b(_al_u2903_o),
    .o(_al_u3057_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(~D*~C))"),
    .INIT(16'h8880))
    _al_u3058 (
    .a(_al_u2884_o),
    .b(_al_u2903_o),
    .c(counter[0]),
    .d(counter[1]),
    .o(_al_u3058_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~B*~(~D*A))"),
    .INIT(16'h0301))
    _al_u3059 (
    .a(_al_u2842_o),
    .b(_al_u3057_o),
    .c(_al_u3058_o),
    .d(counter[0]),
    .o(_al_u3059_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3060 (
    .a(mux16_b15_sel_is_2_o),
    .b(_al_u2922_o),
    .c(_al_u3059_o),
    .o(_al_u3060_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3061 (
    .a(_al_u3060_o),
    .b(_al_u2929_o),
    .o(_al_u3061_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3062 (
    .a(_al_u2886_o),
    .b(_al_u2927_o),
    .o(_al_u3062_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3063 (
    .a(_al_u3062_o),
    .b(_al_u2935_o),
    .o(_al_u3063_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3064 (
    .a(_al_u2897_o),
    .b(_al_u2927_o),
    .o(_al_u3064_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3065 (
    .a(_al_u3061_o),
    .b(_al_u3063_o),
    .c(_al_u3064_o),
    .o(_al_u3065_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u3066 (
    .a(_al_u2913_o),
    .b(_al_u2887_o),
    .c(_al_u2907_o),
    .o(_al_u3066_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u3067 (
    .a(_al_u2982_o),
    .b(_al_u2887_o),
    .o(_al_u3067_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u3068 (
    .a(_al_u3066_o),
    .b(_al_u3067_o),
    .c(_al_u2890_o),
    .o(_al_u3068_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3069 (
    .a(_al_u2938_o),
    .b(_al_u2887_o),
    .o(_al_u3069_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3070 (
    .a(_al_u3069_o),
    .b(_al_u2979_o),
    .o(mux94_b10_sel_is_0_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3071 (
    .a(_al_u2973_o),
    .b(mux94_b10_sel_is_0_o),
    .o(mux97_b15_sel_is_2_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3072 (
    .a(_al_u3065_o),
    .b(_al_u3068_o),
    .c(mux97_b15_sel_is_2_o),
    .o(_al_u3072_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3073 (
    .a(_al_u3072_o),
    .b(_al_u2983_o),
    .o(_al_u3073_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u3074 (
    .a(_al_u2913_o),
    .b(_al_u2969_o),
    .o(_al_u3074_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3075 (
    .a(_al_u3074_o),
    .b(_al_u2990_o),
    .o(_al_u3075_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3076 (
    .a(_al_u2955_o),
    .b(_al_u2969_o),
    .o(_al_u3076_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3077 (
    .a(_al_u2974_o),
    .b(_al_u2969_o),
    .o(_al_u3077_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3078 (
    .a(_al_u3076_o),
    .b(_al_u3077_o),
    .o(_al_u3078_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3079 (
    .a(_al_u3073_o),
    .b(_al_u3075_o),
    .c(_al_u3078_o),
    .o(_al_u3079_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3080 (
    .a(_al_u2993_o),
    .b(_al_u2996_o),
    .o(_al_u3080_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3081 (
    .a(_al_u3080_o),
    .b(_al_u2995_o),
    .o(_al_u3081_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*B))"),
    .INIT(8'ha2))
    _al_u3082 (
    .a(_al_u3081_o),
    .b(_al_u2989_o),
    .c(counter[0]),
    .o(_al_u3082_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3083 (
    .a(_al_u2961_o),
    .b(_al_u2992_o),
    .o(_al_u3083_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3084 (
    .a(_al_u3083_o),
    .b(_al_u3015_o),
    .o(_al_u3084_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3085 (
    .a(_al_u3079_o),
    .b(_al_u3082_o),
    .c(_al_u3084_o),
    .o(_al_u3085_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3086 (
    .a(_al_u2889_o),
    .b(_al_u3010_o),
    .o(_al_u3086_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3087 (
    .a(_al_u3017_o),
    .b(_al_u3086_o),
    .o(mux132_b0_sel_is_0_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3088 (
    .a(_al_u3085_o),
    .b(mux132_b0_sel_is_0_o),
    .c(_al_u3011_o),
    .o(_al_u3088_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3089 (
    .a(_al_u2955_o),
    .b(_al_u3010_o),
    .o(_al_u3089_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3090 (
    .a(_al_u3089_o),
    .b(counter[0]),
    .o(_al_u3090_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3091 (
    .a(_al_u2897_o),
    .b(_al_u3010_o),
    .o(_al_u3091_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3092 (
    .a(_al_u2896_o),
    .b(_al_u3010_o),
    .o(_al_u3092_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3093 (
    .a(_al_u3091_o),
    .b(_al_u3092_o),
    .o(mux135_b11_sel_is_0_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u3094 (
    .a(_al_u3088_o),
    .b(_al_u3090_o),
    .c(mux135_b11_sel_is_0_o),
    .o(_al_u3094_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(~B*~A))"),
    .INIT(8'he0))
    _al_u3095 (
    .a(_al_u2894_o),
    .b(_al_u2901_o),
    .c(_al_u3022_o),
    .o(_al_u3095_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(~B*~A))"),
    .INIT(8'he0))
    _al_u3096 (
    .a(_al_u2931_o),
    .b(_al_u2938_o),
    .c(_al_u3010_o),
    .o(_al_u3096_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u3097 (
    .a(_al_u3094_o),
    .b(_al_u3095_o),
    .c(_al_u3096_o),
    .o(_al_u3097_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    _al_u3098 (
    .a(_al_u3048_o),
    .b(_al_u3033_o),
    .c(_al_u3097_o),
    .o(_al_u3098_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3099 (
    .a(_al_u2938_o),
    .b(_al_u3042_o),
    .o(_al_u3099_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3100 (
    .a(_al_u3098_o),
    .b(_al_u3099_o),
    .o(_al_u3100_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3101 (
    .a(sel1_b1_sel_o),
    .b(state_next[0]),
    .o(n376_lutinv));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3102 (
    .a(_al_u2931_o),
    .b(_al_u3042_o),
    .c(counter[0]),
    .o(_al_u3102_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(B*~(~C*A)))"),
    .INIT(16'h003b))
    _al_u3103 (
    .a(_al_u3100_o),
    .b(n376_lutinv),
    .c(_al_u3102_o),
    .d(n375_lutinv),
    .o(_al_u3103_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3104 (
    .a(_al_u2931_o),
    .b(_al_u3042_o),
    .c(counter[0]),
    .o(_al_u3104_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3105 (
    .a(_al_u3104_o),
    .b(_al_u3099_o),
    .o(mux174_b0_sel_is_0_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3106 (
    .a(mux174_b0_sel_is_0_o),
    .b(_al_u3102_o),
    .o(_al_u3106_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3107 (
    .a(_al_u3106_o),
    .b(n377_lutinv),
    .o(_al_u3107_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C*A))"),
    .INIT(8'hb3))
    _al_u3108 (
    .a(_al_u3051_o),
    .b(_al_u3103_o),
    .c(_al_u3107_o),
    .o(\sel2_b6/or_B6_or_B7_B8_o_o ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*B))"),
    .INIT(8'ha2))
    _al_u3109 (
    .a(n184[0]),
    .b(_al_u2903_o),
    .c(counter[2]),
    .o(_al_u3109_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3110 (
    .a(_al_u2897_o),
    .b(_al_u2903_o),
    .o(_al_u3110_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3111 (
    .a(_al_u3109_o),
    .b(_al_u3110_o),
    .o(_al_u3111_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*~A)"),
    .INIT(8'h04))
    _al_u3112 (
    .a(_al_u3111_o),
    .b(mux14_b11_sel_is_2_o),
    .c(_al_u2908_o),
    .o(_al_u3112_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u3113 (
    .a(_al_u3055_o),
    .b(_al_u3053_o),
    .c(counter[0]),
    .o(mux16_b1_sel_is_0_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    _al_u3114 (
    .a(_al_u3112_o),
    .b(mux16_b1_sel_is_0_o),
    .c(_al_u3053_o),
    .o(n198[2]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3115 (
    .a(_al_u2886_o),
    .b(_al_u2917_o),
    .o(_al_u3115_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3116 (
    .a(_al_u2921_o),
    .b(_al_u3115_o),
    .o(mux19_b2_sel_is_0_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3117 (
    .a(n198[2]),
    .b(mux19_b2_sel_is_0_o),
    .o(n212[2]));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u3118 (
    .a(_al_u3063_o),
    .b(_al_u3064_o),
    .c(_al_u2934_o),
    .o(mux38_b12_sel_is_2_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3119 (
    .a(mux38_b12_sel_is_2_o),
    .b(_al_u2930_o),
    .o(mux38_b1_sel_is_2_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(~D*~(B*A)))"),
    .INIT(16'h0f08))
    _al_u3120 (
    .a(n212[2]),
    .b(mux38_b1_sel_is_2_o),
    .c(_al_u2942_o),
    .d(_al_u3064_o),
    .o(n225[2]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3121 (
    .a(n225[2]),
    .b(mux47_b1_sel_is_2_o),
    .o(_al_u3121_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u3122 (
    .a(_al_u3121_o),
    .b(_al_u2940_o),
    .c(counter[0]),
    .o(_al_u3122_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3123 (
    .a(_al_u2913_o),
    .b(_al_u2982_o),
    .c(_al_u2907_o),
    .o(_al_u3123_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*~B))"),
    .INIT(8'h8a))
    _al_u3124 (
    .a(mux52_b1_sel_is_2_o),
    .b(_al_u3123_o),
    .c(_al_u2944_o),
    .o(mux60_b1_sel_is_2_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3125 (
    .a(mux60_b1_sel_is_2_o),
    .b(_al_u2945_o),
    .o(_al_u3125_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*~B))"),
    .INIT(8'h54))
    _al_u3126 (
    .a(_al_u3122_o),
    .b(_al_u3125_o),
    .c(_al_u2910_o),
    .o(n240[2]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u3127 (
    .a(n240[2]),
    .b(_al_u2938_o),
    .c(_al_u2944_o),
    .o(_al_u3127_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u3128 (
    .a(_al_u3127_o),
    .b(_al_u2901_o),
    .c(_al_u2958_o),
    .o(_al_u3128_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(~B*~A))"),
    .INIT(8'he0))
    _al_u3129 (
    .a(_al_u2885_o),
    .b(_al_u2889_o),
    .c(_al_u2958_o),
    .o(_al_u3129_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u3130 (
    .a(_al_u3129_o),
    .b(_al_u2886_o),
    .c(_al_u2958_o),
    .o(mux68_b1_sel_is_2_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3131 (
    .a(_al_u3128_o),
    .b(mux68_b1_sel_is_2_o),
    .o(_al_u3131_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u3132 (
    .a(_al_u3131_o),
    .b(_al_u2956_o),
    .c(_al_u2958_o),
    .o(_al_u3132_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u3133 (
    .a(_al_u3132_o),
    .b(_al_u2912_o),
    .c(_al_u2958_o),
    .o(_al_u3133_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(~B*~A))"),
    .INIT(8'he0))
    _al_u3134 (
    .a(_al_u2886_o),
    .b(_al_u2894_o),
    .c(_al_u2887_o),
    .o(_al_u3134_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3135 (
    .a(_al_u2840_o),
    .b(_al_u2958_o),
    .c(counter[1]),
    .o(_al_u3135_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u3136 (
    .a(_al_u2902_o),
    .b(_al_u3134_o),
    .c(_al_u3135_o),
    .o(_al_u3136_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*~B))"),
    .INIT(8'ha8))
    _al_u3137 (
    .a(_al_u3133_o),
    .b(_al_u3136_o),
    .c(_al_u2886_o),
    .o(_al_u3137_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*~B))"),
    .INIT(8'h8a))
    _al_u3138 (
    .a(mux94_b10_sel_is_0_o),
    .b(_al_u2913_o),
    .c(_al_u2887_o),
    .o(mux94_b0_sel_is_2_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u3139 (
    .a(_al_u3019_o),
    .b(_al_u2887_o),
    .o(_al_u3139_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3140 (
    .a(_al_u2974_o),
    .b(_al_u2887_o),
    .o(_al_u3140_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*~B*A)"),
    .INIT(16'h0020))
    _al_u3141 (
    .a(mux94_b0_sel_is_2_o),
    .b(_al_u3139_o),
    .c(_al_u2973_o),
    .d(_al_u3140_o),
    .o(mux97_b2_sel_is_2_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3142 (
    .a(_al_u2885_o),
    .b(_al_u2887_o),
    .o(_al_u3142_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3143 (
    .a(_al_u3137_o),
    .b(mux97_b2_sel_is_2_o),
    .c(_al_u3142_o),
    .o(_al_u3143_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3144 (
    .a(_al_u3143_o),
    .b(mux103_b0_sel_is_2_o),
    .o(_al_u3144_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3145 (
    .a(_al_u2896_o),
    .b(_al_u2992_o),
    .o(_al_u3145_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3146 (
    .a(_al_u3145_o),
    .b(_al_u3004_o),
    .o(mux119_b3_sel_is_0_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(~B*~A))"),
    .INIT(8'he0))
    _al_u3147 (
    .a(_al_u2893_o),
    .b(_al_u2889_o),
    .c(_al_u2992_o),
    .o(_al_u3147_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3148 (
    .a(mux119_b3_sel_is_0_o),
    .b(_al_u3147_o),
    .o(mux119_b10_sel_is_2_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3149 (
    .a(mux119_b10_sel_is_2_o),
    .b(_al_u3006_o),
    .o(mux121_b7_sel_is_2_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3150 (
    .a(mux115_b2_sel_is_2_o),
    .b(mux121_b7_sel_is_2_o),
    .c(_al_u3083_o),
    .o(_al_u3150_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3151 (
    .a(_al_u2912_o),
    .b(_al_u2969_o),
    .o(_al_u3151_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3152 (
    .a(_al_u3144_o),
    .b(_al_u3150_o),
    .c(_al_u3151_o),
    .o(_al_u3152_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~B*~(~C*~A))"),
    .INIT(16'h0032))
    _al_u3153 (
    .a(_al_u3152_o),
    .b(_al_u3012_o),
    .c(_al_u3014_o),
    .d(_al_u3015_o),
    .o(_al_u3153_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3154 (
    .a(_al_u3153_o),
    .b(mux132_b0_sel_is_0_o),
    .o(_al_u3154_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3155 (
    .a(_al_u2910_o),
    .b(_al_u3010_o),
    .o(_al_u3155_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3156 (
    .a(_al_u3027_o),
    .b(_al_u3155_o),
    .o(mux140_b5_sel_is_0_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3157 (
    .a(_al_u2974_o),
    .b(_al_u3010_o),
    .o(_al_u3157_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3158 (
    .a(mux140_b5_sel_is_0_o),
    .b(_al_u3157_o),
    .o(mux140_b1_sel_is_2_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3159 (
    .a(mux135_b11_sel_is_0_o),
    .b(_al_u3089_o),
    .o(mux137_b2_sel_is_2_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3160 (
    .a(_al_u2886_o),
    .b(_al_u3022_o),
    .o(_al_u3160_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(~B*~A))"),
    .INIT(8'he0))
    _al_u3161 (
    .a(_al_u2885_o),
    .b(_al_u2889_o),
    .c(_al_u3022_o),
    .o(_al_u3161_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u3162 (
    .a(_al_u3160_o),
    .b(_al_u3095_o),
    .c(_al_u3096_o),
    .d(_al_u3161_o),
    .o(mux148_b3_sel_is_2_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u3163 (
    .a(_al_u3154_o),
    .b(mux140_b1_sel_is_2_o),
    .c(mux137_b2_sel_is_2_o),
    .d(mux148_b3_sel_is_2_o),
    .o(_al_u3163_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3164 (
    .a(_al_u2901_o),
    .b(_al_u3042_o),
    .o(_al_u3164_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3165 (
    .a(_al_u3043_o),
    .b(_al_u3164_o),
    .o(_al_u3165_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3166 (
    .a(_al_u2886_o),
    .b(_al_u3042_o),
    .o(_al_u3166_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3167 (
    .a(_al_u3165_o),
    .b(_al_u3166_o),
    .o(_al_u3167_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3168 (
    .a(mux159_b1_sel_is_2_o),
    .b(_al_u3167_o),
    .o(_al_u3168_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3169 (
    .a(_al_u2885_o),
    .b(_al_u3022_o),
    .o(_al_u3169_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~C*~(~D*A)))"),
    .INIT(16'hc0c8))
    _al_u3170 (
    .a(_al_u3163_o),
    .b(_al_u3168_o),
    .c(_al_u3169_o),
    .d(_al_u3022_o),
    .o(_al_u3170_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u3171 (
    .a(_al_u3170_o),
    .b(_al_u3042_o),
    .c(_al_u2889_o),
    .o(_al_u3171_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3172 (
    .a(_al_u3171_o),
    .b(mux170_b2_sel_is_2_o),
    .o(_al_u3172_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(B*A))"),
    .INIT(8'h07))
    _al_u3173 (
    .a(_al_u2886_o),
    .b(_al_u2903_o),
    .c(_al_u2842_o),
    .o(_al_u3173_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3174 (
    .a(_al_u2893_o),
    .b(_al_u2903_o),
    .o(_al_u3174_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3175 (
    .a(_al_u2955_o),
    .b(_al_u2903_o),
    .o(_al_u3175_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u3176 (
    .a(_al_u3173_o),
    .b(_al_u3174_o),
    .c(_al_u3175_o),
    .o(_al_u3176_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B)*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hc8aa))
    _al_u3177 (
    .a(_al_u3176_o),
    .b(_al_u2913_o),
    .c(_al_u2986_o),
    .d(_al_u2903_o),
    .o(_al_u3177_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D*C*~B))"),
    .INIT(16'h8aaa))
    _al_u3178 (
    .a(mux21_b0_sel_is_0_o),
    .b(_al_u2900_o),
    .c(_al_u2884_o),
    .d(_al_u2917_o),
    .o(mux21_b12_sel_is_2_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3179 (
    .a(_al_u3177_o),
    .b(mux21_b12_sel_is_2_o),
    .o(_al_u3179_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(B*~A))"),
    .INIT(8'h0b))
    _al_u3180 (
    .a(_al_u3179_o),
    .b(_al_u2922_o),
    .c(_al_u2918_o),
    .o(_al_u3180_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u3181 (
    .a(_al_u2957_o),
    .b(_al_u2917_o),
    .o(_al_u3181_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3182 (
    .a(_al_u2897_o),
    .b(_al_u2917_o),
    .o(_al_u3182_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3183 (
    .a(_al_u3181_o),
    .b(_al_u3182_o),
    .o(mux24_b10_sel_is_2_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(A*~(D)*~(C)+A*D*~(C)+~(A)*D*C+A*D*C))"),
    .INIT(16'h04c4))
    _al_u3184 (
    .a(_al_u3180_o),
    .b(mux24_b10_sel_is_2_o),
    .c(_al_u2924_o),
    .d(_al_u2883_o),
    .o(_al_u3184_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3185 (
    .a(_al_u2938_o),
    .b(_al_u2917_o),
    .o(_al_u3185_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3186 (
    .a(_al_u3184_o),
    .b(_al_u3185_o),
    .o(_al_u3186_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*B))"),
    .INIT(8'ha2))
    _al_u3187 (
    .a(_al_u2930_o),
    .b(_al_u2932_o),
    .c(counter[0]),
    .o(mux33_b0_sel_is_2_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3188 (
    .a(_al_u3186_o),
    .b(mux33_b0_sel_is_2_o),
    .o(_al_u3188_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*~B))"),
    .INIT(8'h8a))
    _al_u3189 (
    .a(_al_u3188_o),
    .b(_al_u2889_o),
    .c(_al_u2927_o),
    .o(_al_u3189_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    _al_u3190 (
    .a(_al_u3189_o),
    .b(_al_u2952_o),
    .c(_al_u3064_o),
    .o(_al_u3190_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3191 (
    .a(_al_u3190_o),
    .b(_al_u3068_o),
    .o(_al_u3191_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3192 (
    .a(_al_u3191_o),
    .b(_al_u2970_o),
    .o(_al_u3192_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3193 (
    .a(_al_u3076_o),
    .b(counter[0]),
    .o(_al_u3193_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3194 (
    .a(_al_u2889_o),
    .b(_al_u2969_o),
    .o(_al_u3194_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3195 (
    .a(_al_u2976_o),
    .b(_al_u3194_o),
    .o(_al_u3195_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u3196 (
    .a(_al_u3192_o),
    .b(_al_u3193_o),
    .c(_al_u3195_o),
    .o(_al_u3196_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u3197 (
    .a(_al_u3196_o),
    .b(_al_u2840_o),
    .c(_al_u2969_o),
    .o(_al_u3197_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3198 (
    .a(_al_u3197_o),
    .b(_al_u3001_o),
    .o(_al_u3198_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    _al_u3199 (
    .a(_al_u3198_o),
    .b(_al_u3006_o),
    .c(counter[0]),
    .o(_al_u3199_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u3200 (
    .a(_al_u2840_o),
    .b(_al_u2992_o),
    .c(counter[0]),
    .d(counter[1]),
    .o(_al_u3200_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u3201 (
    .a(_al_u3199_o),
    .b(_al_u3011_o),
    .c(_al_u3200_o),
    .o(_al_u3201_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u3202 (
    .a(_al_u2982_o),
    .b(_al_u3010_o),
    .o(_al_u3202_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3203 (
    .a(_al_u3201_o),
    .b(_al_u3202_o),
    .o(_al_u3203_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u3204 (
    .a(_al_u3203_o),
    .b(_al_u2911_o),
    .c(_al_u3010_o),
    .o(_al_u3204_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(~B*A))"),
    .INIT(8'hd0))
    _al_u3205 (
    .a(_al_u2982_o),
    .b(_al_u2896_o),
    .c(_al_u3022_o),
    .o(_al_u3205_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(~B*~A))"),
    .INIT(8'he0))
    _al_u3206 (
    .a(_al_u2886_o),
    .b(_al_u2894_o),
    .c(_al_u3022_o),
    .o(_al_u3206_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u3207 (
    .a(_al_u3205_o),
    .b(_al_u3206_o),
    .c(_al_u3161_o),
    .o(_al_u3207_o));
  AL_MAP_LUT4 #(
    .EQN("~((B*A)*~(D)*~(C)+(B*A)*D*~(C)+~((B*A))*D*C+(B*A)*D*C)"),
    .INIT(16'h07f7))
    _al_u3208 (
    .a(_al_u3204_o),
    .b(_al_u3207_o),
    .c(_al_u3031_o),
    .d(counter[0]),
    .o(_al_u3208_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3209 (
    .a(_al_u2912_o),
    .b(_al_u3022_o),
    .o(_al_u3209_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3210 (
    .a(_al_u3208_o),
    .b(_al_u3209_o),
    .o(_al_u3210_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3211 (
    .a(_al_u3210_o),
    .b(_al_u3034_o),
    .o(_al_u3211_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    _al_u3212 (
    .a(_al_u2885_o),
    .b(_al_u3042_o),
    .c(_al_u2889_o),
    .o(_al_u3212_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u3213 (
    .a(_al_u3211_o),
    .b(_al_u3036_o),
    .c(_al_u3212_o),
    .o(_al_u3213_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3214 (
    .a(_al_u2897_o),
    .b(_al_u3042_o),
    .o(_al_u3214_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3215 (
    .a(_al_u3213_o),
    .b(_al_u3214_o),
    .o(_al_u3215_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(~C*~B*A))"),
    .INIT(16'hfd00))
    _al_u3216 (
    .a(_al_u2913_o),
    .b(_al_u2938_o),
    .c(_al_u2986_o),
    .d(_al_u3042_o),
    .o(_al_u3216_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u3217 (
    .a(_al_u3215_o),
    .b(_al_u3216_o),
    .c(_al_u3102_o),
    .o(_al_u3217_o));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*~B)*~(C*A))"),
    .INIT(16'hb3a0))
    _al_u3218 (
    .a(_al_u3172_o),
    .b(_al_u3217_o),
    .c(_al_u3107_o),
    .d(n376_lutinv),
    .o(\sel2_b2/or_B6_or_B7_B8_o_o ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3219 (
    .a(_al_u2896_o),
    .b(_al_u2903_o),
    .o(_al_u3219_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3220 (
    .a(_al_u3110_o),
    .b(_al_u3219_o),
    .o(_al_u3220_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*~(D*~C)))"),
    .INIT(16'h2a22))
    _al_u3221 (
    .a(mux15_b15_sel_is_2_o),
    .b(_al_u3220_o),
    .c(_al_u2843_o),
    .d(_al_u3059_o),
    .o(_al_u3221_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*~A))"),
    .INIT(8'h8c))
    _al_u3222 (
    .a(_al_u2911_o),
    .b(_al_u2917_o),
    .c(_al_u2907_o),
    .o(_al_u3222_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~C)*~(~B*~A))"),
    .INIT(16'he0ee))
    _al_u3223 (
    .a(_al_u3221_o),
    .b(_al_u3053_o),
    .c(_al_u3222_o),
    .d(_al_u2917_o),
    .o(_al_u3223_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    _al_u3224 (
    .a(_al_u3223_o),
    .b(mux33_b0_sel_is_2_o),
    .c(_al_u2932_o),
    .o(_al_u3224_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(B*~(~D*~A)))"),
    .INIT(16'h0307))
    _al_u3225 (
    .a(_al_u3224_o),
    .b(mux38_b12_sel_is_2_o),
    .c(_al_u3064_o),
    .d(_al_u2928_o),
    .o(_al_u3225_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3226 (
    .a(_al_u2974_o),
    .b(_al_u2927_o),
    .o(_al_u3226_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(~B*~A))"),
    .INIT(8'he0))
    _al_u3227 (
    .a(_al_u2955_o),
    .b(_al_u2896_o),
    .c(_al_u2927_o),
    .o(_al_u3227_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3228 (
    .a(_al_u3226_o),
    .b(_al_u3227_o),
    .o(mux42_b0_sel_is_2_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*~B))"),
    .INIT(8'h54))
    _al_u3229 (
    .a(_al_u3225_o),
    .b(mux42_b0_sel_is_2_o),
    .c(_al_u2986_o),
    .o(n223[7]));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D*~(~C*~B)))"),
    .INIT(16'h02aa))
    _al_u3230 (
    .a(mux60_b1_sel_is_2_o),
    .b(_al_u2931_o),
    .c(_al_u2938_o),
    .d(_al_u2944_o),
    .o(mux63_b1_sel_is_2_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u3231 (
    .a(_al_u2913_o),
    .b(_al_u2927_o),
    .o(_al_u3231_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*A)"),
    .INIT(16'h0080))
    _al_u3232 (
    .a(mux63_b1_sel_is_2_o),
    .b(mux49_b5_sel_is_0_o),
    .c(mux47_b1_sel_is_2_o),
    .d(_al_u3231_o),
    .o(mux63_b7_sel_is_2_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3233 (
    .a(n223[7]),
    .b(mux63_b7_sel_is_2_o),
    .c(mux67_b0_sel_is_2_o),
    .o(n256[7]));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3234 (
    .a(_al_u3142_o),
    .b(_al_u3134_o),
    .o(mux83_b0_sel_is_2_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3235 (
    .a(_al_u3135_o),
    .b(counter[0]),
    .o(_al_u3235_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3236 (
    .a(_al_u2840_o),
    .b(_al_u2958_o),
    .c(counter[1]),
    .o(_al_u3236_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3237 (
    .a(_al_u3235_o),
    .b(_al_u3236_o),
    .o(_al_u3237_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3238 (
    .a(_al_u3135_o),
    .b(counter[0]),
    .o(_al_u3238_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    _al_u3239 (
    .a(mux83_b0_sel_is_2_o),
    .b(_al_u3237_o),
    .c(_al_u2902_o),
    .d(_al_u3238_o),
    .o(mux83_b7_sel_is_2_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*~A)"),
    .INIT(16'h0004))
    _al_u3240 (
    .a(_al_u3139_o),
    .b(mux83_b7_sel_is_2_o),
    .c(_al_u2975_o),
    .d(_al_u2890_o),
    .o(_al_u3240_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3241 (
    .a(n256[7]),
    .b(_al_u3240_o),
    .o(_al_u3241_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(~B*~A))"),
    .INIT(8'h0e))
    _al_u3242 (
    .a(_al_u3241_o),
    .b(_al_u3069_o),
    .c(_al_u2979_o),
    .o(_al_u3242_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*~B))"),
    .INIT(8'h8a))
    _al_u3243 (
    .a(_al_u3242_o),
    .b(_al_u2883_o),
    .c(_al_u2969_o),
    .o(_al_u3243_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3244 (
    .a(_al_u3193_o),
    .b(_al_u2984_o),
    .o(_al_u3244_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u3245 (
    .a(_al_u3243_o),
    .b(_al_u3244_o),
    .o(_al_u3245_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u3246 (
    .a(_al_u3245_o),
    .b(_al_u2994_o),
    .o(_al_u3246_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3247 (
    .a(_al_u3246_o),
    .b(mux121_b7_sel_is_2_o),
    .o(_al_u3247_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3248 (
    .a(_al_u2931_o),
    .b(_al_u2992_o),
    .c(counter[0]),
    .o(_al_u3248_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*~B))"),
    .INIT(8'h8a))
    _al_u3249 (
    .a(_al_u3247_o),
    .b(_al_u3248_o),
    .c(_al_u3015_o),
    .o(_al_u3249_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    _al_u3250 (
    .a(_al_u3249_o),
    .b(_al_u2894_o),
    .c(_al_u3010_o),
    .o(_al_u3250_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3251 (
    .a(_al_u3250_o),
    .b(_al_u3017_o),
    .o(_al_u3251_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3252 (
    .a(_al_u3089_o),
    .b(counter[0]),
    .o(_al_u3252_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u3253 (
    .a(_al_u3251_o),
    .b(_al_u3252_o),
    .c(_al_u3024_o),
    .o(_al_u3253_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*~A)"),
    .INIT(8'h04))
    _al_u3254 (
    .a(_al_u3253_o),
    .b(mux144_b7_sel_is_2_o),
    .c(_al_u3206_o),
    .o(_al_u3254_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u3255 (
    .a(_al_u3254_o),
    .b(_al_u2897_o),
    .c(_al_u3022_o),
    .o(_al_u3255_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3256 (
    .a(_al_u2961_o),
    .b(_al_u3022_o),
    .o(_al_u3256_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(~A*~(D)*~(B)+~A*D*~(B)+~(~A)*D*B+~A*D*B))"),
    .INIT(16'h020e))
    _al_u3257 (
    .a(_al_u3255_o),
    .b(_al_u3031_o),
    .c(_al_u3256_o),
    .d(counter[0]),
    .o(_al_u3257_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3258 (
    .a(_al_u3038_o),
    .b(_al_u3209_o),
    .o(_al_u3258_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*~A))"),
    .INIT(8'h8c))
    _al_u3259 (
    .a(_al_u3257_o),
    .b(mux159_b1_sel_is_2_o),
    .c(_al_u3258_o),
    .o(_al_u3259_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3260 (
    .a(_al_u3166_o),
    .b(_al_u3212_o),
    .o(_al_u3260_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3261 (
    .a(_al_u3259_o),
    .b(_al_u3260_o),
    .c(_al_u3043_o),
    .o(_al_u3261_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3262 (
    .a(_al_u3261_o),
    .b(mux170_b2_sel_is_2_o),
    .c(_al_u3099_o),
    .o(_al_u3262_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3263 (
    .a(_al_u3262_o),
    .b(n377_lutinv),
    .c(_al_u3102_o),
    .o(_al_u3263_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf131))
    _al_u3264 (
    .a(_al_u2932_o),
    .b(_al_u2924_o),
    .c(counter[0]),
    .d(counter[1]),
    .o(_al_u3264_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3265 (
    .a(_al_u2932_o),
    .b(counter[0]),
    .o(_al_u3265_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    _al_u3266 (
    .a(mux24_b10_sel_is_2_o),
    .b(_al_u3264_o),
    .c(_al_u3265_o),
    .d(_al_u2925_o),
    .o(_al_u3266_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u3267 (
    .a(mux68_b1_sel_is_2_o),
    .b(_al_u2894_o),
    .c(_al_u2958_o),
    .o(mux68_b0_sel_is_2_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3268 (
    .a(_al_u2901_o),
    .b(_al_u2958_o),
    .o(_al_u3268_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u3269 (
    .a(_al_u3268_o),
    .b(_al_u2931_o),
    .c(_al_u2944_o),
    .o(_al_u3269_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3270 (
    .a(mux68_b0_sel_is_2_o),
    .b(_al_u3269_o),
    .o(_al_u3270_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3271 (
    .a(_al_u3266_o),
    .b(mux38_b1_sel_is_2_o),
    .c(_al_u3270_o),
    .o(_al_u3271_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3272 (
    .a(mux83_b0_sel_is_2_o),
    .b(_al_u2958_o),
    .o(_al_u3272_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*(B@A))"),
    .INIT(8'h06))
    _al_u3273 (
    .a(counter[1]),
    .b(counter[2]),
    .c(counter[3]),
    .o(_al_u3273_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*A))"),
    .INIT(8'hc4))
    _al_u3274 (
    .a(_al_u3019_o),
    .b(_al_u2944_o),
    .c(_al_u3273_o),
    .o(_al_u3274_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*B*A)"),
    .INIT(16'h0800))
    _al_u3275 (
    .a(_al_u2952_o),
    .b(_al_u3272_o),
    .c(_al_u3274_o),
    .d(mux21_b12_sel_is_2_o),
    .o(_al_u3275_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*C*D+A*B*C*D)"),
    .INIT(16'ha1b1))
    _al_u3276 (
    .a(_al_u2842_o),
    .b(_al_u3058_o),
    .c(counter[0]),
    .d(_al_u3057_o),
    .o(_al_u3276_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3277 (
    .a(_al_u3220_o),
    .b(_al_u3276_o),
    .o(_al_u3277_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*A)"),
    .INIT(16'h0080))
    _al_u3278 (
    .a(_al_u3271_o),
    .b(_al_u3275_o),
    .c(_al_u3277_o),
    .d(_al_u2902_o),
    .o(_al_u3278_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3279 (
    .a(_al_u3278_o),
    .b(mux97_b15_sel_is_2_o),
    .c(_al_u2978_o),
    .o(_al_u3279_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*B))"),
    .INIT(8'ha2))
    _al_u3280 (
    .a(_al_u3279_o),
    .b(_al_u3076_o),
    .c(counter[0]),
    .o(_al_u3280_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3281 (
    .a(_al_u3280_o),
    .b(_al_u3075_o),
    .o(_al_u3281_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u3282 (
    .a(_al_u3281_o),
    .b(_al_u3048_o),
    .c(_al_u3099_o),
    .o(_al_u3282_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3283 (
    .a(_al_u3282_o),
    .b(_al_u3102_o),
    .o(_al_u3283_o));
  AL_MAP_LUT3 #(
    .EQN("~(~A*~(C*~B))"),
    .INIT(8'hba))
    _al_u3284 (
    .a(_al_u3263_o),
    .b(_al_u3283_o),
    .c(n376_lutinv),
    .o(\sel2_b7/or_B6_or_B7_B8_o_o ));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(D*~(~C*~B)))"),
    .INIT(16'h0155))
    _al_u3285 (
    .a(_al_u2843_o),
    .b(_al_u2894_o),
    .c(_al_u2901_o),
    .d(_al_u2903_o),
    .o(n185[3]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3286 (
    .a(n185[3]),
    .b(_al_u3174_o),
    .o(n187[3]));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u3287 (
    .a(mux14_b11_sel_is_2_o),
    .b(_al_u3055_o),
    .c(_al_u3053_o),
    .o(mux16_b11_sel_is_2_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3288 (
    .a(_al_u2974_o),
    .b(_al_u2903_o),
    .o(_al_u3288_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3289 (
    .a(mux16_b11_sel_is_2_o),
    .b(_al_u3288_o),
    .o(mux16_b0_sel_is_2_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3290 (
    .a(_al_u2955_o),
    .b(_al_u2903_o),
    .c(counter[0]),
    .o(_al_u3290_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(~B*~A))"),
    .INIT(8'he0))
    _al_u3291 (
    .a(_al_u2955_o),
    .b(_al_u2896_o),
    .c(_al_u2903_o),
    .o(_al_u3291_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~C*~(~D*A)))"),
    .INIT(16'hc0c8))
    _al_u3292 (
    .a(n187[3]),
    .b(mux16_b0_sel_is_2_o),
    .c(_al_u3290_o),
    .d(_al_u3291_o),
    .o(_al_u3292_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3293 (
    .a(_al_u3053_o),
    .b(counter[0]),
    .o(_al_u3293_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(~B*~A))"),
    .INIT(8'h0e))
    _al_u3294 (
    .a(_al_u3292_o),
    .b(_al_u3293_o),
    .c(_al_u3115_o),
    .o(n200[3]));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u3295 (
    .a(n200[3]),
    .b(_al_u3181_o),
    .c(_al_u2919_o),
    .o(n206[3]));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3296 (
    .a(_al_u2924_o),
    .b(counter[0]),
    .c(counter[1]),
    .o(_al_u3296_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3297 (
    .a(n206[3]),
    .b(_al_u3296_o),
    .o(n207[3]));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3298 (
    .a(_al_u2932_o),
    .b(_al_u3185_o),
    .o(mux31_b3_sel_is_2_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3299 (
    .a(mux38_b1_sel_is_2_o),
    .b(mux31_b3_sel_is_2_o),
    .o(_al_u3299_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(~C*~(B*A)))"),
    .INIT(16'h00f8))
    _al_u3300 (
    .a(n207[3]),
    .b(_al_u3299_o),
    .c(_al_u3064_o),
    .d(_al_u3227_o),
    .o(_al_u3300_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3301 (
    .a(_al_u3300_o),
    .b(_al_u3231_o),
    .o(_al_u3301_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u3302 (
    .a(_al_u3301_o),
    .b(_al_u2945_o),
    .c(_al_u2940_o),
    .o(_al_u3302_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3303 (
    .a(_al_u2889_o),
    .b(_al_u2958_o),
    .o(_al_u3303_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(D*~(~C*~B)))"),
    .INIT(16'h0155))
    _al_u3304 (
    .a(_al_u3274_o),
    .b(_al_u2885_o),
    .c(_al_u2889_o),
    .d(_al_u2944_o),
    .o(mux61_b0_sel_is_2_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3305 (
    .a(_al_u3270_o),
    .b(mux61_b0_sel_is_2_o),
    .o(mux68_b4_sel_is_2_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(A*~(~D*~C)))"),
    .INIT(16'h1113))
    _al_u3306 (
    .a(_al_u3302_o),
    .b(_al_u2949_o),
    .c(_al_u3303_o),
    .d(mux68_b4_sel_is_2_o),
    .o(_al_u3306_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u3307 (
    .a(_al_u2982_o),
    .b(_al_u2958_o),
    .o(_al_u3307_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(~B*~A))"),
    .INIT(8'he0))
    _al_u3308 (
    .a(_al_u2956_o),
    .b(_al_u2986_o),
    .c(_al_u2958_o),
    .o(_al_u3308_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u3309 (
    .a(_al_u3306_o),
    .b(_al_u3307_o),
    .c(_al_u3308_o),
    .o(_al_u3309_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3310 (
    .a(_al_u2938_o),
    .b(_al_u2958_o),
    .o(_al_u3310_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*~A))"),
    .INIT(8'h32))
    _al_u3311 (
    .a(_al_u3309_o),
    .b(_al_u3310_o),
    .c(_al_u2962_o),
    .o(_al_u3311_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u3312 (
    .a(_al_u3311_o),
    .b(_al_u2902_o),
    .c(_al_u3142_o),
    .o(_al_u3312_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3313 (
    .a(_al_u3312_o),
    .b(_al_u3067_o),
    .o(_al_u3313_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3314 (
    .a(_al_u3313_o),
    .b(_al_u2973_o),
    .c(_al_u2975_o),
    .o(_al_u3314_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3315 (
    .a(_al_u3314_o),
    .b(_al_u3195_o),
    .o(_al_u3315_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3316 (
    .a(_al_u2987_o),
    .b(_al_u3151_o),
    .o(mux107_b0_sel_is_2_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3317 (
    .a(_al_u2897_o),
    .b(_al_u2969_o),
    .o(_al_u3317_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3318 (
    .a(_al_u2984_o),
    .b(_al_u3317_o),
    .o(mux103_b3_sel_is_0_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3319 (
    .a(_al_u3315_o),
    .b(mux107_b0_sel_is_2_o),
    .c(mux103_b3_sel_is_0_o),
    .o(_al_u3319_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3320 (
    .a(_al_u3319_o),
    .b(_al_u2990_o),
    .o(_al_u3320_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(C*~(B*A)))"),
    .INIT(16'h008f))
    _al_u3321 (
    .a(_al_u3320_o),
    .b(_al_u3082_o),
    .c(_al_u2997_o),
    .d(_al_u2998_o),
    .o(_al_u3321_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u3322 (
    .a(_al_u3013_o),
    .b(_al_u2931_o),
    .c(_al_u2992_o),
    .o(_al_u3322_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u3323 (
    .a(_al_u3322_o),
    .b(_al_u2938_o),
    .c(_al_u2992_o),
    .o(mux130_b1_sel_is_2_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3324 (
    .a(_al_u2910_o),
    .b(_al_u2992_o),
    .o(_al_u3324_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u3325 (
    .a(mux122_b11_sel_is_2_o),
    .b(_al_u3324_o),
    .c(_al_u3014_o),
    .o(mux124_b11_sel_is_2_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u3326 (
    .a(mux130_b1_sel_is_2_o),
    .b(mux124_b11_sel_is_2_o),
    .c(mux119_b3_sel_is_0_o),
    .d(mux132_b0_sel_is_0_o),
    .o(mux132_b3_sel_is_2_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3327 (
    .a(_al_u3321_o),
    .b(mux132_b3_sel_is_2_o),
    .o(_al_u3327_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3328 (
    .a(_al_u3327_o),
    .b(mux137_b2_sel_is_2_o),
    .c(_al_u3027_o),
    .o(_al_u3328_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3329 (
    .a(_al_u3328_o),
    .b(mux148_b3_sel_is_2_o),
    .o(_al_u3329_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u3330 (
    .a(_al_u2957_o),
    .b(_al_u3022_o),
    .o(_al_u3330_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3331 (
    .a(_al_u3330_o),
    .b(_al_u3031_o),
    .o(mux153_b3_sel_is_2_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3332 (
    .a(_al_u3329_o),
    .b(mux159_b3_sel_is_2_o),
    .c(mux153_b3_sel_is_2_o),
    .o(_al_u3332_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3333 (
    .a(_al_u3332_o),
    .b(_al_u3043_o),
    .o(_al_u3333_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3334 (
    .a(_al_u2893_o),
    .b(_al_u3042_o),
    .o(_al_u3334_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D*~C*A))"),
    .INIT(16'h3133))
    _al_u3335 (
    .a(_al_u3333_o),
    .b(_al_u3214_o),
    .c(_al_u3334_o),
    .d(mux170_b2_sel_is_2_o),
    .o(_al_u3335_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u3336 (
    .a(_al_u2905_o),
    .b(_al_u2842_o),
    .c(counter[0]),
    .o(_al_u3336_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3337 (
    .a(_al_u3336_o),
    .b(_al_u3052_o),
    .o(_al_u3337_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3338 (
    .a(_al_u3337_o),
    .b(_al_u3115_o),
    .o(_al_u3338_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B*A))"),
    .INIT(8'h70))
    _al_u3339 (
    .a(_al_u2910_o),
    .b(_al_u2917_o),
    .c(_al_u3338_o),
    .o(_al_u3339_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*A))"),
    .INIT(8'hc4))
    _al_u3340 (
    .a(_al_u3339_o),
    .b(mux33_b0_sel_is_2_o),
    .c(_al_u2932_o),
    .o(_al_u3340_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~A*~(D*C))"),
    .INIT(16'h0111))
    _al_u3341 (
    .a(_al_u3340_o),
    .b(_al_u2928_o),
    .c(_al_u2889_o),
    .d(_al_u2927_o),
    .o(_al_u3341_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3342 (
    .a(_al_u3341_o),
    .b(_al_u3068_o),
    .c(mux94_b10_sel_is_0_o),
    .o(_al_u3342_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3343 (
    .a(_al_u3342_o),
    .b(_al_u2971_o),
    .o(_al_u3343_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u3344 (
    .a(_al_u3343_o),
    .b(_al_u2977_o),
    .c(_al_u3194_o),
    .o(_al_u3344_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3345 (
    .a(_al_u3344_o),
    .b(_al_u3151_o),
    .o(_al_u3345_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3346 (
    .a(_al_u3345_o),
    .b(_al_u2994_o),
    .o(_al_u3346_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3347 (
    .a(_al_u2893_o),
    .b(_al_u2992_o),
    .o(_al_u3347_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3348 (
    .a(mux119_b3_sel_is_0_o),
    .b(_al_u3347_o),
    .o(_al_u3348_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3349 (
    .a(_al_u3346_o),
    .b(_al_u3348_o),
    .c(_al_u2995_o),
    .o(_al_u3349_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3350 (
    .a(_al_u3349_o),
    .b(_al_u3200_o),
    .o(_al_u3350_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*~B))"),
    .INIT(8'h8a))
    _al_u3351 (
    .a(_al_u3350_o),
    .b(_al_u2894_o),
    .c(_al_u3010_o),
    .o(_al_u3351_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u3352 (
    .a(_al_u3351_o),
    .b(mux132_b0_sel_is_0_o),
    .o(_al_u3352_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3353 (
    .a(_al_u3352_o),
    .b(mux135_b11_sel_is_0_o),
    .o(_al_u3353_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3354 (
    .a(mux140_b1_sel_is_2_o),
    .b(_al_u3252_o),
    .o(mux140_b11_sel_is_2_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3355 (
    .a(_al_u3353_o),
    .b(mux140_b11_sel_is_2_o),
    .o(_al_u3355_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3356 (
    .a(_al_u3169_o),
    .b(_al_u3160_o),
    .o(_al_u3356_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3357 (
    .a(_al_u3356_o),
    .b(_al_u3095_o),
    .o(mux147_b12_sel_is_2_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3358 (
    .a(_al_u3021_o),
    .b(counter[0]),
    .o(_al_u3358_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3359 (
    .a(mux147_b12_sel_is_2_o),
    .b(_al_u3358_o),
    .o(_al_u3359_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*A))"),
    .INIT(8'hc4))
    _al_u3360 (
    .a(_al_u3355_o),
    .b(_al_u3359_o),
    .c(_al_u3021_o),
    .o(_al_u3360_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3361 (
    .a(_al_u3360_o),
    .b(_al_u3038_o),
    .o(_al_u3361_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3362 (
    .a(_al_u3361_o),
    .b(_al_u3165_o),
    .c(_al_u3036_o),
    .o(_al_u3362_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3363 (
    .a(_al_u3362_o),
    .b(_al_u3050_o),
    .o(_al_u3363_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u3364 (
    .a(_al_u3363_o),
    .b(_al_u2896_o),
    .c(_al_u3042_o),
    .o(_al_u3364_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3365 (
    .a(_al_u3364_o),
    .b(_al_u3216_o),
    .o(_al_u3365_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*A))"),
    .INIT(8'hc4))
    _al_u3366 (
    .a(_al_u3365_o),
    .b(n376_lutinv),
    .c(_al_u3102_o),
    .o(_al_u3366_o));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*~A))"),
    .INIT(8'hdc))
    _al_u3367 (
    .a(_al_u3335_o),
    .b(_al_u3366_o),
    .c(_al_u3107_o),
    .o(\sel2_b3/or_B6_or_B7_B8_o_o ));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3368 (
    .a(_al_u2931_o),
    .b(_al_u2927_o),
    .c(counter[0]),
    .o(_al_u3368_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(~D*~B*A))"),
    .INIT(16'h0f0d))
    _al_u3369 (
    .a(n185[3]),
    .b(_al_u3052_o),
    .c(_al_u3288_o),
    .d(_al_u3057_o),
    .o(_al_u3369_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(~D*~(B*~A)))"),
    .INIT(16'hf040))
    _al_u3370 (
    .a(_al_u3369_o),
    .b(mux14_b11_sel_is_2_o),
    .c(mux16_b1_sel_is_0_o),
    .d(_al_u3053_o),
    .o(n198[4]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3371 (
    .a(mux21_b0_sel_is_0_o),
    .b(mux19_b2_sel_is_0_o),
    .o(_al_u3371_o));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'h47))
    _al_u3372 (
    .a(n198[4]),
    .b(_al_u3371_o),
    .c(_al_u2918_o),
    .o(_al_u3372_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3373 (
    .a(_al_u3372_o),
    .b(_al_u3182_o),
    .o(n204[4]));
  AL_MAP_LUT4 #(
    .EQN("(A*~((D@C))*~(B)+A*(D@C)*~(B)+~(A)*(D@C)*B+A*(D@C)*B)"),
    .INIT(16'h2ee2))
    _al_u3374 (
    .a(n204[4]),
    .b(_al_u2924_o),
    .c(counter[0]),
    .d(counter[1]),
    .o(n209[4]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3375 (
    .a(n209[4]),
    .b(mux31_b3_sel_is_2_o),
    .o(n213[4]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3376 (
    .a(_al_u3063_o),
    .b(_al_u2929_o),
    .o(_al_u3376_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(A*~(D*~C)))"),
    .INIT(16'h4c44))
    _al_u3377 (
    .a(n213[4]),
    .b(_al_u3376_o),
    .c(_al_u3226_o),
    .d(_al_u2927_o),
    .o(_al_u3377_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*C)*~(B*~A))"),
    .INIT(16'hbb0b))
    _al_u3378 (
    .a(_al_u3368_o),
    .b(_al_u3377_o),
    .c(_al_u2944_o),
    .d(_al_u2886_o),
    .o(_al_u3378_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*B))"),
    .INIT(8'ha2))
    _al_u3379 (
    .a(_al_u3378_o),
    .b(_al_u2958_o),
    .c(_al_u2893_o),
    .o(_al_u3379_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u3380 (
    .a(_al_u3379_o),
    .b(_al_u2960_o),
    .c(_al_u3236_o),
    .o(_al_u3380_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*A))"),
    .INIT(8'hc4))
    _al_u3381 (
    .a(_al_u3380_o),
    .b(mux84_b4_sel_is_2_o),
    .c(_al_u3238_o),
    .o(_al_u3381_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(~D*C*~B))"),
    .INIT(16'haa8a))
    _al_u3382 (
    .a(_al_u3381_o),
    .b(_al_u2893_o),
    .c(_al_u2887_o),
    .d(_al_u2884_o),
    .o(_al_u3382_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3383 (
    .a(_al_u3382_o),
    .b(_al_u2970_o),
    .o(_al_u3383_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3384 (
    .a(_al_u3383_o),
    .b(mux103_b3_sel_is_0_o),
    .c(_al_u3194_o),
    .o(_al_u3384_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*~B))"),
    .INIT(8'ha8))
    _al_u3385 (
    .a(_al_u3384_o),
    .b(_al_u3076_o),
    .c(mux107_b0_sel_is_2_o),
    .o(_al_u3385_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(~B*~A))"),
    .INIT(8'he0))
    _al_u3386 (
    .a(_al_u2885_o),
    .b(_al_u2889_o),
    .c(_al_u2992_o),
    .o(_al_u3386_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3387 (
    .a(_al_u3082_o),
    .b(_al_u3348_o),
    .c(_al_u3386_o),
    .o(mux119_b4_sel_is_2_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3388 (
    .a(_al_u3385_o),
    .b(mux119_b4_sel_is_2_o),
    .c(_al_u2990_o),
    .o(_al_u3388_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u3389 (
    .a(_al_u3006_o),
    .b(_al_u3083_o),
    .c(counter[0]),
    .o(mux123_b10_sel_is_2_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(B*A))"),
    .INIT(8'h07))
    _al_u3390 (
    .a(_al_u3388_o),
    .b(mux123_b10_sel_is_2_o),
    .c(_al_u3014_o),
    .o(_al_u3390_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    _al_u3391 (
    .a(_al_u2900_o),
    .b(_al_u2884_o),
    .c(_al_u3010_o),
    .o(_al_u3391_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u3392 (
    .a(_al_u3390_o),
    .b(_al_u3015_o),
    .c(_al_u3391_o),
    .o(_al_u3392_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3393 (
    .a(_al_u3392_o),
    .b(mux137_b2_sel_is_2_o),
    .o(_al_u3393_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u3394 (
    .a(mux148_b3_sel_is_2_o),
    .b(_al_u2893_o),
    .c(_al_u3022_o),
    .o(mux149_b4_sel_is_2_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3395 (
    .a(_al_u3393_o),
    .b(mux149_b4_sel_is_2_o),
    .c(_al_u3027_o),
    .o(_al_u3395_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3396 (
    .a(_al_u3395_o),
    .b(mux153_b3_sel_is_2_o),
    .o(_al_u3396_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~D*~C*A))"),
    .INIT(16'hccc4))
    _al_u3397 (
    .a(_al_u3396_o),
    .b(_al_u3167_o),
    .c(_al_u3036_o),
    .d(_al_u3042_o),
    .o(_al_u3397_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u3398 (
    .a(_al_u2913_o),
    .b(_al_u3042_o),
    .o(_al_u3398_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3399 (
    .a(_al_u3045_o),
    .b(counter[0]),
    .o(_al_u3399_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u3400 (
    .a(_al_u3397_o),
    .b(_al_u3398_o),
    .c(_al_u3399_o),
    .o(_al_u3400_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u3401 (
    .a(mux63_b12_sel_is_2_o),
    .b(_al_u2902_o),
    .c(_al_u3272_o),
    .o(mux83_b12_sel_is_2_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3402 (
    .a(_al_u3336_o),
    .b(_al_u3291_o),
    .o(_al_u3402_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3403 (
    .a(_al_u3266_o),
    .b(mux16_b0_sel_is_2_o),
    .c(_al_u3402_o),
    .o(_al_u3403_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3404 (
    .a(_al_u3403_o),
    .b(_al_u2928_o),
    .o(_al_u3404_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3405 (
    .a(mux83_b12_sel_is_2_o),
    .b(_al_u3404_o),
    .c(_al_u3068_o),
    .o(_al_u3405_o));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    _al_u3406 (
    .a(_al_u3405_o),
    .b(_al_u2973_o),
    .o(_al_u3406_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u3407 (
    .a(_al_u3406_o),
    .b(_al_u3244_o),
    .o(_al_u3407_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3408 (
    .a(_al_u3407_o),
    .b(mux111_b0_sel_is_2_o),
    .c(_al_u3151_o),
    .o(_al_u3408_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u3409 (
    .a(_al_u3408_o),
    .b(_al_u2989_o),
    .c(counter[0]),
    .o(_al_u3409_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u3410 (
    .a(_al_u3409_o),
    .b(_al_u2995_o),
    .c(_al_u2992_o),
    .o(_al_u3410_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(B*~A))"),
    .INIT(8'h0b))
    _al_u3411 (
    .a(_al_u3410_o),
    .b(mux130_b1_sel_is_2_o),
    .c(_al_u3011_o),
    .o(_al_u3411_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3412 (
    .a(_al_u3411_o),
    .b(_al_u3090_o),
    .o(_al_u3412_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3413 (
    .a(_al_u3412_o),
    .b(_al_u3358_o),
    .o(_al_u3413_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(~B*~A))"),
    .INIT(8'he0))
    _al_u3414 (
    .a(_al_u2896_o),
    .b(_al_u2897_o),
    .c(_al_u3022_o),
    .o(_al_u3414_o));
  AL_MAP_LUT4 #(
    .EQN("~((~C*A)*~(D)*~(B)+(~C*A)*D*~(B)+~((~C*A))*D*B+(~C*A)*D*B)"),
    .INIT(16'h31fd))
    _al_u3415 (
    .a(_al_u3413_o),
    .b(_al_u3031_o),
    .c(_al_u3414_o),
    .d(counter[0]),
    .o(_al_u3415_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*~A)"),
    .INIT(8'h04))
    _al_u3416 (
    .a(_al_u3415_o),
    .b(_al_u3258_o),
    .c(_al_u3034_o),
    .o(_al_u3416_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u3417 (
    .a(_al_u3165_o),
    .b(_al_u3166_o),
    .c(_al_u3036_o),
    .o(_al_u3417_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3418 (
    .a(_al_u3416_o),
    .b(_al_u3417_o),
    .o(_al_u3418_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    _al_u3419 (
    .a(_al_u2893_o),
    .b(_al_u3042_o),
    .c(_al_u2889_o),
    .o(_al_u3419_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3420 (
    .a(_al_u3418_o),
    .b(_al_u3419_o),
    .o(_al_u3420_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3421 (
    .a(_al_u3048_o),
    .b(_al_u3045_o),
    .o(_al_u3421_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3422 (
    .a(_al_u3420_o),
    .b(_al_u3106_o),
    .c(_al_u3421_o),
    .o(_al_u3422_o));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*~B)*~(C*~A))"),
    .INIT(16'h7350))
    _al_u3423 (
    .a(_al_u3400_o),
    .b(_al_u3422_o),
    .c(_al_u3107_o),
    .d(n376_lutinv),
    .o(\sel2_b4/or_B6_or_B7_B8_o_o ));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u3424 (
    .a(_al_u2842_o),
    .b(_al_u3058_o),
    .c(_al_u2900_o),
    .o(_al_u3424_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*~A)"),
    .INIT(8'h04))
    _al_u3425 (
    .a(_al_u3290_o),
    .b(_al_u3424_o),
    .c(_al_u3110_o),
    .o(_al_u3425_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3426 (
    .a(_al_u2912_o),
    .b(_al_u2903_o),
    .o(_al_u3426_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3427 (
    .a(_al_u3425_o),
    .b(_al_u3426_o),
    .o(_al_u3427_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*A*~(~D*~C))"),
    .INIT(16'h2220))
    _al_u3428 (
    .a(_al_u3427_o),
    .b(_al_u2921_o),
    .c(counter[0]),
    .d(_al_u3109_o),
    .o(_al_u3428_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*B))"),
    .INIT(8'ha2))
    _al_u3429 (
    .a(_al_u3428_o),
    .b(_al_u3222_o),
    .c(counter[0]),
    .o(_al_u3429_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3430 (
    .a(_al_u3429_o),
    .b(_al_u2930_o),
    .c(_al_u2925_o),
    .o(_al_u3430_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3431 (
    .a(_al_u3430_o),
    .b(_al_u2935_o),
    .o(_al_u3431_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3432 (
    .a(_al_u2897_o),
    .b(_al_u2927_o),
    .o(_al_u3432_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(~B*~(~D*C)))"),
    .INIT(16'h88a8))
    _al_u3433 (
    .a(_al_u3431_o),
    .b(_al_u2950_o),
    .c(mux83_b12_sel_is_2_o),
    .d(_al_u3432_o),
    .o(_al_u3433_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u3434 (
    .a(_al_u3142_o),
    .b(_al_u2886_o),
    .c(_al_u2958_o),
    .o(_al_u3434_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(A*~(~D*C)))"),
    .INIT(16'h44c4))
    _al_u3435 (
    .a(_al_u3433_o),
    .b(_al_u3434_o),
    .c(_al_u2887_o),
    .d(_al_u2896_o),
    .o(_al_u3435_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3436 (
    .a(_al_u3435_o),
    .b(_al_u3140_o),
    .o(_al_u3436_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3437 (
    .a(_al_u2910_o),
    .b(_al_u2887_o),
    .o(_al_u3437_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u3438 (
    .a(_al_u3436_o),
    .b(_al_u2979_o),
    .c(_al_u3437_o),
    .o(_al_u3438_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*~A)"),
    .INIT(8'h04))
    _al_u3439 (
    .a(_al_u3438_o),
    .b(_al_u2973_o),
    .c(_al_u2976_o),
    .o(_al_u3439_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3440 (
    .a(_al_u2893_o),
    .b(_al_u2969_o),
    .o(_al_u3440_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3441 (
    .a(_al_u3439_o),
    .b(_al_u3440_o),
    .o(_al_u3441_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u3442 (
    .a(_al_u3075_o),
    .b(_al_u2989_o),
    .c(_al_u3077_o),
    .o(_al_u3442_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3443 (
    .a(_al_u3441_o),
    .b(_al_u3442_o),
    .c(_al_u2984_o),
    .o(_al_u3443_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3444 (
    .a(_al_u3443_o),
    .b(_al_u3001_o),
    .o(_al_u3444_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u3445 (
    .a(_al_u3006_o),
    .b(_al_u3083_o),
    .c(counter[0]),
    .o(_al_u3445_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3446 (
    .a(_al_u3444_o),
    .b(_al_u3445_o),
    .c(_al_u3004_o),
    .o(_al_u3446_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3447 (
    .a(_al_u3446_o),
    .b(_al_u3248_o),
    .o(_al_u3447_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u3448 (
    .a(_al_u3447_o),
    .b(_al_u3092_o),
    .c(_al_u3086_o),
    .o(_al_u3448_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3449 (
    .a(_al_u3448_o),
    .b(_al_u3157_o),
    .o(_al_u3449_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u3450 (
    .a(_al_u3449_o),
    .b(_al_u3358_o),
    .c(_al_u3155_o),
    .o(_al_u3450_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3451 (
    .a(_al_u3450_o),
    .b(_al_u3161_o),
    .o(_al_u3451_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3452 (
    .a(_al_u3451_o),
    .b(_al_u3258_o),
    .c(_al_u3031_o),
    .o(_al_u3452_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3453 (
    .a(_al_u3452_o),
    .b(_al_u3033_o),
    .o(_al_u3453_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u3454 (
    .a(_al_u3453_o),
    .b(_al_u3166_o),
    .c(_al_u3164_o),
    .o(_al_u3454_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3455 (
    .a(_al_u3454_o),
    .b(_al_u3334_o),
    .o(_al_u3455_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(~B*~(D*A)))"),
    .INIT(16'he0c0))
    _al_u3456 (
    .a(_al_u2955_o),
    .b(_al_u2896_o),
    .c(_al_u3042_o),
    .d(counter[0]),
    .o(_al_u3456_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u3457 (
    .a(_al_u3455_o),
    .b(_al_u3048_o),
    .c(_al_u3456_o),
    .o(_al_u3457_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3458 (
    .a(_al_u3457_o),
    .b(_al_u3099_o),
    .o(_al_u3458_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u3459 (
    .a(_al_u3111_o),
    .b(_al_u3175_o),
    .c(_al_u3290_o),
    .o(_al_u3459_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3460 (
    .a(_al_u3459_o),
    .b(mux16_b0_sel_is_2_o),
    .c(_al_u3115_o),
    .o(n200[0]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3461 (
    .a(n200[0]),
    .b(mux21_b0_sel_is_0_o),
    .o(n203[0]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(~D*~C*A))"),
    .INIT(16'h3331))
    _al_u3462 (
    .a(n203[0]),
    .b(_al_u2924_o),
    .c(_al_u2925_o),
    .d(_al_u3222_o),
    .o(_al_u3462_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u3463 (
    .a(_al_u3462_o),
    .b(mux33_b0_sel_is_2_o),
    .o(n214[0]));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3464 (
    .a(n214[0]),
    .b(mux49_b0_sel_is_2_o),
    .c(_al_u2934_o),
    .o(_al_u3464_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3465 (
    .a(_al_u3464_o),
    .b(mux61_b0_sel_is_2_o),
    .o(_al_u3465_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3466 (
    .a(_al_u2897_o),
    .b(_al_u2958_o),
    .o(_al_u3466_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3467 (
    .a(_al_u3465_o),
    .b(mux68_b0_sel_is_2_o),
    .c(_al_u3466_o),
    .o(_al_u3467_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3468 (
    .a(_al_u3467_o),
    .b(_al_u2960_o),
    .o(_al_u3468_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(~B*~A))"),
    .INIT(8'he0))
    _al_u3469 (
    .a(_al_u2910_o),
    .b(_al_u2912_o),
    .c(_al_u2958_o),
    .o(_al_u3469_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u3470 (
    .a(_al_u3468_o),
    .b(_al_u3469_o),
    .c(_al_u3238_o),
    .o(_al_u3470_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3471 (
    .a(_al_u3470_o),
    .b(mux87_b0_sel_is_2_o),
    .o(_al_u3471_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(~D*~C*~B))"),
    .INIT(16'haaa8))
    _al_u3472 (
    .a(_al_u3471_o),
    .b(_al_u3140_o),
    .c(mux97_b2_sel_is_2_o),
    .d(_al_u2894_o),
    .o(_al_u3472_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3473 (
    .a(_al_u3472_o),
    .b(mux103_b0_sel_is_2_o),
    .c(mux107_b0_sel_is_2_o),
    .o(_al_u3473_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3474 (
    .a(_al_u3473_o),
    .b(mux111_b0_sel_is_2_o),
    .o(_al_u3474_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3475 (
    .a(_al_u3474_o),
    .b(_al_u2999_o),
    .c(mux119_b3_sel_is_0_o),
    .o(_al_u3475_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~B*~A)*~(D)*~(C)+~(~B*~A)*D*~(C)+~(~(~B*~A))*D*C+~(~B*~A)*D*C)"),
    .INIT(16'hfe0e))
    _al_u3476 (
    .a(_al_u3475_o),
    .b(_al_u3145_o),
    .c(_al_u3006_o),
    .d(counter[0]),
    .o(_al_u3476_o));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'h47))
    _al_u3477 (
    .a(_al_u3476_o),
    .b(mux130_b6_sel_is_2_o),
    .c(_al_u3011_o),
    .o(_al_u3477_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u3478 (
    .a(mux132_b0_sel_is_0_o),
    .b(_al_u3202_o),
    .c(_al_u3092_o),
    .o(mux135_b0_sel_is_2_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u3479 (
    .a(mux135_b0_sel_is_2_o),
    .b(_al_u2911_o),
    .c(_al_u3010_o),
    .o(mux139_b0_sel_is_2_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    _al_u3480 (
    .a(_al_u3477_o),
    .b(_al_u3359_o),
    .c(mux139_b0_sel_is_2_o),
    .o(_al_u3480_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(~B*~A))"),
    .INIT(8'he0))
    _al_u3481 (
    .a(_al_u2956_o),
    .b(_al_u2892_o),
    .c(_al_u3022_o),
    .o(_al_u3481_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*~A))"),
    .INIT(8'h23))
    _al_u3482 (
    .a(_al_u3480_o),
    .b(_al_u3481_o),
    .c(_al_u3356_o),
    .o(_al_u3482_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3483 (
    .a(_al_u3038_o),
    .b(_al_u3256_o),
    .o(mux156_b0_sel_is_2_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3484 (
    .a(mux158_b11_sel_is_0_o),
    .b(mux156_b0_sel_is_2_o),
    .o(_al_u3484_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(~C*~(B*A)))"),
    .INIT(16'h00f8))
    _al_u3485 (
    .a(_al_u3482_o),
    .b(_al_u3484_o),
    .c(_al_u3033_o),
    .d(_al_u3036_o),
    .o(_al_u3485_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3486 (
    .a(_al_u3485_o),
    .b(_al_u3260_o),
    .o(_al_u3486_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3487 (
    .a(_al_u3486_o),
    .b(mux169_b0_sel_is_2_o),
    .c(mux174_b0_sel_is_0_o),
    .o(_al_u3487_o));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'h47))
    _al_u3488 (
    .a(_al_u3487_o),
    .b(n377_lutinv),
    .c(n378_lutinv),
    .o(_al_u3488_o));
  AL_MAP_LUT4 #(
    .EQN("~(B*~(C*~(~D*A)))"),
    .INIT(16'hf373))
    _al_u3489 (
    .a(_al_u3458_o),
    .b(_al_u3488_o),
    .c(n376_lutinv),
    .d(_al_u3102_o),
    .o(\sel2_b0/or_or_B4_B5_o_or_B6__o ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    _al_u3490 (
    .a(_al_u2909_o),
    .b(mux16_b11_sel_is_2_o),
    .c(_al_u2986_o),
    .o(n198[5]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3491 (
    .a(n198[5]),
    .b(mux19_b2_sel_is_0_o),
    .o(n201[5]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u3492 (
    .a(_al_u2982_o),
    .b(_al_u2917_o),
    .o(_al_u3492_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u3493 (
    .a(n201[5]),
    .b(_al_u3181_o),
    .c(_al_u3492_o),
    .o(n206[5]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3494 (
    .a(n206[5]),
    .b(_al_u3296_o),
    .o(n212[5]));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(B*A))"),
    .INIT(8'h07))
    _al_u3495 (
    .a(n212[5]),
    .b(mux38_b1_sel_is_2_o),
    .c(_al_u3432_o),
    .o(_al_u3495_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*~A)"),
    .INIT(16'h4000))
    _al_u3496 (
    .a(_al_u3274_o),
    .b(mux49_b5_sel_is_0_o),
    .c(mux52_b1_sel_is_2_o),
    .d(_al_u3269_o),
    .o(_al_u3496_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*~A)"),
    .INIT(8'h04))
    _al_u3497 (
    .a(_al_u3495_o),
    .b(_al_u3496_o),
    .c(_al_u2942_o),
    .o(_al_u3497_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*~A))"),
    .INIT(8'h32))
    _al_u3498 (
    .a(_al_u3497_o),
    .b(_al_u2965_o),
    .c(_al_u3268_o),
    .o(_al_u3498_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3499 (
    .a(_al_u3498_o),
    .b(mux75_b5_sel_is_2_o),
    .c(_al_u3307_o),
    .o(_al_u3499_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3500 (
    .a(_al_u3499_o),
    .b(_al_u3238_o),
    .o(_al_u3500_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3501 (
    .a(_al_u3500_o),
    .b(mux85_b0_sel_is_2_o),
    .o(_al_u3501_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3502 (
    .a(_al_u3501_o),
    .b(mux97_b15_sel_is_2_o),
    .c(_al_u3066_o),
    .o(_al_u3502_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3503 (
    .a(_al_u3502_o),
    .b(_al_u3195_o),
    .c(_al_u3440_o),
    .o(_al_u3503_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u3504 (
    .a(_al_u3503_o),
    .b(_al_u3076_o),
    .c(counter[0]),
    .o(_al_u3504_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*~A)"),
    .INIT(8'h04))
    _al_u3505 (
    .a(_al_u3504_o),
    .b(mux111_b0_sel_is_2_o),
    .c(_al_u3151_o),
    .o(_al_u3505_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3506 (
    .a(_al_u2989_o),
    .b(counter[0]),
    .o(_al_u3506_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(A*~(D*B)))"),
    .INIT(16'h0d05))
    _al_u3507 (
    .a(_al_u3505_o),
    .b(_al_u3080_o),
    .c(_al_u3506_o),
    .d(_al_u2992_o),
    .o(_al_u3507_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3508 (
    .a(_al_u3507_o),
    .b(_al_u3391_o),
    .o(_al_u3508_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3509 (
    .a(_al_u3089_o),
    .b(_al_u3092_o),
    .o(mux137_b5_sel_is_2_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3510 (
    .a(_al_u3508_o),
    .b(mux137_b5_sel_is_2_o),
    .o(_al_u3510_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3511 (
    .a(mux140_b5_sel_is_0_o),
    .b(_al_u3022_o),
    .o(_al_u3511_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3512 (
    .a(_al_u3511_o),
    .b(_al_u3096_o),
    .o(mux159_b5_sel_is_2_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3513 (
    .a(_al_u3510_o),
    .b(mux159_b5_sel_is_2_o),
    .c(_al_u3212_o),
    .o(_al_u3513_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3514 (
    .a(_al_u3513_o),
    .b(_al_u3456_o),
    .o(_al_u3514_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*~B))"),
    .INIT(8'h8a))
    _al_u3515 (
    .a(_al_u3514_o),
    .b(_al_u3399_o),
    .c(_al_u3216_o),
    .o(_al_u3515_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~A*~(D*C)))"),
    .INIT(16'hc888))
    _al_u3516 (
    .a(_al_u3515_o),
    .b(_al_u3107_o),
    .c(_al_u2910_o),
    .d(_al_u3042_o),
    .o(_al_u3516_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3517 (
    .a(_al_u3174_o),
    .b(_al_u3058_o),
    .o(_al_u3517_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3518 (
    .a(_al_u3266_o),
    .b(_al_u3517_o),
    .o(_al_u3518_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u3519 (
    .a(_al_u3518_o),
    .b(_al_u2928_o),
    .c(_al_u2934_o),
    .o(_al_u3519_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3520 (
    .a(_al_u3519_o),
    .b(_al_u3068_o),
    .o(_al_u3520_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    _al_u3521 (
    .a(_al_u3076_o),
    .b(_al_u2984_o),
    .c(_al_u3520_o),
    .o(_al_u3521_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3522 (
    .a(_al_u3521_o),
    .b(_al_u3075_o),
    .c(_al_u2989_o),
    .o(_al_u3522_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3523 (
    .a(_al_u3522_o),
    .b(_al_u3386_o),
    .o(_al_u3523_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u3524 (
    .a(_al_u3523_o),
    .b(_al_u3013_o),
    .c(_al_u3084_o),
    .d(mux132_b0_sel_is_0_o),
    .o(_al_u3524_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3525 (
    .a(_al_u3524_o),
    .b(_al_u3092_o),
    .o(_al_u3525_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3526 (
    .a(_al_u3525_o),
    .b(mux140_b11_sel_is_2_o),
    .o(_al_u3526_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    _al_u3527 (
    .a(_al_u3526_o),
    .b(mux156_b0_sel_is_2_o),
    .c(_al_u3031_o),
    .d(_al_u3414_o),
    .o(_al_u3527_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3528 (
    .a(_al_u3527_o),
    .b(_al_u3417_o),
    .c(_al_u3050_o),
    .o(_al_u3528_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    _al_u3529 (
    .a(_al_u3216_o),
    .b(_al_u3102_o),
    .c(_al_u3528_o),
    .o(_al_u3529_o));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~A*~(C*~B))"),
    .INIT(16'hffba))
    _al_u3530 (
    .a(_al_u3516_o),
    .b(_al_u3529_o),
    .c(n376_lutinv),
    .d(n375_lutinv),
    .o(\sel2_b5/or_B6_or_B7_B8_o_o ));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(~B*~(~C*~A)))"),
    .INIT(16'h00cd))
    _al_u3531 (
    .a(_al_u3109_o),
    .b(_al_u3052_o),
    .c(_al_u3219_o),
    .d(_al_u3288_o),
    .o(_al_u3531_o));
  AL_MAP_LUT3 #(
    .EQN("(~(A)*~(B)*~(C)+A*~(B)*~(C)+A*B*~(C)+~(A)*~(B)*C+A*B*C)"),
    .INIT(8'h9b))
    _al_u3532 (
    .a(_al_u3531_o),
    .b(mux14_b11_sel_is_2_o),
    .c(_al_u3053_o),
    .o(_al_u3532_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*~A))"),
    .INIT(8'h32))
    _al_u3533 (
    .a(_al_u3532_o),
    .b(_al_u2921_o),
    .c(_al_u2917_o),
    .o(_al_u3533_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3534 (
    .a(_al_u3533_o),
    .b(_al_u3264_o),
    .c(_al_u3182_o),
    .o(_al_u3534_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    _al_u3535 (
    .a(_al_u3534_o),
    .b(mux38_b1_sel_is_2_o),
    .c(mux42_b0_sel_is_2_o),
    .o(n223[1]));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3536 (
    .a(n223[1]),
    .b(mux47_b1_sel_is_2_o),
    .c(_al_u2946_o),
    .o(_al_u3536_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3537 (
    .a(_al_u3536_o),
    .b(mux63_b1_sel_is_2_o),
    .o(_al_u3537_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3538 (
    .a(_al_u3537_o),
    .b(mux68_b1_sel_is_2_o),
    .c(_al_u3466_o),
    .o(_al_u3538_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u3539 (
    .a(_al_u3538_o),
    .b(_al_u2912_o),
    .c(_al_u2958_o),
    .o(_al_u3539_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3540 (
    .a(_al_u3310_o),
    .b(_al_u3235_o),
    .o(_al_u3540_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3541 (
    .a(_al_u3539_o),
    .b(_al_u3540_o),
    .o(_al_u3541_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3542 (
    .a(_al_u3541_o),
    .b(_al_u2902_o),
    .o(_al_u3542_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u3543 (
    .a(_al_u3542_o),
    .b(_al_u3139_o),
    .c(_al_u3142_o),
    .o(_al_u3543_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3544 (
    .a(_al_u3543_o),
    .b(mux94_b0_sel_is_2_o),
    .o(_al_u3544_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*A*~(~D*C))"),
    .INIT(16'h2202))
    _al_u3545 (
    .a(_al_u3544_o),
    .b(_al_u2971_o),
    .c(_al_u2969_o),
    .d(_al_u2981_o),
    .o(_al_u3545_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~A*~(D*C))"),
    .INIT(16'h0111))
    _al_u3546 (
    .a(_al_u3545_o),
    .b(_al_u3193_o),
    .c(mux107_b0_sel_is_2_o),
    .d(_al_u3074_o),
    .o(_al_u3546_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3547 (
    .a(_al_u3546_o),
    .b(_al_u2996_o),
    .o(_al_u3547_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3548 (
    .a(_al_u3547_o),
    .b(_al_u3386_o),
    .o(_al_u3548_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3549 (
    .a(_al_u3548_o),
    .b(mux124_b11_sel_is_2_o),
    .c(_al_u3004_o),
    .o(_al_u3549_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3550 (
    .a(mux130_b1_sel_is_2_o),
    .b(mux132_b0_sel_is_0_o),
    .c(_al_u3202_o),
    .o(_al_u3550_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(B*~(~C*~A)))"),
    .INIT(16'h0037))
    _al_u3551 (
    .a(_al_u3549_o),
    .b(_al_u3550_o),
    .c(_al_u3324_o),
    .d(_al_u3091_o),
    .o(_al_u3551_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u3552 (
    .a(mux140_b1_sel_is_2_o),
    .b(_al_u2938_o),
    .c(_al_u3010_o),
    .o(mux141_b1_sel_is_2_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~C*~(D*~A)))"),
    .INIT(16'hc4c0))
    _al_u3553 (
    .a(_al_u3551_o),
    .b(mux141_b1_sel_is_2_o),
    .c(_al_u3252_o),
    .d(mux137_b5_sel_is_2_o),
    .o(_al_u3553_o));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'h47))
    _al_u3554 (
    .a(_al_u3553_o),
    .b(_al_u3359_o),
    .c(_al_u3169_o),
    .o(_al_u3554_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(~B*~A))"),
    .INIT(8'he0))
    _al_u3555 (
    .a(_al_u2893_o),
    .b(_al_u2889_o),
    .c(_al_u3022_o),
    .o(_al_u3555_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u3556 (
    .a(_al_u3554_o),
    .b(_al_u3330_o),
    .c(_al_u3555_o),
    .o(_al_u3556_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3557 (
    .a(_al_u3556_o),
    .b(mux159_b1_sel_is_2_o),
    .o(_al_u3557_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u3558 (
    .a(_al_u3260_o),
    .b(_al_u3214_o),
    .c(_al_u3334_o),
    .o(mux166_b1_sel_is_2_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u3559 (
    .a(_al_u3048_o),
    .b(_al_u3045_o),
    .c(counter[0]),
    .o(_al_u3559_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3560 (
    .a(_al_u3557_o),
    .b(mux166_b1_sel_is_2_o),
    .c(_al_u3559_o),
    .o(_al_u3560_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u3561 (
    .a(_al_u2986_o),
    .b(_al_u3057_o),
    .c(_al_u2903_o),
    .o(mux12_b9_sel_is_2_o_neg_lutinv));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3562 (
    .a(mux12_b9_sel_is_2_o_neg_lutinv),
    .b(_al_u2914_o),
    .o(mux16_b9_sel_is_2_o_neg_lutinv));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*~(D*C)))"),
    .INIT(16'ha222))
    _al_u3563 (
    .a(_al_u3371_o),
    .b(mux16_b9_sel_is_2_o_neg_lutinv),
    .c(mux16_b1_sel_is_0_o),
    .d(_al_u2917_o),
    .o(_al_u3563_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*B))"),
    .INIT(8'ha2))
    _al_u3564 (
    .a(_al_u3563_o),
    .b(_al_u2917_o),
    .c(_al_u2907_o),
    .o(_al_u3564_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u3565 (
    .a(_al_u2910_o),
    .b(_al_u3564_o),
    .o(_al_u3565_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~D*~(~C*A)))"),
    .INIT(16'hcc08))
    _al_u3566 (
    .a(_al_u3565_o),
    .b(mux37_b6_sel_is_2_o),
    .c(_al_u3265_o),
    .d(_al_u2927_o),
    .o(_al_u3566_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*~A)"),
    .INIT(8'h04))
    _al_u3567 (
    .a(_al_u3566_o),
    .b(_al_u3496_o),
    .c(_al_u2965_o),
    .o(_al_u3567_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    _al_u3568 (
    .a(_al_u2970_o),
    .b(_al_u2972_o),
    .c(_al_u3567_o),
    .o(_al_u3568_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3569 (
    .a(_al_u3568_o),
    .b(_al_u2976_o),
    .o(_al_u3569_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*~B))"),
    .INIT(8'h8a))
    _al_u3570 (
    .a(_al_u3244_o),
    .b(_al_u2982_o),
    .c(_al_u2969_o),
    .o(mux104_b11_sel_is_2_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3571 (
    .a(_al_u3569_o),
    .b(mux104_b11_sel_is_2_o),
    .o(_al_u3571_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3572 (
    .a(_al_u3571_o),
    .b(_al_u2990_o),
    .o(_al_u3572_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3573 (
    .a(_al_u3572_o),
    .b(_al_u2993_o),
    .o(_al_u3573_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3574 (
    .a(_al_u3573_o),
    .b(_al_u3001_o),
    .c(_al_u3147_o),
    .o(_al_u3574_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3575 (
    .a(_al_u3574_o),
    .b(mux122_b11_sel_is_2_o),
    .o(_al_u3575_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u3576 (
    .a(_al_u3575_o),
    .b(_al_u2938_o),
    .c(_al_u2992_o),
    .o(_al_u3576_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3577 (
    .a(_al_u3576_o),
    .b(mux137_b2_sel_is_2_o),
    .c(_al_u3017_o),
    .o(_al_u3577_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u3578 (
    .a(_al_u3577_o),
    .b(_al_u3090_o),
    .c(_al_u3096_o),
    .o(_al_u3578_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3579 (
    .a(_al_u3578_o),
    .b(_al_u3160_o),
    .o(_al_u3579_o));
  AL_MAP_LUT4 #(
    .EQN("~(A*~(B)*~((D*C))+A*B*~((D*C))+~(A)*B*(D*C)+A*B*(D*C))"),
    .INIT(16'h3555))
    _al_u3580 (
    .a(_al_u3579_o),
    .b(_al_u2883_o),
    .c(_al_u2892_o),
    .d(_al_u3022_o),
    .o(_al_u3580_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u3581 (
    .a(_al_u3580_o),
    .b(_al_u3040_o),
    .c(_al_u3031_o),
    .o(_al_u3581_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3582 (
    .a(_al_u3581_o),
    .b(_al_u3168_o),
    .o(_al_u3582_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3583 (
    .a(_al_u3582_o),
    .b(_al_u3334_o),
    .o(_al_u3583_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u3584 (
    .a(_al_u3583_o),
    .b(_al_u2961_o),
    .c(_al_u3042_o),
    .o(_al_u3584_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B*A))"),
    .INIT(8'h70))
    _al_u3585 (
    .a(_al_u3584_o),
    .b(_al_u3106_o),
    .c(n376_lutinv),
    .o(_al_u3585_o));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    _al_u3586 (
    .a(_al_u3560_o),
    .b(_al_u3585_o),
    .c(_al_u3107_o),
    .o(\sel2_b1/or_B6_or_B7_B8_o_o ));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add0/u0  (
    .a(divider2[0]),
    .b(1'b1),
    .c(\add0/c0 ),
    .o({\add0/c1 ,n0[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add0/u1  (
    .a(divider2[1]),
    .b(1'b0),
    .c(\add0/c1 ),
    .o({\add0/c2 ,n0[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add0/u2  (
    .a(divider2[2]),
    .b(1'b0),
    .c(\add0/c2 ),
    .o({\add0/c3 ,n0[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add0/u3  (
    .a(divider2[3]),
    .b(1'b0),
    .c(\add0/c3 ),
    .o({\add0/c4 ,n0[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add0/u4  (
    .a(divider2[4]),
    .b(1'b0),
    .c(\add0/c4 ),
    .o({\add0/c5 ,n0[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add0/u5  (
    .a(divider2[5]),
    .b(1'b0),
    .c(\add0/c5 ),
    .o({\add0/c6 ,n0[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add0/u6  (
    .a(divider2[6]),
    .b(1'b0),
    .c(\add0/c6 ),
    .o({\add0/c7 ,n0[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add0/u7  (
    .a(divider2[7]),
    .b(1'b0),
    .c(\add0/c7 ),
    .o({\add0/c8 ,n0[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add0/u8  (
    .a(divider2[8]),
    .b(1'b0),
    .c(\add0/c8 ),
    .o({open_n0,n0[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \add0/ucin  (
    .a(1'b0),
    .o({\add0/c0 ,open_n3}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add1/u0  (
    .a(cnt[0]),
    .b(1'b1),
    .c(\add1/c0 ),
    .o({\add1/c1 ,n371[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add1/u1  (
    .a(cnt[1]),
    .b(1'b0),
    .c(\add1/c1 ),
    .o({\add1/c2 ,n371[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add1/u2  (
    .a(cnt[2]),
    .b(1'b0),
    .c(\add1/c2 ),
    .o({\add1/c3 ,n371[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add1/u3  (
    .a(cnt[3]),
    .b(1'b0),
    .c(\add1/c3 ),
    .o({\add1/c4 ,n371[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add1/u4  (
    .a(cnt[4]),
    .b(1'b0),
    .c(\add1/c4 ),
    .o({\add1/c5 ,n371[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add1/u5  (
    .a(cnt[5]),
    .b(1'b0),
    .c(\add1/c5 ),
    .o({\add1/c6 ,n371[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add1/u6  (
    .a(cnt[6]),
    .b(1'b0),
    .c(\add1/c6 ),
    .o({\add1/c7 ,n371[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add1/u7  (
    .a(cnt[7]),
    .b(1'b0),
    .c(\add1/c7 ),
    .o({open_n4,n371[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \add1/ucin  (
    .a(1'b0),
    .o({\add1/c0 ,open_n7}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add2/u0  (
    .a(counter[0]),
    .b(1'b1),
    .c(\add2/c0 ),
    .o({\add2/c1 ,n372[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add2/u1  (
    .a(counter[1]),
    .b(1'b0),
    .c(\add2/c1 ),
    .o({\add2/c2 ,n372[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add2/u2  (
    .a(counter[2]),
    .b(1'b0),
    .c(\add2/c2 ),
    .o({\add2/c3 ,n372[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add2/u3  (
    .a(counter[3]),
    .b(1'b0),
    .c(\add2/c3 ),
    .o({\add2/c4 ,n372[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add2/u4  (
    .a(counter[4]),
    .b(1'b0),
    .c(\add2/c4 ),
    .o({\add2/c5 ,n372[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add2/u5  (
    .a(counter[5]),
    .b(1'b0),
    .c(\add2/c5 ),
    .o({\add2/c6 ,n372[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add2/u6  (
    .a(counter[6]),
    .b(1'b0),
    .c(\add2/c6 ),
    .o({\add2/c7 ,n372[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add2/u7  (
    .a(counter[7]),
    .b(1'b0),
    .c(\add2/c7 ),
    .o({open_n8,n372[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \add2/ucin  (
    .a(1'b0),
    .o({\add2/c0 ,open_n11}));
  reg_ar_as_w1 bus_write_reg (
    .clk(divider2[8]),
    .d(n366),
    .en(1'b1),
    .reset(~reset_n),
    .set(1'b0),
    .q(bus_write));  // sources/rtl/camera_init.v(389)
  reg_ar_as_w1 ready_reg (
    .clk(clk),
    .d(n382),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(ready));  // sources/rtl/camera_init.v(265)
  reg_ar_as_w1 reg0_b0 (
    .clk(divider2[8]),
    .d(sel1_b0_sel_o),
    .en(1'b1),
    .reset(~reset_n),
    .set(1'b0),
    .q(reg_address[0]));  // sources/rtl/camera_init.v(389)
  reg_ar_as_w1 reg0_b1 (
    .clk(divider2[8]),
    .d(sel1_b1_sel_o),
    .en(1'b1),
    .reset(~reset_n),
    .set(1'b0),
    .q(reg_address[1]));  // sources/rtl/camera_init.v(389)
  reg_ar_as_w1 reg1_b0 (
    .clk(divider2[8]),
    .d(\sel2_b0/or_or_B4_B5_o_or_B6__o ),
    .en(1'b1),
    .reset(~reset_n),
    .set(1'b0),
    .q(data_in_bus[0]));  // sources/rtl/camera_init.v(389)
  reg_ar_as_w1 reg1_b1 (
    .clk(divider2[8]),
    .d(\sel2_b1/or_B6_or_B7_B8_o_o ),
    .en(1'b1),
    .reset(~reset_n),
    .set(1'b0),
    .q(data_in_bus[1]));  // sources/rtl/camera_init.v(389)
  reg_ar_as_w1 reg1_b2 (
    .clk(divider2[8]),
    .d(\sel2_b2/or_B6_or_B7_B8_o_o ),
    .en(1'b1),
    .reset(~reset_n),
    .set(1'b0),
    .q(data_in_bus[2]));  // sources/rtl/camera_init.v(389)
  reg_ar_as_w1 reg1_b3 (
    .clk(divider2[8]),
    .d(\sel2_b3/or_B6_or_B7_B8_o_o ),
    .en(1'b1),
    .reset(~reset_n),
    .set(1'b0),
    .q(data_in_bus[3]));  // sources/rtl/camera_init.v(389)
  reg_ar_as_w1 reg1_b4 (
    .clk(divider2[8]),
    .d(\sel2_b4/or_B6_or_B7_B8_o_o ),
    .en(1'b1),
    .reset(~reset_n),
    .set(1'b0),
    .q(data_in_bus[4]));  // sources/rtl/camera_init.v(389)
  reg_ar_as_w1 reg1_b5 (
    .clk(divider2[8]),
    .d(\sel2_b5/or_B6_or_B7_B8_o_o ),
    .en(1'b1),
    .reset(~reset_n),
    .set(1'b0),
    .q(data_in_bus[5]));  // sources/rtl/camera_init.v(389)
  reg_ar_as_w1 reg1_b6 (
    .clk(divider2[8]),
    .d(\sel2_b6/or_B6_or_B7_B8_o_o ),
    .en(1'b1),
    .reset(~reset_n),
    .set(1'b0),
    .q(data_in_bus[6]));  // sources/rtl/camera_init.v(389)
  reg_ar_as_w1 reg1_b7 (
    .clk(divider2[8]),
    .d(\sel2_b7/or_B6_or_B7_B8_o_o ),
    .en(1'b1),
    .reset(~reset_n),
    .set(1'b0),
    .q(data_in_bus[7]));  // sources/rtl/camera_init.v(389)
  reg_ar_as_w1 reg2_b0 (
    .clk(divider2[8]),
    .d(n374[0]),
    .en(n380),
    .reset(~reset_n),
    .set(1'b0),
    .q(counter[0]));  // sources/rtl/camera_init.v(389)
  reg_ar_as_w1 reg2_b1 (
    .clk(divider2[8]),
    .d(n374[1]),
    .en(n380),
    .reset(~reset_n),
    .set(1'b0),
    .q(counter[1]));  // sources/rtl/camera_init.v(389)
  reg_ar_as_w1 reg2_b2 (
    .clk(divider2[8]),
    .d(n374[2]),
    .en(n380),
    .reset(~reset_n),
    .set(1'b0),
    .q(counter[2]));  // sources/rtl/camera_init.v(389)
  reg_ar_as_w1 reg2_b3 (
    .clk(divider2[8]),
    .d(n374[3]),
    .en(n380),
    .reset(~reset_n),
    .set(1'b0),
    .q(counter[3]));  // sources/rtl/camera_init.v(389)
  reg_ar_as_w1 reg2_b4 (
    .clk(divider2[8]),
    .d(n374[4]),
    .en(n380),
    .reset(~reset_n),
    .set(1'b0),
    .q(counter[4]));  // sources/rtl/camera_init.v(389)
  reg_ar_as_w1 reg2_b5 (
    .clk(divider2[8]),
    .d(n374[5]),
    .en(n380),
    .reset(~reset_n),
    .set(1'b0),
    .q(counter[5]));  // sources/rtl/camera_init.v(389)
  reg_ar_as_w1 reg2_b6 (
    .clk(divider2[8]),
    .d(n374[6]),
    .en(n380),
    .reset(~reset_n),
    .set(1'b0),
    .q(counter[6]));  // sources/rtl/camera_init.v(389)
  reg_ar_as_w1 reg2_b7 (
    .clk(divider2[8]),
    .d(n374[7]),
    .en(n380),
    .reset(~reset_n),
    .set(1'b0),
    .q(counter[7]));  // sources/rtl/camera_init.v(389)
  reg_ar_as_w1 reg3_b0 (
    .clk(divider2[8]),
    .d(n371[0]),
    .en(mux181_b0_sel_is_2_o),
    .reset(1'b0),
    .set(1'b0),
    .q(cnt[0]));  // sources/rtl/camera_init.v(389)
  reg_ar_as_w1 reg3_b1 (
    .clk(divider2[8]),
    .d(n371[1]),
    .en(mux181_b0_sel_is_2_o),
    .reset(1'b0),
    .set(1'b0),
    .q(cnt[1]));  // sources/rtl/camera_init.v(389)
  reg_ar_as_w1 reg3_b2 (
    .clk(divider2[8]),
    .d(n371[2]),
    .en(mux181_b0_sel_is_2_o),
    .reset(1'b0),
    .set(1'b0),
    .q(cnt[2]));  // sources/rtl/camera_init.v(389)
  reg_ar_as_w1 reg3_b3 (
    .clk(divider2[8]),
    .d(n371[3]),
    .en(mux181_b0_sel_is_2_o),
    .reset(1'b0),
    .set(1'b0),
    .q(cnt[3]));  // sources/rtl/camera_init.v(389)
  reg_ar_as_w1 reg3_b4 (
    .clk(divider2[8]),
    .d(n371[4]),
    .en(mux181_b0_sel_is_2_o),
    .reset(1'b0),
    .set(1'b0),
    .q(cnt[4]));  // sources/rtl/camera_init.v(389)
  reg_ar_as_w1 reg3_b5 (
    .clk(divider2[8]),
    .d(n371[5]),
    .en(mux181_b0_sel_is_2_o),
    .reset(1'b0),
    .set(1'b0),
    .q(cnt[5]));  // sources/rtl/camera_init.v(389)
  reg_ar_as_w1 reg3_b6 (
    .clk(divider2[8]),
    .d(n371[6]),
    .en(mux181_b0_sel_is_2_o),
    .reset(1'b0),
    .set(1'b0),
    .q(cnt[6]));  // sources/rtl/camera_init.v(389)
  reg_ar_as_w1 reg3_b7 (
    .clk(divider2[8]),
    .d(n371[7]),
    .en(mux181_b0_sel_is_2_o),
    .reset(1'b0),
    .set(1'b0),
    .q(cnt[7]));  // sources/rtl/camera_init.v(389)
  reg_ar_as_w1 reg4_b0 (
    .clk(clk),
    .d(n0[0]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(divider2[0]));  // sources/rtl/camera_init.v(72)
  reg_ar_as_w1 reg4_b1 (
    .clk(clk),
    .d(n0[1]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(divider2[1]));  // sources/rtl/camera_init.v(72)
  reg_ar_as_w1 reg4_b2 (
    .clk(clk),
    .d(n0[2]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(divider2[2]));  // sources/rtl/camera_init.v(72)
  reg_ar_as_w1 reg4_b3 (
    .clk(clk),
    .d(n0[3]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(divider2[3]));  // sources/rtl/camera_init.v(72)
  reg_ar_as_w1 reg4_b4 (
    .clk(clk),
    .d(n0[4]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(divider2[4]));  // sources/rtl/camera_init.v(72)
  reg_ar_as_w1 reg4_b5 (
    .clk(clk),
    .d(n0[5]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(divider2[5]));  // sources/rtl/camera_init.v(72)
  reg_ar_as_w1 reg4_b6 (
    .clk(clk),
    .d(n0[6]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(divider2[6]));  // sources/rtl/camera_init.v(72)
  reg_ar_as_w1 reg4_b7 (
    .clk(clk),
    .d(n0[7]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(divider2[7]));  // sources/rtl/camera_init.v(72)
  reg_ar_as_w1 reg4_b8 (
    .clk(clk),
    .d(n0[8]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(divider2[8]));  // sources/rtl/camera_init.v(72)
  reg_ar_as_w1 reg5_b0 (
    .clk(divider2[8]),
    .d(n369[0]),
    .en(1'b1),
    .reset(1'b0),
    .set(~reset_n),
    .q(state_next[0]));  // sources/rtl/camera_init.v(311)
  reg_ar_as_w1 reg5_b1 (
    .clk(divider2[8]),
    .d(n369[1]),
    .en(1'b1),
    .reset(1'b0),
    .set(~reset_n),
    .q(state_next[1]));  // sources/rtl/camera_init.v(311)
  reg_ar_as_w1 reg5_b2 (
    .clk(divider2[8]),
    .d(n369[2]),
    .en(1'b1),
    .reset(~reset_n),
    .set(1'b0),
    .q(state_next[2]));  // sources/rtl/camera_init.v(311)
  reg_ar_as_w1 reg5_b3 (
    .clk(divider2[8]),
    .d(n369[3]),
    .en(1'b1),
    .reset(1'b0),
    .set(~reset_n),
    .q(state_next[3]));  // sources/rtl/camera_init.v(311)
  reg_ar_as_w1 reg5_b4 (
    .clk(divider2[8]),
    .d(n369[4]),
    .en(1'b1),
    .reset(~reset_n),
    .set(1'b0),
    .q(state_next[4]));  // sources/rtl/camera_init.v(311)
  reg_ar_as_w1 reg5_b5 (
    .clk(divider2[8]),
    .d(n369[5]),
    .en(1'b1),
    .reset(~reset_n),
    .set(1'b0),
    .q(n369[5]));  // sources/rtl/camera_init.v(311)
  reg_ar_as_w1 reg5_b6 (
    .clk(divider2[8]),
    .d(n369[6]),
    .en(1'b1),
    .reset(~reset_n),
    .set(1'b0),
    .q(n369[6]));  // sources/rtl/camera_init.v(311)
  reg_ar_as_w1 reg5_b7 (
    .clk(divider2[8]),
    .d(n369[7]),
    .en(1'b1),
    .reset(~reset_n),
    .set(1'b0),
    .q(n369[7]));  // sources/rtl/camera_init.v(311)
  i2c_module u_i2c_write (
    .address({1'b0,reg_address[1:0]}),
    .clk(clk),
    .reset_n(reset_n),
    .sda_in(sda_in),
    .write(bus_write),
    .writedata(data_in_bus),
    .ready(ready_out),
    .scl_out(scl),
    .sda(sda),
    .sda_oe(sda_oe),
    .success_out(success_out));  // sources/rtl/camera_init.v(48)

endmodule 

module reg_ar_as_w1
  (
  clk,
  d,
  en,
  reset,
  set,
  q
  );

  input clk;
  input d;
  input en;
  input reset;
  input set;
  output q;

  parameter REGSET = "RESET";
  wire enout;

  AL_MUX u_en0 (
    .i0(q),
    .i1(d),
    .sel(en),
    .o(enout));
  AL_DFF #(
    .INI((REGSET == "SET") ? 1'b1 : 1'b0))
    u_seq0 (
    .clk(clk),
    .d(enout),
    .reset(reset),
    .set(set),
    .q(q));

endmodule 

module \lcd_sync(IMG_Y=1)   // sources/rtl/lcd_sync.v(14)
  (
  clk,
  rest_n,
  addr,
  hsync_cnt,
  img_ack,
  lcd_clk,
  lcd_de,
  lcd_hsync,
  lcd_pwm,
  lcd_vsync,
  vsync_cnt
  );

  input clk;  // sources/rtl/lcd_sync.v(23)
  input rest_n;  // sources/rtl/lcd_sync.v(24)
  output [15:0] addr;  // sources/rtl/lcd_sync.v(33)
  output [10:0] hsync_cnt;  // sources/rtl/lcd_sync.v(30)
  output img_ack;  // sources/rtl/lcd_sync.v(32)
  output lcd_clk;  // sources/rtl/lcd_sync.v(25)
  output lcd_de;  // sources/rtl/lcd_sync.v(29)
  output lcd_hsync;  // sources/rtl/lcd_sync.v(27)
  output lcd_pwm;  // sources/rtl/lcd_sync.v(26)
  output lcd_vsync;  // sources/rtl/lcd_sync.v(28)
  output [10:0] vsync_cnt;  // sources/rtl/lcd_sync.v(31)

  parameter IMG_H = 164;
  parameter IMG_W = 200;
  parameter IMG_X = 0;
  parameter IMG_Y = 1;
  // localparam TFT_H = 640;
  // localparam TFT_V = 480;
  // localparam TH = 800;
  // localparam THB = 160;
  // localparam TV = 525;
  // localparam TVB = 45;
  wire [10:0] n10;
  wire [10:0] n2;
  wire [11:0] n24;
  wire [12:0] n28;
  wire [6:0] n29;
  wire [10:0] n3;
  wire [10:0] n30;
  wire [39:0] n32;
  wire [15:0] n34;
  wire [10:0] n8;
  wire _al_u25_o;
  wire _al_u26_o;
  wire _al_u27_o;
  wire _al_u40_o;
  wire _al_u41_o;
  wire _al_u42_o;
  wire \add0/c0 ;
  wire \add0/c1 ;
  wire \add0/c10 ;
  wire \add0/c2 ;
  wire \add0/c3 ;
  wire \add0/c4 ;
  wire \add0/c5 ;
  wire \add0/c6 ;
  wire \add0/c7 ;
  wire \add0/c8 ;
  wire \add0/c9 ;
  wire \add1/c0 ;
  wire \add1/c1 ;
  wire \add1/c10 ;
  wire \add1/c2 ;
  wire \add1/c3 ;
  wire \add1/c4 ;
  wire \add1/c5 ;
  wire \add1/c6 ;
  wire \add1/c7 ;
  wire \add1/c8 ;
  wire \add1/c9 ;
  wire lt0_c0;
  wire lt0_c1;
  wire lt0_c10;
  wire lt0_c11;
  wire lt0_c2;
  wire lt0_c3;
  wire lt0_c4;
  wire lt0_c5;
  wire lt0_c6;
  wire lt0_c7;
  wire lt0_c8;
  wire lt0_c9;
  wire lt10_2_c0;
  wire lt10_2_c1;
  wire lt10_2_c10;
  wire lt10_2_c11;
  wire lt10_2_c12;
  wire lt10_2_c2;
  wire lt10_2_c3;
  wire lt10_2_c4;
  wire lt10_2_c5;
  wire lt10_2_c6;
  wire lt10_2_c7;
  wire lt10_2_c8;
  wire lt10_2_c9;
  wire lt1_c0;
  wire lt1_c1;
  wire lt1_c10;
  wire lt1_c11;
  wire lt1_c2;
  wire lt1_c3;
  wire lt1_c4;
  wire lt1_c5;
  wire lt1_c6;
  wire lt1_c7;
  wire lt1_c8;
  wire lt1_c9;
  wire lt2_c0;
  wire lt2_c1;
  wire lt2_c10;
  wire lt2_c11;
  wire lt2_c2;
  wire lt2_c3;
  wire lt2_c4;
  wire lt2_c5;
  wire lt2_c6;
  wire lt2_c7;
  wire lt2_c8;
  wire lt2_c9;
  wire lt3_c0;
  wire lt3_c1;
  wire lt3_c10;
  wire lt3_c11;
  wire lt3_c2;
  wire lt3_c3;
  wire lt3_c4;
  wire lt3_c5;
  wire lt3_c6;
  wire lt3_c7;
  wire lt3_c8;
  wire lt3_c9;
  wire lt4_c0;
  wire lt4_c1;
  wire lt4_c10;
  wire lt4_c11;
  wire lt4_c2;
  wire lt4_c3;
  wire lt4_c4;
  wire lt4_c5;
  wire lt4_c6;
  wire lt4_c7;
  wire lt4_c8;
  wire lt4_c9;
  wire lt5_c0;
  wire lt5_c1;
  wire lt5_c10;
  wire lt5_c11;
  wire lt5_c2;
  wire lt5_c3;
  wire lt5_c4;
  wire lt5_c5;
  wire lt5_c6;
  wire lt5_c7;
  wire lt5_c8;
  wire lt5_c9;
  wire lt6_c0;
  wire lt6_c1;
  wire lt6_c10;
  wire lt6_c11;
  wire lt6_c2;
  wire lt6_c3;
  wire lt6_c4;
  wire lt6_c5;
  wire lt6_c6;
  wire lt6_c7;
  wire lt6_c8;
  wire lt6_c9;
  wire lt7_c0;
  wire lt7_c1;
  wire lt7_c10;
  wire lt7_c11;
  wire lt7_c2;
  wire lt7_c3;
  wire lt7_c4;
  wire lt7_c5;
  wire lt7_c6;
  wire lt7_c7;
  wire lt7_c8;
  wire lt7_c9;
  wire lt8_2_c0;
  wire lt8_2_c1;
  wire lt8_2_c10;
  wire lt8_2_c11;
  wire lt8_2_c12;
  wire lt8_2_c2;
  wire lt8_2_c3;
  wire lt8_2_c4;
  wire lt8_2_c5;
  wire lt8_2_c6;
  wire lt8_2_c7;
  wire lt8_2_c8;
  wire lt8_2_c9;
  wire lt9_2_c0;
  wire lt9_2_c1;
  wire lt9_2_c10;
  wire lt9_2_c11;
  wire lt9_2_c12;
  wire lt9_2_c2;
  wire lt9_2_c3;
  wire lt9_2_c4;
  wire lt9_2_c5;
  wire lt9_2_c6;
  wire lt9_2_c7;
  wire lt9_2_c8;
  wire lt9_2_c9;
  wire n11;
  wire n12;
  wire n13;
  wire n14;
  wire n15;
  wire n16;
  wire n18;
  wire n1_lutinv;
  wire n20;
  wire n22;
  wire n25;
  wire n26;
  wire n4_lutinv;
  wire \sub0/c0 ;
  wire \sub0/c1 ;
  wire \sub0/c2 ;
  wire \sub0/c3 ;
  wire \sub0/c4 ;
  wire \sub0/c5 ;
  wire \sub0/c6 ;
  wire \sub1/c0 ;
  wire \sub1/c1 ;
  wire \sub1/c10 ;
  wire \sub1/c11 ;
  wire \sub1/c2 ;
  wire \sub1/c3 ;
  wire \sub1/c4 ;
  wire \sub1/c5 ;
  wire \sub1/c6 ;
  wire \sub1/c7 ;
  wire \sub1/c8 ;
  wire \sub1/c9 ;
  wire \sub4_sub5/c0 ;
  wire \sub4_sub5/c1 ;
  wire \sub4_sub5/c10 ;
  wire \sub4_sub5/c2 ;
  wire \sub4_sub5/c3 ;
  wire \sub4_sub5/c4 ;
  wire \sub4_sub5/c5 ;
  wire \sub4_sub5/c6 ;
  wire \sub4_sub5/c7 ;
  wire \sub4_sub5/c8 ;
  wire \sub4_sub5/c9 ;
  wire \u2/c0 ;
  wire \u2/c1 ;
  wire \u2/c10 ;
  wire \u2/c11 ;
  wire \u2/c12 ;
  wire \u2/c2 ;
  wire \u2/c3 ;
  wire \u2/c4 ;
  wire \u2/c5 ;
  wire \u2/c6 ;
  wire \u2/c7 ;
  wire \u2/c8 ;
  wire \u2/c9 ;

  assign lcd_pwm = rest_n;
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u10 (
    .a(img_ack),
    .b(n28[5]),
    .o(n34[8]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u11 (
    .a(img_ack),
    .b(n28[4]),
    .o(n34[7]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u12 (
    .a(img_ack),
    .b(n28[3]),
    .o(n34[6]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u13 (
    .a(img_ack),
    .b(n28[2]),
    .o(n34[5]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u14 (
    .a(img_ack),
    .b(n28[1]),
    .o(n34[4]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u15 (
    .a(img_ack),
    .b(n28[0]),
    .o(n34[3]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u16 (
    .a(img_ack),
    .b(hsync_cnt[2]),
    .o(n34[2]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u17 (
    .a(img_ack),
    .b(n28[12]),
    .o(n34[15]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u18 (
    .a(img_ack),
    .b(n28[11]),
    .o(n34[14]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u19 (
    .a(img_ack),
    .b(n28[10]),
    .o(n34[13]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u20 (
    .a(img_ack),
    .b(n28[9]),
    .o(n34[12]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u21 (
    .a(img_ack),
    .b(n28[8]),
    .o(n34[11]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u22 (
    .a(img_ack),
    .b(n28[7]),
    .o(n34[10]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u23 (
    .a(img_ack),
    .b(hsync_cnt[1]),
    .o(n34[1]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u24 (
    .a(img_ack),
    .b(hsync_cnt[0]),
    .o(n34[0]));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    _al_u25 (
    .a(hsync_cnt[7]),
    .b(hsync_cnt[8]),
    .c(hsync_cnt[9]),
    .o(_al_u25_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*~B*~A)"),
    .INIT(16'h0010))
    _al_u26 (
    .a(hsync_cnt[3]),
    .b(hsync_cnt[4]),
    .c(hsync_cnt[5]),
    .d(hsync_cnt[6]),
    .o(_al_u26_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u27 (
    .a(hsync_cnt[0]),
    .b(hsync_cnt[1]),
    .c(hsync_cnt[10]),
    .d(hsync_cnt[2]),
    .o(_al_u27_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u28 (
    .a(_al_u25_o),
    .b(_al_u26_o),
    .c(_al_u27_o),
    .o(n1_lutinv));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u29 (
    .a(n1_lutinv),
    .b(n2[9]),
    .o(n3[9]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u30 (
    .a(n1_lutinv),
    .b(n2[8]),
    .o(n3[8]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u31 (
    .a(n1_lutinv),
    .b(n2[7]),
    .o(n3[7]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u32 (
    .a(n1_lutinv),
    .b(n2[6]),
    .o(n3[6]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u33 (
    .a(n1_lutinv),
    .b(n2[5]),
    .o(n3[5]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u34 (
    .a(n1_lutinv),
    .b(n2[4]),
    .o(n3[4]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u35 (
    .a(n1_lutinv),
    .b(n2[3]),
    .o(n3[3]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u36 (
    .a(n1_lutinv),
    .b(n2[2]),
    .o(n3[2]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u37 (
    .a(n1_lutinv),
    .b(n2[10]),
    .o(n3[10]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u38 (
    .a(n1_lutinv),
    .b(n2[1]),
    .o(n3[1]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u39 (
    .a(n1_lutinv),
    .b(n2[0]),
    .o(n3[0]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u4 (
    .a(n11),
    .b(n12),
    .o(lcd_hsync));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    _al_u40 (
    .a(vsync_cnt[7]),
    .b(vsync_cnt[8]),
    .c(vsync_cnt[9]),
    .o(_al_u40_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*A)"),
    .INIT(16'h0002))
    _al_u41 (
    .a(vsync_cnt[3]),
    .b(vsync_cnt[4]),
    .c(vsync_cnt[5]),
    .d(vsync_cnt[6]),
    .o(_al_u41_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*A)"),
    .INIT(16'h0200))
    _al_u42 (
    .a(vsync_cnt[0]),
    .b(vsync_cnt[1]),
    .c(vsync_cnt[10]),
    .d(vsync_cnt[2]),
    .o(_al_u42_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u43 (
    .a(_al_u40_o),
    .b(_al_u41_o),
    .c(_al_u42_o),
    .o(n4_lutinv));
  AL_MAP_LUT4 #(
    .EQN("(D*~((C*~B))*~(A)+D*(C*~B)*~(A)+~(D)*(C*~B)*A+D*(C*~B)*A)"),
    .INIT(16'h7520))
    _al_u44 (
    .a(n1_lutinv),
    .b(n4_lutinv),
    .c(n8[9]),
    .d(vsync_cnt[9]),
    .o(n10[9]));
  AL_MAP_LUT4 #(
    .EQN("(D*~((C*~B))*~(A)+D*(C*~B)*~(A)+~(D)*(C*~B)*A+D*(C*~B)*A)"),
    .INIT(16'h7520))
    _al_u45 (
    .a(n1_lutinv),
    .b(n4_lutinv),
    .c(n8[8]),
    .d(vsync_cnt[8]),
    .o(n10[8]));
  AL_MAP_LUT4 #(
    .EQN("(D*~((C*~B))*~(A)+D*(C*~B)*~(A)+~(D)*(C*~B)*A+D*(C*~B)*A)"),
    .INIT(16'h7520))
    _al_u46 (
    .a(n1_lutinv),
    .b(n4_lutinv),
    .c(n8[7]),
    .d(vsync_cnt[7]),
    .o(n10[7]));
  AL_MAP_LUT4 #(
    .EQN("(D*~((C*~B))*~(A)+D*(C*~B)*~(A)+~(D)*(C*~B)*A+D*(C*~B)*A)"),
    .INIT(16'h7520))
    _al_u47 (
    .a(n1_lutinv),
    .b(n4_lutinv),
    .c(n8[6]),
    .d(vsync_cnt[6]),
    .o(n10[6]));
  AL_MAP_LUT4 #(
    .EQN("(D*~((C*~B))*~(A)+D*(C*~B)*~(A)+~(D)*(C*~B)*A+D*(C*~B)*A)"),
    .INIT(16'h7520))
    _al_u48 (
    .a(n1_lutinv),
    .b(n4_lutinv),
    .c(n8[5]),
    .d(vsync_cnt[5]),
    .o(n10[5]));
  AL_MAP_LUT4 #(
    .EQN("(D*~((C*~B))*~(A)+D*(C*~B)*~(A)+~(D)*(C*~B)*A+D*(C*~B)*A)"),
    .INIT(16'h7520))
    _al_u49 (
    .a(n1_lutinv),
    .b(n4_lutinv),
    .c(n8[4]),
    .d(vsync_cnt[4]),
    .o(n10[4]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u5 (
    .a(n13),
    .b(n14),
    .o(lcd_vsync));
  AL_MAP_LUT4 #(
    .EQN("(D*~((C*~B))*~(A)+D*(C*~B)*~(A)+~(D)*(C*~B)*A+D*(C*~B)*A)"),
    .INIT(16'h7520))
    _al_u50 (
    .a(n1_lutinv),
    .b(n4_lutinv),
    .c(n8[3]),
    .d(vsync_cnt[3]),
    .o(n10[3]));
  AL_MAP_LUT4 #(
    .EQN("(D*~((C*~B))*~(A)+D*(C*~B)*~(A)+~(D)*(C*~B)*A+D*(C*~B)*A)"),
    .INIT(16'h7520))
    _al_u51 (
    .a(n1_lutinv),
    .b(n4_lutinv),
    .c(n8[2]),
    .d(vsync_cnt[2]),
    .o(n10[2]));
  AL_MAP_LUT4 #(
    .EQN("(D*~((C*~B))*~(A)+D*(C*~B)*~(A)+~(D)*(C*~B)*A+D*(C*~B)*A)"),
    .INIT(16'h7520))
    _al_u52 (
    .a(n1_lutinv),
    .b(n4_lutinv),
    .c(n8[10]),
    .d(vsync_cnt[10]),
    .o(n10[10]));
  AL_MAP_LUT4 #(
    .EQN("(D*~((C*~B))*~(A)+D*(C*~B)*~(A)+~(D)*(C*~B)*A+D*(C*~B)*A)"),
    .INIT(16'h7520))
    _al_u53 (
    .a(n1_lutinv),
    .b(n4_lutinv),
    .c(n8[1]),
    .d(vsync_cnt[1]),
    .o(n10[1]));
  AL_MAP_LUT4 #(
    .EQN("(D*~((C*~B))*~(A)+D*(C*~B)*~(A)+~(D)*(C*~B)*A+D*(C*~B)*A)"),
    .INIT(16'h7520))
    _al_u54 (
    .a(n1_lutinv),
    .b(n4_lutinv),
    .c(n8[0]),
    .d(vsync_cnt[0]),
    .o(n10[0]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u6 (
    .a(clk),
    .b(lcd_pwm),
    .o(lcd_clk));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u7 (
    .a(n15),
    .b(n16),
    .c(n18),
    .d(n20),
    .o(lcd_de));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u8 (
    .a(lcd_de),
    .b(n26),
    .c(n22),
    .d(n25),
    .o(img_ack));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u9 (
    .a(img_ack),
    .b(n28[6]),
    .o(n34[9]));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add0/u0  (
    .a(hsync_cnt[0]),
    .b(1'b1),
    .c(\add0/c0 ),
    .o({\add0/c1 ,n2[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add0/u1  (
    .a(hsync_cnt[1]),
    .b(1'b0),
    .c(\add0/c1 ),
    .o({\add0/c2 ,n2[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add0/u10  (
    .a(hsync_cnt[10]),
    .b(1'b0),
    .c(\add0/c10 ),
    .o({open_n0,n2[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add0/u2  (
    .a(hsync_cnt[2]),
    .b(1'b0),
    .c(\add0/c2 ),
    .o({\add0/c3 ,n2[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add0/u3  (
    .a(hsync_cnt[3]),
    .b(1'b0),
    .c(\add0/c3 ),
    .o({\add0/c4 ,n2[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add0/u4  (
    .a(hsync_cnt[4]),
    .b(1'b0),
    .c(\add0/c4 ),
    .o({\add0/c5 ,n2[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add0/u5  (
    .a(hsync_cnt[5]),
    .b(1'b0),
    .c(\add0/c5 ),
    .o({\add0/c6 ,n2[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add0/u6  (
    .a(hsync_cnt[6]),
    .b(1'b0),
    .c(\add0/c6 ),
    .o({\add0/c7 ,n2[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add0/u7  (
    .a(hsync_cnt[7]),
    .b(1'b0),
    .c(\add0/c7 ),
    .o({\add0/c8 ,n2[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add0/u8  (
    .a(hsync_cnt[8]),
    .b(1'b0),
    .c(\add0/c8 ),
    .o({\add0/c9 ,n2[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add0/u9  (
    .a(hsync_cnt[9]),
    .b(1'b0),
    .c(\add0/c9 ),
    .o({\add0/c10 ,n2[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \add0/ucin  (
    .a(1'b0),
    .o({\add0/c0 ,open_n3}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add1/u0  (
    .a(vsync_cnt[0]),
    .b(1'b1),
    .c(\add1/c0 ),
    .o({\add1/c1 ,n8[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add1/u1  (
    .a(vsync_cnt[1]),
    .b(1'b0),
    .c(\add1/c1 ),
    .o({\add1/c2 ,n8[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add1/u10  (
    .a(vsync_cnt[10]),
    .b(1'b0),
    .c(\add1/c10 ),
    .o({open_n4,n8[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add1/u2  (
    .a(vsync_cnt[2]),
    .b(1'b0),
    .c(\add1/c2 ),
    .o({\add1/c3 ,n8[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add1/u3  (
    .a(vsync_cnt[3]),
    .b(1'b0),
    .c(\add1/c3 ),
    .o({\add1/c4 ,n8[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add1/u4  (
    .a(vsync_cnt[4]),
    .b(1'b0),
    .c(\add1/c4 ),
    .o({\add1/c5 ,n8[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add1/u5  (
    .a(vsync_cnt[5]),
    .b(1'b0),
    .c(\add1/c5 ),
    .o({\add1/c6 ,n8[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add1/u6  (
    .a(vsync_cnt[6]),
    .b(1'b0),
    .c(\add1/c6 ),
    .o({\add1/c7 ,n8[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add1/u7  (
    .a(vsync_cnt[7]),
    .b(1'b0),
    .c(\add1/c7 ),
    .o({\add1/c8 ,n8[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add1/u8  (
    .a(vsync_cnt[8]),
    .b(1'b0),
    .c(\add1/c8 ),
    .o({\add1/c9 ,n8[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add1/u9  (
    .a(vsync_cnt[9]),
    .b(1'b0),
    .c(\add1/c9 ),
    .o({\add1/c10 ,n8[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \add1/ucin  (
    .a(1'b0),
    .o({\add1/c0 ,open_n7}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt0_0 (
    .a(1'b0),
    .b(hsync_cnt[0]),
    .c(lt0_c0),
    .o({lt0_c1,open_n8}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt0_1 (
    .a(1'b0),
    .b(hsync_cnt[1]),
    .c(lt0_c1),
    .o({lt0_c2,open_n9}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt0_10 (
    .a(1'b0),
    .b(hsync_cnt[10]),
    .c(lt0_c10),
    .o({lt0_c11,open_n10}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt0_2 (
    .a(1'b0),
    .b(hsync_cnt[2]),
    .c(lt0_c2),
    .o({lt0_c3,open_n11}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt0_3 (
    .a(1'b0),
    .b(hsync_cnt[3]),
    .c(lt0_c3),
    .o({lt0_c4,open_n12}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt0_4 (
    .a(1'b1),
    .b(hsync_cnt[4]),
    .c(lt0_c4),
    .o({lt0_c5,open_n13}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt0_5 (
    .a(1'b0),
    .b(hsync_cnt[5]),
    .c(lt0_c5),
    .o({lt0_c6,open_n14}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt0_6 (
    .a(1'b0),
    .b(hsync_cnt[6]),
    .c(lt0_c6),
    .o({lt0_c7,open_n15}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt0_7 (
    .a(1'b0),
    .b(hsync_cnt[7]),
    .c(lt0_c7),
    .o({lt0_c8,open_n16}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt0_8 (
    .a(1'b0),
    .b(hsync_cnt[8]),
    .c(lt0_c8),
    .o({lt0_c9,open_n17}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt0_9 (
    .a(1'b0),
    .b(hsync_cnt[9]),
    .c(lt0_c9),
    .o({lt0_c10,open_n18}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    lt0_cin (
    .a(1'b1),
    .o({lt0_c0,open_n21}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt0_cout (
    .a(1'b0),
    .b(1'b1),
    .c(lt0_c11),
    .o({open_n22,n11}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt10_2_0 (
    .a(n24[0]),
    .b(1'b1),
    .c(lt10_2_c0),
    .o({lt10_2_c1,open_n23}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt10_2_1 (
    .a(n24[1]),
    .b(1'b0),
    .c(lt10_2_c1),
    .o({lt10_2_c2,open_n24}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt10_2_10 (
    .a(n24[10]),
    .b(1'b0),
    .c(lt10_2_c10),
    .o({lt10_2_c11,open_n25}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt10_2_11 (
    .a(n24[11]),
    .b(1'b0),
    .c(lt10_2_c11),
    .o({lt10_2_c12,open_n26}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt10_2_2 (
    .a(n24[2]),
    .b(1'b1),
    .c(lt10_2_c2),
    .o({lt10_2_c3,open_n27}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt10_2_3 (
    .a(n24[3]),
    .b(1'b0),
    .c(lt10_2_c3),
    .o({lt10_2_c4,open_n28}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt10_2_4 (
    .a(n24[4]),
    .b(1'b0),
    .c(lt10_2_c4),
    .o({lt10_2_c5,open_n29}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt10_2_5 (
    .a(n24[5]),
    .b(1'b1),
    .c(lt10_2_c5),
    .o({lt10_2_c6,open_n30}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt10_2_6 (
    .a(n24[6]),
    .b(1'b0),
    .c(lt10_2_c6),
    .o({lt10_2_c7,open_n31}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt10_2_7 (
    .a(n24[7]),
    .b(1'b1),
    .c(lt10_2_c7),
    .o({lt10_2_c8,open_n32}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt10_2_8 (
    .a(n24[8]),
    .b(1'b0),
    .c(lt10_2_c8),
    .o({lt10_2_c9,open_n33}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt10_2_9 (
    .a(n24[9]),
    .b(1'b0),
    .c(lt10_2_c9),
    .o({lt10_2_c10,open_n34}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    lt10_2_cin (
    .a(1'b0),
    .o({lt10_2_c0,open_n37}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt10_2_cout (
    .a(1'b0),
    .b(1'b1),
    .c(lt10_2_c12),
    .o({open_n38,n26}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt1_0 (
    .a(hsync_cnt[0]),
    .b(1'b0),
    .c(lt1_c0),
    .o({lt1_c1,open_n39}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt1_1 (
    .a(hsync_cnt[1]),
    .b(1'b0),
    .c(lt1_c1),
    .o({lt1_c2,open_n40}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt1_10 (
    .a(hsync_cnt[10]),
    .b(1'b0),
    .c(lt1_c10),
    .o({lt1_c11,open_n41}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt1_2 (
    .a(hsync_cnt[2]),
    .b(1'b0),
    .c(lt1_c2),
    .o({lt1_c3,open_n42}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt1_3 (
    .a(hsync_cnt[3]),
    .b(1'b0),
    .c(lt1_c3),
    .o({lt1_c4,open_n43}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt1_4 (
    .a(hsync_cnt[4]),
    .b(1'b1),
    .c(lt1_c4),
    .o({lt1_c5,open_n44}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt1_5 (
    .a(hsync_cnt[5]),
    .b(1'b1),
    .c(lt1_c5),
    .o({lt1_c6,open_n45}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt1_6 (
    .a(hsync_cnt[6]),
    .b(1'b1),
    .c(lt1_c6),
    .o({lt1_c7,open_n46}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt1_7 (
    .a(hsync_cnt[7]),
    .b(1'b0),
    .c(lt1_c7),
    .o({lt1_c8,open_n47}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt1_8 (
    .a(hsync_cnt[8]),
    .b(1'b0),
    .c(lt1_c8),
    .o({lt1_c9,open_n48}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt1_9 (
    .a(hsync_cnt[9]),
    .b(1'b0),
    .c(lt1_c9),
    .o({lt1_c10,open_n49}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    lt1_cin (
    .a(1'b0),
    .o({lt1_c0,open_n52}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt1_cout (
    .a(1'b0),
    .b(1'b1),
    .c(lt1_c11),
    .o({open_n53,n12}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt2_0 (
    .a(1'b0),
    .b(vsync_cnt[0]),
    .c(lt2_c0),
    .o({lt2_c1,open_n54}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt2_1 (
    .a(1'b1),
    .b(vsync_cnt[1]),
    .c(lt2_c1),
    .o({lt2_c2,open_n55}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt2_10 (
    .a(1'b0),
    .b(vsync_cnt[10]),
    .c(lt2_c10),
    .o({lt2_c11,open_n56}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt2_2 (
    .a(1'b0),
    .b(vsync_cnt[2]),
    .c(lt2_c2),
    .o({lt2_c3,open_n57}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt2_3 (
    .a(1'b1),
    .b(vsync_cnt[3]),
    .c(lt2_c3),
    .o({lt2_c4,open_n58}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt2_4 (
    .a(1'b0),
    .b(vsync_cnt[4]),
    .c(lt2_c4),
    .o({lt2_c5,open_n59}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt2_5 (
    .a(1'b0),
    .b(vsync_cnt[5]),
    .c(lt2_c5),
    .o({lt2_c6,open_n60}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt2_6 (
    .a(1'b0),
    .b(vsync_cnt[6]),
    .c(lt2_c6),
    .o({lt2_c7,open_n61}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt2_7 (
    .a(1'b0),
    .b(vsync_cnt[7]),
    .c(lt2_c7),
    .o({lt2_c8,open_n62}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt2_8 (
    .a(1'b0),
    .b(vsync_cnt[8]),
    .c(lt2_c8),
    .o({lt2_c9,open_n63}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt2_9 (
    .a(1'b0),
    .b(vsync_cnt[9]),
    .c(lt2_c9),
    .o({lt2_c10,open_n64}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    lt2_cin (
    .a(1'b1),
    .o({lt2_c0,open_n67}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt2_cout (
    .a(1'b0),
    .b(1'b1),
    .c(lt2_c11),
    .o({open_n68,n13}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt3_0 (
    .a(vsync_cnt[0]),
    .b(1'b0),
    .c(lt3_c0),
    .o({lt3_c1,open_n69}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt3_1 (
    .a(vsync_cnt[1]),
    .b(1'b0),
    .c(lt3_c1),
    .o({lt3_c2,open_n70}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt3_10 (
    .a(vsync_cnt[10]),
    .b(1'b0),
    .c(lt3_c10),
    .o({lt3_c11,open_n71}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt3_2 (
    .a(vsync_cnt[2]),
    .b(1'b1),
    .c(lt3_c2),
    .o({lt3_c3,open_n72}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt3_3 (
    .a(vsync_cnt[3]),
    .b(1'b1),
    .c(lt3_c3),
    .o({lt3_c4,open_n73}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt3_4 (
    .a(vsync_cnt[4]),
    .b(1'b0),
    .c(lt3_c4),
    .o({lt3_c5,open_n74}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt3_5 (
    .a(vsync_cnt[5]),
    .b(1'b0),
    .c(lt3_c5),
    .o({lt3_c6,open_n75}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt3_6 (
    .a(vsync_cnt[6]),
    .b(1'b0),
    .c(lt3_c6),
    .o({lt3_c7,open_n76}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt3_7 (
    .a(vsync_cnt[7]),
    .b(1'b0),
    .c(lt3_c7),
    .o({lt3_c8,open_n77}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt3_8 (
    .a(vsync_cnt[8]),
    .b(1'b0),
    .c(lt3_c8),
    .o({lt3_c9,open_n78}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt3_9 (
    .a(vsync_cnt[9]),
    .b(1'b0),
    .c(lt3_c9),
    .o({lt3_c10,open_n79}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    lt3_cin (
    .a(1'b0),
    .o({lt3_c0,open_n82}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt3_cout (
    .a(1'b0),
    .b(1'b1),
    .c(lt3_c11),
    .o({open_n83,n14}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt4_0 (
    .a(1'b0),
    .b(hsync_cnt[0]),
    .c(lt4_c0),
    .o({lt4_c1,open_n84}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt4_1 (
    .a(1'b0),
    .b(hsync_cnt[1]),
    .c(lt4_c1),
    .o({lt4_c2,open_n85}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt4_10 (
    .a(1'b0),
    .b(hsync_cnt[10]),
    .c(lt4_c10),
    .o({lt4_c11,open_n86}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt4_2 (
    .a(1'b0),
    .b(hsync_cnt[2]),
    .c(lt4_c2),
    .o({lt4_c3,open_n87}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt4_3 (
    .a(1'b0),
    .b(hsync_cnt[3]),
    .c(lt4_c3),
    .o({lt4_c4,open_n88}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt4_4 (
    .a(1'b0),
    .b(hsync_cnt[4]),
    .c(lt4_c4),
    .o({lt4_c5,open_n89}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt4_5 (
    .a(1'b1),
    .b(hsync_cnt[5]),
    .c(lt4_c5),
    .o({lt4_c6,open_n90}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt4_6 (
    .a(1'b0),
    .b(hsync_cnt[6]),
    .c(lt4_c6),
    .o({lt4_c7,open_n91}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt4_7 (
    .a(1'b1),
    .b(hsync_cnt[7]),
    .c(lt4_c7),
    .o({lt4_c8,open_n92}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt4_8 (
    .a(1'b0),
    .b(hsync_cnt[8]),
    .c(lt4_c8),
    .o({lt4_c9,open_n93}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt4_9 (
    .a(1'b0),
    .b(hsync_cnt[9]),
    .c(lt4_c9),
    .o({lt4_c10,open_n94}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    lt4_cin (
    .a(1'b1),
    .o({lt4_c0,open_n97}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt4_cout (
    .a(1'b0),
    .b(1'b1),
    .c(lt4_c11),
    .o({open_n98,n15}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt5_0 (
    .a(hsync_cnt[0]),
    .b(1'b0),
    .c(lt5_c0),
    .o({lt5_c1,open_n99}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt5_1 (
    .a(hsync_cnt[1]),
    .b(1'b0),
    .c(lt5_c1),
    .o({lt5_c2,open_n100}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt5_10 (
    .a(hsync_cnt[10]),
    .b(1'b0),
    .c(lt5_c10),
    .o({lt5_c11,open_n101}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt5_2 (
    .a(hsync_cnt[2]),
    .b(1'b0),
    .c(lt5_c2),
    .o({lt5_c3,open_n102}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt5_3 (
    .a(hsync_cnt[3]),
    .b(1'b0),
    .c(lt5_c3),
    .o({lt5_c4,open_n103}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt5_4 (
    .a(hsync_cnt[4]),
    .b(1'b0),
    .c(lt5_c4),
    .o({lt5_c5,open_n104}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt5_5 (
    .a(hsync_cnt[5]),
    .b(1'b1),
    .c(lt5_c5),
    .o({lt5_c6,open_n105}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt5_6 (
    .a(hsync_cnt[6]),
    .b(1'b0),
    .c(lt5_c6),
    .o({lt5_c7,open_n106}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt5_7 (
    .a(hsync_cnt[7]),
    .b(1'b0),
    .c(lt5_c7),
    .o({lt5_c8,open_n107}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt5_8 (
    .a(hsync_cnt[8]),
    .b(1'b1),
    .c(lt5_c8),
    .o({lt5_c9,open_n108}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt5_9 (
    .a(hsync_cnt[9]),
    .b(1'b1),
    .c(lt5_c9),
    .o({lt5_c10,open_n109}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    lt5_cin (
    .a(1'b1),
    .o({lt5_c0,open_n112}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt5_cout (
    .a(1'b0),
    .b(1'b1),
    .c(lt5_c11),
    .o({open_n113,n16}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt6_0 (
    .a(1'b1),
    .b(vsync_cnt[0]),
    .c(lt6_c0),
    .o({lt6_c1,open_n114}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt6_1 (
    .a(1'b0),
    .b(vsync_cnt[1]),
    .c(lt6_c1),
    .o({lt6_c2,open_n115}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt6_10 (
    .a(1'b0),
    .b(vsync_cnt[10]),
    .c(lt6_c10),
    .o({lt6_c11,open_n116}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt6_2 (
    .a(1'b1),
    .b(vsync_cnt[2]),
    .c(lt6_c2),
    .o({lt6_c3,open_n117}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt6_3 (
    .a(1'b1),
    .b(vsync_cnt[3]),
    .c(lt6_c3),
    .o({lt6_c4,open_n118}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt6_4 (
    .a(1'b0),
    .b(vsync_cnt[4]),
    .c(lt6_c4),
    .o({lt6_c5,open_n119}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt6_5 (
    .a(1'b1),
    .b(vsync_cnt[5]),
    .c(lt6_c5),
    .o({lt6_c6,open_n120}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt6_6 (
    .a(1'b0),
    .b(vsync_cnt[6]),
    .c(lt6_c6),
    .o({lt6_c7,open_n121}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt6_7 (
    .a(1'b0),
    .b(vsync_cnt[7]),
    .c(lt6_c7),
    .o({lt6_c8,open_n122}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt6_8 (
    .a(1'b0),
    .b(vsync_cnt[8]),
    .c(lt6_c8),
    .o({lt6_c9,open_n123}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt6_9 (
    .a(1'b0),
    .b(vsync_cnt[9]),
    .c(lt6_c9),
    .o({lt6_c10,open_n124}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    lt6_cin (
    .a(1'b1),
    .o({lt6_c0,open_n127}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt6_cout (
    .a(1'b0),
    .b(1'b1),
    .c(lt6_c11),
    .o({open_n128,n18}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt7_0 (
    .a(vsync_cnt[0]),
    .b(1'b1),
    .c(lt7_c0),
    .o({lt7_c1,open_n129}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt7_1 (
    .a(vsync_cnt[1]),
    .b(1'b0),
    .c(lt7_c1),
    .o({lt7_c2,open_n130}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt7_10 (
    .a(vsync_cnt[10]),
    .b(1'b0),
    .c(lt7_c10),
    .o({lt7_c11,open_n131}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt7_2 (
    .a(vsync_cnt[2]),
    .b(1'b1),
    .c(lt7_c2),
    .o({lt7_c3,open_n132}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt7_3 (
    .a(vsync_cnt[3]),
    .b(1'b1),
    .c(lt7_c3),
    .o({lt7_c4,open_n133}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt7_4 (
    .a(vsync_cnt[4]),
    .b(1'b0),
    .c(lt7_c4),
    .o({lt7_c5,open_n134}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt7_5 (
    .a(vsync_cnt[5]),
    .b(1'b0),
    .c(lt7_c5),
    .o({lt7_c6,open_n135}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt7_6 (
    .a(vsync_cnt[6]),
    .b(1'b0),
    .c(lt7_c6),
    .o({lt7_c7,open_n136}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt7_7 (
    .a(vsync_cnt[7]),
    .b(1'b0),
    .c(lt7_c7),
    .o({lt7_c8,open_n137}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt7_8 (
    .a(vsync_cnt[8]),
    .b(1'b0),
    .c(lt7_c8),
    .o({lt7_c9,open_n138}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt7_9 (
    .a(vsync_cnt[9]),
    .b(1'b1),
    .c(lt7_c9),
    .o({lt7_c10,open_n139}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    lt7_cin (
    .a(1'b0),
    .o({lt7_c0,open_n142}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt7_cout (
    .a(1'b0),
    .b(1'b1),
    .c(lt7_c11),
    .o({open_n143,n20}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt8_2_0 (
    .a(hsync_cnt[0]),
    .b(1'b0),
    .c(lt8_2_c0),
    .o({lt8_2_c1,open_n144}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt8_2_1 (
    .a(hsync_cnt[1]),
    .b(1'b0),
    .c(lt8_2_c1),
    .o({lt8_2_c2,open_n145}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt8_2_10 (
    .a(n29[5]),
    .b(1'b0),
    .c(lt8_2_c10),
    .o({lt8_2_c11,open_n146}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt8_2_11 (
    .a(n29[6]),
    .b(1'b0),
    .c(lt8_2_c11),
    .o({lt8_2_c12,open_n147}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt8_2_2 (
    .a(hsync_cnt[2]),
    .b(1'b0),
    .c(lt8_2_c2),
    .o({lt8_2_c3,open_n148}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt8_2_3 (
    .a(hsync_cnt[3]),
    .b(1'b1),
    .c(lt8_2_c3),
    .o({lt8_2_c4,open_n149}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt8_2_4 (
    .a(hsync_cnt[4]),
    .b(1'b0),
    .c(lt8_2_c4),
    .o({lt8_2_c5,open_n150}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt8_2_5 (
    .a(n29[0]),
    .b(1'b0),
    .c(lt8_2_c5),
    .o({lt8_2_c6,open_n151}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt8_2_6 (
    .a(n29[1]),
    .b(1'b1),
    .c(lt8_2_c6),
    .o({lt8_2_c7,open_n152}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt8_2_7 (
    .a(n29[2]),
    .b(1'b1),
    .c(lt8_2_c7),
    .o({lt8_2_c8,open_n153}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt8_2_8 (
    .a(n29[3]),
    .b(1'b0),
    .c(lt8_2_c8),
    .o({lt8_2_c9,open_n154}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt8_2_9 (
    .a(n29[4]),
    .b(1'b0),
    .c(lt8_2_c9),
    .o({lt8_2_c10,open_n155}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    lt8_2_cin (
    .a(1'b0),
    .o({lt8_2_c0,open_n158}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt8_2_cout (
    .a(1'b0),
    .b(1'b1),
    .c(lt8_2_c12),
    .o({open_n159,n22}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt9_2_0 (
    .a(1'b1),
    .b(n24[0]),
    .c(lt9_2_c0),
    .o({lt9_2_c1,open_n160}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt9_2_1 (
    .a(1'b0),
    .b(n24[1]),
    .c(lt9_2_c1),
    .o({lt9_2_c2,open_n161}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt9_2_10 (
    .a(1'b0),
    .b(n24[10]),
    .c(lt9_2_c10),
    .o({lt9_2_c11,open_n162}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt9_2_11 (
    .a(1'b0),
    .b(n24[11]),
    .c(lt9_2_c11),
    .o({lt9_2_c12,open_n163}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt9_2_2 (
    .a(1'b0),
    .b(n24[2]),
    .c(lt9_2_c2),
    .o({lt9_2_c3,open_n164}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt9_2_3 (
    .a(1'b0),
    .b(n24[3]),
    .c(lt9_2_c3),
    .o({lt9_2_c4,open_n165}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt9_2_4 (
    .a(1'b0),
    .b(n24[4]),
    .c(lt9_2_c4),
    .o({lt9_2_c5,open_n166}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt9_2_5 (
    .a(1'b0),
    .b(n24[5]),
    .c(lt9_2_c5),
    .o({lt9_2_c6,open_n167}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt9_2_6 (
    .a(1'b0),
    .b(n24[6]),
    .c(lt9_2_c6),
    .o({lt9_2_c7,open_n168}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt9_2_7 (
    .a(1'b0),
    .b(n24[7]),
    .c(lt9_2_c7),
    .o({lt9_2_c8,open_n169}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt9_2_8 (
    .a(1'b0),
    .b(n24[8]),
    .c(lt9_2_c8),
    .o({lt9_2_c9,open_n170}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt9_2_9 (
    .a(1'b0),
    .b(n24[9]),
    .c(lt9_2_c9),
    .o({lt9_2_c10,open_n171}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    lt9_2_cin (
    .a(1'b1),
    .o({lt9_2_c0,open_n174}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt9_2_cout (
    .a(1'b0),
    .b(1'b1),
    .c(lt9_2_c12),
    .o({open_n175,n25}));
  EG_PHY_MULT18 #(
    .INPUTREGA("DISABLE"),
    .INPUTREGB("DISABLE"),
    .MODE("MULT18X18C"),
    .OUTPUTREG("DISABLE"),
    .SIGNEDAMUX("0"),
    .SIGNEDBMUX("0"))
    mult0_ (
    .a({5'b00000,n30[10],n30,vsync_cnt[0]}),
    .b(18'b000000000000011001),
    .p({open_n259,open_n260,open_n261,open_n262,open_n263,open_n264,open_n265,open_n266,open_n267,open_n268,open_n269,open_n270,open_n271,open_n272,open_n273,open_n274,open_n275,open_n276,open_n277,open_n278,open_n279,open_n280,open_n281,n32[15:3]}));
  reg_ar_as_w1 reg0_b0 (
    .clk(clk),
    .d(n10[0]),
    .en(1'b1),
    .reset(~lcd_pwm),
    .set(1'b0),
    .q(vsync_cnt[0]));  // sources/rtl/lcd_sync.v(71)
  reg_ar_as_w1 reg0_b1 (
    .clk(clk),
    .d(n10[1]),
    .en(1'b1),
    .reset(~lcd_pwm),
    .set(1'b0),
    .q(vsync_cnt[1]));  // sources/rtl/lcd_sync.v(71)
  reg_ar_as_w1 reg0_b10 (
    .clk(clk),
    .d(n10[10]),
    .en(1'b1),
    .reset(~lcd_pwm),
    .set(1'b0),
    .q(vsync_cnt[10]));  // sources/rtl/lcd_sync.v(71)
  reg_ar_as_w1 reg0_b2 (
    .clk(clk),
    .d(n10[2]),
    .en(1'b1),
    .reset(~lcd_pwm),
    .set(1'b0),
    .q(vsync_cnt[2]));  // sources/rtl/lcd_sync.v(71)
  reg_ar_as_w1 reg0_b3 (
    .clk(clk),
    .d(n10[3]),
    .en(1'b1),
    .reset(~lcd_pwm),
    .set(1'b0),
    .q(vsync_cnt[3]));  // sources/rtl/lcd_sync.v(71)
  reg_ar_as_w1 reg0_b4 (
    .clk(clk),
    .d(n10[4]),
    .en(1'b1),
    .reset(~lcd_pwm),
    .set(1'b0),
    .q(vsync_cnt[4]));  // sources/rtl/lcd_sync.v(71)
  reg_ar_as_w1 reg0_b5 (
    .clk(clk),
    .d(n10[5]),
    .en(1'b1),
    .reset(~lcd_pwm),
    .set(1'b0),
    .q(vsync_cnt[5]));  // sources/rtl/lcd_sync.v(71)
  reg_ar_as_w1 reg0_b6 (
    .clk(clk),
    .d(n10[6]),
    .en(1'b1),
    .reset(~lcd_pwm),
    .set(1'b0),
    .q(vsync_cnt[6]));  // sources/rtl/lcd_sync.v(71)
  reg_ar_as_w1 reg0_b7 (
    .clk(clk),
    .d(n10[7]),
    .en(1'b1),
    .reset(~lcd_pwm),
    .set(1'b0),
    .q(vsync_cnt[7]));  // sources/rtl/lcd_sync.v(71)
  reg_ar_as_w1 reg0_b8 (
    .clk(clk),
    .d(n10[8]),
    .en(1'b1),
    .reset(~lcd_pwm),
    .set(1'b0),
    .q(vsync_cnt[8]));  // sources/rtl/lcd_sync.v(71)
  reg_ar_as_w1 reg0_b9 (
    .clk(clk),
    .d(n10[9]),
    .en(1'b1),
    .reset(~lcd_pwm),
    .set(1'b0),
    .q(vsync_cnt[9]));  // sources/rtl/lcd_sync.v(71)
  reg_ar_as_w1 reg1_b0 (
    .clk(clk),
    .d(n34[0]),
    .en(1'b1),
    .reset(~lcd_pwm),
    .set(1'b0),
    .q(addr[0]));  // sources/rtl/lcd_sync.v(95)
  reg_ar_as_w1 reg1_b1 (
    .clk(clk),
    .d(n34[1]),
    .en(1'b1),
    .reset(~lcd_pwm),
    .set(1'b0),
    .q(addr[1]));  // sources/rtl/lcd_sync.v(95)
  reg_ar_as_w1 reg1_b10 (
    .clk(clk),
    .d(n34[10]),
    .en(1'b1),
    .reset(~lcd_pwm),
    .set(1'b0),
    .q(addr[10]));  // sources/rtl/lcd_sync.v(95)
  reg_ar_as_w1 reg1_b11 (
    .clk(clk),
    .d(n34[11]),
    .en(1'b1),
    .reset(~lcd_pwm),
    .set(1'b0),
    .q(addr[11]));  // sources/rtl/lcd_sync.v(95)
  reg_ar_as_w1 reg1_b12 (
    .clk(clk),
    .d(n34[12]),
    .en(1'b1),
    .reset(~lcd_pwm),
    .set(1'b0),
    .q(addr[12]));  // sources/rtl/lcd_sync.v(95)
  reg_ar_as_w1 reg1_b13 (
    .clk(clk),
    .d(n34[13]),
    .en(1'b1),
    .reset(~lcd_pwm),
    .set(1'b0),
    .q(addr[13]));  // sources/rtl/lcd_sync.v(95)
  reg_ar_as_w1 reg1_b14 (
    .clk(clk),
    .d(n34[14]),
    .en(1'b1),
    .reset(~lcd_pwm),
    .set(1'b0),
    .q(addr[14]));  // sources/rtl/lcd_sync.v(95)
  reg_ar_as_w1 reg1_b15 (
    .clk(clk),
    .d(n34[15]),
    .en(1'b1),
    .reset(~lcd_pwm),
    .set(1'b0),
    .q(addr[15]));  // sources/rtl/lcd_sync.v(95)
  reg_ar_as_w1 reg1_b2 (
    .clk(clk),
    .d(n34[2]),
    .en(1'b1),
    .reset(~lcd_pwm),
    .set(1'b0),
    .q(addr[2]));  // sources/rtl/lcd_sync.v(95)
  reg_ar_as_w1 reg1_b3 (
    .clk(clk),
    .d(n34[3]),
    .en(1'b1),
    .reset(~lcd_pwm),
    .set(1'b0),
    .q(addr[3]));  // sources/rtl/lcd_sync.v(95)
  reg_ar_as_w1 reg1_b4 (
    .clk(clk),
    .d(n34[4]),
    .en(1'b1),
    .reset(~lcd_pwm),
    .set(1'b0),
    .q(addr[4]));  // sources/rtl/lcd_sync.v(95)
  reg_ar_as_w1 reg1_b5 (
    .clk(clk),
    .d(n34[5]),
    .en(1'b1),
    .reset(~lcd_pwm),
    .set(1'b0),
    .q(addr[5]));  // sources/rtl/lcd_sync.v(95)
  reg_ar_as_w1 reg1_b6 (
    .clk(clk),
    .d(n34[6]),
    .en(1'b1),
    .reset(~lcd_pwm),
    .set(1'b0),
    .q(addr[6]));  // sources/rtl/lcd_sync.v(95)
  reg_ar_as_w1 reg1_b7 (
    .clk(clk),
    .d(n34[7]),
    .en(1'b1),
    .reset(~lcd_pwm),
    .set(1'b0),
    .q(addr[7]));  // sources/rtl/lcd_sync.v(95)
  reg_ar_as_w1 reg1_b8 (
    .clk(clk),
    .d(n34[8]),
    .en(1'b1),
    .reset(~lcd_pwm),
    .set(1'b0),
    .q(addr[8]));  // sources/rtl/lcd_sync.v(95)
  reg_ar_as_w1 reg1_b9 (
    .clk(clk),
    .d(n34[9]),
    .en(1'b1),
    .reset(~lcd_pwm),
    .set(1'b0),
    .q(addr[9]));  // sources/rtl/lcd_sync.v(95)
  reg_ar_as_w1 reg2_b0 (
    .clk(clk),
    .d(n3[0]),
    .en(1'b1),
    .reset(~lcd_pwm),
    .set(1'b0),
    .q(hsync_cnt[0]));  // sources/rtl/lcd_sync.v(61)
  reg_ar_as_w1 reg2_b1 (
    .clk(clk),
    .d(n3[1]),
    .en(1'b1),
    .reset(~lcd_pwm),
    .set(1'b0),
    .q(hsync_cnt[1]));  // sources/rtl/lcd_sync.v(61)
  reg_ar_as_w1 reg2_b10 (
    .clk(clk),
    .d(n3[10]),
    .en(1'b1),
    .reset(~lcd_pwm),
    .set(1'b0),
    .q(hsync_cnt[10]));  // sources/rtl/lcd_sync.v(61)
  reg_ar_as_w1 reg2_b2 (
    .clk(clk),
    .d(n3[2]),
    .en(1'b1),
    .reset(~lcd_pwm),
    .set(1'b0),
    .q(hsync_cnt[2]));  // sources/rtl/lcd_sync.v(61)
  reg_ar_as_w1 reg2_b3 (
    .clk(clk),
    .d(n3[3]),
    .en(1'b1),
    .reset(~lcd_pwm),
    .set(1'b0),
    .q(hsync_cnt[3]));  // sources/rtl/lcd_sync.v(61)
  reg_ar_as_w1 reg2_b4 (
    .clk(clk),
    .d(n3[4]),
    .en(1'b1),
    .reset(~lcd_pwm),
    .set(1'b0),
    .q(hsync_cnt[4]));  // sources/rtl/lcd_sync.v(61)
  reg_ar_as_w1 reg2_b5 (
    .clk(clk),
    .d(n3[5]),
    .en(1'b1),
    .reset(~lcd_pwm),
    .set(1'b0),
    .q(hsync_cnt[5]));  // sources/rtl/lcd_sync.v(61)
  reg_ar_as_w1 reg2_b6 (
    .clk(clk),
    .d(n3[6]),
    .en(1'b1),
    .reset(~lcd_pwm),
    .set(1'b0),
    .q(hsync_cnt[6]));  // sources/rtl/lcd_sync.v(61)
  reg_ar_as_w1 reg2_b7 (
    .clk(clk),
    .d(n3[7]),
    .en(1'b1),
    .reset(~lcd_pwm),
    .set(1'b0),
    .q(hsync_cnt[7]));  // sources/rtl/lcd_sync.v(61)
  reg_ar_as_w1 reg2_b8 (
    .clk(clk),
    .d(n3[8]),
    .en(1'b1),
    .reset(~lcd_pwm),
    .set(1'b0),
    .q(hsync_cnt[8]));  // sources/rtl/lcd_sync.v(61)
  reg_ar_as_w1 reg2_b9 (
    .clk(clk),
    .d(n3[9]),
    .en(1'b1),
    .reset(~lcd_pwm),
    .set(1'b0),
    .q(hsync_cnt[9]));  // sources/rtl/lcd_sync.v(61)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \sub0/u0  (
    .a(hsync_cnt[5]),
    .b(1'b1),
    .c(\sub0/c0 ),
    .o({\sub0/c1 ,n29[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \sub0/u1  (
    .a(hsync_cnt[6]),
    .b(1'b0),
    .c(\sub0/c1 ),
    .o({\sub0/c2 ,n29[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \sub0/u2  (
    .a(hsync_cnt[7]),
    .b(1'b1),
    .c(\sub0/c2 ),
    .o({\sub0/c3 ,n29[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \sub0/u3  (
    .a(hsync_cnt[8]),
    .b(1'b0),
    .c(\sub0/c3 ),
    .o({\sub0/c4 ,n29[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \sub0/u4  (
    .a(hsync_cnt[9]),
    .b(1'b0),
    .c(\sub0/c4 ),
    .o({\sub0/c5 ,n29[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \sub0/u5  (
    .a(hsync_cnt[10]),
    .b(1'b0),
    .c(\sub0/c5 ),
    .o({\sub0/c6 ,n29[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    \sub0/ucin  (
    .a(1'b0),
    .o({\sub0/c0 ,open_n284}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \sub0/ucout  (
    .c(\sub0/c6 ),
    .o({open_n287,n29[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \sub1/u0  (
    .a(vsync_cnt[0]),
    .b(1'b1),
    .c(\sub1/c0 ),
    .o({\sub1/c1 ,n24[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \sub1/u1  (
    .a(vsync_cnt[1]),
    .b(1'b0),
    .c(\sub1/c1 ),
    .o({\sub1/c2 ,n24[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \sub1/u10  (
    .a(vsync_cnt[10]),
    .b(1'b0),
    .c(\sub1/c10 ),
    .o({\sub1/c11 ,n24[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \sub1/u2  (
    .a(vsync_cnt[2]),
    .b(1'b1),
    .c(\sub1/c2 ),
    .o({\sub1/c3 ,n24[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \sub1/u3  (
    .a(vsync_cnt[3]),
    .b(1'b1),
    .c(\sub1/c3 ),
    .o({\sub1/c4 ,n24[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \sub1/u4  (
    .a(vsync_cnt[4]),
    .b(1'b0),
    .c(\sub1/c4 ),
    .o({\sub1/c5 ,n24[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \sub1/u5  (
    .a(vsync_cnt[5]),
    .b(1'b1),
    .c(\sub1/c5 ),
    .o({\sub1/c6 ,n24[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \sub1/u6  (
    .a(vsync_cnt[6]),
    .b(1'b0),
    .c(\sub1/c6 ),
    .o({\sub1/c7 ,n24[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \sub1/u7  (
    .a(vsync_cnt[7]),
    .b(1'b0),
    .c(\sub1/c7 ),
    .o({\sub1/c8 ,n24[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \sub1/u8  (
    .a(vsync_cnt[8]),
    .b(1'b0),
    .c(\sub1/c8 ),
    .o({\sub1/c9 ,n24[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \sub1/u9  (
    .a(vsync_cnt[9]),
    .b(1'b0),
    .c(\sub1/c9 ),
    .o({\sub1/c10 ,n24[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    \sub1/ucin  (
    .a(1'b0),
    .o({\sub1/c0 ,open_n290}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \sub1/ucout  (
    .c(\sub1/c11 ),
    .o({open_n293,n24[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \sub4_sub5/u0  (
    .a(vsync_cnt[1]),
    .b(1'b1),
    .c(\sub4_sub5/c0 ),
    .o({\sub4_sub5/c1 ,n30[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \sub4_sub5/u1  (
    .a(vsync_cnt[2]),
    .b(1'b1),
    .c(\sub4_sub5/c1 ),
    .o({\sub4_sub5/c2 ,n30[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \sub4_sub5/u2  (
    .a(vsync_cnt[3]),
    .b(1'b1),
    .c(\sub4_sub5/c2 ),
    .o({\sub4_sub5/c3 ,n30[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \sub4_sub5/u3  (
    .a(vsync_cnt[4]),
    .b(1'b0),
    .c(\sub4_sub5/c3 ),
    .o({\sub4_sub5/c4 ,n30[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \sub4_sub5/u4  (
    .a(vsync_cnt[5]),
    .b(1'b1),
    .c(\sub4_sub5/c4 ),
    .o({\sub4_sub5/c5 ,n30[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \sub4_sub5/u5  (
    .a(vsync_cnt[6]),
    .b(1'b0),
    .c(\sub4_sub5/c5 ),
    .o({\sub4_sub5/c6 ,n30[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \sub4_sub5/u6  (
    .a(vsync_cnt[7]),
    .b(1'b0),
    .c(\sub4_sub5/c6 ),
    .o({\sub4_sub5/c7 ,n30[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \sub4_sub5/u7  (
    .a(vsync_cnt[8]),
    .b(1'b0),
    .c(\sub4_sub5/c7 ),
    .o({\sub4_sub5/c8 ,n30[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \sub4_sub5/u8  (
    .a(vsync_cnt[9]),
    .b(1'b0),
    .c(\sub4_sub5/c8 ),
    .o({\sub4_sub5/c9 ,n30[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \sub4_sub5/u9  (
    .a(vsync_cnt[10]),
    .b(1'b0),
    .c(\sub4_sub5/c9 ),
    .o({\sub4_sub5/c10 ,n30[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    \sub4_sub5/ucin  (
    .a(1'b0),
    .o({\sub4_sub5/c0 ,open_n296}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \sub4_sub5/ucout  (
    .c(\sub4_sub5/c10 ),
    .o({open_n299,n30[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2/u0  (
    .a(hsync_cnt[3]),
    .b(n32[3]),
    .c(\u2/c0 ),
    .o({\u2/c1 ,n28[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2/u1  (
    .a(hsync_cnt[4]),
    .b(n32[4]),
    .c(\u2/c1 ),
    .o({\u2/c2 ,n28[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2/u10  (
    .a(n29[6]),
    .b(n32[13]),
    .c(\u2/c10 ),
    .o({\u2/c11 ,n28[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2/u11  (
    .a(n29[6]),
    .b(n32[14]),
    .c(\u2/c11 ),
    .o({\u2/c12 ,n28[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2/u12  (
    .a(n29[6]),
    .b(n32[15]),
    .c(\u2/c12 ),
    .o({open_n300,n28[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2/u2  (
    .a(n29[0]),
    .b(n32[5]),
    .c(\u2/c2 ),
    .o({\u2/c3 ,n28[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2/u3  (
    .a(n29[1]),
    .b(n32[6]),
    .c(\u2/c3 ),
    .o({\u2/c4 ,n28[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2/u4  (
    .a(n29[2]),
    .b(n32[7]),
    .c(\u2/c4 ),
    .o({\u2/c5 ,n28[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2/u5  (
    .a(n29[3]),
    .b(n32[8]),
    .c(\u2/c5 ),
    .o({\u2/c6 ,n28[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2/u6  (
    .a(n29[4]),
    .b(n32[9]),
    .c(\u2/c6 ),
    .o({\u2/c7 ,n28[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2/u7  (
    .a(n29[5]),
    .b(n32[10]),
    .c(\u2/c7 ),
    .o({\u2/c8 ,n28[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2/u8  (
    .a(n29[6]),
    .b(n32[11]),
    .c(\u2/c8 ),
    .o({\u2/c9 ,n28[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2/u9  (
    .a(n29[6]),
    .b(n32[12]),
    .c(\u2/c9 ),
    .o({\u2/c10 ,n28[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2/ucin  (
    .a(1'b0),
    .o({\u2/c0 ,open_n303}));

endmodule 

module reg_sr_as_w1
  (
  clk,
  d,
  en,
  reset,
  set,
  q
  );

  input clk;
  input d;
  input en;
  input reset;
  input set;
  output q;

  parameter REGSET = "RESET";
  wire enout;
  wire resetout;

  AL_MUX u_en0 (
    .i0(q),
    .i1(d),
    .sel(en),
    .o(enout));
  AL_MUX u_reset0 (
    .i0(enout),
    .i1(1'b0),
    .sel(reset),
    .o(resetout));
  AL_DFF #(
    .INI((REGSET == "SET") ? 1'b1 : 1'b0))
    u_seq0 (
    .clk(clk),
    .d(resetout),
    .reset(1'b0),
    .set(set),
    .q(q));

endmodule 

module i2c_module  // sources/rtl/i2c_module.v(2)
  (
  address,
  clk,
  reset_n,
  sda_in,
  write,
  writedata,
  ready,
  scl_out,
  sda,
  sda_oe,
  success_out
  );

  input [2:0] address;  // sources/rtl/i2c_module.v(14)
  input clk;  // sources/rtl/i2c_module.v(3)
  input reset_n;  // sources/rtl/i2c_module.v(4)
  input sda_in;  // sources/rtl/i2c_module.v(7)
  input write;  // sources/rtl/i2c_module.v(13)
  input [7:0] writedata;  // sources/rtl/i2c_module.v(12)
  output ready;  // sources/rtl/i2c_module.v(16)
  output scl_out;  // sources/rtl/i2c_module.v(10)
  output sda;  // sources/rtl/i2c_module.v(8)
  output sda_oe;  // sources/rtl/i2c_module.v(6)
  output success_out;  // sources/rtl/i2c_module.v(17)

  // localparam STATE_ADDRESS_ACK = 10;
  // localparam STATE_ADDRESS_BIT_1 = 2;
  // localparam STATE_ADDRESS_BIT_2 = 3;
  // localparam STATE_ADDRESS_BIT_3 = 4;
  // localparam STATE_ADDRESS_BIT_4 = 5;
  // localparam STATE_ADDRESS_BIT_5 = 6;
  // localparam STATE_ADDRESS_BIT_6 = 7;
  // localparam STATE_ADDRESS_BIT_7 = 8;
  // localparam STATE_ADDRESS_BIT_8 = 9;
  // localparam STATE_ADDRESS_START = 1;
  // localparam STATE_ADDRESS_START_2 = 111;
  // localparam STATE_ADDRESS_START_3 = 112;
  // localparam STATE_DATA_ACK = 28;
  // localparam STATE_DATA_BIT_1 = 20;
  // localparam STATE_DATA_BIT_2 = 21;
  // localparam STATE_DATA_BIT_3 = 22;
  // localparam STATE_DATA_BIT_4 = 23;
  // localparam STATE_DATA_BIT_5 = 24;
  // localparam STATE_DATA_BIT_6 = 25;
  // localparam STATE_DATA_BIT_7 = 26;
  // localparam STATE_DATA_BIT_8 = 27;
  // localparam STATE_IDLE = 0;
  // localparam STATE_REG_ACK = 19;
  // localparam STATE_REG_BIT_1 = 11;
  // localparam STATE_REG_BIT_2 = 12;
  // localparam STATE_REG_BIT_3 = 13;
  // localparam STATE_REG_BIT_4 = 14;
  // localparam STATE_REG_BIT_5 = 15;
  // localparam STATE_REG_BIT_6 = 16;
  // localparam STATE_REG_BIT_7 = 17;
  // localparam STATE_REG_BIT_8 = 18;
  // localparam STATE_STOP = 29;
  // localparam STATE_STOP_1 = 30;
  // localparam STATE_STOP_2 = 31;
  // localparam STATE_TRANSIT_1 = 102;
  // localparam STATE_TRANSIT_2 = 192;
  wire [7:0] control_reg;  // sources/rtl/i2c_module.v(85)
  wire [7:0] divider2;  // sources/rtl/i2c_module.v(71)
  wire [7:0] n1;
  wire [7:0] n99;
  wire  \sel0_b0/B1 ;
  wire  \sel0_b0/B35 ;
  wire  \sel0_b1/B10 ;
  wire  \sel0_b1/B23 ;
  wire  \sel0_b2/B11 ;
  wire  \sel0_b2/B12 ;
  wire  \sel0_b2/B20 ;
  wire  \sel0_b2/B21 ;
  wire  \sel0_b2/B29 ;
  wire  \sel0_b2/B3 ;
  wire  \sel0_b2/B4 ;
  wire  \sel0_b3/B22 ;
  wire  \sel0_b3/B26 ;
  wire  \sel0_b3/B8 ;
  wire  \sel0_b4/B16 ;
  wire  \sel0_b4/B17 ;
  wire  \sel0_b4/B9 ;
  wire  \sel0_b5/B34 ;
  wire  \sel1/B33 ;
  wire  \sel5/B3 ;
  wire [7:0] slave_address;  // sources/rtl/i2c_module.v(86)
  wire [7:0] slave_data_1;  // sources/rtl/i2c_module.v(88)
  wire [7:0] slave_reg_address;  // sources/rtl/i2c_module.v(87)
  wire [7:0] state_next;  // sources/rtl/i2c_module.v(21)
  wire _al_u108_o;
  wire _al_u109_o;
  wire _al_u113_o;
  wire _al_u114_o;
  wire _al_u115_o;
  wire _al_u117_o;
  wire _al_u121_o;
  wire _al_u122_o;
  wire _al_u123_o;
  wire _al_u126_o;
  wire _al_u127_o;
  wire _al_u129_o;
  wire _al_u131_o;
  wire _al_u132_o;
  wire _al_u133_o;
  wire _al_u134_o;
  wire _al_u135_o;
  wire _al_u136_o;
  wire _al_u138_o;
  wire _al_u139_o;
  wire _al_u141_o;
  wire _al_u142_o;
  wire _al_u143_o;
  wire _al_u144_o;
  wire _al_u145_o;
  wire _al_u146_o;
  wire _al_u147_o;
  wire _al_u149_o;
  wire _al_u150_o;
  wire _al_u151_o;
  wire _al_u153_o;
  wire _al_u154_o;
  wire _al_u155_o;
  wire _al_u156_o;
  wire _al_u157_o;
  wire _al_u158_o;
  wire _al_u160_o;
  wire _al_u161_o;
  wire _al_u164_o;
  wire _al_u165_o;
  wire _al_u166_o;
  wire _al_u168_o;
  wire _al_u170_o;
  wire _al_u171_o;
  wire _al_u172_o;
  wire _al_u175_o;
  wire _al_u176_o;
  wire _al_u177_o;
  wire _al_u180_o;
  wire _al_u181_o;
  wire _al_u183_o;
  wire _al_u185_o;
  wire _al_u186_o;
  wire _al_u187_o;
  wire _al_u189_o;
  wire _al_u193_o;
  wire _al_u194_o;
  wire _al_u195_o;
  wire _al_u196_o;
  wire _al_u197_o;
  wire _al_u198_o;
  wire _al_u200_o;
  wire _al_u202_o;
  wire _al_u203_o;
  wire _al_u205_o;
  wire _al_u206_o;
  wire _al_u207_o;
  wire _al_u208_o;
  wire _al_u209_o;
  wire _al_u210_o;
  wire _al_u211_o;
  wire _al_u212_o;
  wire _al_u213_o;
  wire _al_u214_o;
  wire _al_u215_o;
  wire _al_u216_o;
  wire _al_u217_o;
  wire _al_u219_o;
  wire _al_u221_o;
  wire _al_u222_o;
  wire _al_u223_o;
  wire _al_u224_o;
  wire _al_u226_o;
  wire _al_u227_o;
  wire _al_u228_o;
  wire _al_u229_o;
  wire _al_u231_o;
  wire _al_u232_o;
  wire _al_u233_o;
  wire _al_u234_o;
  wire _al_u235_o;
  wire _al_u236_o;
  wire _al_u238_o;
  wire _al_u239_o;
  wire _al_u241_o;
  wire _al_u243_o;
  wire _al_u244_o;
  wire _al_u245_o;
  wire _al_u246_o;
  wire _al_u247_o;
  wire _al_u248_o;
  wire _al_u249_o;
  wire _al_u250_o;
  wire _al_u251_o;
  wire _al_u253_o;
  wire _al_u255_o;
  wire _al_u258_o;
  wire _al_u259_o;
  wire _al_u260_o;
  wire _al_u261_o;
  wire _al_u263_o;
  wire _al_u264_o;
  wire _al_u265_o;
  wire _al_u266_o;
  wire _al_u268_o;
  wire _al_u269_o;
  wire _al_u272_o;
  wire _al_u273_o;
  wire _al_u274_o;
  wire _al_u276_o;
  wire _al_u277_o;
  wire _al_u278_o;
  wire _al_u280_o;
  wire _al_u281_o;
  wire _al_u282_o;
  wire _al_u283_o;
  wire _al_u284_o;
  wire _al_u285_o;
  wire _al_u286_o;
  wire _al_u287_o;
  wire _al_u288_o;
  wire _al_u289_o;
  wire _al_u290_o;
  wire _al_u291_o;
  wire _al_u292_o;
  wire _al_u294_o;
  wire _al_u295_o;
  wire _al_u296_o;
  wire _al_u297_o;
  wire _al_u298_o;
  wire _al_u299_o;
  wire _al_u300_o;
  wire _al_u301_o;
  wire _al_u302_o;
  wire _al_u303_o;
  wire _al_u304_o;
  wire _al_u305_o;
  wire _al_u308_o;
  wire _al_u309_o;
  wire _al_u311_o;
  wire _al_u312_o;
  wire ack_ok;  // sources/rtl/i2c_module.v(143)
  wire \add0/c0 ;
  wire \add0/c1 ;
  wire \add0/c2 ;
  wire \add0/c3 ;
  wire \add0/c4 ;
  wire \add0/c5 ;
  wire \add0/c6 ;
  wire \add0/c7 ;
  wire clk_div_neg;
  wire mux4_b0_sel_is_3_o;
  wire mux5_b0_sel_is_3_o;
  wire mux6_b0_sel_is_3_o;
  wire mux7_b0_sel_is_3_o;
  wire mux9_b0_sel_is_0_o;
  wire n106_lutinv;
  wire n107_lutinv;
  wire n146_lutinv;
  wire n155_lutinv;
  wire n158_lutinv;
  wire n164_lutinv;
  wire n168_lutinv;
  wire n169_lutinv;
  wire n180_lutinv;
  wire n181_lutinv;
  wire n183_lutinv;
  wire n184;
  wire n186;
  wire n188;
  wire n190;
  wire n191_lutinv;
  wire n192;
  wire n194;
  wire n2;
  wire n20;
  wire n28;
  wire n29;
  wire n33;
  wire n80_lutinv;
  wire n81_lutinv;
  wire n88_lutinv;
  wire n94_lutinv;
  wire scl_out_pad;  // sources/rtl/i2c_module.v(10)
  wire scl_output_enable;  // sources/rtl/i2c_module.v(120)
  wire scl_output_zero;  // sources/rtl/i2c_module.v(121)
  wire \sel0_b3/or_or_B13_B14_o_or_B_o_lutinv ;
  wire success;  // sources/rtl/i2c_module.v(141)

  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u104 (
    .a(address[1]),
    .b(address[0]),
    .c(write),
    .o(mux4_b0_sel_is_3_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    _al_u105 (
    .a(address[1]),
    .b(address[0]),
    .c(write),
    .o(mux6_b0_sel_is_3_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    _al_u106 (
    .a(address[1]),
    .b(address[0]),
    .c(write),
    .o(mux7_b0_sel_is_3_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u107 (
    .a(address[1]),
    .b(address[0]),
    .c(write),
    .o(mux5_b0_sel_is_3_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u108 (
    .a(state_next[4]),
    .b(state_next[5]),
    .c(state_next[6]),
    .d(state_next[7]),
    .o(_al_u108_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u109 (
    .a(state_next[0]),
    .b(state_next[1]),
    .c(state_next[2]),
    .d(state_next[3]),
    .o(_al_u109_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u110 (
    .a(_al_u108_o),
    .b(_al_u109_o),
    .o(n146_lutinv));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u111 (
    .a(n146_lutinv),
    .b(reset_n),
    .o(mux9_b0_sel_is_0_o));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'h47))
    _al_u112 (
    .a(scl_out_pad),
    .b(scl_output_enable),
    .c(scl_output_zero),
    .o(n20));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*A)"),
    .INIT(16'h0002))
    _al_u113 (
    .a(state_next[4]),
    .b(state_next[5]),
    .c(state_next[6]),
    .d(state_next[7]),
    .o(_al_u113_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u114 (
    .a(state_next[0]),
    .b(state_next[1]),
    .o(_al_u114_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u115 (
    .a(state_next[2]),
    .b(state_next[3]),
    .o(_al_u115_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u116 (
    .a(_al_u113_o),
    .b(_al_u114_o),
    .c(_al_u115_o),
    .o(\sel0_b2/B3 ));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*A)"),
    .INIT(16'h0002))
    _al_u117 (
    .a(state_next[0]),
    .b(state_next[1]),
    .c(state_next[2]),
    .d(state_next[3]),
    .o(_al_u117_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u118 (
    .a(_al_u108_o),
    .b(_al_u117_o),
    .o(\sel0_b0/B35 ));
  AL_MAP_LUT4 #(
    .EQN("~(~(C*~B)*~(D*A))"),
    .INIT(16'hba30))
    _al_u119 (
    .a(\sel0_b2/B3 ),
    .b(\sel0_b0/B35 ),
    .c(success_out),
    .d(success),
    .o(n33));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    _al_u120 (
    .a(_al_u113_o),
    .b(_al_u115_o),
    .c(state_next[0]),
    .d(state_next[1]),
    .o(\sel0_b2/B4 ));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*B*~A)"),
    .INIT(16'h0400))
    _al_u121 (
    .a(state_next[0]),
    .b(state_next[1]),
    .c(state_next[2]),
    .d(state_next[3]),
    .o(_al_u121_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    _al_u122 (
    .a(state_next[0]),
    .b(state_next[1]),
    .c(state_next[2]),
    .d(state_next[3]),
    .o(_al_u122_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u123 (
    .a(_al_u108_o),
    .b(_al_u113_o),
    .c(_al_u121_o),
    .d(_al_u122_o),
    .o(_al_u123_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~(B*~A))"),
    .INIT(16'h0b00))
    _al_u124 (
    .a(\sel0_b2/B4 ),
    .b(_al_u123_o),
    .c(sda_in),
    .d(n28),
    .o(n29));
  AL_MAP_LUT4 #(
    .EQN("(B*A*(D@C))"),
    .INIT(16'h0880))
    _al_u125 (
    .a(_al_u108_o),
    .b(_al_u115_o),
    .c(state_next[0]),
    .d(state_next[1]),
    .o(n88_lutinv));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u126 (
    .a(state_next[2]),
    .b(state_next[3]),
    .o(_al_u126_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u127 (
    .a(state_next[0]),
    .b(state_next[1]),
    .o(_al_u127_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u128 (
    .a(_al_u108_o),
    .b(_al_u126_o),
    .c(_al_u127_o),
    .o(\sel0_b3/B22 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u129 (
    .a(state_next[0]),
    .b(state_next[1]),
    .o(_al_u129_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u130 (
    .a(_al_u129_o),
    .b(_al_u108_o),
    .c(_al_u115_o),
    .o(\sel0_b2/B21 ));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u131 (
    .a(n88_lutinv),
    .b(\sel0_b3/B22 ),
    .c(\sel0_b2/B21 ),
    .o(_al_u131_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*~A)"),
    .INIT(16'h0100))
    _al_u132 (
    .a(state_next[0]),
    .b(state_next[1]),
    .c(state_next[2]),
    .d(state_next[3]),
    .o(_al_u132_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*A)"),
    .INIT(16'h0080))
    _al_u133 (
    .a(state_next[0]),
    .b(state_next[1]),
    .c(state_next[2]),
    .d(state_next[3]),
    .o(_al_u133_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u134 (
    .a(state_next[0]),
    .b(state_next[1]),
    .c(state_next[3]),
    .o(_al_u134_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(~D*~C*~B))"),
    .INIT(16'haaa8))
    _al_u135 (
    .a(_al_u108_o),
    .b(_al_u132_o),
    .c(_al_u133_o),
    .d(_al_u134_o),
    .o(_al_u135_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*~B*~A)"),
    .INIT(16'h0010))
    _al_u136 (
    .a(state_next[0]),
    .b(state_next[1]),
    .c(state_next[2]),
    .d(state_next[3]),
    .o(_al_u136_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*~B))"),
    .INIT(8'ha8))
    _al_u137 (
    .a(_al_u108_o),
    .b(_al_u122_o),
    .c(_al_u136_o),
    .o(n80_lutinv));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*~A)"),
    .INIT(16'h0040))
    _al_u138 (
    .a(state_next[0]),
    .b(state_next[1]),
    .c(state_next[2]),
    .d(state_next[3]),
    .o(_al_u138_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*~B*A)"),
    .INIT(16'h0020))
    _al_u139 (
    .a(state_next[0]),
    .b(state_next[1]),
    .c(state_next[2]),
    .d(state_next[3]),
    .o(_al_u139_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*~B))"),
    .INIT(8'ha8))
    _al_u140 (
    .a(_al_u108_o),
    .b(_al_u138_o),
    .c(_al_u139_o),
    .o(n81_lutinv));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*~A)"),
    .INIT(16'h0004))
    _al_u141 (
    .a(state_next[0]),
    .b(state_next[1]),
    .c(state_next[2]),
    .d(state_next[3]),
    .o(_al_u141_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*A)"),
    .INIT(16'h0080))
    _al_u142 (
    .a(state_next[4]),
    .b(state_next[5]),
    .c(state_next[6]),
    .d(state_next[7]),
    .o(_al_u142_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*C)*~(B*A))"),
    .INIT(16'h0777))
    _al_u143 (
    .a(_al_u108_o),
    .b(_al_u141_o),
    .c(_al_u109_o),
    .d(_al_u142_o),
    .o(_al_u143_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*~A)"),
    .INIT(16'h0100))
    _al_u144 (
    .a(_al_u135_o),
    .b(n80_lutinv),
    .c(n81_lutinv),
    .d(_al_u143_o),
    .o(_al_u144_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*~A)"),
    .INIT(16'h1000))
    _al_u145 (
    .a(state_next[4]),
    .b(state_next[5]),
    .c(state_next[6]),
    .d(state_next[7]),
    .o(_al_u145_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*C)*~(B*A))"),
    .INIT(16'h0777))
    _al_u146 (
    .a(_al_u113_o),
    .b(_al_u139_o),
    .c(_al_u109_o),
    .d(_al_u145_o),
    .o(_al_u146_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*~B))"),
    .INIT(8'ha8))
    _al_u147 (
    .a(_al_u113_o),
    .b(_al_u136_o),
    .c(_al_u138_o),
    .o(_al_u147_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u148 (
    .a(_al_u113_o),
    .b(_al_u117_o),
    .o(\sel0_b4/B16 ));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u149 (
    .a(state_next[0]),
    .b(state_next[1]),
    .c(state_next[2]),
    .d(state_next[3]),
    .o(_al_u149_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u150 (
    .a(_al_u108_o),
    .b(_al_u113_o),
    .c(_al_u109_o),
    .d(_al_u149_o),
    .o(_al_u150_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*A)"),
    .INIT(16'h0200))
    _al_u151 (
    .a(_al_u146_o),
    .b(_al_u147_o),
    .c(\sel0_b4/B16 ),
    .d(_al_u150_o),
    .o(_al_u151_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u152 (
    .a(_al_u113_o),
    .b(_al_u133_o),
    .o(\sel0_b4/B9 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u153 (
    .a(_al_u113_o),
    .b(_al_u126_o),
    .o(_al_u153_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*~A)"),
    .INIT(16'h0040))
    _al_u154 (
    .a(state_next[4]),
    .b(state_next[5]),
    .c(state_next[6]),
    .d(state_next[7]),
    .o(_al_u154_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u155 (
    .a(_al_u113_o),
    .b(_al_u138_o),
    .c(_al_u141_o),
    .d(_al_u154_o),
    .o(_al_u155_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    _al_u156 (
    .a(\sel0_b4/B9 ),
    .b(_al_u153_o),
    .c(_al_u155_o),
    .o(_al_u156_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u157 (
    .a(_al_u131_o),
    .b(_al_u144_o),
    .c(_al_u151_o),
    .d(_al_u156_o),
    .o(_al_u157_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*~A)"),
    .INIT(16'h4000))
    _al_u158 (
    .a(state_next[0]),
    .b(state_next[1]),
    .c(state_next[2]),
    .d(state_next[3]),
    .o(_al_u158_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u159 (
    .a(_al_u113_o),
    .b(_al_u158_o),
    .o(n180_lutinv));
  EG_PHY_PAD #(
    //.LOCATION("D16"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u16 (
    .do({open_n1,open_n2,open_n3,scl_out_pad}),
    .opad(scl_out));  // sources/rtl/i2c_module.v(10)
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u160 (
    .a(\sel0_b0/B35 ),
    .b(n180_lutinv),
    .o(_al_u160_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~(B*A))"),
    .INIT(16'h7000))
    _al_u161 (
    .a(_al_u157_o),
    .b(_al_u160_o),
    .c(n28),
    .d(scl_output_zero),
    .o(_al_u161_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u162 (
    .a(_al_u113_o),
    .b(_al_u149_o),
    .o(n181_lutinv));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u163 (
    .a(_al_u149_o),
    .b(_al_u154_o),
    .o(\sel0_b5/B34 ));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(~D*~(~C*~A)))"),
    .INIT(16'h3301))
    _al_u164 (
    .a(\sel0_b2/B3 ),
    .b(n181_lutinv),
    .c(\sel0_b5/B34 ),
    .d(n28),
    .o(_al_u164_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u165 (
    .a(_al_u164_o),
    .b(\sel0_b5/B34 ),
    .c(scl_output_zero),
    .o(_al_u165_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*C)*~(B*~A))"),
    .INIT(16'hbb0b))
    _al_u166 (
    .a(\sel0_b2/B4 ),
    .b(_al_u123_o),
    .c(n28),
    .d(scl_output_zero),
    .o(_al_u166_o));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~B*~A)"),
    .INIT(8'hfe))
    _al_u167 (
    .a(_al_u161_o),
    .b(_al_u165_o),
    .c(_al_u166_o),
    .o(n194));
  AL_MAP_LUT4 #(
    .EQN("(~(D*C)*~(B*A))"),
    .INIT(16'h0777))
    _al_u168 (
    .a(_al_u108_o),
    .b(_al_u121_o),
    .c(_al_u138_o),
    .d(_al_u154_o),
    .o(_al_u168_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*~B))"),
    .INIT(8'ha8))
    _al_u169 (
    .a(_al_u113_o),
    .b(_al_u122_o),
    .c(_al_u141_o),
    .o(n94_lutinv));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*~B*~A)"),
    .INIT(16'h0010))
    _al_u170 (
    .a(\sel0_b4/B9 ),
    .b(_al_u153_o),
    .c(_al_u168_o),
    .d(n94_lutinv),
    .o(_al_u170_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u171 (
    .a(_al_u131_o),
    .b(_al_u144_o),
    .c(_al_u151_o),
    .d(_al_u170_o),
    .o(_al_u171_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~(B*A))"),
    .INIT(16'h7000))
    _al_u172 (
    .a(_al_u171_o),
    .b(_al_u160_o),
    .c(n28),
    .d(success),
    .o(_al_u172_o));
  AL_MAP_LUT4 #(
    .EQN("(A*(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C))"),
    .INIT(16'ha808))
    _al_u173 (
    .a(\sel0_b2/B4 ),
    .b(ack_ok),
    .c(n28),
    .d(success),
    .o(\sel5/B3 ));
  AL_MAP_LUT4 #(
    .EQN("~(~C*~A*~(D*~B))"),
    .INIT(16'hfbfa))
    _al_u174 (
    .a(_al_u172_o),
    .b(_al_u164_o),
    .c(\sel5/B3 ),
    .d(success),
    .o(n192));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*~A)"),
    .INIT(8'h04))
    _al_u175 (
    .a(\sel0_b0/B35 ),
    .b(_al_u123_o),
    .c(n180_lutinv),
    .o(_al_u175_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(A*~(C*~B)))"),
    .INIT(16'h7500))
    _al_u176 (
    .a(_al_u164_o),
    .b(_al_u175_o),
    .c(n28),
    .d(scl_output_enable),
    .o(_al_u176_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(B*~(~D*~C)))"),
    .INIT(16'h1115))
    _al_u177 (
    .a(_al_u176_o),
    .b(\sel0_b2/B4 ),
    .c(ack_ok),
    .d(n28),
    .o(_al_u177_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*C)*~(B*A))"),
    .INIT(16'h7707))
    _al_u178 (
    .a(_al_u177_o),
    .b(_al_u157_o),
    .c(n28),
    .d(scl_output_enable),
    .o(n188));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u179 (
    .a(_al_u113_o),
    .b(_al_u115_o),
    .o(n191_lutinv));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u180 (
    .a(n191_lutinv),
    .b(\sel0_b5/B34 ),
    .o(_al_u180_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u181 (
    .a(_al_u171_o),
    .b(_al_u180_o),
    .o(_al_u181_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u182 (
    .a(_al_u113_o),
    .b(_al_u122_o),
    .o(n168_lutinv));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u183 (
    .a(n168_lutinv),
    .b(ack_ok),
    .o(_al_u183_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((~B*~A))+C*D*~((~B*~A))+~(C)*D*(~B*~A)+C*D*(~B*~A))"),
    .INIT(16'hf1e0))
    _al_u184 (
    .a(_al_u181_o),
    .b(n28),
    .c(state_next[7]),
    .d(_al_u183_o),
    .o(n99[7]));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*~A)"),
    .INIT(8'h04))
    _al_u185 (
    .a(_al_u123_o),
    .b(ack_ok),
    .c(n28),
    .o(_al_u185_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(B)*~(A)+~C*B*~(A)+~(~C)*B*A+~C*B*A)"),
    .INIT(8'h8d))
    _al_u186 (
    .a(\sel0_b0/B35 ),
    .b(n28),
    .c(_al_u185_o),
    .o(_al_u186_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u187 (
    .a(\sel0_b5/B34 ),
    .b(_al_u186_o),
    .o(_al_u187_o));
  AL_MAP_LUT4 #(
    .EQN("~(D*~(B*~(~C*~A)))"),
    .INIT(16'hc8ff))
    _al_u188 (
    .a(_al_u181_o),
    .b(state_next[6]),
    .c(n28),
    .d(_al_u187_o),
    .o(n99[6]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u189 (
    .a(_al_u186_o),
    .b(state_next[5]),
    .o(_al_u189_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(~D*~C*~A))"),
    .INIT(16'h3332))
    _al_u190 (
    .a(_al_u181_o),
    .b(_al_u189_o),
    .c(n28),
    .d(state_next[3]),
    .o(n99[5]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u191 (
    .a(_al_u109_o),
    .b(_al_u145_o),
    .o(n169_lutinv));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u192 (
    .a(_al_u113_o),
    .b(_al_u109_o),
    .o(\sel0_b4/B17 ));
  AL_MAP_LUT4 #(
    .EQN("(A*~(~D*~C*~B))"),
    .INIT(16'haaa8))
    _al_u193 (
    .a(_al_u113_o),
    .b(_al_u117_o),
    .c(_al_u139_o),
    .d(_al_u141_o),
    .o(_al_u193_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u194 (
    .a(n169_lutinv),
    .b(_al_u147_o),
    .c(\sel0_b4/B17 ),
    .d(_al_u193_o),
    .o(_al_u194_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*A)"),
    .INIT(16'h0002))
    _al_u195 (
    .a(_al_u194_o),
    .b(\sel0_b2/B4 ),
    .c(\sel0_b4/B9 ),
    .d(_al_u153_o),
    .o(_al_u195_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u196 (
    .a(\sel0_b2/B3 ),
    .b(\sel0_b5/B34 ),
    .o(_al_u196_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h7735))
    _al_u197 (
    .a(_al_u195_o),
    .b(_al_u196_o),
    .c(n28),
    .d(state_next[4]),
    .o(_al_u197_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u198 (
    .a(_al_u123_o),
    .b(ack_ok),
    .c(n28),
    .o(_al_u198_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u199 (
    .a(_al_u108_o),
    .b(_al_u149_o),
    .o(n164_lutinv));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u200 (
    .a(n180_lutinv),
    .b(n164_lutinv),
    .c(n28),
    .o(_al_u200_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u201 (
    .a(_al_u113_o),
    .b(_al_u149_o),
    .c(n28),
    .o(\sel0_b0/B1 ));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*~A)"),
    .INIT(8'h04))
    _al_u202 (
    .a(_al_u198_o),
    .b(_al_u200_o),
    .c(\sel0_b0/B1 ),
    .o(_al_u202_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hd151))
    _al_u203 (
    .a(_al_u202_o),
    .b(n28),
    .c(state_next[4]),
    .d(state_next[5]),
    .o(_al_u203_o));
  AL_MAP_LUT4 #(
    .EQN("~(~C*~B*~(D*A))"),
    .INIT(16'hfefc))
    _al_u204 (
    .a(_al_u181_o),
    .b(_al_u197_o),
    .c(_al_u203_o),
    .d(state_next[4]),
    .o(n99[4]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*C)*~(B*A))"),
    .INIT(16'h0777))
    _al_u205 (
    .a(_al_u108_o),
    .b(_al_u134_o),
    .c(_al_u138_o),
    .d(_al_u154_o),
    .o(_al_u205_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*~B))"),
    .INIT(8'h8a))
    _al_u206 (
    .a(_al_u126_o),
    .b(state_next[0]),
    .c(state_next[1]),
    .o(_al_u206_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*~B*~A)"),
    .INIT(16'h0010))
    _al_u207 (
    .a(n88_lutinv),
    .b(\sel0_b2/B21 ),
    .c(_al_u205_o),
    .d(_al_u206_o),
    .o(_al_u207_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u208 (
    .a(_al_u207_o),
    .b(\sel0_b2/B4 ),
    .c(_al_u153_o),
    .o(_al_u208_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u209 (
    .a(_al_u208_o),
    .b(n28),
    .c(state_next[3]),
    .o(_al_u209_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(~B*~A))"),
    .INIT(8'he0))
    _al_u210 (
    .a(n180_lutinv),
    .b(n164_lutinv),
    .c(n28),
    .o(_al_u210_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*B))"),
    .INIT(8'ha2))
    _al_u211 (
    .a(_al_u198_o),
    .b(n28),
    .c(state_next[3]),
    .o(_al_u211_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u212 (
    .a(\sel0_b2/B3 ),
    .b(\sel0_b4/B9 ),
    .c(n28),
    .o(_al_u212_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*~B))"),
    .INIT(8'ha8))
    _al_u213 (
    .a(_al_u108_o),
    .b(_al_u117_o),
    .c(_al_u133_o),
    .o(_al_u213_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u214 (
    .a(_al_u213_o),
    .b(n28),
    .o(_al_u214_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(~B*~A))"),
    .INIT(8'h0e))
    _al_u215 (
    .a(n181_lutinv),
    .b(\sel0_b5/B34 ),
    .c(n28),
    .o(_al_u215_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u216 (
    .a(_al_u212_o),
    .b(_al_u214_o),
    .c(_al_u215_o),
    .o(_al_u216_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    _al_u217 (
    .a(_al_u210_o),
    .b(_al_u211_o),
    .c(_al_u216_o),
    .o(_al_u217_o));
  AL_MAP_LUT4 #(
    .EQN("~(C*~B*~(D*A))"),
    .INIT(16'hefcf))
    _al_u218 (
    .a(_al_u181_o),
    .b(_al_u209_o),
    .c(_al_u217_o),
    .d(state_next[3]),
    .o(n99[3]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u219 (
    .a(_al_u146_o),
    .b(_al_u147_o),
    .o(_al_u219_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u220 (
    .a(_al_u108_o),
    .b(_al_u121_o),
    .o(n158_lutinv));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u221 (
    .a(\sel0_b0/B35 ),
    .b(n158_lutinv),
    .c(n80_lutinv),
    .d(n81_lutinv),
    .o(_al_u221_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u222 (
    .a(_al_u126_o),
    .b(_al_u127_o),
    .o(_al_u222_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u223 (
    .a(\sel0_b2/B4 ),
    .b(_al_u222_o),
    .c(_al_u113_o),
    .o(_al_u223_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u224 (
    .a(_al_u131_o),
    .b(_al_u219_o),
    .c(_al_u221_o),
    .d(_al_u223_o),
    .o(_al_u224_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u225 (
    .a(n168_lutinv),
    .b(ack_ok),
    .c(n28),
    .o(\sel0_b3/or_or_B13_B14_o_or_B_o_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(~D*C*B))"),
    .INIT(16'h5515))
    _al_u226 (
    .a(\sel0_b2/B3 ),
    .b(n28),
    .c(state_next[2]),
    .d(state_next[0]),
    .o(_al_u226_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    _al_u227 (
    .a(\sel0_b3/or_or_B13_B14_o_or_B_o_lutinv ),
    .b(_al_u215_o),
    .c(_al_u226_o),
    .o(_al_u227_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    _al_u228 (
    .a(_al_u224_o),
    .b(_al_u227_o),
    .c(n28),
    .o(_al_u228_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u229 (
    .a(n28),
    .b(_al_u180_o),
    .o(_al_u229_o));
  AL_MAP_LUT4 #(
    .EQN("~(B*~(D*~(~C*~A)))"),
    .INIT(16'hfb33))
    _al_u230 (
    .a(_al_u181_o),
    .b(_al_u228_o),
    .c(_al_u229_o),
    .d(state_next[2]),
    .o(n99[2]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u231 (
    .a(n81_lutinv),
    .b(_al_u143_o),
    .o(_al_u231_o));
  AL_MAP_LUT3 #(
    .EQN("(A*(C@B))"),
    .INIT(8'h28))
    _al_u232 (
    .a(_al_u153_o),
    .b(state_next[0]),
    .c(state_next[1]),
    .o(_al_u232_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(~C*~B*A))"),
    .INIT(16'h00fd))
    _al_u233 (
    .a(_al_u231_o),
    .b(_al_u232_o),
    .c(\sel0_b0/B35 ),
    .d(n28),
    .o(_al_u233_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u234 (
    .a(\sel0_b2/B3 ),
    .b(n180_lutinv),
    .o(_al_u234_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*C)*~(B*~A))"),
    .INIT(16'h0bbb))
    _al_u235 (
    .a(_al_u234_o),
    .b(n28),
    .c(_al_u108_o),
    .d(_al_u185_o),
    .o(_al_u235_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u236 (
    .a(n88_lutinv),
    .b(_al_u205_o),
    .o(_al_u236_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u237 (
    .a(_al_u113_o),
    .b(_al_u138_o),
    .o(\sel0_b1/B10 ));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(~C*~B*A))"),
    .INIT(16'h00fd))
    _al_u238 (
    .a(_al_u236_o),
    .b(\sel0_b1/B10 ),
    .c(_al_u193_o),
    .d(n28),
    .o(_al_u238_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*~A)"),
    .INIT(16'h0004))
    _al_u239 (
    .a(_al_u233_o),
    .b(_al_u235_o),
    .c(_al_u238_o),
    .d(_al_u215_o),
    .o(_al_u239_o));
  AL_MAP_LUT4 #(
    .EQN("~(B*~(C*~(~D*~A)))"),
    .INIT(16'hf3b3))
    _al_u240 (
    .a(_al_u181_o),
    .b(_al_u239_o),
    .c(state_next[1]),
    .d(_al_u229_o),
    .o(n99[1]));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u241 (
    .a(\sel0_b2/B4 ),
    .b(_al_u153_o),
    .c(state_next[0]),
    .o(_al_u241_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u242 (
    .a(_al_u108_o),
    .b(_al_u132_o),
    .o(\sel0_b3/B26 ));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u243 (
    .a(\sel0_b2/B21 ),
    .b(\sel0_b3/B26 ),
    .c(_al_u147_o),
    .o(_al_u243_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*~B))"),
    .INIT(8'ha8))
    _al_u244 (
    .a(_al_u108_o),
    .b(_al_u136_o),
    .c(_al_u138_o),
    .o(_al_u244_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*~B))"),
    .INIT(8'ha8))
    _al_u245 (
    .a(_al_u108_o),
    .b(_al_u158_o),
    .c(_al_u141_o),
    .o(_al_u245_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*~A)"),
    .INIT(16'h0004))
    _al_u246 (
    .a(\sel0_b4/B17 ),
    .b(_al_u155_o),
    .c(_al_u244_o),
    .d(_al_u245_o),
    .o(_al_u246_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*~A)"),
    .INIT(16'h4000))
    _al_u247 (
    .a(_al_u198_o),
    .b(_al_u241_o),
    .c(_al_u243_o),
    .d(_al_u246_o),
    .o(_al_u247_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~(~B*~A))"),
    .INIT(16'h0e00))
    _al_u248 (
    .a(n191_lutinv),
    .b(\sel0_b5/B34 ),
    .c(n28),
    .d(state_next[0]),
    .o(_al_u248_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u249 (
    .a(_al_u248_o),
    .b(n146_lutinv),
    .c(control_reg[0]),
    .o(_al_u249_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u250 (
    .a(n28),
    .b(state_next[0]),
    .o(_al_u250_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~C*~(~D*A)))"),
    .INIT(16'hc0c8))
    _al_u251 (
    .a(_al_u247_o),
    .b(_al_u249_o),
    .c(_al_u250_o),
    .d(_al_u229_o),
    .o(_al_u251_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C*A))"),
    .INIT(8'hb3))
    _al_u252 (
    .a(_al_u181_o),
    .b(_al_u251_o),
    .c(state_next[0]),
    .o(n99[0]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u253 (
    .a(_al_u115_o),
    .b(state_next[0]),
    .o(_al_u253_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u254 (
    .a(n28),
    .b(ready),
    .o(n107_lutinv));
  AL_MAP_LUT4 #(
    .EQN("(D*~(~C*~B*A))"),
    .INIT(16'hfd00))
    _al_u255 (
    .a(_al_u171_o),
    .b(\sel0_b0/B35 ),
    .c(_al_u253_o),
    .d(n107_lutinv),
    .o(_al_u255_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u256 (
    .a(_al_u171_o),
    .b(_al_u180_o),
    .c(\sel0_b0/B35 ),
    .o(n183_lutinv));
  AL_MAP_LUT4 #(
    .EQN("~(~B*~A*~(D*~C))"),
    .INIT(16'hefee))
    _al_u257 (
    .a(_al_u255_o),
    .b(n183_lutinv),
    .c(_al_u164_o),
    .d(ready),
    .o(n190));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u258 (
    .a(n80_lutinv),
    .b(_al_u150_o),
    .o(_al_u258_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u259 (
    .a(_al_u219_o),
    .b(_al_u232_o),
    .c(_al_u258_o),
    .o(_al_u259_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u260 (
    .a(_al_u117_o),
    .b(_al_u133_o),
    .o(_al_u260_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    _al_u261 (
    .a(_al_u253_o),
    .b(_al_u168_o),
    .c(_al_u260_o),
    .o(_al_u261_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u262 (
    .a(_al_u113_o),
    .b(_al_u132_o),
    .o(\sel0_b3/B8 ));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u263 (
    .a(n168_lutinv),
    .b(\sel0_b3/B26 ),
    .c(\sel0_b3/B8 ),
    .o(_al_u263_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u264 (
    .a(_al_u131_o),
    .b(_al_u231_o),
    .c(_al_u261_o),
    .d(_al_u263_o),
    .o(_al_u264_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(B*A))"),
    .INIT(8'h07))
    _al_u265 (
    .a(_al_u259_o),
    .b(_al_u264_o),
    .c(n28),
    .o(_al_u265_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf5d0))
    _al_u266 (
    .a(_al_u196_o),
    .b(n181_lutinv),
    .c(sda_oe),
    .d(n28),
    .o(_al_u266_o));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~B*~A)"),
    .INIT(8'hfe))
    _al_u267 (
    .a(n183_lutinv),
    .b(_al_u265_o),
    .c(_al_u266_o),
    .o(n186));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u268 (
    .a(n28),
    .b(slave_address[7]),
    .o(_al_u268_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u269 (
    .a(_al_u268_o),
    .b(_al_u142_o),
    .o(_al_u269_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u270 (
    .a(_al_u108_o),
    .b(_al_u114_o),
    .c(_al_u115_o),
    .o(\sel0_b2/B20 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u271 (
    .a(_al_u108_o),
    .b(_al_u139_o),
    .o(\sel0_b2/B29 ));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u272 (
    .a(n28),
    .b(slave_address[3]),
    .o(_al_u272_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u273 (
    .a(n28),
    .b(slave_reg_address[4]),
    .o(_al_u273_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u274 (
    .a(\sel0_b2/B20 ),
    .b(\sel0_b2/B29 ),
    .c(_al_u272_o),
    .d(_al_u273_o),
    .o(_al_u274_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u275 (
    .a(_al_u138_o),
    .b(_al_u154_o),
    .o(\sel0_b1/B23 ));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u276 (
    .a(n28),
    .b(slave_address[2]),
    .o(_al_u276_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u277 (
    .a(_al_u108_o),
    .b(_al_u138_o),
    .c(_al_u276_o),
    .o(_al_u277_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D*~C*A))"),
    .INIT(16'h3133))
    _al_u278 (
    .a(\sel0_b1/B23 ),
    .b(_al_u277_o),
    .c(n28),
    .d(slave_reg_address[7]),
    .o(_al_u278_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u279 (
    .a(_al_u113_o),
    .b(_al_u139_o),
    .o(\sel0_b2/B11 ));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u280 (
    .a(n28),
    .b(slave_data_1[5]),
    .o(_al_u280_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u281 (
    .a(n28),
    .b(slave_data_1[4]),
    .o(_al_u281_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u282 (
    .a(\sel0_b2/B11 ),
    .b(\sel0_b1/B10 ),
    .c(_al_u280_o),
    .d(_al_u281_o),
    .o(_al_u282_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*~A)"),
    .INIT(16'h4000))
    _al_u283 (
    .a(_al_u269_o),
    .b(_al_u274_o),
    .c(_al_u278_o),
    .d(_al_u282_o),
    .o(_al_u283_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u284 (
    .a(n28),
    .b(slave_address[0]),
    .o(_al_u284_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u285 (
    .a(\sel0_b3/B26 ),
    .b(_al_u284_o),
    .o(_al_u285_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u286 (
    .a(n28),
    .b(slave_reg_address[3]),
    .o(_al_u286_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u287 (
    .a(n28),
    .b(slave_address[6]),
    .o(_al_u287_o));
  AL_MAP_LUT4 #(
    .EQN("~((D*B)*~(A)*~(C)+(D*B)*A*~(C)+~((D*B))*A*C+(D*B)*A*C)"),
    .INIT(16'h535f))
    _al_u288 (
    .a(_al_u286_o),
    .b(_al_u287_o),
    .c(_al_u158_o),
    .d(_al_u245_o),
    .o(_al_u288_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u289 (
    .a(_al_u114_o),
    .b(n28),
    .c(slave_data_1[1]),
    .o(_al_u289_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u290 (
    .a(n28),
    .b(slave_data_1[2]),
    .o(_al_u290_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u291 (
    .a(_al_u153_o),
    .b(\sel0_b3/B8 ),
    .c(_al_u289_o),
    .d(_al_u290_o),
    .o(_al_u291_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    _al_u292 (
    .a(_al_u285_o),
    .b(_al_u288_o),
    .c(_al_u291_o),
    .o(_al_u292_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u293 (
    .a(\sel0_b5/B34 ),
    .b(n28),
    .c(sda),
    .o(\sel1/B33 ));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u294 (
    .a(_al_u283_o),
    .b(_al_u292_o),
    .c(\sel1/B33 ),
    .o(_al_u294_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u295 (
    .a(_al_u108_o),
    .b(_al_u122_o),
    .c(slave_address[5]),
    .o(_al_u295_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u296 (
    .a(_al_u108_o),
    .b(_al_u136_o),
    .c(slave_address[4]),
    .o(_al_u296_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~B*~(D*A))"),
    .INIT(16'h0103))
    _al_u297 (
    .a(\sel0_b3/B22 ),
    .b(_al_u295_o),
    .c(_al_u296_o),
    .d(slave_reg_address[6]),
    .o(_al_u297_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(A*~(D*B)))"),
    .INIT(16'h0d05))
    _al_u298 (
    .a(_al_u297_o),
    .b(\sel0_b2/B21 ),
    .c(n28),
    .d(slave_reg_address[5]),
    .o(_al_u298_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u299 (
    .a(\sel0_b4/B16 ),
    .b(\sel0_b4/B9 ),
    .c(slave_reg_address[0]),
    .d(slave_data_1[3]),
    .o(_al_u299_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(~B*~(~C*A)))"),
    .INIT(16'hce00))
    _al_u300 (
    .a(\sel0_b2/B3 ),
    .b(n181_lutinv),
    .c(n28),
    .d(sda),
    .o(_al_u300_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u301 (
    .a(_al_u121_o),
    .b(n28),
    .c(slave_data_1[0]),
    .o(_al_u301_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u302 (
    .a(_al_u153_o),
    .b(_al_u301_o),
    .o(_al_u302_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~B*~(~D*~A))"),
    .INIT(16'h0302))
    _al_u303 (
    .a(_al_u299_o),
    .b(_al_u300_o),
    .c(_al_u302_o),
    .d(n28),
    .o(_al_u303_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u304 (
    .a(n180_lutinv),
    .b(\sel0_b4/B17 ),
    .c(slave_reg_address[1]),
    .o(_al_u304_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u305 (
    .a(n169_lutinv),
    .b(n164_lutinv),
    .c(slave_reg_address[2]),
    .d(slave_data_1[7]),
    .o(_al_u305_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u306 (
    .a(_al_u108_o),
    .b(_al_u133_o),
    .o(n155_lutinv));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u307 (
    .a(_al_u113_o),
    .b(_al_u136_o),
    .o(\sel0_b2/B12 ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u308 (
    .a(n155_lutinv),
    .b(\sel0_b2/B12 ),
    .c(slave_address[1]),
    .d(slave_data_1[6]),
    .o(_al_u308_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(C*B*A))"),
    .INIT(16'h007f))
    _al_u309 (
    .a(_al_u304_o),
    .b(_al_u305_o),
    .c(_al_u308_o),
    .d(n28),
    .o(_al_u309_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u310 (
    .a(n28),
    .b(sda),
    .o(n106_lutinv));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u311 (
    .a(n106_lutinv),
    .b(_al_u196_o),
    .o(_al_u311_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*~A)"),
    .INIT(16'h0004))
    _al_u312 (
    .a(_al_u298_o),
    .b(_al_u303_o),
    .c(_al_u309_o),
    .d(_al_u311_o),
    .o(_al_u312_o));
  AL_MAP_LUT3 #(
    .EQN("~(C*B*~A)"),
    .INIT(8'hbf))
    _al_u313 (
    .a(n183_lutinv),
    .b(_al_u294_o),
    .c(_al_u312_o),
    .o(n184));
  AL_MAP_LUT1 #(
    .EQN("(~A)"),
    .INIT(2'h1))
    _al_u314 (
    .a(reset_n),
    .o(n2));
  AL_MAP_LUT1 #(
    .EQN("(~A)"),
    .INIT(2'h1))
    _al_u315 (
    .a(n28),
    .o(clk_div_neg));
  reg_ar_as_w1 ack_ok_reg (
    .clk(divider2[7]),
    .d(n29),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(ack_ok));  // sources/rtl/i2c_module.v(153)
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add0/u0  (
    .a(divider2[0]),
    .b(1'b1),
    .c(\add0/c0 ),
    .o({\add0/c1 ,n1[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add0/u1  (
    .a(divider2[1]),
    .b(1'b0),
    .c(\add0/c1 ),
    .o({\add0/c2 ,n1[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add0/u2  (
    .a(divider2[2]),
    .b(1'b0),
    .c(\add0/c2 ),
    .o({\add0/c3 ,n1[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add0/u3  (
    .a(divider2[3]),
    .b(1'b0),
    .c(\add0/c3 ),
    .o({\add0/c4 ,n1[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add0/u4  (
    .a(divider2[4]),
    .b(1'b0),
    .c(\add0/c4 ),
    .o({\add0/c5 ,n1[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add0/u5  (
    .a(divider2[5]),
    .b(1'b0),
    .c(\add0/c5 ),
    .o({\add0/c6 ,n1[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add0/u6  (
    .a(divider2[6]),
    .b(1'b0),
    .c(\add0/c6 ),
    .o({\add0/c7 ,n1[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add0/u7  (
    .a(divider2[7]),
    .b(1'b0),
    .c(\add0/c7 ),
    .o({open_n17,n1[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \add0/ucin  (
    .a(1'b0),
    .o({\add0/c0 ,open_n20}));
  reg_ar_as_w1 clk_div_reg (
    .clk(divider2[7]),
    .d(clk_div_neg),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(n28));  // sources/rtl/i2c_module.v(76)
  reg_ar_ss_w1 ready_reg (
    .clk(~divider2[7]),
    .d(n190),
    .en(1'b1),
    .reset(1'b0),
    .set(~reset_n),
    .q(ready));  // sources/rtl/i2c_module.v(1066)
  reg_ar_as_w1 reg0_b0 (
    .clk(clk),
    .d(n1[0]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(divider2[0]));  // sources/rtl/i2c_module.v(81)
  reg_ar_as_w1 reg0_b1 (
    .clk(clk),
    .d(n1[1]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(divider2[1]));  // sources/rtl/i2c_module.v(81)
  reg_ar_as_w1 reg0_b2 (
    .clk(clk),
    .d(n1[2]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(divider2[2]));  // sources/rtl/i2c_module.v(81)
  reg_ar_as_w1 reg0_b3 (
    .clk(clk),
    .d(n1[3]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(divider2[3]));  // sources/rtl/i2c_module.v(81)
  reg_ar_as_w1 reg0_b4 (
    .clk(clk),
    .d(n1[4]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(divider2[4]));  // sources/rtl/i2c_module.v(81)
  reg_ar_as_w1 reg0_b5 (
    .clk(clk),
    .d(n1[5]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(divider2[5]));  // sources/rtl/i2c_module.v(81)
  reg_ar_as_w1 reg0_b6 (
    .clk(clk),
    .d(n1[6]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(divider2[6]));  // sources/rtl/i2c_module.v(81)
  reg_ar_as_w1 reg0_b7 (
    .clk(clk),
    .d(n1[7]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(divider2[7]));  // sources/rtl/i2c_module.v(81)
  reg_sr_as_w1 reg1_b0 (
    .clk(clk),
    .d(writedata[0]),
    .en(mux7_b0_sel_is_3_o),
    .reset(~mux9_b0_sel_is_0_o),
    .set(1'b0),
    .q(control_reg[0]));  // sources/rtl/i2c_module.v(117)
  reg_sr_as_w1 reg2_b0 (
    .clk(clk),
    .d(writedata[0]),
    .en(mux6_b0_sel_is_3_o),
    .reset(n2),
    .set(1'b0),
    .q(slave_address[0]));  // sources/rtl/i2c_module.v(117)
  reg_sr_as_w1 reg2_b1 (
    .clk(clk),
    .d(writedata[1]),
    .en(mux6_b0_sel_is_3_o),
    .reset(n2),
    .set(1'b0),
    .q(slave_address[1]));  // sources/rtl/i2c_module.v(117)
  reg_sr_as_w1 reg2_b2 (
    .clk(clk),
    .d(writedata[2]),
    .en(mux6_b0_sel_is_3_o),
    .reset(n2),
    .set(1'b0),
    .q(slave_address[2]));  // sources/rtl/i2c_module.v(117)
  reg_sr_as_w1 reg2_b3 (
    .clk(clk),
    .d(writedata[3]),
    .en(mux6_b0_sel_is_3_o),
    .reset(n2),
    .set(1'b0),
    .q(slave_address[3]));  // sources/rtl/i2c_module.v(117)
  reg_sr_as_w1 reg2_b4 (
    .clk(clk),
    .d(writedata[4]),
    .en(mux6_b0_sel_is_3_o),
    .reset(n2),
    .set(1'b0),
    .q(slave_address[4]));  // sources/rtl/i2c_module.v(117)
  reg_sr_as_w1 reg2_b5 (
    .clk(clk),
    .d(writedata[5]),
    .en(mux6_b0_sel_is_3_o),
    .reset(n2),
    .set(1'b0),
    .q(slave_address[5]));  // sources/rtl/i2c_module.v(117)
  reg_sr_as_w1 reg2_b6 (
    .clk(clk),
    .d(writedata[6]),
    .en(mux6_b0_sel_is_3_o),
    .reset(n2),
    .set(1'b0),
    .q(slave_address[6]));  // sources/rtl/i2c_module.v(117)
  reg_sr_as_w1 reg2_b7 (
    .clk(clk),
    .d(writedata[7]),
    .en(mux6_b0_sel_is_3_o),
    .reset(n2),
    .set(1'b0),
    .q(slave_address[7]));  // sources/rtl/i2c_module.v(117)
  reg_sr_as_w1 reg3_b0 (
    .clk(clk),
    .d(writedata[0]),
    .en(mux5_b0_sel_is_3_o),
    .reset(n2),
    .set(1'b0),
    .q(slave_reg_address[0]));  // sources/rtl/i2c_module.v(117)
  reg_sr_as_w1 reg3_b1 (
    .clk(clk),
    .d(writedata[1]),
    .en(mux5_b0_sel_is_3_o),
    .reset(n2),
    .set(1'b0),
    .q(slave_reg_address[1]));  // sources/rtl/i2c_module.v(117)
  reg_sr_as_w1 reg3_b2 (
    .clk(clk),
    .d(writedata[2]),
    .en(mux5_b0_sel_is_3_o),
    .reset(n2),
    .set(1'b0),
    .q(slave_reg_address[2]));  // sources/rtl/i2c_module.v(117)
  reg_sr_as_w1 reg3_b3 (
    .clk(clk),
    .d(writedata[3]),
    .en(mux5_b0_sel_is_3_o),
    .reset(n2),
    .set(1'b0),
    .q(slave_reg_address[3]));  // sources/rtl/i2c_module.v(117)
  reg_sr_as_w1 reg3_b4 (
    .clk(clk),
    .d(writedata[4]),
    .en(mux5_b0_sel_is_3_o),
    .reset(n2),
    .set(1'b0),
    .q(slave_reg_address[4]));  // sources/rtl/i2c_module.v(117)
  reg_sr_as_w1 reg3_b5 (
    .clk(clk),
    .d(writedata[5]),
    .en(mux5_b0_sel_is_3_o),
    .reset(n2),
    .set(1'b0),
    .q(slave_reg_address[5]));  // sources/rtl/i2c_module.v(117)
  reg_sr_as_w1 reg3_b6 (
    .clk(clk),
    .d(writedata[6]),
    .en(mux5_b0_sel_is_3_o),
    .reset(n2),
    .set(1'b0),
    .q(slave_reg_address[6]));  // sources/rtl/i2c_module.v(117)
  reg_sr_as_w1 reg3_b7 (
    .clk(clk),
    .d(writedata[7]),
    .en(mux5_b0_sel_is_3_o),
    .reset(n2),
    .set(1'b0),
    .q(slave_reg_address[7]));  // sources/rtl/i2c_module.v(117)
  reg_sr_as_w1 reg4_b0 (
    .clk(clk),
    .d(writedata[0]),
    .en(mux4_b0_sel_is_3_o),
    .reset(n2),
    .set(1'b0),
    .q(slave_data_1[0]));  // sources/rtl/i2c_module.v(117)
  reg_sr_as_w1 reg4_b1 (
    .clk(clk),
    .d(writedata[1]),
    .en(mux4_b0_sel_is_3_o),
    .reset(n2),
    .set(1'b0),
    .q(slave_data_1[1]));  // sources/rtl/i2c_module.v(117)
  reg_sr_as_w1 reg4_b2 (
    .clk(clk),
    .d(writedata[2]),
    .en(mux4_b0_sel_is_3_o),
    .reset(n2),
    .set(1'b0),
    .q(slave_data_1[2]));  // sources/rtl/i2c_module.v(117)
  reg_sr_as_w1 reg4_b3 (
    .clk(clk),
    .d(writedata[3]),
    .en(mux4_b0_sel_is_3_o),
    .reset(n2),
    .set(1'b0),
    .q(slave_data_1[3]));  // sources/rtl/i2c_module.v(117)
  reg_sr_as_w1 reg4_b4 (
    .clk(clk),
    .d(writedata[4]),
    .en(mux4_b0_sel_is_3_o),
    .reset(n2),
    .set(1'b0),
    .q(slave_data_1[4]));  // sources/rtl/i2c_module.v(117)
  reg_sr_as_w1 reg4_b5 (
    .clk(clk),
    .d(writedata[5]),
    .en(mux4_b0_sel_is_3_o),
    .reset(n2),
    .set(1'b0),
    .q(slave_data_1[5]));  // sources/rtl/i2c_module.v(117)
  reg_sr_as_w1 reg4_b6 (
    .clk(clk),
    .d(writedata[6]),
    .en(mux4_b0_sel_is_3_o),
    .reset(n2),
    .set(1'b0),
    .q(slave_data_1[6]));  // sources/rtl/i2c_module.v(117)
  reg_sr_as_w1 reg4_b7 (
    .clk(clk),
    .d(writedata[7]),
    .en(mux4_b0_sel_is_3_o),
    .reset(n2),
    .set(1'b0),
    .q(slave_data_1[7]));  // sources/rtl/i2c_module.v(117)
  reg_sr_as_w1 reg5_b0 (
    .clk(~divider2[7]),
    .d(n99[0]),
    .en(1'b1),
    .reset(n2),
    .set(1'b0),
    .q(state_next[0]));  // sources/rtl/i2c_module.v(510)
  reg_sr_as_w1 reg5_b1 (
    .clk(~divider2[7]),
    .d(n99[1]),
    .en(1'b1),
    .reset(n2),
    .set(1'b0),
    .q(state_next[1]));  // sources/rtl/i2c_module.v(510)
  reg_sr_as_w1 reg5_b2 (
    .clk(~divider2[7]),
    .d(n99[2]),
    .en(1'b1),
    .reset(n2),
    .set(1'b0),
    .q(state_next[2]));  // sources/rtl/i2c_module.v(510)
  reg_sr_as_w1 reg5_b3 (
    .clk(~divider2[7]),
    .d(n99[3]),
    .en(1'b1),
    .reset(n2),
    .set(1'b0),
    .q(state_next[3]));  // sources/rtl/i2c_module.v(510)
  reg_sr_as_w1 reg5_b4 (
    .clk(~divider2[7]),
    .d(n99[4]),
    .en(1'b1),
    .reset(n2),
    .set(1'b0),
    .q(state_next[4]));  // sources/rtl/i2c_module.v(510)
  reg_sr_as_w1 reg5_b5 (
    .clk(~divider2[7]),
    .d(n99[5]),
    .en(1'b1),
    .reset(n2),
    .set(1'b0),
    .q(state_next[5]));  // sources/rtl/i2c_module.v(510)
  reg_sr_as_w1 reg5_b6 (
    .clk(~divider2[7]),
    .d(n99[6]),
    .en(1'b1),
    .reset(n2),
    .set(1'b0),
    .q(state_next[6]));  // sources/rtl/i2c_module.v(510)
  reg_sr_as_w1 reg5_b7 (
    .clk(~divider2[7]),
    .d(n99[7]),
    .en(1'b1),
    .reset(n2),
    .set(1'b0),
    .q(state_next[7]));  // sources/rtl/i2c_module.v(510)
  reg_ar_as_w1 scl_out_reg (
    .clk(divider2[7]),
    .d(n20),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(scl_out_pad));  // sources/rtl/i2c_module.v(137)
  reg_sr_as_w1 scl_output_enable_reg (
    .clk(~divider2[7]),
    .d(n188),
    .en(1'b1),
    .reset(~reset_n),
    .set(1'b0),
    .q(scl_output_enable));  // sources/rtl/i2c_module.v(1066)
  reg_ar_as_w1 scl_output_zero_reg (
    .clk(~divider2[7]),
    .d(n194),
    .en(~n2),
    .reset(1'b0),
    .set(1'b0),
    .q(scl_output_zero));  // sources/rtl/i2c_module.v(1066)
  reg_ar_ss_w1 sda_oe_reg (
    .clk(~divider2[7]),
    .d(n186),
    .en(1'b1),
    .reset(1'b0),
    .set(~reset_n),
    .q(sda_oe));  // sources/rtl/i2c_module.v(1066)
  reg_ar_ss_w1 sda_reg (
    .clk(~divider2[7]),
    .d(n184),
    .en(1'b1),
    .reset(1'b0),
    .set(~reset_n),
    .q(sda));  // sources/rtl/i2c_module.v(1066)
  reg_ar_as_w1 success_out_reg (
    .clk(~divider2[7]),
    .d(n33),
    .en(n28),
    .reset(1'b0),
    .set(1'b0),
    .q(success_out));  // sources/rtl/i2c_module.v(167)
  reg_sr_as_w1 success_reg (
    .clk(~divider2[7]),
    .d(n192),
    .en(1'b1),
    .reset(~reset_n),
    .set(1'b0),
    .q(success));  // sources/rtl/i2c_module.v(1066)

endmodule 

module reg_ar_ss_w1
  (
  clk,
  d,
  en,
  reset,
  set,
  q
  );

  input clk;
  input d;
  input en;
  input reset;
  input set;
  output q;

  parameter REGSET = "RESET";
  wire enout;
  wire setout;

  AL_MUX u_en0 (
    .i0(q),
    .i1(d),
    .sel(en),
    .o(enout));
  AL_DFF #(
    .INI((REGSET == "SET") ? 1'b1 : 1'b0))
    u_seq0 (
    .clk(clk),
    .d(setout),
    .reset(reset),
    .set(1'b0),
    .q(q));
  AL_MUX u_set0 (
    .i0(enout),
    .i1(1'b1),
    .sel(set),
    .o(setout));

endmodule 

module AL_MUX
  (
  input i0,
  input i1,
  input sel,
  output o
  );

  wire not_sel, sel_i0, sel_i1;
  not u0 (not_sel, sel);
  and u1 (sel_i1, sel, i1);
  and u2 (sel_i0, not_sel, i0);
  or u3 (o, sel_i1, sel_i0);

endmodule

module AL_DFF
  (
  input reset,
  input set,
  input clk,
  input d,
  output reg q
  );

  parameter INI = 1'b0;

  always @(posedge reset or posedge set or posedge clk)
  begin
    if (reset)
      q <= 1'b0;
    else if (set)
      q <= 1'b1;
    else
      q <= d;
  end

endmodule

