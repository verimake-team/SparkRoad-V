`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company:        anlogic
// Engineer:       liguang
// 
// Create Date:    14:07:14 11/19/2014 
// Design Name: 
// Module Name:    DP_1024X8_1024X8
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments:  
//
//////////////////////////////////////////////////////////////////////////////////
module DP_1024X8_1024X8 (DataInA, DataInB, AddressA, AddressB, ClockA, ClockB, WrA, WrB, ResetA, ResetB, QA, QB);
    input wire [7:0] DataInA;
    input wire [7:0] DataInB;
    input wire [9:0] AddressA;
    input wire [9:0] AddressB;
    input wire ClockA;
    input wire ClockB;
    input wire WrA;
    input wire WrB;
    input wire ResetA;
    input wire ResetB;
    output wire [7:0] QA;
    output wire [7:0] QB;

    wire [8:0] doa_0,dob_0;
    
    AL_PHY_BRAM  RAM_01 (
        .dia({1'b0,DataInA[7:0]}),
        .addra({AddressA,3'b111}),
        .cea(1'b1), 
        .ocea(1'b1),
        .clka(ClockA),
        .wea(WrA),
        .csa(3'b111),
        .rsta(ResetA),
        .dib({1'b0,DataInB[7:0]}),
        .addrb({AddressB,3'b111}),
        .ceb(1'b1), 
        .oceb(1'b1), 
        .clkb(ClockB), 
        .web(WrB), 
        .csb(3'b111),
        .rstb(ResetB),
        .doa(doa_0), 
        .dob(dob_0));

    defparam RAM_01.DATA_WIDTH_A = "9" ; // 1, 2, 4, 9, 18
    defparam RAM_01.DATA_WIDTH_B = "9" ; // 1, 2, 4, 9, 18    
    defparam RAM_01.INIT_1F = 256'h543210FEDCBA9876BA9876543210FEDCBA9876543210FEDCBA9876543210FEDC;
    defparam RAM_01.INIT_1E = 256'hFEDCBA9876543210FEDCBA9876543210543210FEDCBA9876543210FEDCBA9876;
    defparam RAM_01.INIT_1D = 256'hFEDCBA9876543210FEDCBA9876543210FEDCBA9876543210FEDCBA9876543210;
    defparam RAM_01.INIT_1C = 256'hBA9876543210FEDC543210FEDCBA9876543210FEDCBA9876543210FEDCBA9876;
    defparam RAM_01.INIT_1B = 256'hFEDCBA9876543210FEDCBA9876543210BA9876543210FEDCBA9876543210FEDC;
    defparam RAM_01.INIT_1A = 256'h543210FEDCBA9876543210FEDCBA9876543210FEDCBA9876FEDCBA9876543210;
    defparam RAM_01.INIT_19 = 256'hFEDCBA9876543210BA9876543210FEDCBA9876543210FEDCBA9876543210FEDC;
    defparam RAM_01.INIT_18 = 256'h543210FEDCBA9876543210FEDCBA9876FEDCBA9876543210FEDCBA9876543210;
    defparam RAM_01.INIT_17 = 256'hBA9876543210FEDCBA9876543210FEDCBA9876543210FEDC543210FEDCBA9876;
    defparam RAM_01.INIT_16 = 256'h543210FEDCBA9876FEDCBA9876543210FEDCBA9876543210FEDCBA9876543210;
    defparam RAM_01.INIT_15 = 256'hBA9876543210FEDCBA9876543210FEDC543210FEDCBA9876543210FEDCBA9876;
    defparam RAM_01.INIT_14 = 256'hFEDCBA9876543210FEDCBA9876543210FEDCBA9876543210BA9876543210FEDC;
    defparam RAM_01.INIT_13 = 256'hBA9876543210FEDC543210FEDCBA9876543210FEDCBA9876543210FEDCBA9876;
    defparam RAM_01.INIT_12 = 256'hFEDCBA9876543210FEDCBA9876543210BA9876543210FEDCBA9876543210FEDC;
    defparam RAM_01.INIT_11 = 256'h543210FEDCBA9876543210FEDCBA9876543210FEDCBA9876FEDCBA9876543210;
    defparam RAM_01.INIT_10 = 256'hFEDCBA9876543210BA9876543210FEDCBA9876543210FEDCBA9876543210FEDC;
    defparam RAM_01.INIT_0F = 256'h543210FEDCBA9876543210FEDCBA9876FEDCBA9876543210FEDCBA9876543210;
    defparam RAM_01.INIT_0E = 256'hBA9876543210FEDCBA9876543210FEDCBA9876543210FEDC543210FEDCBA9876;
    defparam RAM_01.INIT_0D = 256'h543210FEDCBA9876FEDCBA9876543210FEDCBA9876543210FEDCBA9876543210;
    defparam RAM_01.INIT_0C = 256'hBA9876543210FEDCBA9876543210FEDC543210FEDCBA9876543210FEDCBA9876;
    defparam RAM_01.INIT_0B = 256'hFEDCBA9876543210FEDCBA9876543210FEDCBA9876543210BA9876543210FEDC;
    defparam RAM_01.INIT_0A = 256'hBA9876543210FEDC543210FEDCBA9876543210FEDCBA9876543210FEDCBA9876;
    defparam RAM_01.INIT_09 = 256'hFEDCBA9876543210FEDCBA9876543210BA9876543210FEDCBA9876543210FEDC;
    defparam RAM_01.INIT_08 = 256'h543210FEDCBA9876543210FEDCBA9876543210FEDCBA9876FEDCBA9876543210;
    defparam RAM_01.INIT_07 = 256'hFEDCBA9876543210BA9876543210FEDCBA9876543210FEDCBA9876543210FEDC;
    defparam RAM_01.INIT_06 = 256'h543210FEDCBA9876543210FEDCBA9876FEDCBA9876543210FEDCBA9876543210;
    defparam RAM_01.INIT_05 = 256'hBA9876543210FEDCBA9876543210FEDCBA9876543210FEDC543210FEDCBA9876;
    defparam RAM_01.INIT_04 = 256'h543210FEDCBA9876FEDCBA9876543210FEDCBA9876543210FEDCBA9876543210;
    defparam RAM_01.INIT_03 = 256'hBA9876543210FEDCBA9876543210FEDC543210FEDCBA9876543210FEDCBA9876;
    defparam RAM_01.INIT_02 = 256'hFEDCBA9876543210FEDCBA9876543210FEDCBA9876543210BA9876543210FEDC;
    defparam RAM_01.INIT_01 = 256'hBA9876543210FEDC543210FEDCBA9876543210FEDCBA9876543210FEDCBA9876;
    defparam RAM_01.INIT_00 = 256'hFEDCBA9876543210FEDCBA9876543210BA9876543210FEDCBA9876543210FEDC;
 //  defparam RAM_01.INIT_FILE    = "tt.mif";
    
    assign QA = doa_0[7:0];
    assign QB = dob_0[7:0];

endmodule