// 译码模块宏定义

`define null_cmd         0
`define wt_a_cmd         1
`define wt_b_cmd         2
`define wt_c_cmd         3
`define wt_d_cmd         4
`define wt_a_rt_cmd      5
`define wt_b_rt_cmd      6
`define wt_c_rt_cmd      7
`define wt_d_rt_cmd      8
`define wt_a_bt_cmd      9
`define wt_b_bt_cmd      10
`define wt_c_bt_cmd      11
`define wt_d_bt_cmd      12
`define wt_pc_cmd        13
`define wt_timer_cmd     14  
`define ex_alua_cmd      15
`define ex_alub_cmd      16
`define ex_aluc_cmd      17
`define ex_alud_cmd      18
`define ex_alue_cmd      19
`define ex_aluf_cmd      20
`define ex_alug_cmd      21
`define ex_aluh_cmd      22
`define ex_alui_cmd      23
`define ex_aluj_cmd      24
`define ex_aluk_cmd      25
`define wt_bus_cmd       26
`define rd_bus_cmd       27
`define rd_ram_cmd       28
`define wt_ram_a_cmd     29
`define wt_ram_b_cmd     30
`define wt_ram_c_cmd     31
`define wt_ram_alu0_cmd  32
`define wt_ram_alu1_cmd  33
`define wt_ram_alu2_cmd  34
`define wt_ram_alu3_cmd  35
`define wt_ram_alu4_cmd  36
`define wt_ram_alu5_cmd  37
`define wt_ram_alu6_cmd  38 
`define dbg_info_cmd     39
