// Verilog netlist created by TD v4.6.12906
// Mon Jul 29 11:23:12 2019

`timescale 1ns / 1ps
module camera  // sources/rtl/test_camera.v(2)
  (
  CLK_IN,
  CSI_D,
  CSI_HREF,
  CSI_PCLK,
  CSI_VSYNC,
  RST_N,
  B,
  CSI_PWDN,
  CSI_RST,
  CSI_SOIC,
  CSI_XCLK,
  G,
  LCD_CLK,
  LCD_DEN,
  LCD_HSYNC,
  LCD_PWM,
  LCD_VSYNC,
  OD,
  R,
  TESTA,
  TESTB,
  TESTC,
  TESTD,
  TESTE,
  TESTF,
  CSI_SOID
  );

  input CLK_IN;  // sources/rtl/test_camera.v(4)
  input [7:0] CSI_D;  // sources/rtl/test_camera.v(15)
  input CSI_HREF;  // sources/rtl/test_camera.v(9)
  input CSI_PCLK;  // sources/rtl/test_camera.v(7)
  input CSI_VSYNC;  // sources/rtl/test_camera.v(10)
  input RST_N;  // sources/rtl/test_camera.v(5)
  output [7:0] B;  // sources/rtl/test_camera.v(19)
  output CSI_PWDN;  // sources/rtl/test_camera.v(11)
  output CSI_RST;  // sources/rtl/test_camera.v(12)
  output CSI_SOIC;  // sources/rtl/test_camera.v(13)
  output CSI_XCLK;  // sources/rtl/test_camera.v(8)
  output [7:0] G;  // sources/rtl/test_camera.v(18)
  output LCD_CLK;  // sources/rtl/test_camera.v(20)
  output LCD_DEN;  // sources/rtl/test_camera.v(23)
  output LCD_HSYNC;  // sources/rtl/test_camera.v(21)
  output LCD_PWM;  // sources/rtl/test_camera.v(24)
  output LCD_VSYNC;  // sources/rtl/test_camera.v(22)
  output [0:7] OD;  // sources/rtl/test_camera.v(32)
  output [7:0] R;  // sources/rtl/test_camera.v(17)
  output TESTA;  // sources/rtl/test_camera.v(26)
  output TESTB;  // sources/rtl/test_camera.v(27)
  output TESTC;  // sources/rtl/test_camera.v(28)
  output TESTD;  // sources/rtl/test_camera.v(29)
  output TESTE;  // sources/rtl/test_camera.v(30)
  output TESTF;  // sources/rtl/test_camera.v(31)
  inout CSI_SOID;  // sources/rtl/test_camera.v(14)

  wire [7:0] B_pad;  // sources/rtl/test_camera.v(19)
  wire [7:0] G_pad;  // sources/rtl/test_camera.v(18)
  wire [0:7] OD_pad;  // sources/rtl/test_camera.v(32)
  wire [7:0] R_pad;  // sources/rtl/test_camera.v(17)
  wire [19:0] camera_addr;  // sources/rtl/test_camera.v(103)
  wire [15:0] camera_wrdat;  // sources/rtl/test_camera.v(102)
  wire [15:0] lcd_rdaddr;  // sources/rtl/test_camera.v(77)
  wire [0:6] lcd_rdaddr_piped;
  wire [0:6] lcd_rdaddr_piped_piped;
  wire [15:0] \u_cameraReader/current_pixel ;  // sources/rtl/cameraReader.v(40)
  wire [19:0] \u_cameraReader/n21 ;
  wire [19:0] \u_cameraReader/n8 ;
  wire [19:0] \u_cameraReader/n9 ;
  wire [19:0] \u_cameraReader/pixel_counter ;  // sources/rtl/cameraReader.v(19)
  wire [7:0] \u_cameraReader/subpixel ;  // sources/rtl/cameraReader.v(39)
  wire CLK_IN_pad;  // sources/rtl/test_camera.v(4)
  wire CSI_PCLK_pad;  // sources/rtl/test_camera.v(7)
  wire CSI_RST_pad;  // sources/rtl/test_camera.v(12)
  wire CSI_RST_pad_neg;
  wire CSI_VSYNC_pad;  // sources/rtl/test_camera.v(10)
  wire CSI_XCLK_pad;  // sources/rtl/test_camera.v(8)
  wire LCD_CLK_pad;  // sources/rtl/test_camera.v(20)
  wire LCD_DEN_pad;  // sources/rtl/test_camera.v(23)
  wire LCD_HSYNC_pad;  // sources/rtl/test_camera.v(21)
  wire LCD_PWM_pad;  // sources/rtl/test_camera.v(24)
  wire LCD_VSYNC_pad;  // sources/rtl/test_camera.v(22)
  wire TESTA_pad;  // sources/rtl/test_camera.v(26)
  wire TESTB_pad;  // sources/rtl/test_camera.v(27)
  wire _al_u461_o;
  wire _al_u471_o;
  wire _al_u477_o;
  wire _al_u498_o;
  wire _al_u499_o;
  wire _al_u500_o;
  wire _al_u501_o;
  wire _al_u502_o;
  wire _al_u503_o;
  wire _al_u504_o;
  wire _al_u505_o;
  wire _al_u506_o;
  wire _al_u507_o;
  wire _al_u508_o;
  wire _al_u509_o;
  wire _al_u510_o;
  wire _al_u511_o;
  wire _al_u512_o;
  wire _al_u513_o;
  wire _al_u514_o;
  wire _al_u515_o;
  wire _al_u516_o;
  wire _al_u517_o;
  wire _al_u518_o;
  wire _al_u519_o;
  wire _al_u520_o;
  wire _al_u521_o;
  wire _al_u522_o;
  wire _al_u523_o;
  wire _al_u524_o;
  wire _al_u526_o;
  wire _al_u527_o;
  wire _al_u528_o;
  wire _al_u529_o;
  wire _al_u530_o;
  wire _al_u531_o;
  wire _al_u532_o;
  wire _al_u533_o;
  wire _al_u534_o;
  wire _al_u535_o;
  wire _al_u536_o;
  wire _al_u537_o;
  wire _al_u538_o;
  wire _al_u539_o;
  wire _al_u540_o;
  wire _al_u541_o;
  wire _al_u542_o;
  wire _al_u543_o;
  wire _al_u544_o;
  wire _al_u545_o;
  wire _al_u546_o;
  wire _al_u547_o;
  wire _al_u548_o;
  wire _al_u549_o;
  wire _al_u550_o;
  wire _al_u551_o;
  wire _al_u552_o;
  wire _al_u554_o;
  wire _al_u555_o;
  wire _al_u556_o;
  wire _al_u557_o;
  wire _al_u558_o;
  wire _al_u559_o;
  wire _al_u560_o;
  wire _al_u561_o;
  wire _al_u562_o;
  wire _al_u563_o;
  wire _al_u564_o;
  wire _al_u565_o;
  wire _al_u566_o;
  wire _al_u567_o;
  wire _al_u568_o;
  wire _al_u569_o;
  wire _al_u570_o;
  wire _al_u571_o;
  wire _al_u572_o;
  wire _al_u573_o;
  wire _al_u574_o;
  wire _al_u575_o;
  wire _al_u576_o;
  wire _al_u577_o;
  wire _al_u578_o;
  wire _al_u579_o;
  wire _al_u580_o;
  wire _al_u582_o;
  wire _al_u583_o;
  wire _al_u584_o;
  wire _al_u585_o;
  wire _al_u586_o;
  wire _al_u587_o;
  wire _al_u588_o;
  wire _al_u589_o;
  wire _al_u590_o;
  wire _al_u591_o;
  wire _al_u592_o;
  wire _al_u593_o;
  wire _al_u594_o;
  wire _al_u595_o;
  wire _al_u596_o;
  wire _al_u597_o;
  wire _al_u598_o;
  wire _al_u599_o;
  wire _al_u600_o;
  wire _al_u601_o;
  wire _al_u602_o;
  wire _al_u603_o;
  wire _al_u604_o;
  wire _al_u605_o;
  wire _al_u606_o;
  wire _al_u607_o;
  wire _al_u608_o;
  wire _al_u610_o;
  wire _al_u611_o;
  wire _al_u612_o;
  wire _al_u613_o;
  wire _al_u614_o;
  wire _al_u615_o;
  wire _al_u616_o;
  wire _al_u617_o;
  wire _al_u618_o;
  wire _al_u619_o;
  wire _al_u620_o;
  wire _al_u621_o;
  wire _al_u622_o;
  wire _al_u623_o;
  wire _al_u624_o;
  wire _al_u625_o;
  wire _al_u626_o;
  wire _al_u627_o;
  wire _al_u628_o;
  wire _al_u629_o;
  wire _al_u630_o;
  wire _al_u631_o;
  wire _al_u632_o;
  wire _al_u633_o;
  wire _al_u634_o;
  wire _al_u635_o;
  wire _al_u636_o;
  wire _al_u638_o;
  wire _al_u639_o;
  wire _al_u640_o;
  wire _al_u641_o;
  wire _al_u642_o;
  wire _al_u643_o;
  wire _al_u644_o;
  wire _al_u645_o;
  wire _al_u646_o;
  wire _al_u647_o;
  wire _al_u648_o;
  wire _al_u649_o;
  wire _al_u650_o;
  wire _al_u651_o;
  wire _al_u652_o;
  wire _al_u653_o;
  wire _al_u654_o;
  wire _al_u655_o;
  wire _al_u656_o;
  wire _al_u657_o;
  wire _al_u658_o;
  wire _al_u659_o;
  wire _al_u660_o;
  wire _al_u661_o;
  wire _al_u662_o;
  wire _al_u663_o;
  wire _al_u664_o;
  wire _al_u666_o;
  wire _al_u667_o;
  wire _al_u668_o;
  wire _al_u669_o;
  wire _al_u670_o;
  wire _al_u671_o;
  wire _al_u672_o;
  wire _al_u673_o;
  wire _al_u674_o;
  wire _al_u675_o;
  wire _al_u676_o;
  wire _al_u677_o;
  wire _al_u678_o;
  wire _al_u679_o;
  wire _al_u680_o;
  wire _al_u681_o;
  wire _al_u682_o;
  wire _al_u683_o;
  wire _al_u684_o;
  wire _al_u685_o;
  wire _al_u686_o;
  wire _al_u687_o;
  wire _al_u688_o;
  wire _al_u689_o;
  wire _al_u690_o;
  wire _al_u691_o;
  wire _al_u692_o;
  wire _al_u694_o;
  wire _al_u695_o;
  wire _al_u696_o;
  wire _al_u697_o;
  wire _al_u698_o;
  wire _al_u699_o;
  wire _al_u700_o;
  wire _al_u701_o;
  wire _al_u702_o;
  wire _al_u703_o;
  wire _al_u704_o;
  wire _al_u705_o;
  wire _al_u706_o;
  wire _al_u707_o;
  wire _al_u708_o;
  wire _al_u709_o;
  wire _al_u710_o;
  wire _al_u711_o;
  wire _al_u712_o;
  wire _al_u713_o;
  wire _al_u714_o;
  wire _al_u715_o;
  wire _al_u716_o;
  wire _al_u717_o;
  wire _al_u718_o;
  wire _al_u719_o;
  wire _al_u720_o;
  wire _al_u722_o;
  wire _al_u723_o;
  wire _al_u724_o;
  wire _al_u725_o;
  wire _al_u726_o;
  wire _al_u727_o;
  wire _al_u728_o;
  wire _al_u729_o;
  wire _al_u730_o;
  wire _al_u731_o;
  wire _al_u732_o;
  wire _al_u733_o;
  wire _al_u734_o;
  wire _al_u735_o;
  wire _al_u736_o;
  wire _al_u737_o;
  wire _al_u738_o;
  wire _al_u739_o;
  wire _al_u740_o;
  wire _al_u741_o;
  wire _al_u742_o;
  wire _al_u743_o;
  wire _al_u744_o;
  wire _al_u745_o;
  wire _al_u746_o;
  wire _al_u747_o;
  wire _al_u748_o;
  wire _al_u750_o;
  wire _al_u751_o;
  wire _al_u752_o;
  wire _al_u754_o;
  wire _al_u755_o;
  wire _al_u756_o;
  wire _al_u758_o;
  wire _al_u759_o;
  wire _al_u760_o;
  wire _al_u762_o;
  wire _al_u763_o;
  wire _al_u764_o;
  wire _al_u766_o;
  wire _al_u767_o;
  wire _al_u768_o;
  wire _al_u770_o;
  wire _al_u771_o;
  wire _al_u772_o;
  wire _al_u774_o;
  wire _al_u775_o;
  wire _al_u776_o;
  wire \and_Ncamera_addr[11]_o_and_camera_wrreq ;
  wire \and_Ncamera_addr[12]_o ;
  wire \and_Ncamera_addr[12]_o_al_n197 ;
  wire \and_Ncamera_addr[12]_o_al_n228 ;
  wire \and_Ncamera_addr[12]_o_al_n260 ;
  wire \and_Nlcd_rdaddr[11]__o_and_lcd_rden ;
  wire \and_Nlcd_rdaddr[12]__o ;
  wire \and_Nlcd_rdaddr[12]__o_al_n200 ;
  wire \and_Nlcd_rdaddr[12]__o_al_n231 ;
  wire \and_Nlcd_rdaddr[12]__o_al_n263 ;
  wire \and_camera_addr[12]__o ;
  wire \and_camera_addr[12]__o_al_n213 ;
  wire \and_camera_addr[12]__o_al_n244 ;
  wire \and_camera_addr[12]__o_al_n276 ;
  wire \and_lcd_rdaddr[12]_N_o ;
  wire \and_lcd_rdaddr[12]_N_o_al_n247 ;
  wire \and_lcd_rdaddr[12]_l_o ;
  wire \and_lcd_rdaddr[12]_l_o_al_n279 ;
  wire camera_wrreq;  // sources/rtl/test_camera.v(101)
  wire clk_cam;  // sources/rtl/test_camera.v(36)
  wire clk_lcd;  // sources/rtl/test_camera.v(35)
  wire clk_sccb;  // sources/rtl/test_camera.v(37)
  wire lcd_rden;  // sources/rtl/test_camera.v(75)
  wire \pll/clk0_buf ;  // al_ip/ip_pll.v(34)
  wire sda;  // sources/rtl/test_camera.v(49)
  wire sda_oe;  // sources/rtl/test_camera.v(48)
  wire \u_cameraReader/add0/c0 ;
  wire \u_cameraReader/add0/c1 ;
  wire \u_cameraReader/add0/c10 ;
  wire \u_cameraReader/add0/c11 ;
  wire \u_cameraReader/add0/c12 ;
  wire \u_cameraReader/add0/c13 ;
  wire \u_cameraReader/add0/c14 ;
  wire \u_cameraReader/add0/c15 ;
  wire \u_cameraReader/add0/c16 ;
  wire \u_cameraReader/add0/c17 ;
  wire \u_cameraReader/add0/c18 ;
  wire \u_cameraReader/add0/c19 ;
  wire \u_cameraReader/add0/c2 ;
  wire \u_cameraReader/add0/c3 ;
  wire \u_cameraReader/add0/c4 ;
  wire \u_cameraReader/add0/c5 ;
  wire \u_cameraReader/add0/c6 ;
  wire \u_cameraReader/add0/c7 ;
  wire \u_cameraReader/add0/c8 ;
  wire \u_cameraReader/add0/c9 ;
  wire \u_cameraReader/add1/c0 ;
  wire \u_cameraReader/add1/c1 ;
  wire \u_cameraReader/add1/c10 ;
  wire \u_cameraReader/add1/c11 ;
  wire \u_cameraReader/add1/c12 ;
  wire \u_cameraReader/add1/c13 ;
  wire \u_cameraReader/add1/c14 ;
  wire \u_cameraReader/add1/c15 ;
  wire \u_cameraReader/add1/c2 ;
  wire \u_cameraReader/add1/c3 ;
  wire \u_cameraReader/add1/c4 ;
  wire \u_cameraReader/add1/c5 ;
  wire \u_cameraReader/add1/c6 ;
  wire \u_cameraReader/add1/c7 ;
  wire \u_cameraReader/add1/c8 ;
  wire \u_cameraReader/add1/c9 ;
  wire \u_cameraReader/lt0_c0 ;
  wire \u_cameraReader/lt0_c1 ;
  wire \u_cameraReader/lt0_c10 ;
  wire \u_cameraReader/lt0_c11 ;
  wire \u_cameraReader/lt0_c12 ;
  wire \u_cameraReader/lt0_c13 ;
  wire \u_cameraReader/lt0_c14 ;
  wire \u_cameraReader/lt0_c15 ;
  wire \u_cameraReader/lt0_c16 ;
  wire \u_cameraReader/lt0_c17 ;
  wire \u_cameraReader/lt0_c18 ;
  wire \u_cameraReader/lt0_c19 ;
  wire \u_cameraReader/lt0_c2 ;
  wire \u_cameraReader/lt0_c20 ;
  wire \u_cameraReader/lt0_c3 ;
  wire \u_cameraReader/lt0_c4 ;
  wire \u_cameraReader/lt0_c5 ;
  wire \u_cameraReader/lt0_c6 ;
  wire \u_cameraReader/lt0_c7 ;
  wire \u_cameraReader/lt0_c8 ;
  wire \u_cameraReader/lt0_c9 ;
  wire \u_cameraReader/mux12_b0_sel_is_2_o ;
  wire \u_cameraReader/mux14_b0_sel_is_2_o ;
  wire \u_cameraReader/mux15_b0_sel_is_2_o ;
  wire \u_cameraReader/mux6_b0_sel_is_1_o ;
  wire \u_cameraReader/n1 ;
  wire \u_cameraReader/n2 ;
  wire \u_cameraReader/n29 ;
  wire \u_cameraReader/vsync_passed ;  // sources/rtl/cameraReader.v(23)
  wire \u_cameraReader/vsync_passed_d ;
  wire \u_cameraReader/wrclk1 ;  // sources/rtl/cameraReader.v(26)
  wire \u_cameraReader/write_pixel ;  // sources/rtl/cameraReader.v(24)
  wire \uimg/inst_dob_i0_000 ;
  wire \uimg/inst_dob_i0_001 ;
  wire \uimg/inst_dob_i0_002 ;
  wire \uimg/inst_dob_i0_003 ;
  wire \uimg/inst_dob_i0_004 ;
  wire \uimg/inst_dob_i0_005 ;
  wire \uimg/inst_dob_i0_006 ;
  wire \uimg/inst_dob_i0_007 ;
  wire \uimg/inst_dob_i0_008 ;
  wire \uimg/inst_dob_i0_009 ;
  wire \uimg/inst_dob_i0_010 ;
  wire \uimg/inst_dob_i0_011 ;
  wire \uimg/inst_dob_i0_012 ;
  wire \uimg/inst_dob_i0_013 ;
  wire \uimg/inst_dob_i0_014 ;
  wire \uimg/inst_dob_i0_015 ;
  wire \uimg/inst_dob_i10_000 ;
  wire \uimg/inst_dob_i10_001 ;
  wire \uimg/inst_dob_i10_002 ;
  wire \uimg/inst_dob_i10_003 ;
  wire \uimg/inst_dob_i10_004 ;
  wire \uimg/inst_dob_i10_005 ;
  wire \uimg/inst_dob_i10_006 ;
  wire \uimg/inst_dob_i10_007 ;
  wire \uimg/inst_dob_i10_008 ;
  wire \uimg/inst_dob_i12_000 ;
  wire \uimg/inst_dob_i12_001 ;
  wire \uimg/inst_dob_i12_002 ;
  wire \uimg/inst_dob_i12_003 ;
  wire \uimg/inst_dob_i12_004 ;
  wire \uimg/inst_dob_i12_005 ;
  wire \uimg/inst_dob_i12_006 ;
  wire \uimg/inst_dob_i12_007 ;
  wire \uimg/inst_dob_i12_008 ;
  wire \uimg/inst_dob_i14_000 ;
  wire \uimg/inst_dob_i14_001 ;
  wire \uimg/inst_dob_i14_002 ;
  wire \uimg/inst_dob_i14_003 ;
  wire \uimg/inst_dob_i14_004 ;
  wire \uimg/inst_dob_i14_005 ;
  wire \uimg/inst_dob_i14_006 ;
  wire \uimg/inst_dob_i14_007 ;
  wire \uimg/inst_dob_i14_008 ;
  wire \uimg/inst_dob_i16_000 ;
  wire \uimg/inst_dob_i16_001 ;
  wire \uimg/inst_dob_i16_002 ;
  wire \uimg/inst_dob_i16_003 ;
  wire \uimg/inst_dob_i16_004 ;
  wire \uimg/inst_dob_i16_005 ;
  wire \uimg/inst_dob_i16_006 ;
  wire \uimg/inst_dob_i16_007 ;
  wire \uimg/inst_dob_i16_008 ;
  wire \uimg/inst_dob_i16_009 ;
  wire \uimg/inst_dob_i16_010 ;
  wire \uimg/inst_dob_i16_011 ;
  wire \uimg/inst_dob_i16_012 ;
  wire \uimg/inst_dob_i16_013 ;
  wire \uimg/inst_dob_i16_014 ;
  wire \uimg/inst_dob_i16_015 ;
  wire \uimg/inst_dob_i18_000 ;
  wire \uimg/inst_dob_i18_001 ;
  wire \uimg/inst_dob_i18_002 ;
  wire \uimg/inst_dob_i18_003 ;
  wire \uimg/inst_dob_i18_004 ;
  wire \uimg/inst_dob_i18_005 ;
  wire \uimg/inst_dob_i18_006 ;
  wire \uimg/inst_dob_i18_007 ;
  wire \uimg/inst_dob_i18_008 ;
  wire \uimg/inst_dob_i20_000 ;
  wire \uimg/inst_dob_i20_001 ;
  wire \uimg/inst_dob_i20_002 ;
  wire \uimg/inst_dob_i20_003 ;
  wire \uimg/inst_dob_i20_004 ;
  wire \uimg/inst_dob_i20_005 ;
  wire \uimg/inst_dob_i20_006 ;
  wire \uimg/inst_dob_i20_007 ;
  wire \uimg/inst_dob_i20_008 ;
  wire \uimg/inst_dob_i22_000 ;
  wire \uimg/inst_dob_i22_001 ;
  wire \uimg/inst_dob_i22_002 ;
  wire \uimg/inst_dob_i22_003 ;
  wire \uimg/inst_dob_i22_004 ;
  wire \uimg/inst_dob_i22_005 ;
  wire \uimg/inst_dob_i22_006 ;
  wire \uimg/inst_dob_i22_007 ;
  wire \uimg/inst_dob_i22_008 ;
  wire \uimg/inst_dob_i24_000 ;
  wire \uimg/inst_dob_i24_001 ;
  wire \uimg/inst_dob_i24_002 ;
  wire \uimg/inst_dob_i24_003 ;
  wire \uimg/inst_dob_i24_004 ;
  wire \uimg/inst_dob_i24_005 ;
  wire \uimg/inst_dob_i24_006 ;
  wire \uimg/inst_dob_i24_007 ;
  wire \uimg/inst_dob_i24_008 ;
  wire \uimg/inst_dob_i26_000 ;
  wire \uimg/inst_dob_i26_001 ;
  wire \uimg/inst_dob_i26_002 ;
  wire \uimg/inst_dob_i26_003 ;
  wire \uimg/inst_dob_i26_004 ;
  wire \uimg/inst_dob_i26_005 ;
  wire \uimg/inst_dob_i26_006 ;
  wire \uimg/inst_dob_i26_007 ;
  wire \uimg/inst_dob_i26_008 ;
  wire \uimg/inst_dob_i28_000 ;
  wire \uimg/inst_dob_i28_001 ;
  wire \uimg/inst_dob_i28_002 ;
  wire \uimg/inst_dob_i28_003 ;
  wire \uimg/inst_dob_i28_004 ;
  wire \uimg/inst_dob_i28_005 ;
  wire \uimg/inst_dob_i28_006 ;
  wire \uimg/inst_dob_i28_007 ;
  wire \uimg/inst_dob_i28_008 ;
  wire \uimg/inst_dob_i2_000 ;
  wire \uimg/inst_dob_i2_001 ;
  wire \uimg/inst_dob_i2_002 ;
  wire \uimg/inst_dob_i2_003 ;
  wire \uimg/inst_dob_i2_004 ;
  wire \uimg/inst_dob_i2_005 ;
  wire \uimg/inst_dob_i2_006 ;
  wire \uimg/inst_dob_i2_007 ;
  wire \uimg/inst_dob_i2_008 ;
  wire \uimg/inst_dob_i30_000 ;
  wire \uimg/inst_dob_i30_001 ;
  wire \uimg/inst_dob_i30_002 ;
  wire \uimg/inst_dob_i30_003 ;
  wire \uimg/inst_dob_i30_004 ;
  wire \uimg/inst_dob_i30_005 ;
  wire \uimg/inst_dob_i30_006 ;
  wire \uimg/inst_dob_i30_007 ;
  wire \uimg/inst_dob_i30_008 ;
  wire \uimg/inst_dob_i32_000 ;
  wire \uimg/inst_dob_i32_001 ;
  wire \uimg/inst_dob_i32_002 ;
  wire \uimg/inst_dob_i32_003 ;
  wire \uimg/inst_dob_i32_004 ;
  wire \uimg/inst_dob_i32_005 ;
  wire \uimg/inst_dob_i32_006 ;
  wire \uimg/inst_dob_i32_007 ;
  wire \uimg/inst_dob_i32_008 ;
  wire \uimg/inst_dob_i32_009 ;
  wire \uimg/inst_dob_i32_010 ;
  wire \uimg/inst_dob_i32_011 ;
  wire \uimg/inst_dob_i32_012 ;
  wire \uimg/inst_dob_i32_013 ;
  wire \uimg/inst_dob_i32_014 ;
  wire \uimg/inst_dob_i32_015 ;
  wire \uimg/inst_dob_i34_000 ;
  wire \uimg/inst_dob_i34_001 ;
  wire \uimg/inst_dob_i34_002 ;
  wire \uimg/inst_dob_i34_003 ;
  wire \uimg/inst_dob_i34_004 ;
  wire \uimg/inst_dob_i34_005 ;
  wire \uimg/inst_dob_i34_006 ;
  wire \uimg/inst_dob_i34_007 ;
  wire \uimg/inst_dob_i34_008 ;
  wire \uimg/inst_dob_i36_000 ;
  wire \uimg/inst_dob_i36_001 ;
  wire \uimg/inst_dob_i36_002 ;
  wire \uimg/inst_dob_i36_003 ;
  wire \uimg/inst_dob_i36_004 ;
  wire \uimg/inst_dob_i36_005 ;
  wire \uimg/inst_dob_i36_006 ;
  wire \uimg/inst_dob_i36_007 ;
  wire \uimg/inst_dob_i36_008 ;
  wire \uimg/inst_dob_i38_000 ;
  wire \uimg/inst_dob_i38_001 ;
  wire \uimg/inst_dob_i38_002 ;
  wire \uimg/inst_dob_i38_003 ;
  wire \uimg/inst_dob_i38_004 ;
  wire \uimg/inst_dob_i38_005 ;
  wire \uimg/inst_dob_i38_006 ;
  wire \uimg/inst_dob_i38_007 ;
  wire \uimg/inst_dob_i38_008 ;
  wire \uimg/inst_dob_i40_000 ;
  wire \uimg/inst_dob_i40_001 ;
  wire \uimg/inst_dob_i40_002 ;
  wire \uimg/inst_dob_i40_003 ;
  wire \uimg/inst_dob_i40_004 ;
  wire \uimg/inst_dob_i40_005 ;
  wire \uimg/inst_dob_i40_006 ;
  wire \uimg/inst_dob_i40_007 ;
  wire \uimg/inst_dob_i40_008 ;
  wire \uimg/inst_dob_i42_000 ;
  wire \uimg/inst_dob_i42_001 ;
  wire \uimg/inst_dob_i42_002 ;
  wire \uimg/inst_dob_i42_003 ;
  wire \uimg/inst_dob_i42_004 ;
  wire \uimg/inst_dob_i42_005 ;
  wire \uimg/inst_dob_i42_006 ;
  wire \uimg/inst_dob_i42_007 ;
  wire \uimg/inst_dob_i42_008 ;
  wire \uimg/inst_dob_i44_000 ;
  wire \uimg/inst_dob_i44_001 ;
  wire \uimg/inst_dob_i44_002 ;
  wire \uimg/inst_dob_i44_003 ;
  wire \uimg/inst_dob_i44_004 ;
  wire \uimg/inst_dob_i44_005 ;
  wire \uimg/inst_dob_i44_006 ;
  wire \uimg/inst_dob_i44_007 ;
  wire \uimg/inst_dob_i44_008 ;
  wire \uimg/inst_dob_i46_000 ;
  wire \uimg/inst_dob_i46_001 ;
  wire \uimg/inst_dob_i46_002 ;
  wire \uimg/inst_dob_i46_003 ;
  wire \uimg/inst_dob_i46_004 ;
  wire \uimg/inst_dob_i46_005 ;
  wire \uimg/inst_dob_i46_006 ;
  wire \uimg/inst_dob_i46_007 ;
  wire \uimg/inst_dob_i46_008 ;
  wire \uimg/inst_dob_i48_000 ;
  wire \uimg/inst_dob_i48_001 ;
  wire \uimg/inst_dob_i48_002 ;
  wire \uimg/inst_dob_i48_003 ;
  wire \uimg/inst_dob_i48_004 ;
  wire \uimg/inst_dob_i48_005 ;
  wire \uimg/inst_dob_i48_006 ;
  wire \uimg/inst_dob_i48_007 ;
  wire \uimg/inst_dob_i48_008 ;
  wire \uimg/inst_dob_i48_009 ;
  wire \uimg/inst_dob_i48_010 ;
  wire \uimg/inst_dob_i48_011 ;
  wire \uimg/inst_dob_i48_012 ;
  wire \uimg/inst_dob_i48_013 ;
  wire \uimg/inst_dob_i48_014 ;
  wire \uimg/inst_dob_i48_015 ;
  wire \uimg/inst_dob_i4_000 ;
  wire \uimg/inst_dob_i4_001 ;
  wire \uimg/inst_dob_i4_002 ;
  wire \uimg/inst_dob_i4_003 ;
  wire \uimg/inst_dob_i4_004 ;
  wire \uimg/inst_dob_i4_005 ;
  wire \uimg/inst_dob_i4_006 ;
  wire \uimg/inst_dob_i4_007 ;
  wire \uimg/inst_dob_i4_008 ;
  wire \uimg/inst_dob_i50_000 ;
  wire \uimg/inst_dob_i50_001 ;
  wire \uimg/inst_dob_i50_002 ;
  wire \uimg/inst_dob_i50_003 ;
  wire \uimg/inst_dob_i50_004 ;
  wire \uimg/inst_dob_i50_005 ;
  wire \uimg/inst_dob_i50_006 ;
  wire \uimg/inst_dob_i50_007 ;
  wire \uimg/inst_dob_i50_008 ;
  wire \uimg/inst_dob_i52_000 ;
  wire \uimg/inst_dob_i52_001 ;
  wire \uimg/inst_dob_i52_002 ;
  wire \uimg/inst_dob_i52_003 ;
  wire \uimg/inst_dob_i52_004 ;
  wire \uimg/inst_dob_i52_005 ;
  wire \uimg/inst_dob_i52_006 ;
  wire \uimg/inst_dob_i52_007 ;
  wire \uimg/inst_dob_i52_008 ;
  wire \uimg/inst_dob_i54_000 ;
  wire \uimg/inst_dob_i54_001 ;
  wire \uimg/inst_dob_i54_002 ;
  wire \uimg/inst_dob_i54_003 ;
  wire \uimg/inst_dob_i54_004 ;
  wire \uimg/inst_dob_i54_005 ;
  wire \uimg/inst_dob_i54_006 ;
  wire \uimg/inst_dob_i54_007 ;
  wire \uimg/inst_dob_i54_008 ;
  wire \uimg/inst_dob_i56_000 ;
  wire \uimg/inst_dob_i56_001 ;
  wire \uimg/inst_dob_i56_002 ;
  wire \uimg/inst_dob_i56_003 ;
  wire \uimg/inst_dob_i56_004 ;
  wire \uimg/inst_dob_i56_005 ;
  wire \uimg/inst_dob_i56_006 ;
  wire \uimg/inst_dob_i56_007 ;
  wire \uimg/inst_dob_i56_008 ;
  wire \uimg/inst_dob_i58_000 ;
  wire \uimg/inst_dob_i58_001 ;
  wire \uimg/inst_dob_i58_002 ;
  wire \uimg/inst_dob_i58_003 ;
  wire \uimg/inst_dob_i58_004 ;
  wire \uimg/inst_dob_i58_005 ;
  wire \uimg/inst_dob_i58_006 ;
  wire \uimg/inst_dob_i58_007 ;
  wire \uimg/inst_dob_i58_008 ;
  wire \uimg/inst_dob_i60_000 ;
  wire \uimg/inst_dob_i60_001 ;
  wire \uimg/inst_dob_i60_002 ;
  wire \uimg/inst_dob_i60_003 ;
  wire \uimg/inst_dob_i60_004 ;
  wire \uimg/inst_dob_i60_005 ;
  wire \uimg/inst_dob_i60_006 ;
  wire \uimg/inst_dob_i60_007 ;
  wire \uimg/inst_dob_i60_008 ;
  wire \uimg/inst_dob_i62_000 ;
  wire \uimg/inst_dob_i62_001 ;
  wire \uimg/inst_dob_i62_002 ;
  wire \uimg/inst_dob_i62_003 ;
  wire \uimg/inst_dob_i62_004 ;
  wire \uimg/inst_dob_i62_005 ;
  wire \uimg/inst_dob_i62_006 ;
  wire \uimg/inst_dob_i62_007 ;
  wire \uimg/inst_dob_i62_008 ;
  wire \uimg/inst_dob_i64_000 ;
  wire \uimg/inst_dob_i64_001 ;
  wire \uimg/inst_dob_i64_002 ;
  wire \uimg/inst_dob_i64_003 ;
  wire \uimg/inst_dob_i64_004 ;
  wire \uimg/inst_dob_i64_005 ;
  wire \uimg/inst_dob_i64_006 ;
  wire \uimg/inst_dob_i64_007 ;
  wire \uimg/inst_dob_i64_008 ;
  wire \uimg/inst_dob_i64_009 ;
  wire \uimg/inst_dob_i64_010 ;
  wire \uimg/inst_dob_i64_011 ;
  wire \uimg/inst_dob_i64_012 ;
  wire \uimg/inst_dob_i64_013 ;
  wire \uimg/inst_dob_i64_014 ;
  wire \uimg/inst_dob_i64_015 ;
  wire \uimg/inst_dob_i6_000 ;
  wire \uimg/inst_dob_i6_001 ;
  wire \uimg/inst_dob_i6_002 ;
  wire \uimg/inst_dob_i6_003 ;
  wire \uimg/inst_dob_i6_004 ;
  wire \uimg/inst_dob_i6_005 ;
  wire \uimg/inst_dob_i6_006 ;
  wire \uimg/inst_dob_i6_007 ;
  wire \uimg/inst_dob_i6_008 ;
  wire \uimg/inst_dob_i8_000 ;
  wire \uimg/inst_dob_i8_001 ;
  wire \uimg/inst_dob_i8_002 ;
  wire \uimg/inst_dob_i8_003 ;
  wire \uimg/inst_dob_i8_004 ;
  wire \uimg/inst_dob_i8_005 ;
  wire \uimg/inst_dob_i8_006 ;
  wire \uimg/inst_dob_i8_007 ;
  wire \uimg/inst_dob_i8_008 ;

  assign TESTD = TESTC;
  assign TESTE = TESTC;
  assign TESTF = TESTC;
  AL_MAP_LUT1 #(
    //.LOCATION("VIRTUALIO"),
    .EQN("a"),
    .INIT(2'h2))
    LCD_DEN_vio (
    .a(LCD_DEN_pad),
    .o(LCD_DEN));
  AL_MAP_LUT1 #(
    //.LOCATION("VIRTUALIO"),
    .EQN("a"),
    .INIT(2'h2))
    LCD_PWM_vio (
    .a(LCD_PWM_pad),
    .o(LCD_PWM));
  AL_MAP_LUT1 #(
    //.LOCATION("VIRTUALIO"),
    .EQN("a"),
    .INIT(2'h2))
    TESTC_vio (
    .a(1'b0),
    .o(TESTC));
  EG_PHY_PAD #(
    //.LOCATION("C1"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("FAST"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u171 (
    .do({open_n1,open_n2,open_n3,B_pad[7]}),
    .opad(B[7]));  // sources/rtl/test_camera.v(19)
  EG_PHY_PAD #(
    //.LOCATION("D1"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("FAST"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u172 (
    .do({open_n18,open_n19,open_n20,B_pad[6]}),
    .opad(B[6]));  // sources/rtl/test_camera.v(19)
  EG_PHY_PAD #(
    //.LOCATION("E2"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("FAST"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u173 (
    .do({open_n35,open_n36,open_n37,B_pad[5]}),
    .opad(B[5]));  // sources/rtl/test_camera.v(19)
  EG_PHY_PAD #(
    //.LOCATION("G3"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("FAST"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u174 (
    .do({open_n52,open_n53,open_n54,B_pad[4]}),
    .opad(B[4]));  // sources/rtl/test_camera.v(19)
  EG_PHY_PAD #(
    //.LOCATION("E1"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("FAST"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u175 (
    .do({open_n69,open_n70,open_n71,B_pad[3]}),
    .opad(B[3]));  // sources/rtl/test_camera.v(19)
  EG_PHY_PAD #(
    //.LOCATION("F2"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("FAST"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u176 (
    .do({open_n86,open_n87,open_n88,1'b0}),
    .opad(B[2]));  // sources/rtl/test_camera.v(19)
  EG_PHY_PAD #(
    //.LOCATION("F1"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("FAST"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u177 (
    .do({open_n103,open_n104,open_n105,1'b0}),
    .opad(B[1]));  // sources/rtl/test_camera.v(19)
  EG_PHY_PAD #(
    //.LOCATION("G1"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("FAST"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u178 (
    .do({open_n120,open_n121,open_n122,1'b0}),
    .opad(B[0]));  // sources/rtl/test_camera.v(19)
  EG_PHY_PAD #(
    //.LOCATION("K14"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u179 (
    .ipad(CLK_IN),
    .di(CLK_IN_pad));  // sources/rtl/test_camera.v(4)
  EG_PHY_PAD #(
    //.LOCATION("H13"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS33"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u180 (
    .ipad(CSI_D[7]),
    .di(OD_pad[0]));  // sources/rtl/test_camera.v(15)
  EG_PHY_PAD #(
    //.LOCATION("G16"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS33"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u181 (
    .ipad(CSI_D[6]),
    .di(OD_pad[1]));  // sources/rtl/test_camera.v(15)
  EG_PHY_PAD #(
    //.LOCATION("H16"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS33"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u182 (
    .ipad(CSI_D[5]),
    .di(OD_pad[2]));  // sources/rtl/test_camera.v(15)
  EG_PHY_PAD #(
    //.LOCATION("G14"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS33"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u183 (
    .ipad(CSI_D[4]),
    .di(OD_pad[3]));  // sources/rtl/test_camera.v(15)
  EG_PHY_PAD #(
    //.LOCATION("K15"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS33"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u184 (
    .ipad(CSI_D[3]),
    .di(OD_pad[4]));  // sources/rtl/test_camera.v(15)
  EG_PHY_PAD #(
    //.LOCATION("K16"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS33"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u185 (
    .ipad(CSI_D[2]),
    .di(OD_pad[5]));  // sources/rtl/test_camera.v(15)
  EG_PHY_PAD #(
    //.LOCATION("J16"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS33"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u186 (
    .ipad(CSI_D[1]),
    .di(OD_pad[6]));  // sources/rtl/test_camera.v(15)
  EG_PHY_PAD #(
    //.LOCATION("H15"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS33"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u187 (
    .ipad(CSI_D[0]),
    .di(OD_pad[7]));  // sources/rtl/test_camera.v(15)
  EG_PHY_PAD #(
    //.LOCATION("F15"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u188 (
    .ipad(CSI_HREF),
    .di(\u_cameraReader/n2 ));  // sources/rtl/test_camera.v(9)
  EG_PHY_PAD #(
    //.LOCATION("K12"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u189 (
    .ipad(CSI_PCLK),
    .di(CSI_PCLK_pad));  // sources/rtl/test_camera.v(7)
  EG_PHY_PAD #(
    //.LOCATION("F14"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u190 (
    .do({open_n324,open_n325,open_n326,1'b0}),
    .opad(CSI_PWDN));  // sources/rtl/test_camera.v(11)
  EG_PHY_PAD #(
    //.LOCATION("F13"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u191 (
    .do({open_n341,open_n342,open_n343,CSI_RST_pad}),
    .opad(CSI_RST));  // sources/rtl/test_camera.v(12)
  EG_PHY_PAD #(
    //.LOCATION("D16"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u192 (
    .do({open_n358,open_n359,open_n360,TESTB_pad}),
    .opad(CSI_SOIC));  // sources/rtl/test_camera.v(13)
  EG_PHY_PAD #(
    //.LOCATION("D14"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("BI"),
    .TSMUX("INV"))
    _al_u193 (
    .do({open_n375,open_n376,open_n377,sda}),
    .ts(sda_oe),
    .di(TESTA_pad),
    .bpad(CSI_SOID));  // sources/rtl/test_camera.v(63)
  EG_PHY_PAD #(
    //.LOCATION("E15"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u194 (
    .ipad(CSI_VSYNC),
    .di(CSI_VSYNC_pad));  // sources/rtl/test_camera.v(10)
  EG_PHY_PAD #(
    //.LOCATION("J12"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u195 (
    .do({open_n407,open_n408,open_n409,CSI_XCLK_pad}),
    .opad(CSI_XCLK));  // sources/rtl/test_camera.v(8)
  EG_PHY_PAD #(
    //.LOCATION("H5"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u196 (
    .do({open_n424,open_n425,open_n426,G_pad[7]}),
    .opad(G[7]));  // sources/rtl/test_camera.v(18)
  EG_PHY_PAD #(
    //.LOCATION("H1"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u197 (
    .do({open_n441,open_n442,open_n443,G_pad[6]}),
    .opad(G[6]));  // sources/rtl/test_camera.v(18)
  EG_PHY_PAD #(
    //.LOCATION("J6"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u198 (
    .do({open_n458,open_n459,open_n460,G_pad[5]}),
    .opad(G[5]));  // sources/rtl/test_camera.v(18)
  EG_PHY_PAD #(
    //.LOCATION("H3"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u199 (
    .do({open_n475,open_n476,open_n477,G_pad[4]}),
    .opad(G[4]));  // sources/rtl/test_camera.v(18)
  EG_PHY_PAD #(
    //.LOCATION("J1"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u200 (
    .do({open_n492,open_n493,open_n494,G_pad[3]}),
    .opad(G[3]));  // sources/rtl/test_camera.v(18)
  EG_PHY_PAD #(
    //.LOCATION("K1"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u201 (
    .do({open_n509,open_n510,open_n511,G_pad[2]}),
    .opad(G[2]));  // sources/rtl/test_camera.v(18)
  EG_PHY_PAD #(
    //.LOCATION("K2"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u202 (
    .do({open_n526,open_n527,open_n528,1'b0}),
    .opad(G[1]));  // sources/rtl/test_camera.v(18)
  EG_PHY_PAD #(
    //.LOCATION("L1"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u203 (
    .do({open_n543,open_n544,open_n545,1'b0}),
    .opad(G[0]));  // sources/rtl/test_camera.v(18)
  EG_PHY_PAD #(
    //.LOCATION("H2"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u204 (
    .do({open_n560,open_n561,open_n562,LCD_CLK_pad}),
    .opad(LCD_CLK));  // sources/rtl/test_camera.v(20)
  EG_PHY_PAD #(
    //.LOCATION("J3"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u205 (
    .do({open_n577,open_n578,open_n579,LCD_HSYNC_pad}),
    .opad(LCD_HSYNC));  // sources/rtl/test_camera.v(21)
  EG_PHY_PAD #(
    //.LOCATION("J4"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u206 (
    .do({open_n594,open_n595,open_n596,LCD_VSYNC_pad}),
    .opad(LCD_VSYNC));  // sources/rtl/test_camera.v(22)
  EG_PHY_PAD #(
    //.LOCATION("A7"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u207 (
    .do({open_n611,open_n612,open_n613,OD_pad[0]}),
    .opad(OD[0]));  // sources/rtl/test_camera.v(32)
  EG_PHY_PAD #(
    //.LOCATION("A8"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u208 (
    .do({open_n628,open_n629,open_n630,OD_pad[1]}),
    .opad(OD[1]));  // sources/rtl/test_camera.v(32)
  EG_PHY_PAD #(
    //.LOCATION("A10"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u209 (
    .do({open_n645,open_n646,open_n647,OD_pad[2]}),
    .opad(OD[2]));  // sources/rtl/test_camera.v(32)
  EG_PHY_PAD #(
    //.LOCATION("A6"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u210 (
    .do({open_n662,open_n663,open_n664,OD_pad[3]}),
    .opad(OD[3]));  // sources/rtl/test_camera.v(32)
  EG_PHY_PAD #(
    //.LOCATION("A4"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u211 (
    .do({open_n679,open_n680,open_n681,OD_pad[4]}),
    .opad(OD[4]));  // sources/rtl/test_camera.v(32)
  EG_PHY_PAD #(
    //.LOCATION("A12"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u212 (
    .do({open_n696,open_n697,open_n698,OD_pad[5]}),
    .opad(OD[5]));  // sources/rtl/test_camera.v(32)
  EG_PHY_PAD #(
    //.LOCATION("E8"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u213 (
    .do({open_n713,open_n714,open_n715,OD_pad[6]}),
    .opad(OD[6]));  // sources/rtl/test_camera.v(32)
  EG_PHY_PAD #(
    //.LOCATION("A14"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u214 (
    .do({open_n730,open_n731,open_n732,OD_pad[7]}),
    .opad(OD[7]));  // sources/rtl/test_camera.v(32)
  EG_PHY_PAD #(
    //.LOCATION("L5"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u215 (
    .do({open_n747,open_n748,open_n749,R_pad[7]}),
    .opad(R[7]));  // sources/rtl/test_camera.v(17)
  EG_PHY_PAD #(
    //.LOCATION("L3"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u216 (
    .do({open_n764,open_n765,open_n766,R_pad[6]}),
    .opad(R[6]));  // sources/rtl/test_camera.v(17)
  EG_PHY_PAD #(
    //.LOCATION("M2"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u217 (
    .do({open_n781,open_n782,open_n783,R_pad[5]}),
    .opad(R[5]));  // sources/rtl/test_camera.v(17)
  EG_PHY_PAD #(
    //.LOCATION("M1"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u218 (
    .do({open_n798,open_n799,open_n800,R_pad[4]}),
    .opad(R[4]));  // sources/rtl/test_camera.v(17)
  EG_PHY_PAD #(
    //.LOCATION("L4"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u219 (
    .do({open_n815,open_n816,open_n817,R_pad[3]}),
    .opad(R[3]));  // sources/rtl/test_camera.v(17)
  EG_PHY_PAD #(
    //.LOCATION("K5"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u220 (
    .do({open_n832,open_n833,open_n834,1'b0}),
    .opad(R[2]));  // sources/rtl/test_camera.v(17)
  EG_PHY_PAD #(
    //.LOCATION("K3"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u221 (
    .do({open_n849,open_n850,open_n851,1'b0}),
    .opad(R[1]));  // sources/rtl/test_camera.v(17)
  EG_PHY_PAD #(
    //.LOCATION("K6"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u222 (
    .do({open_n866,open_n867,open_n868,1'b0}),
    .opad(R[0]));  // sources/rtl/test_camera.v(17)
  EG_PHY_PAD #(
    //.LOCATION("G11"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u223 (
    .ipad(RST_N),
    .di(CSI_RST_pad));  // sources/rtl/test_camera.v(5)
  EG_PHY_PAD #(
    //.LOCATION("A5"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u224 (
    .do({open_n900,open_n901,open_n902,TESTA_pad}),
    .opad(TESTA));  // sources/rtl/test_camera.v(26)
  EG_PHY_PAD #(
    //.LOCATION("A9"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u225 (
    .do({open_n917,open_n918,open_n919,TESTB_pad}),
    .opad(TESTB));  // sources/rtl/test_camera.v(27)
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*A)"),
    .INIT(16'h0080))
    _al_u454 (
    .a(camera_addr[12]),
    .b(camera_addr[13]),
    .c(camera_addr[14]),
    .d(camera_addr[15]),
    .o(\and_camera_addr[12]__o_al_n276 ));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*~B*A)"),
    .INIT(16'h0020))
    _al_u455 (
    .a(camera_addr[12]),
    .b(camera_addr[13]),
    .c(camera_addr[14]),
    .d(camera_addr[15]),
    .o(\and_camera_addr[12]__o_al_n244 ));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    _al_u456 (
    .a(camera_addr[12]),
    .b(camera_addr[13]),
    .c(camera_addr[14]),
    .d(camera_addr[15]),
    .o(\and_camera_addr[12]__o_al_n213 ));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*A)"),
    .INIT(16'h0002))
    _al_u457 (
    .a(camera_addr[12]),
    .b(camera_addr[13]),
    .c(camera_addr[14]),
    .d(camera_addr[15]),
    .o(\and_camera_addr[12]__o ));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*~A)"),
    .INIT(16'h0040))
    _al_u458 (
    .a(camera_addr[12]),
    .b(camera_addr[13]),
    .c(camera_addr[14]),
    .d(camera_addr[15]),
    .o(\and_Ncamera_addr[12]_o_al_n260 ));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*~B*~A)"),
    .INIT(16'h0010))
    _al_u459 (
    .a(camera_addr[12]),
    .b(camera_addr[13]),
    .c(camera_addr[14]),
    .d(camera_addr[15]),
    .o(\and_Ncamera_addr[12]_o_al_n228 ));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*~A)"),
    .INIT(16'h0004))
    _al_u460 (
    .a(camera_addr[12]),
    .b(camera_addr[13]),
    .c(camera_addr[14]),
    .d(camera_addr[15]),
    .o(\and_Ncamera_addr[12]_o_al_n197 ));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u461 (
    .a(camera_addr[12]),
    .b(camera_addr[13]),
    .c(camera_addr[14]),
    .o(_al_u461_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u462 (
    .a(_al_u461_o),
    .b(camera_addr[15]),
    .o(\and_Ncamera_addr[12]_o ));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*~A)"),
    .INIT(16'h4000))
    _al_u463 (
    .a(lcd_rdaddr[15]),
    .b(lcd_rdaddr[14]),
    .c(lcd_rdaddr[13]),
    .d(lcd_rdaddr[12]),
    .o(\and_lcd_rdaddr[12]_l_o_al_n279 ));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*~A)"),
    .INIT(16'h1000))
    _al_u464 (
    .a(lcd_rdaddr[15]),
    .b(lcd_rdaddr[14]),
    .c(lcd_rdaddr[13]),
    .d(lcd_rdaddr[12]),
    .o(\and_lcd_rdaddr[12]_l_o ));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*B*~A)"),
    .INIT(16'h0400))
    _al_u465 (
    .a(lcd_rdaddr[15]),
    .b(lcd_rdaddr[14]),
    .c(lcd_rdaddr[13]),
    .d(lcd_rdaddr[12]),
    .o(\and_lcd_rdaddr[12]_N_o_al_n247 ));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*~A)"),
    .INIT(16'h0100))
    _al_u466 (
    .a(lcd_rdaddr[15]),
    .b(lcd_rdaddr[14]),
    .c(lcd_rdaddr[13]),
    .d(lcd_rdaddr[12]),
    .o(\and_lcd_rdaddr[12]_N_o ));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*~A)"),
    .INIT(16'h0040))
    _al_u467 (
    .a(lcd_rdaddr[15]),
    .b(lcd_rdaddr[14]),
    .c(lcd_rdaddr[13]),
    .d(lcd_rdaddr[12]),
    .o(\and_Nlcd_rdaddr[12]__o_al_n263 ));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*~A)"),
    .INIT(16'h0004))
    _al_u468 (
    .a(lcd_rdaddr[15]),
    .b(lcd_rdaddr[14]),
    .c(lcd_rdaddr[13]),
    .d(lcd_rdaddr[12]),
    .o(\and_Nlcd_rdaddr[12]__o_al_n231 ));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*~B*~A)"),
    .INIT(16'h0010))
    _al_u469 (
    .a(lcd_rdaddr[15]),
    .b(lcd_rdaddr[14]),
    .c(lcd_rdaddr[13]),
    .d(lcd_rdaddr[12]),
    .o(\and_Nlcd_rdaddr[12]__o_al_n200 ));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u470 (
    .a(lcd_rdaddr[15]),
    .b(lcd_rdaddr[14]),
    .c(lcd_rdaddr[13]),
    .d(lcd_rdaddr[12]),
    .o(\and_Nlcd_rdaddr[12]__o ));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*A)"),
    .INIT(16'h0200))
    _al_u471 (
    .a(lcd_rdaddr[15]),
    .b(lcd_rdaddr[14]),
    .c(lcd_rdaddr[11]),
    .d(lcd_rden),
    .o(_al_u471_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u472 (
    .a(_al_u471_o),
    .b(lcd_rdaddr[13]),
    .c(lcd_rdaddr[12]),
    .o(\and_Nlcd_rdaddr[11]__o_and_lcd_rden ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u473 (
    .a(CSI_RST_pad),
    .b(clk_cam),
    .o(CSI_XCLK_pad));
  AL_MAP_LUT2 #(
    .EQN("~(~B*A)"),
    .INIT(4'hd))
    _al_u474 (
    .a(CSI_VSYNC_pad),
    .b(\u_cameraReader/vsync_passed ),
    .o(\u_cameraReader/vsync_passed_d ));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u475 (
    .a(\u_cameraReader/n29 ),
    .b(\u_cameraReader/wrclk1 ),
    .c(\u_cameraReader/write_pixel ),
    .o(camera_wrreq));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*B*A)"),
    .INIT(16'h0800))
    _al_u476 (
    .a(_al_u461_o),
    .b(camera_wrreq),
    .c(camera_addr[11]),
    .d(camera_addr[15]),
    .o(\and_Ncamera_addr[11]_o_and_camera_wrreq ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u477 (
    .a(\u_cameraReader/n2 ),
    .b(\u_cameraReader/vsync_passed ),
    .o(_al_u477_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u478 (
    .a(_al_u477_o),
    .b(\u_cameraReader/pixel_counter [0]),
    .o(\u_cameraReader/mux6_b0_sel_is_1_o ));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u479 (
    .a(\u_cameraReader/mux6_b0_sel_is_1_o ),
    .b(CSI_VSYNC_pad),
    .c(\u_cameraReader/n9 [9]),
    .d(camera_addr[9]),
    .o(\u_cameraReader/n21 [9]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u480 (
    .a(\u_cameraReader/mux6_b0_sel_is_1_o ),
    .b(CSI_VSYNC_pad),
    .c(\u_cameraReader/n9 [8]),
    .d(camera_addr[8]),
    .o(\u_cameraReader/n21 [8]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u481 (
    .a(\u_cameraReader/mux6_b0_sel_is_1_o ),
    .b(CSI_VSYNC_pad),
    .c(\u_cameraReader/n9 [7]),
    .d(camera_addr[7]),
    .o(\u_cameraReader/n21 [7]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u482 (
    .a(\u_cameraReader/mux6_b0_sel_is_1_o ),
    .b(CSI_VSYNC_pad),
    .c(\u_cameraReader/n9 [6]),
    .d(camera_addr[6]),
    .o(\u_cameraReader/n21 [6]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u483 (
    .a(\u_cameraReader/mux6_b0_sel_is_1_o ),
    .b(CSI_VSYNC_pad),
    .c(\u_cameraReader/n9 [5]),
    .d(camera_addr[5]),
    .o(\u_cameraReader/n21 [5]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u484 (
    .a(\u_cameraReader/mux6_b0_sel_is_1_o ),
    .b(CSI_VSYNC_pad),
    .c(\u_cameraReader/n9 [4]),
    .d(camera_addr[4]),
    .o(\u_cameraReader/n21 [4]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u485 (
    .a(\u_cameraReader/mux6_b0_sel_is_1_o ),
    .b(CSI_VSYNC_pad),
    .c(\u_cameraReader/n9 [3]),
    .d(camera_addr[3]),
    .o(\u_cameraReader/n21 [3]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u486 (
    .a(\u_cameraReader/mux6_b0_sel_is_1_o ),
    .b(CSI_VSYNC_pad),
    .c(\u_cameraReader/n9 [2]),
    .d(camera_addr[2]),
    .o(\u_cameraReader/n21 [2]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u487 (
    .a(\u_cameraReader/mux6_b0_sel_is_1_o ),
    .b(CSI_VSYNC_pad),
    .c(\u_cameraReader/n9 [1]),
    .d(camera_addr[1]),
    .o(\u_cameraReader/n21 [1]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u488 (
    .a(\u_cameraReader/mux6_b0_sel_is_1_o ),
    .b(CSI_VSYNC_pad),
    .c(\u_cameraReader/n9 [15]),
    .d(camera_addr[15]),
    .o(\u_cameraReader/n21 [15]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u489 (
    .a(\u_cameraReader/mux6_b0_sel_is_1_o ),
    .b(CSI_VSYNC_pad),
    .c(\u_cameraReader/n9 [14]),
    .d(camera_addr[14]),
    .o(\u_cameraReader/n21 [14]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u490 (
    .a(\u_cameraReader/mux6_b0_sel_is_1_o ),
    .b(CSI_VSYNC_pad),
    .c(\u_cameraReader/n9 [13]),
    .d(camera_addr[13]),
    .o(\u_cameraReader/n21 [13]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u491 (
    .a(\u_cameraReader/mux6_b0_sel_is_1_o ),
    .b(CSI_VSYNC_pad),
    .c(\u_cameraReader/n9 [12]),
    .d(camera_addr[12]),
    .o(\u_cameraReader/n21 [12]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u492 (
    .a(\u_cameraReader/mux6_b0_sel_is_1_o ),
    .b(CSI_VSYNC_pad),
    .c(\u_cameraReader/n9 [11]),
    .d(camera_addr[11]),
    .o(\u_cameraReader/n21 [11]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u493 (
    .a(\u_cameraReader/mux6_b0_sel_is_1_o ),
    .b(CSI_VSYNC_pad),
    .c(\u_cameraReader/n9 [10]),
    .d(camera_addr[10]),
    .o(\u_cameraReader/n21 [10]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u494 (
    .a(\u_cameraReader/mux6_b0_sel_is_1_o ),
    .b(CSI_VSYNC_pad),
    .c(\u_cameraReader/n9 [0]),
    .d(camera_addr[0]),
    .o(\u_cameraReader/n21 [0]));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u495 (
    .a(\u_cameraReader/mux6_b0_sel_is_1_o ),
    .b(CSI_VSYNC_pad),
    .c(CSI_RST_pad),
    .o(\u_cameraReader/mux15_b0_sel_is_2_o ));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*A)"),
    .INIT(16'h0080))
    _al_u496 (
    .a(_al_u477_o),
    .b(CSI_VSYNC_pad),
    .c(CSI_RST_pad),
    .d(\u_cameraReader/pixel_counter [0]),
    .o(\u_cameraReader/mux14_b0_sel_is_2_o ));
  AL_MAP_LUT4 #(
    .EQN("(C*B*~(~D*~A))"),
    .INIT(16'hc080))
    _al_u497 (
    .a(_al_u477_o),
    .b(CSI_VSYNC_pad),
    .c(CSI_RST_pad),
    .d(\u_cameraReader/write_pixel ),
    .o(\u_cameraReader/mux12_b0_sel_is_2_o ));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u498 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(\uimg/inst_dob_i4_008 ),
    .c(\uimg/inst_dob_i6_008 ),
    .o(_al_u498_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u499 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(\uimg/inst_dob_i0_008 ),
    .c(\uimg/inst_dob_i2_008 ),
    .o(_al_u499_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'h00ac))
    _al_u500 (
    .a(_al_u498_o),
    .b(_al_u499_o),
    .c(lcd_rdaddr_piped_piped[2]),
    .d(lcd_rdaddr_piped_piped[3]),
    .o(_al_u500_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u501 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(lcd_rdaddr_piped_piped[2]),
    .c(\uimg/inst_dob_i12_008 ),
    .d(\uimg/inst_dob_i14_008 ),
    .o(_al_u501_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h3210))
    _al_u502 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(lcd_rdaddr_piped_piped[2]),
    .c(\uimg/inst_dob_i8_008 ),
    .d(\uimg/inst_dob_i10_008 ),
    .o(_al_u502_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(C*~B*~A))"),
    .INIT(16'h00ef))
    _al_u503 (
    .a(_al_u501_o),
    .b(_al_u502_o),
    .c(lcd_rdaddr_piped_piped[3]),
    .d(lcd_rdaddr_piped_piped[4]),
    .o(_al_u503_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u504 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(\uimg/inst_dob_i28_008 ),
    .c(\uimg/inst_dob_i30_008 ),
    .o(_al_u504_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u505 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(\uimg/inst_dob_i24_008 ),
    .c(\uimg/inst_dob_i26_008 ),
    .o(_al_u505_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'hac00))
    _al_u506 (
    .a(_al_u504_o),
    .b(_al_u505_o),
    .c(lcd_rdaddr_piped_piped[2]),
    .d(lcd_rdaddr_piped_piped[3]),
    .o(_al_u506_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u507 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(lcd_rdaddr_piped_piped[2]),
    .c(\uimg/inst_dob_i20_008 ),
    .d(\uimg/inst_dob_i22_008 ),
    .o(_al_u507_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h3210))
    _al_u508 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(lcd_rdaddr_piped_piped[2]),
    .c(\uimg/inst_dob_i16_008 ),
    .d(\uimg/inst_dob_i18_008 ),
    .o(_al_u508_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(~C*~B*~A))"),
    .INIT(16'hfe00))
    _al_u509 (
    .a(_al_u507_o),
    .b(_al_u508_o),
    .c(lcd_rdaddr_piped_piped[3]),
    .d(lcd_rdaddr_piped_piped[4]),
    .o(_al_u509_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~C)*~(B*~A))"),
    .INIT(16'hb0bb))
    _al_u510 (
    .a(_al_u500_o),
    .b(_al_u503_o),
    .c(_al_u506_o),
    .d(_al_u509_o),
    .o(_al_u510_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u511 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(\uimg/inst_dob_i36_008 ),
    .c(\uimg/inst_dob_i38_008 ),
    .o(_al_u511_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u512 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(\uimg/inst_dob_i32_008 ),
    .c(\uimg/inst_dob_i34_008 ),
    .o(_al_u512_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'h00ac))
    _al_u513 (
    .a(_al_u511_o),
    .b(_al_u512_o),
    .c(lcd_rdaddr_piped_piped[2]),
    .d(lcd_rdaddr_piped_piped[3]),
    .o(_al_u513_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u514 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(lcd_rdaddr_piped_piped[2]),
    .c(\uimg/inst_dob_i44_008 ),
    .d(\uimg/inst_dob_i46_008 ),
    .o(_al_u514_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h3210))
    _al_u515 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(lcd_rdaddr_piped_piped[2]),
    .c(\uimg/inst_dob_i40_008 ),
    .d(\uimg/inst_dob_i42_008 ),
    .o(_al_u515_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(C*~B*~A))"),
    .INIT(16'h00ef))
    _al_u516 (
    .a(_al_u514_o),
    .b(_al_u515_o),
    .c(lcd_rdaddr_piped_piped[3]),
    .d(lcd_rdaddr_piped_piped[4]),
    .o(_al_u516_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u517 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(\uimg/inst_dob_i52_008 ),
    .c(\uimg/inst_dob_i54_008 ),
    .o(_al_u517_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u518 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(\uimg/inst_dob_i48_008 ),
    .c(\uimg/inst_dob_i50_008 ),
    .o(_al_u518_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'h00ac))
    _al_u519 (
    .a(_al_u517_o),
    .b(_al_u518_o),
    .c(lcd_rdaddr_piped_piped[2]),
    .d(lcd_rdaddr_piped_piped[3]),
    .o(_al_u519_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h3210))
    _al_u520 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(lcd_rdaddr_piped_piped[2]),
    .c(\uimg/inst_dob_i56_008 ),
    .d(\uimg/inst_dob_i58_008 ),
    .o(_al_u520_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u521 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(lcd_rdaddr_piped_piped[2]),
    .c(\uimg/inst_dob_i60_008 ),
    .d(\uimg/inst_dob_i62_008 ),
    .o(_al_u521_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C*~B*~A))"),
    .INIT(16'hef00))
    _al_u522 (
    .a(_al_u520_o),
    .b(_al_u521_o),
    .c(lcd_rdaddr_piped_piped[3]),
    .d(lcd_rdaddr_piped_piped[4]),
    .o(_al_u522_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~C)*~(B*~A))"),
    .INIT(16'hb0bb))
    _al_u523 (
    .a(_al_u513_o),
    .b(_al_u516_o),
    .c(_al_u519_o),
    .d(_al_u522_o),
    .o(_al_u523_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h00ca))
    _al_u524 (
    .a(_al_u510_o),
    .b(_al_u523_o),
    .c(lcd_rdaddr_piped_piped[5]),
    .d(lcd_rdaddr_piped_piped[6]),
    .o(_al_u524_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*~(~D*B))"),
    .INIT(16'h5010))
    _al_u525 (
    .a(_al_u524_o),
    .b(lcd_rdaddr_piped_piped[6]),
    .c(lcd_rden),
    .d(\uimg/inst_dob_i64_008 ),
    .o(G_pad[5]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u526 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(\uimg/inst_dob_i8_007 ),
    .c(\uimg/inst_dob_i10_007 ),
    .o(_al_u526_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u527 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(\uimg/inst_dob_i12_007 ),
    .c(\uimg/inst_dob_i14_007 ),
    .o(_al_u527_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'hca00))
    _al_u528 (
    .a(_al_u526_o),
    .b(_al_u527_o),
    .c(lcd_rdaddr_piped_piped[2]),
    .d(lcd_rdaddr_piped_piped[3]),
    .o(_al_u528_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u529 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(lcd_rdaddr_piped_piped[2]),
    .c(\uimg/inst_dob_i4_007 ),
    .d(\uimg/inst_dob_i6_007 ),
    .o(_al_u529_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h3210))
    _al_u530 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(lcd_rdaddr_piped_piped[2]),
    .c(\uimg/inst_dob_i0_007 ),
    .d(\uimg/inst_dob_i2_007 ),
    .o(_al_u530_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(~C*~B*~A))"),
    .INIT(16'h00fe))
    _al_u531 (
    .a(_al_u529_o),
    .b(_al_u530_o),
    .c(lcd_rdaddr_piped_piped[3]),
    .d(lcd_rdaddr_piped_piped[4]),
    .o(_al_u531_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u532 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(\uimg/inst_dob_i20_007 ),
    .c(\uimg/inst_dob_i22_007 ),
    .o(_al_u532_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u533 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(\uimg/inst_dob_i16_007 ),
    .c(\uimg/inst_dob_i18_007 ),
    .o(_al_u533_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'h00ac))
    _al_u534 (
    .a(_al_u532_o),
    .b(_al_u533_o),
    .c(lcd_rdaddr_piped_piped[2]),
    .d(lcd_rdaddr_piped_piped[3]),
    .o(_al_u534_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h3210))
    _al_u535 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(lcd_rdaddr_piped_piped[2]),
    .c(\uimg/inst_dob_i24_007 ),
    .d(\uimg/inst_dob_i26_007 ),
    .o(_al_u535_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u536 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(lcd_rdaddr_piped_piped[2]),
    .c(\uimg/inst_dob_i28_007 ),
    .d(\uimg/inst_dob_i30_007 ),
    .o(_al_u536_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C*~B*~A))"),
    .INIT(16'hef00))
    _al_u537 (
    .a(_al_u535_o),
    .b(_al_u536_o),
    .c(lcd_rdaddr_piped_piped[3]),
    .d(lcd_rdaddr_piped_piped[4]),
    .o(_al_u537_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~C)*~(B*~A))"),
    .INIT(16'hb0bb))
    _al_u538 (
    .a(_al_u528_o),
    .b(_al_u531_o),
    .c(_al_u534_o),
    .d(_al_u537_o),
    .o(_al_u538_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u539 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(\uimg/inst_dob_i40_007 ),
    .c(\uimg/inst_dob_i42_007 ),
    .o(_al_u539_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u540 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(\uimg/inst_dob_i44_007 ),
    .c(\uimg/inst_dob_i46_007 ),
    .o(_al_u540_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'hca00))
    _al_u541 (
    .a(_al_u539_o),
    .b(_al_u540_o),
    .c(lcd_rdaddr_piped_piped[2]),
    .d(lcd_rdaddr_piped_piped[3]),
    .o(_al_u541_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u542 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(lcd_rdaddr_piped_piped[2]),
    .c(\uimg/inst_dob_i36_007 ),
    .d(\uimg/inst_dob_i38_007 ),
    .o(_al_u542_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h3210))
    _al_u543 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(lcd_rdaddr_piped_piped[2]),
    .c(\uimg/inst_dob_i32_007 ),
    .d(\uimg/inst_dob_i34_007 ),
    .o(_al_u543_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(~C*~B*~A))"),
    .INIT(16'h00fe))
    _al_u544 (
    .a(_al_u542_o),
    .b(_al_u543_o),
    .c(lcd_rdaddr_piped_piped[3]),
    .d(lcd_rdaddr_piped_piped[4]),
    .o(_al_u544_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u545 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(\uimg/inst_dob_i52_007 ),
    .c(\uimg/inst_dob_i54_007 ),
    .o(_al_u545_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u546 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(\uimg/inst_dob_i48_007 ),
    .c(\uimg/inst_dob_i50_007 ),
    .o(_al_u546_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'h00ac))
    _al_u547 (
    .a(_al_u545_o),
    .b(_al_u546_o),
    .c(lcd_rdaddr_piped_piped[2]),
    .d(lcd_rdaddr_piped_piped[3]),
    .o(_al_u547_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h3210))
    _al_u548 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(lcd_rdaddr_piped_piped[2]),
    .c(\uimg/inst_dob_i56_007 ),
    .d(\uimg/inst_dob_i58_007 ),
    .o(_al_u548_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u549 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(lcd_rdaddr_piped_piped[2]),
    .c(\uimg/inst_dob_i60_007 ),
    .d(\uimg/inst_dob_i62_007 ),
    .o(_al_u549_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C*~B*~A))"),
    .INIT(16'hef00))
    _al_u550 (
    .a(_al_u548_o),
    .b(_al_u549_o),
    .c(lcd_rdaddr_piped_piped[3]),
    .d(lcd_rdaddr_piped_piped[4]),
    .o(_al_u550_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~C)*~(B*~A))"),
    .INIT(16'hb0bb))
    _al_u551 (
    .a(_al_u541_o),
    .b(_al_u544_o),
    .c(_al_u547_o),
    .d(_al_u550_o),
    .o(_al_u551_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h00ca))
    _al_u552 (
    .a(_al_u538_o),
    .b(_al_u551_o),
    .c(lcd_rdaddr_piped_piped[5]),
    .d(lcd_rdaddr_piped_piped[6]),
    .o(_al_u552_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*~(~D*B))"),
    .INIT(16'h5010))
    _al_u553 (
    .a(_al_u552_o),
    .b(lcd_rdaddr_piped_piped[6]),
    .c(lcd_rden),
    .d(\uimg/inst_dob_i64_007 ),
    .o(G_pad[4]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u554 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(\uimg/inst_dob_i36_006 ),
    .c(\uimg/inst_dob_i38_006 ),
    .o(_al_u554_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u555 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(\uimg/inst_dob_i32_006 ),
    .c(\uimg/inst_dob_i34_006 ),
    .o(_al_u555_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'h00ac))
    _al_u556 (
    .a(_al_u554_o),
    .b(_al_u555_o),
    .c(lcd_rdaddr_piped_piped[2]),
    .d(lcd_rdaddr_piped_piped[3]),
    .o(_al_u556_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u557 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(lcd_rdaddr_piped_piped[2]),
    .c(\uimg/inst_dob_i44_006 ),
    .d(\uimg/inst_dob_i46_006 ),
    .o(_al_u557_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h3210))
    _al_u558 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(lcd_rdaddr_piped_piped[2]),
    .c(\uimg/inst_dob_i40_006 ),
    .d(\uimg/inst_dob_i42_006 ),
    .o(_al_u558_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(C*~B*~A))"),
    .INIT(16'h00ef))
    _al_u559 (
    .a(_al_u557_o),
    .b(_al_u558_o),
    .c(lcd_rdaddr_piped_piped[3]),
    .d(lcd_rdaddr_piped_piped[4]),
    .o(_al_u559_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u560 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(\uimg/inst_dob_i52_006 ),
    .c(\uimg/inst_dob_i54_006 ),
    .o(_al_u560_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u561 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(\uimg/inst_dob_i48_006 ),
    .c(\uimg/inst_dob_i50_006 ),
    .o(_al_u561_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'h00ac))
    _al_u562 (
    .a(_al_u560_o),
    .b(_al_u561_o),
    .c(lcd_rdaddr_piped_piped[2]),
    .d(lcd_rdaddr_piped_piped[3]),
    .o(_al_u562_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u563 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(lcd_rdaddr_piped_piped[2]),
    .c(\uimg/inst_dob_i60_006 ),
    .d(\uimg/inst_dob_i62_006 ),
    .o(_al_u563_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h3210))
    _al_u564 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(lcd_rdaddr_piped_piped[2]),
    .c(\uimg/inst_dob_i56_006 ),
    .d(\uimg/inst_dob_i58_006 ),
    .o(_al_u564_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C*~B*~A))"),
    .INIT(16'hef00))
    _al_u565 (
    .a(_al_u563_o),
    .b(_al_u564_o),
    .c(lcd_rdaddr_piped_piped[3]),
    .d(lcd_rdaddr_piped_piped[4]),
    .o(_al_u565_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~C)*~(B*~A))"),
    .INIT(16'hb0bb))
    _al_u566 (
    .a(_al_u556_o),
    .b(_al_u559_o),
    .c(_al_u562_o),
    .d(_al_u565_o),
    .o(_al_u566_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u567 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(\uimg/inst_dob_i4_006 ),
    .c(\uimg/inst_dob_i6_006 ),
    .o(_al_u567_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u568 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(\uimg/inst_dob_i0_006 ),
    .c(\uimg/inst_dob_i2_006 ),
    .o(_al_u568_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'h00ac))
    _al_u569 (
    .a(_al_u567_o),
    .b(_al_u568_o),
    .c(lcd_rdaddr_piped_piped[2]),
    .d(lcd_rdaddr_piped_piped[3]),
    .o(_al_u569_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u570 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(lcd_rdaddr_piped_piped[2]),
    .c(\uimg/inst_dob_i12_006 ),
    .d(\uimg/inst_dob_i14_006 ),
    .o(_al_u570_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h3210))
    _al_u571 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(lcd_rdaddr_piped_piped[2]),
    .c(\uimg/inst_dob_i8_006 ),
    .d(\uimg/inst_dob_i10_006 ),
    .o(_al_u571_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(C*~B*~A))"),
    .INIT(16'h00ef))
    _al_u572 (
    .a(_al_u570_o),
    .b(_al_u571_o),
    .c(lcd_rdaddr_piped_piped[3]),
    .d(lcd_rdaddr_piped_piped[4]),
    .o(_al_u572_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u573 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(\uimg/inst_dob_i28_006 ),
    .c(\uimg/inst_dob_i30_006 ),
    .o(_al_u573_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u574 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(\uimg/inst_dob_i24_006 ),
    .c(\uimg/inst_dob_i26_006 ),
    .o(_al_u574_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'hac00))
    _al_u575 (
    .a(_al_u573_o),
    .b(_al_u574_o),
    .c(lcd_rdaddr_piped_piped[2]),
    .d(lcd_rdaddr_piped_piped[3]),
    .o(_al_u575_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u576 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(lcd_rdaddr_piped_piped[2]),
    .c(\uimg/inst_dob_i20_006 ),
    .d(\uimg/inst_dob_i22_006 ),
    .o(_al_u576_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h3210))
    _al_u577 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(lcd_rdaddr_piped_piped[2]),
    .c(\uimg/inst_dob_i16_006 ),
    .d(\uimg/inst_dob_i18_006 ),
    .o(_al_u577_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(~C*~B*~A))"),
    .INIT(16'hfe00))
    _al_u578 (
    .a(_al_u576_o),
    .b(_al_u577_o),
    .c(lcd_rdaddr_piped_piped[3]),
    .d(lcd_rdaddr_piped_piped[4]),
    .o(_al_u578_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~C)*~(B*~A))"),
    .INIT(16'hb0bb))
    _al_u579 (
    .a(_al_u569_o),
    .b(_al_u572_o),
    .c(_al_u575_o),
    .d(_al_u578_o),
    .o(_al_u579_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'h00ac))
    _al_u580 (
    .a(_al_u566_o),
    .b(_al_u579_o),
    .c(lcd_rdaddr_piped_piped[5]),
    .d(lcd_rdaddr_piped_piped[6]),
    .o(_al_u580_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*~(~D*B))"),
    .INIT(16'h5010))
    _al_u581 (
    .a(_al_u580_o),
    .b(lcd_rdaddr_piped_piped[6]),
    .c(lcd_rden),
    .d(\uimg/inst_dob_i64_006 ),
    .o(G_pad[3]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u582 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(\uimg/inst_dob_i4_005 ),
    .c(\uimg/inst_dob_i6_005 ),
    .o(_al_u582_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u583 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(\uimg/inst_dob_i0_005 ),
    .c(\uimg/inst_dob_i2_005 ),
    .o(_al_u583_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'h00ac))
    _al_u584 (
    .a(_al_u582_o),
    .b(_al_u583_o),
    .c(lcd_rdaddr_piped_piped[2]),
    .d(lcd_rdaddr_piped_piped[3]),
    .o(_al_u584_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u585 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(lcd_rdaddr_piped_piped[2]),
    .c(\uimg/inst_dob_i12_005 ),
    .d(\uimg/inst_dob_i14_005 ),
    .o(_al_u585_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h3210))
    _al_u586 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(lcd_rdaddr_piped_piped[2]),
    .c(\uimg/inst_dob_i8_005 ),
    .d(\uimg/inst_dob_i10_005 ),
    .o(_al_u586_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(C*~B*~A))"),
    .INIT(16'h00ef))
    _al_u587 (
    .a(_al_u585_o),
    .b(_al_u586_o),
    .c(lcd_rdaddr_piped_piped[3]),
    .d(lcd_rdaddr_piped_piped[4]),
    .o(_al_u587_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u588 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(\uimg/inst_dob_i28_005 ),
    .c(\uimg/inst_dob_i30_005 ),
    .o(_al_u588_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u589 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(\uimg/inst_dob_i24_005 ),
    .c(\uimg/inst_dob_i26_005 ),
    .o(_al_u589_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'hac00))
    _al_u590 (
    .a(_al_u588_o),
    .b(_al_u589_o),
    .c(lcd_rdaddr_piped_piped[2]),
    .d(lcd_rdaddr_piped_piped[3]),
    .o(_al_u590_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u591 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(lcd_rdaddr_piped_piped[2]),
    .c(\uimg/inst_dob_i20_005 ),
    .d(\uimg/inst_dob_i22_005 ),
    .o(_al_u591_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h3210))
    _al_u592 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(lcd_rdaddr_piped_piped[2]),
    .c(\uimg/inst_dob_i16_005 ),
    .d(\uimg/inst_dob_i18_005 ),
    .o(_al_u592_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(~C*~B*~A))"),
    .INIT(16'hfe00))
    _al_u593 (
    .a(_al_u591_o),
    .b(_al_u592_o),
    .c(lcd_rdaddr_piped_piped[3]),
    .d(lcd_rdaddr_piped_piped[4]),
    .o(_al_u593_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~C)*~(B*~A))"),
    .INIT(16'hb0bb))
    _al_u594 (
    .a(_al_u584_o),
    .b(_al_u587_o),
    .c(_al_u590_o),
    .d(_al_u593_o),
    .o(_al_u594_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u595 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(\uimg/inst_dob_i36_005 ),
    .c(\uimg/inst_dob_i38_005 ),
    .o(_al_u595_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u596 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(\uimg/inst_dob_i32_005 ),
    .c(\uimg/inst_dob_i34_005 ),
    .o(_al_u596_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'h00ac))
    _al_u597 (
    .a(_al_u595_o),
    .b(_al_u596_o),
    .c(lcd_rdaddr_piped_piped[2]),
    .d(lcd_rdaddr_piped_piped[3]),
    .o(_al_u597_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u598 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(lcd_rdaddr_piped_piped[2]),
    .c(\uimg/inst_dob_i44_005 ),
    .d(\uimg/inst_dob_i46_005 ),
    .o(_al_u598_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h3210))
    _al_u599 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(lcd_rdaddr_piped_piped[2]),
    .c(\uimg/inst_dob_i40_005 ),
    .d(\uimg/inst_dob_i42_005 ),
    .o(_al_u599_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(C*~B*~A))"),
    .INIT(16'h00ef))
    _al_u600 (
    .a(_al_u598_o),
    .b(_al_u599_o),
    .c(lcd_rdaddr_piped_piped[3]),
    .d(lcd_rdaddr_piped_piped[4]),
    .o(_al_u600_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u601 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(\uimg/inst_dob_i60_005 ),
    .c(\uimg/inst_dob_i62_005 ),
    .o(_al_u601_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u602 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(\uimg/inst_dob_i56_005 ),
    .c(\uimg/inst_dob_i58_005 ),
    .o(_al_u602_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'hac00))
    _al_u603 (
    .a(_al_u601_o),
    .b(_al_u602_o),
    .c(lcd_rdaddr_piped_piped[2]),
    .d(lcd_rdaddr_piped_piped[3]),
    .o(_al_u603_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u604 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(lcd_rdaddr_piped_piped[2]),
    .c(\uimg/inst_dob_i52_005 ),
    .d(\uimg/inst_dob_i54_005 ),
    .o(_al_u604_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h3210))
    _al_u605 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(lcd_rdaddr_piped_piped[2]),
    .c(\uimg/inst_dob_i48_005 ),
    .d(\uimg/inst_dob_i50_005 ),
    .o(_al_u605_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(~C*~B*~A))"),
    .INIT(16'hfe00))
    _al_u606 (
    .a(_al_u604_o),
    .b(_al_u605_o),
    .c(lcd_rdaddr_piped_piped[3]),
    .d(lcd_rdaddr_piped_piped[4]),
    .o(_al_u606_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~C)*~(B*~A))"),
    .INIT(16'hb0bb))
    _al_u607 (
    .a(_al_u597_o),
    .b(_al_u600_o),
    .c(_al_u603_o),
    .d(_al_u606_o),
    .o(_al_u607_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h00ca))
    _al_u608 (
    .a(_al_u594_o),
    .b(_al_u607_o),
    .c(lcd_rdaddr_piped_piped[5]),
    .d(lcd_rdaddr_piped_piped[6]),
    .o(_al_u608_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*~(~D*B))"),
    .INIT(16'h5010))
    _al_u609 (
    .a(_al_u608_o),
    .b(lcd_rdaddr_piped_piped[6]),
    .c(lcd_rden),
    .d(\uimg/inst_dob_i64_005 ),
    .o(G_pad[2]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u610 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(\uimg/inst_dob_i4_004 ),
    .c(\uimg/inst_dob_i6_004 ),
    .o(_al_u610_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u611 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(\uimg/inst_dob_i0_004 ),
    .c(\uimg/inst_dob_i2_004 ),
    .o(_al_u611_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'h00ac))
    _al_u612 (
    .a(_al_u610_o),
    .b(_al_u611_o),
    .c(lcd_rdaddr_piped_piped[2]),
    .d(lcd_rdaddr_piped_piped[3]),
    .o(_al_u612_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u613 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(lcd_rdaddr_piped_piped[2]),
    .c(\uimg/inst_dob_i12_004 ),
    .d(\uimg/inst_dob_i14_004 ),
    .o(_al_u613_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h3210))
    _al_u614 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(lcd_rdaddr_piped_piped[2]),
    .c(\uimg/inst_dob_i8_004 ),
    .d(\uimg/inst_dob_i10_004 ),
    .o(_al_u614_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(C*~B*~A))"),
    .INIT(16'h00ef))
    _al_u615 (
    .a(_al_u613_o),
    .b(_al_u614_o),
    .c(lcd_rdaddr_piped_piped[3]),
    .d(lcd_rdaddr_piped_piped[4]),
    .o(_al_u615_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u616 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(\uimg/inst_dob_i28_004 ),
    .c(\uimg/inst_dob_i30_004 ),
    .o(_al_u616_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u617 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(\uimg/inst_dob_i24_004 ),
    .c(\uimg/inst_dob_i26_004 ),
    .o(_al_u617_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'hac00))
    _al_u618 (
    .a(_al_u616_o),
    .b(_al_u617_o),
    .c(lcd_rdaddr_piped_piped[2]),
    .d(lcd_rdaddr_piped_piped[3]),
    .o(_al_u618_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u619 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(lcd_rdaddr_piped_piped[2]),
    .c(\uimg/inst_dob_i20_004 ),
    .d(\uimg/inst_dob_i22_004 ),
    .o(_al_u619_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h3210))
    _al_u620 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(lcd_rdaddr_piped_piped[2]),
    .c(\uimg/inst_dob_i16_004 ),
    .d(\uimg/inst_dob_i18_004 ),
    .o(_al_u620_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(~C*~B*~A))"),
    .INIT(16'hfe00))
    _al_u621 (
    .a(_al_u619_o),
    .b(_al_u620_o),
    .c(lcd_rdaddr_piped_piped[3]),
    .d(lcd_rdaddr_piped_piped[4]),
    .o(_al_u621_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~C)*~(B*~A))"),
    .INIT(16'hb0bb))
    _al_u622 (
    .a(_al_u612_o),
    .b(_al_u615_o),
    .c(_al_u618_o),
    .d(_al_u621_o),
    .o(_al_u622_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u623 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(\uimg/inst_dob_i40_004 ),
    .c(\uimg/inst_dob_i42_004 ),
    .o(_al_u623_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u624 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(\uimg/inst_dob_i44_004 ),
    .c(\uimg/inst_dob_i46_004 ),
    .o(_al_u624_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'hca00))
    _al_u625 (
    .a(_al_u623_o),
    .b(_al_u624_o),
    .c(lcd_rdaddr_piped_piped[2]),
    .d(lcd_rdaddr_piped_piped[3]),
    .o(_al_u625_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u626 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(lcd_rdaddr_piped_piped[2]),
    .c(\uimg/inst_dob_i36_004 ),
    .d(\uimg/inst_dob_i38_004 ),
    .o(_al_u626_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h3210))
    _al_u627 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(lcd_rdaddr_piped_piped[2]),
    .c(\uimg/inst_dob_i32_004 ),
    .d(\uimg/inst_dob_i34_004 ),
    .o(_al_u627_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(~C*~B*~A))"),
    .INIT(16'h00fe))
    _al_u628 (
    .a(_al_u626_o),
    .b(_al_u627_o),
    .c(lcd_rdaddr_piped_piped[3]),
    .d(lcd_rdaddr_piped_piped[4]),
    .o(_al_u628_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u629 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(\uimg/inst_dob_i60_004 ),
    .c(\uimg/inst_dob_i62_004 ),
    .o(_al_u629_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u630 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(\uimg/inst_dob_i56_004 ),
    .c(\uimg/inst_dob_i58_004 ),
    .o(_al_u630_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'hac00))
    _al_u631 (
    .a(_al_u629_o),
    .b(_al_u630_o),
    .c(lcd_rdaddr_piped_piped[2]),
    .d(lcd_rdaddr_piped_piped[3]),
    .o(_al_u631_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u632 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(lcd_rdaddr_piped_piped[2]),
    .c(\uimg/inst_dob_i52_004 ),
    .d(\uimg/inst_dob_i54_004 ),
    .o(_al_u632_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h3210))
    _al_u633 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(lcd_rdaddr_piped_piped[2]),
    .c(\uimg/inst_dob_i48_004 ),
    .d(\uimg/inst_dob_i50_004 ),
    .o(_al_u633_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(~C*~B*~A))"),
    .INIT(16'hfe00))
    _al_u634 (
    .a(_al_u632_o),
    .b(_al_u633_o),
    .c(lcd_rdaddr_piped_piped[3]),
    .d(lcd_rdaddr_piped_piped[4]),
    .o(_al_u634_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~C)*~(B*~A))"),
    .INIT(16'hb0bb))
    _al_u635 (
    .a(_al_u625_o),
    .b(_al_u628_o),
    .c(_al_u631_o),
    .d(_al_u634_o),
    .o(_al_u635_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h00ca))
    _al_u636 (
    .a(_al_u622_o),
    .b(_al_u635_o),
    .c(lcd_rdaddr_piped_piped[5]),
    .d(lcd_rdaddr_piped_piped[6]),
    .o(_al_u636_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*~(~D*B))"),
    .INIT(16'h5010))
    _al_u637 (
    .a(_al_u636_o),
    .b(lcd_rdaddr_piped_piped[6]),
    .c(lcd_rden),
    .d(\uimg/inst_dob_i64_004 ),
    .o(B_pad[7]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u638 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(lcd_rdaddr_piped_piped[2]),
    .c(\uimg/inst_dob_i56_003 ),
    .d(\uimg/inst_dob_i58_003 ),
    .o(_al_u638_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h048c))
    _al_u639 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(lcd_rdaddr_piped_piped[2]),
    .c(\uimg/inst_dob_i60_003 ),
    .d(\uimg/inst_dob_i62_003 ),
    .o(_al_u639_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u640 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(lcd_rdaddr_piped_piped[2]),
    .c(\uimg/inst_dob_i48_003 ),
    .d(\uimg/inst_dob_i50_003 ),
    .o(_al_u640_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h048c))
    _al_u641 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(lcd_rdaddr_piped_piped[2]),
    .c(\uimg/inst_dob_i52_003 ),
    .d(\uimg/inst_dob_i54_003 ),
    .o(_al_u641_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u642 (
    .a(_al_u640_o),
    .b(_al_u641_o),
    .c(lcd_rdaddr_piped_piped[3]),
    .o(_al_u642_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(D*~C*~B))"),
    .INIT(16'h5455))
    _al_u643 (
    .a(_al_u642_o),
    .b(_al_u638_o),
    .c(_al_u639_o),
    .d(lcd_rdaddr_piped_piped[3]),
    .o(_al_u643_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u644 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(lcd_rdaddr_piped_piped[2]),
    .c(\uimg/inst_dob_i40_003 ),
    .d(\uimg/inst_dob_i42_003 ),
    .o(_al_u644_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h048c))
    _al_u645 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(lcd_rdaddr_piped_piped[2]),
    .c(\uimg/inst_dob_i44_003 ),
    .d(\uimg/inst_dob_i46_003 ),
    .o(_al_u645_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u646 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(lcd_rdaddr_piped_piped[2]),
    .c(\uimg/inst_dob_i32_003 ),
    .d(\uimg/inst_dob_i34_003 ),
    .o(_al_u646_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h048c))
    _al_u647 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(lcd_rdaddr_piped_piped[2]),
    .c(\uimg/inst_dob_i36_003 ),
    .d(\uimg/inst_dob_i38_003 ),
    .o(_al_u647_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u648 (
    .a(_al_u646_o),
    .b(_al_u647_o),
    .c(lcd_rdaddr_piped_piped[3]),
    .o(_al_u648_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(D*~C*~B))"),
    .INIT(16'h5455))
    _al_u649 (
    .a(_al_u648_o),
    .b(_al_u644_o),
    .c(_al_u645_o),
    .d(lcd_rdaddr_piped_piped[3]),
    .o(_al_u649_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'hac00))
    _al_u650 (
    .a(_al_u643_o),
    .b(_al_u649_o),
    .c(lcd_rdaddr_piped_piped[4]),
    .d(lcd_rdaddr_piped_piped[5]),
    .o(_al_u650_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u651 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(lcd_rdaddr_piped_piped[2]),
    .c(\uimg/inst_dob_i24_003 ),
    .d(\uimg/inst_dob_i26_003 ),
    .o(_al_u651_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h048c))
    _al_u652 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(lcd_rdaddr_piped_piped[2]),
    .c(\uimg/inst_dob_i28_003 ),
    .d(\uimg/inst_dob_i30_003 ),
    .o(_al_u652_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u653 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(lcd_rdaddr_piped_piped[2]),
    .c(\uimg/inst_dob_i16_003 ),
    .d(\uimg/inst_dob_i18_003 ),
    .o(_al_u653_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h048c))
    _al_u654 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(lcd_rdaddr_piped_piped[2]),
    .c(\uimg/inst_dob_i20_003 ),
    .d(\uimg/inst_dob_i22_003 ),
    .o(_al_u654_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u655 (
    .a(_al_u653_o),
    .b(_al_u654_o),
    .c(lcd_rdaddr_piped_piped[3]),
    .o(_al_u655_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(D*~C*~B))"),
    .INIT(16'h5455))
    _al_u656 (
    .a(_al_u655_o),
    .b(_al_u651_o),
    .c(_al_u652_o),
    .d(lcd_rdaddr_piped_piped[3]),
    .o(_al_u656_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u657 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(lcd_rdaddr_piped_piped[2]),
    .c(\uimg/inst_dob_i8_003 ),
    .d(\uimg/inst_dob_i10_003 ),
    .o(_al_u657_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h048c))
    _al_u658 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(lcd_rdaddr_piped_piped[2]),
    .c(\uimg/inst_dob_i12_003 ),
    .d(\uimg/inst_dob_i14_003 ),
    .o(_al_u658_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u659 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(lcd_rdaddr_piped_piped[2]),
    .c(\uimg/inst_dob_i0_003 ),
    .d(\uimg/inst_dob_i2_003 ),
    .o(_al_u659_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h048c))
    _al_u660 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(lcd_rdaddr_piped_piped[2]),
    .c(\uimg/inst_dob_i4_003 ),
    .d(\uimg/inst_dob_i6_003 ),
    .o(_al_u660_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u661 (
    .a(_al_u659_o),
    .b(_al_u660_o),
    .c(lcd_rdaddr_piped_piped[3]),
    .o(_al_u661_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(D*~C*~B))"),
    .INIT(16'h5455))
    _al_u662 (
    .a(_al_u661_o),
    .b(_al_u657_o),
    .c(_al_u658_o),
    .d(lcd_rdaddr_piped_piped[3]),
    .o(_al_u662_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'h00ac))
    _al_u663 (
    .a(_al_u656_o),
    .b(_al_u662_o),
    .c(lcd_rdaddr_piped_piped[4]),
    .d(lcd_rdaddr_piped_piped[5]),
    .o(_al_u663_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*A))"),
    .INIT(8'hc4))
    _al_u664 (
    .a(lcd_rdaddr_piped_piped[6]),
    .b(lcd_rden),
    .c(\uimg/inst_dob_i64_003 ),
    .o(_al_u664_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(~D*~(~B*~A)))"),
    .INIT(16'hf010))
    _al_u665 (
    .a(_al_u650_o),
    .b(_al_u663_o),
    .c(_al_u664_o),
    .d(lcd_rdaddr_piped_piped[6]),
    .o(B_pad[6]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u666 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(\uimg/inst_dob_i36_002 ),
    .c(\uimg/inst_dob_i38_002 ),
    .o(_al_u666_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u667 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(\uimg/inst_dob_i32_002 ),
    .c(\uimg/inst_dob_i34_002 ),
    .o(_al_u667_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'h00ac))
    _al_u668 (
    .a(_al_u666_o),
    .b(_al_u667_o),
    .c(lcd_rdaddr_piped_piped[2]),
    .d(lcd_rdaddr_piped_piped[3]),
    .o(_al_u668_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u669 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(lcd_rdaddr_piped_piped[2]),
    .c(\uimg/inst_dob_i44_002 ),
    .d(\uimg/inst_dob_i46_002 ),
    .o(_al_u669_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h3210))
    _al_u670 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(lcd_rdaddr_piped_piped[2]),
    .c(\uimg/inst_dob_i40_002 ),
    .d(\uimg/inst_dob_i42_002 ),
    .o(_al_u670_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(C*~B*~A))"),
    .INIT(16'h00ef))
    _al_u671 (
    .a(_al_u669_o),
    .b(_al_u670_o),
    .c(lcd_rdaddr_piped_piped[3]),
    .d(lcd_rdaddr_piped_piped[4]),
    .o(_al_u671_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u672 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(\uimg/inst_dob_i52_002 ),
    .c(\uimg/inst_dob_i54_002 ),
    .o(_al_u672_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u673 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(\uimg/inst_dob_i48_002 ),
    .c(\uimg/inst_dob_i50_002 ),
    .o(_al_u673_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'h00ac))
    _al_u674 (
    .a(_al_u672_o),
    .b(_al_u673_o),
    .c(lcd_rdaddr_piped_piped[2]),
    .d(lcd_rdaddr_piped_piped[3]),
    .o(_al_u674_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h3210))
    _al_u675 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(lcd_rdaddr_piped_piped[2]),
    .c(\uimg/inst_dob_i56_002 ),
    .d(\uimg/inst_dob_i58_002 ),
    .o(_al_u675_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u676 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(lcd_rdaddr_piped_piped[2]),
    .c(\uimg/inst_dob_i60_002 ),
    .d(\uimg/inst_dob_i62_002 ),
    .o(_al_u676_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C*~B*~A))"),
    .INIT(16'hef00))
    _al_u677 (
    .a(_al_u675_o),
    .b(_al_u676_o),
    .c(lcd_rdaddr_piped_piped[3]),
    .d(lcd_rdaddr_piped_piped[4]),
    .o(_al_u677_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~C)*~(B*~A))"),
    .INIT(16'hb0bb))
    _al_u678 (
    .a(_al_u668_o),
    .b(_al_u671_o),
    .c(_al_u674_o),
    .d(_al_u677_o),
    .o(_al_u678_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u679 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(\uimg/inst_dob_i8_002 ),
    .c(\uimg/inst_dob_i10_002 ),
    .o(_al_u679_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u680 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(\uimg/inst_dob_i12_002 ),
    .c(\uimg/inst_dob_i14_002 ),
    .o(_al_u680_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'hca00))
    _al_u681 (
    .a(_al_u679_o),
    .b(_al_u680_o),
    .c(lcd_rdaddr_piped_piped[2]),
    .d(lcd_rdaddr_piped_piped[3]),
    .o(_al_u681_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u682 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(lcd_rdaddr_piped_piped[2]),
    .c(\uimg/inst_dob_i4_002 ),
    .d(\uimg/inst_dob_i6_002 ),
    .o(_al_u682_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h3210))
    _al_u683 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(lcd_rdaddr_piped_piped[2]),
    .c(\uimg/inst_dob_i0_002 ),
    .d(\uimg/inst_dob_i2_002 ),
    .o(_al_u683_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(~C*~B*~A))"),
    .INIT(16'h00fe))
    _al_u684 (
    .a(_al_u682_o),
    .b(_al_u683_o),
    .c(lcd_rdaddr_piped_piped[3]),
    .d(lcd_rdaddr_piped_piped[4]),
    .o(_al_u684_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u685 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(\uimg/inst_dob_i20_002 ),
    .c(\uimg/inst_dob_i22_002 ),
    .o(_al_u685_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u686 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(\uimg/inst_dob_i16_002 ),
    .c(\uimg/inst_dob_i18_002 ),
    .o(_al_u686_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'h00ac))
    _al_u687 (
    .a(_al_u685_o),
    .b(_al_u686_o),
    .c(lcd_rdaddr_piped_piped[2]),
    .d(lcd_rdaddr_piped_piped[3]),
    .o(_al_u687_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h3210))
    _al_u688 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(lcd_rdaddr_piped_piped[2]),
    .c(\uimg/inst_dob_i24_002 ),
    .d(\uimg/inst_dob_i26_002 ),
    .o(_al_u688_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u689 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(lcd_rdaddr_piped_piped[2]),
    .c(\uimg/inst_dob_i28_002 ),
    .d(\uimg/inst_dob_i30_002 ),
    .o(_al_u689_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C*~B*~A))"),
    .INIT(16'hef00))
    _al_u690 (
    .a(_al_u688_o),
    .b(_al_u689_o),
    .c(lcd_rdaddr_piped_piped[3]),
    .d(lcd_rdaddr_piped_piped[4]),
    .o(_al_u690_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~C)*~(B*~A))"),
    .INIT(16'hb0bb))
    _al_u691 (
    .a(_al_u681_o),
    .b(_al_u684_o),
    .c(_al_u687_o),
    .d(_al_u690_o),
    .o(_al_u691_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'h00ac))
    _al_u692 (
    .a(_al_u678_o),
    .b(_al_u691_o),
    .c(lcd_rdaddr_piped_piped[5]),
    .d(lcd_rdaddr_piped_piped[6]),
    .o(_al_u692_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*~(~D*B))"),
    .INIT(16'h5010))
    _al_u693 (
    .a(_al_u692_o),
    .b(lcd_rdaddr_piped_piped[6]),
    .c(lcd_rden),
    .d(\uimg/inst_dob_i64_002 ),
    .o(B_pad[5]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u694 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(lcd_rdaddr_piped_piped[2]),
    .c(\uimg/inst_dob_i56_001 ),
    .d(\uimg/inst_dob_i58_001 ),
    .o(_al_u694_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h048c))
    _al_u695 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(lcd_rdaddr_piped_piped[2]),
    .c(\uimg/inst_dob_i60_001 ),
    .d(\uimg/inst_dob_i62_001 ),
    .o(_al_u695_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u696 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(lcd_rdaddr_piped_piped[2]),
    .c(\uimg/inst_dob_i48_001 ),
    .d(\uimg/inst_dob_i50_001 ),
    .o(_al_u696_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h048c))
    _al_u697 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(lcd_rdaddr_piped_piped[2]),
    .c(\uimg/inst_dob_i52_001 ),
    .d(\uimg/inst_dob_i54_001 ),
    .o(_al_u697_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u698 (
    .a(_al_u696_o),
    .b(_al_u697_o),
    .c(lcd_rdaddr_piped_piped[3]),
    .o(_al_u698_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(D*~C*~B))"),
    .INIT(16'h5455))
    _al_u699 (
    .a(_al_u698_o),
    .b(_al_u694_o),
    .c(_al_u695_o),
    .d(lcd_rdaddr_piped_piped[3]),
    .o(_al_u699_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u700 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(lcd_rdaddr_piped_piped[2]),
    .c(\uimg/inst_dob_i40_001 ),
    .d(\uimg/inst_dob_i42_001 ),
    .o(_al_u700_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h048c))
    _al_u701 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(lcd_rdaddr_piped_piped[2]),
    .c(\uimg/inst_dob_i44_001 ),
    .d(\uimg/inst_dob_i46_001 ),
    .o(_al_u701_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u702 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(lcd_rdaddr_piped_piped[2]),
    .c(\uimg/inst_dob_i32_001 ),
    .d(\uimg/inst_dob_i34_001 ),
    .o(_al_u702_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h048c))
    _al_u703 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(lcd_rdaddr_piped_piped[2]),
    .c(\uimg/inst_dob_i36_001 ),
    .d(\uimg/inst_dob_i38_001 ),
    .o(_al_u703_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u704 (
    .a(_al_u702_o),
    .b(_al_u703_o),
    .c(lcd_rdaddr_piped_piped[3]),
    .o(_al_u704_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(D*~C*~B))"),
    .INIT(16'h5455))
    _al_u705 (
    .a(_al_u704_o),
    .b(_al_u700_o),
    .c(_al_u701_o),
    .d(lcd_rdaddr_piped_piped[3]),
    .o(_al_u705_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'hac00))
    _al_u706 (
    .a(_al_u699_o),
    .b(_al_u705_o),
    .c(lcd_rdaddr_piped_piped[4]),
    .d(lcd_rdaddr_piped_piped[5]),
    .o(_al_u706_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u707 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(lcd_rdaddr_piped_piped[2]),
    .c(\uimg/inst_dob_i24_001 ),
    .d(\uimg/inst_dob_i26_001 ),
    .o(_al_u707_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h048c))
    _al_u708 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(lcd_rdaddr_piped_piped[2]),
    .c(\uimg/inst_dob_i28_001 ),
    .d(\uimg/inst_dob_i30_001 ),
    .o(_al_u708_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u709 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(lcd_rdaddr_piped_piped[2]),
    .c(\uimg/inst_dob_i16_001 ),
    .d(\uimg/inst_dob_i18_001 ),
    .o(_al_u709_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h048c))
    _al_u710 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(lcd_rdaddr_piped_piped[2]),
    .c(\uimg/inst_dob_i20_001 ),
    .d(\uimg/inst_dob_i22_001 ),
    .o(_al_u710_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u711 (
    .a(_al_u709_o),
    .b(_al_u710_o),
    .c(lcd_rdaddr_piped_piped[3]),
    .o(_al_u711_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(D*~C*~B))"),
    .INIT(16'h5455))
    _al_u712 (
    .a(_al_u711_o),
    .b(_al_u707_o),
    .c(_al_u708_o),
    .d(lcd_rdaddr_piped_piped[3]),
    .o(_al_u712_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u713 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(lcd_rdaddr_piped_piped[2]),
    .c(\uimg/inst_dob_i8_001 ),
    .d(\uimg/inst_dob_i10_001 ),
    .o(_al_u713_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h048c))
    _al_u714 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(lcd_rdaddr_piped_piped[2]),
    .c(\uimg/inst_dob_i12_001 ),
    .d(\uimg/inst_dob_i14_001 ),
    .o(_al_u714_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u715 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(lcd_rdaddr_piped_piped[2]),
    .c(\uimg/inst_dob_i0_001 ),
    .d(\uimg/inst_dob_i2_001 ),
    .o(_al_u715_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h048c))
    _al_u716 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(lcd_rdaddr_piped_piped[2]),
    .c(\uimg/inst_dob_i4_001 ),
    .d(\uimg/inst_dob_i6_001 ),
    .o(_al_u716_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u717 (
    .a(_al_u715_o),
    .b(_al_u716_o),
    .c(lcd_rdaddr_piped_piped[3]),
    .o(_al_u717_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(D*~C*~B))"),
    .INIT(16'h5455))
    _al_u718 (
    .a(_al_u717_o),
    .b(_al_u713_o),
    .c(_al_u714_o),
    .d(lcd_rdaddr_piped_piped[3]),
    .o(_al_u718_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'h00ac))
    _al_u719 (
    .a(_al_u712_o),
    .b(_al_u718_o),
    .c(lcd_rdaddr_piped_piped[4]),
    .d(lcd_rdaddr_piped_piped[5]),
    .o(_al_u719_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*A))"),
    .INIT(8'hc4))
    _al_u720 (
    .a(lcd_rdaddr_piped_piped[6]),
    .b(lcd_rden),
    .c(\uimg/inst_dob_i64_001 ),
    .o(_al_u720_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(~D*~(~B*~A)))"),
    .INIT(16'hf010))
    _al_u721 (
    .a(_al_u706_o),
    .b(_al_u719_o),
    .c(_al_u720_o),
    .d(lcd_rdaddr_piped_piped[6]),
    .o(B_pad[4]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u722 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(\uimg/inst_dob_i36_000 ),
    .c(\uimg/inst_dob_i38_000 ),
    .o(_al_u722_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u723 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(\uimg/inst_dob_i32_000 ),
    .c(\uimg/inst_dob_i34_000 ),
    .o(_al_u723_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'h00ac))
    _al_u724 (
    .a(_al_u722_o),
    .b(_al_u723_o),
    .c(lcd_rdaddr_piped_piped[2]),
    .d(lcd_rdaddr_piped_piped[3]),
    .o(_al_u724_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u725 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(lcd_rdaddr_piped_piped[2]),
    .c(\uimg/inst_dob_i44_000 ),
    .d(\uimg/inst_dob_i46_000 ),
    .o(_al_u725_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h3210))
    _al_u726 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(lcd_rdaddr_piped_piped[2]),
    .c(\uimg/inst_dob_i40_000 ),
    .d(\uimg/inst_dob_i42_000 ),
    .o(_al_u726_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(C*~B*~A))"),
    .INIT(16'h00ef))
    _al_u727 (
    .a(_al_u725_o),
    .b(_al_u726_o),
    .c(lcd_rdaddr_piped_piped[3]),
    .d(lcd_rdaddr_piped_piped[4]),
    .o(_al_u727_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u728 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(\uimg/inst_dob_i52_000 ),
    .c(\uimg/inst_dob_i54_000 ),
    .o(_al_u728_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u729 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(\uimg/inst_dob_i48_000 ),
    .c(\uimg/inst_dob_i50_000 ),
    .o(_al_u729_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'h00ac))
    _al_u730 (
    .a(_al_u728_o),
    .b(_al_u729_o),
    .c(lcd_rdaddr_piped_piped[2]),
    .d(lcd_rdaddr_piped_piped[3]),
    .o(_al_u730_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h3210))
    _al_u731 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(lcd_rdaddr_piped_piped[2]),
    .c(\uimg/inst_dob_i56_000 ),
    .d(\uimg/inst_dob_i58_000 ),
    .o(_al_u731_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u732 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(lcd_rdaddr_piped_piped[2]),
    .c(\uimg/inst_dob_i60_000 ),
    .d(\uimg/inst_dob_i62_000 ),
    .o(_al_u732_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C*~B*~A))"),
    .INIT(16'hef00))
    _al_u733 (
    .a(_al_u731_o),
    .b(_al_u732_o),
    .c(lcd_rdaddr_piped_piped[3]),
    .d(lcd_rdaddr_piped_piped[4]),
    .o(_al_u733_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~C)*~(B*~A))"),
    .INIT(16'hb0bb))
    _al_u734 (
    .a(_al_u724_o),
    .b(_al_u727_o),
    .c(_al_u730_o),
    .d(_al_u733_o),
    .o(_al_u734_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u735 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(\uimg/inst_dob_i4_000 ),
    .c(\uimg/inst_dob_i6_000 ),
    .o(_al_u735_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u736 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(\uimg/inst_dob_i0_000 ),
    .c(\uimg/inst_dob_i2_000 ),
    .o(_al_u736_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'h00ac))
    _al_u737 (
    .a(_al_u735_o),
    .b(_al_u736_o),
    .c(lcd_rdaddr_piped_piped[2]),
    .d(lcd_rdaddr_piped_piped[3]),
    .o(_al_u737_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u738 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(lcd_rdaddr_piped_piped[2]),
    .c(\uimg/inst_dob_i12_000 ),
    .d(\uimg/inst_dob_i14_000 ),
    .o(_al_u738_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h3210))
    _al_u739 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(lcd_rdaddr_piped_piped[2]),
    .c(\uimg/inst_dob_i8_000 ),
    .d(\uimg/inst_dob_i10_000 ),
    .o(_al_u739_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(C*~B*~A))"),
    .INIT(16'h00ef))
    _al_u740 (
    .a(_al_u738_o),
    .b(_al_u739_o),
    .c(lcd_rdaddr_piped_piped[3]),
    .d(lcd_rdaddr_piped_piped[4]),
    .o(_al_u740_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u741 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(\uimg/inst_dob_i28_000 ),
    .c(\uimg/inst_dob_i30_000 ),
    .o(_al_u741_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u742 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(\uimg/inst_dob_i24_000 ),
    .c(\uimg/inst_dob_i26_000 ),
    .o(_al_u742_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'hac00))
    _al_u743 (
    .a(_al_u741_o),
    .b(_al_u742_o),
    .c(lcd_rdaddr_piped_piped[2]),
    .d(lcd_rdaddr_piped_piped[3]),
    .o(_al_u743_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u744 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(lcd_rdaddr_piped_piped[2]),
    .c(\uimg/inst_dob_i20_000 ),
    .d(\uimg/inst_dob_i22_000 ),
    .o(_al_u744_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h3210))
    _al_u745 (
    .a(lcd_rdaddr_piped_piped[1]),
    .b(lcd_rdaddr_piped_piped[2]),
    .c(\uimg/inst_dob_i16_000 ),
    .d(\uimg/inst_dob_i18_000 ),
    .o(_al_u745_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(~C*~B*~A))"),
    .INIT(16'hfe00))
    _al_u746 (
    .a(_al_u744_o),
    .b(_al_u745_o),
    .c(lcd_rdaddr_piped_piped[3]),
    .d(lcd_rdaddr_piped_piped[4]),
    .o(_al_u746_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~C)*~(B*~A))"),
    .INIT(16'hb0bb))
    _al_u747 (
    .a(_al_u737_o),
    .b(_al_u740_o),
    .c(_al_u743_o),
    .d(_al_u746_o),
    .o(_al_u747_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'h00ac))
    _al_u748 (
    .a(_al_u734_o),
    .b(_al_u747_o),
    .c(lcd_rdaddr_piped_piped[5]),
    .d(lcd_rdaddr_piped_piped[6]),
    .o(_al_u748_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*~(~D*B))"),
    .INIT(16'h5010))
    _al_u749 (
    .a(_al_u748_o),
    .b(lcd_rdaddr_piped_piped[6]),
    .c(lcd_rden),
    .d(\uimg/inst_dob_i64_000 ),
    .o(B_pad[3]));
  AL_MAP_LUT4 #(
    .EQN("(~B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h3210))
    _al_u750 (
    .a(lcd_rdaddr_piped_piped[4]),
    .b(lcd_rdaddr_piped_piped[5]),
    .c(\uimg/inst_dob_i0_015 ),
    .d(\uimg/inst_dob_i16_015 ),
    .o(_al_u750_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u751 (
    .a(lcd_rdaddr_piped_piped[4]),
    .b(lcd_rdaddr_piped_piped[5]),
    .c(\uimg/inst_dob_i32_015 ),
    .d(\uimg/inst_dob_i48_015 ),
    .o(_al_u751_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*A))"),
    .INIT(8'hc4))
    _al_u752 (
    .a(lcd_rdaddr_piped_piped[6]),
    .b(lcd_rden),
    .c(\uimg/inst_dob_i64_015 ),
    .o(_al_u752_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(~D*~B*~A))"),
    .INIT(16'hf0e0))
    _al_u753 (
    .a(_al_u750_o),
    .b(_al_u751_o),
    .c(_al_u752_o),
    .d(lcd_rdaddr_piped_piped[6]),
    .o(R_pad[7]));
  AL_MAP_LUT4 #(
    .EQN("(~B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h3210))
    _al_u754 (
    .a(lcd_rdaddr_piped_piped[4]),
    .b(lcd_rdaddr_piped_piped[5]),
    .c(\uimg/inst_dob_i0_014 ),
    .d(\uimg/inst_dob_i16_014 ),
    .o(_al_u754_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u755 (
    .a(lcd_rdaddr_piped_piped[4]),
    .b(lcd_rdaddr_piped_piped[5]),
    .c(\uimg/inst_dob_i32_014 ),
    .d(\uimg/inst_dob_i48_014 ),
    .o(_al_u755_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*A))"),
    .INIT(8'hc4))
    _al_u756 (
    .a(lcd_rdaddr_piped_piped[6]),
    .b(lcd_rden),
    .c(\uimg/inst_dob_i64_014 ),
    .o(_al_u756_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(~D*~B*~A))"),
    .INIT(16'hf0e0))
    _al_u757 (
    .a(_al_u754_o),
    .b(_al_u755_o),
    .c(_al_u756_o),
    .d(lcd_rdaddr_piped_piped[6]),
    .o(R_pad[6]));
  AL_MAP_LUT4 #(
    .EQN("(~B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h3210))
    _al_u758 (
    .a(lcd_rdaddr_piped_piped[4]),
    .b(lcd_rdaddr_piped_piped[5]),
    .c(\uimg/inst_dob_i0_013 ),
    .d(\uimg/inst_dob_i16_013 ),
    .o(_al_u758_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u759 (
    .a(lcd_rdaddr_piped_piped[4]),
    .b(lcd_rdaddr_piped_piped[5]),
    .c(\uimg/inst_dob_i32_013 ),
    .d(\uimg/inst_dob_i48_013 ),
    .o(_al_u759_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*A))"),
    .INIT(8'hc4))
    _al_u760 (
    .a(lcd_rdaddr_piped_piped[6]),
    .b(lcd_rden),
    .c(\uimg/inst_dob_i64_013 ),
    .o(_al_u760_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(~D*~B*~A))"),
    .INIT(16'hf0e0))
    _al_u761 (
    .a(_al_u758_o),
    .b(_al_u759_o),
    .c(_al_u760_o),
    .d(lcd_rdaddr_piped_piped[6]),
    .o(R_pad[5]));
  AL_MAP_LUT4 #(
    .EQN("(~B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h3210))
    _al_u762 (
    .a(lcd_rdaddr_piped_piped[4]),
    .b(lcd_rdaddr_piped_piped[5]),
    .c(\uimg/inst_dob_i0_012 ),
    .d(\uimg/inst_dob_i16_012 ),
    .o(_al_u762_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u763 (
    .a(lcd_rdaddr_piped_piped[4]),
    .b(lcd_rdaddr_piped_piped[5]),
    .c(\uimg/inst_dob_i32_012 ),
    .d(\uimg/inst_dob_i48_012 ),
    .o(_al_u763_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*A))"),
    .INIT(8'hc4))
    _al_u764 (
    .a(lcd_rdaddr_piped_piped[6]),
    .b(lcd_rden),
    .c(\uimg/inst_dob_i64_012 ),
    .o(_al_u764_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(~D*~B*~A))"),
    .INIT(16'hf0e0))
    _al_u765 (
    .a(_al_u762_o),
    .b(_al_u763_o),
    .c(_al_u764_o),
    .d(lcd_rdaddr_piped_piped[6]),
    .o(R_pad[4]));
  AL_MAP_LUT4 #(
    .EQN("(~B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h3210))
    _al_u766 (
    .a(lcd_rdaddr_piped_piped[4]),
    .b(lcd_rdaddr_piped_piped[5]),
    .c(\uimg/inst_dob_i0_011 ),
    .d(\uimg/inst_dob_i16_011 ),
    .o(_al_u766_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u767 (
    .a(lcd_rdaddr_piped_piped[4]),
    .b(lcd_rdaddr_piped_piped[5]),
    .c(\uimg/inst_dob_i32_011 ),
    .d(\uimg/inst_dob_i48_011 ),
    .o(_al_u767_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*A))"),
    .INIT(8'hc4))
    _al_u768 (
    .a(lcd_rdaddr_piped_piped[6]),
    .b(lcd_rden),
    .c(\uimg/inst_dob_i64_011 ),
    .o(_al_u768_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(~D*~B*~A))"),
    .INIT(16'hf0e0))
    _al_u769 (
    .a(_al_u766_o),
    .b(_al_u767_o),
    .c(_al_u768_o),
    .d(lcd_rdaddr_piped_piped[6]),
    .o(R_pad[3]));
  AL_MAP_LUT4 #(
    .EQN("(~B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h3210))
    _al_u770 (
    .a(lcd_rdaddr_piped_piped[4]),
    .b(lcd_rdaddr_piped_piped[5]),
    .c(\uimg/inst_dob_i0_010 ),
    .d(\uimg/inst_dob_i16_010 ),
    .o(_al_u770_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u771 (
    .a(lcd_rdaddr_piped_piped[4]),
    .b(lcd_rdaddr_piped_piped[5]),
    .c(\uimg/inst_dob_i32_010 ),
    .d(\uimg/inst_dob_i48_010 ),
    .o(_al_u771_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*A))"),
    .INIT(8'hc4))
    _al_u772 (
    .a(lcd_rdaddr_piped_piped[6]),
    .b(lcd_rden),
    .c(\uimg/inst_dob_i64_010 ),
    .o(_al_u772_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(~D*~B*~A))"),
    .INIT(16'hf0e0))
    _al_u773 (
    .a(_al_u770_o),
    .b(_al_u771_o),
    .c(_al_u772_o),
    .d(lcd_rdaddr_piped_piped[6]),
    .o(G_pad[7]));
  AL_MAP_LUT4 #(
    .EQN("(~B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h3210))
    _al_u774 (
    .a(lcd_rdaddr_piped_piped[4]),
    .b(lcd_rdaddr_piped_piped[5]),
    .c(\uimg/inst_dob_i0_009 ),
    .d(\uimg/inst_dob_i16_009 ),
    .o(_al_u774_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u775 (
    .a(lcd_rdaddr_piped_piped[4]),
    .b(lcd_rdaddr_piped_piped[5]),
    .c(\uimg/inst_dob_i32_009 ),
    .d(\uimg/inst_dob_i48_009 ),
    .o(_al_u775_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*A))"),
    .INIT(8'hc4))
    _al_u776 (
    .a(lcd_rdaddr_piped_piped[6]),
    .b(lcd_rden),
    .c(\uimg/inst_dob_i64_009 ),
    .o(_al_u776_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(~D*~B*~A))"),
    .INIT(16'hf0e0))
    _al_u777 (
    .a(_al_u774_o),
    .b(_al_u775_o),
    .c(_al_u776_o),
    .d(lcd_rdaddr_piped_piped[6]),
    .o(G_pad[6]));
  AL_MAP_LUT1 #(
    .EQN("(~A)"),
    .INIT(2'h1))
    _al_u778 (
    .a(CSI_RST_pad),
    .o(CSI_RST_pad_neg));
  AL_MAP_LUT1 #(
    .EQN("(~A)"),
    .INIT(2'h1))
    _al_u779 (
    .a(\u_cameraReader/wrclk1 ),
    .o(\u_cameraReader/n1 ));
  EG_PHY_CONFIG #(
    .DONE_PERSISTN("ENABLE"),
    .INIT_PERSISTN("ENABLE"),
    .JTAG_PERSISTN("DISABLE"),
    .PROGRAMN_PERSISTN("DISABLE"))
    config_inst ();
  reg_sr_as_w1 lcd_rdaddr_pipe_b0 (
    .clk(clk_lcd),
    .d(lcd_rdaddr[9]),
    .en(lcd_rden),
    .reset(CSI_RST_pad_neg),
    .set(1'b0),
    .q(lcd_rdaddr_piped[0]));
  reg_sr_as_w1 lcd_rdaddr_pipe_b1 (
    .clk(clk_lcd),
    .d(lcd_rdaddr[10]),
    .en(lcd_rden),
    .reset(CSI_RST_pad_neg),
    .set(1'b0),
    .q(lcd_rdaddr_piped[1]));
  reg_sr_as_w1 lcd_rdaddr_pipe_b2 (
    .clk(clk_lcd),
    .d(lcd_rdaddr[11]),
    .en(lcd_rden),
    .reset(CSI_RST_pad_neg),
    .set(1'b0),
    .q(lcd_rdaddr_piped[2]));
  reg_sr_as_w1 lcd_rdaddr_pipe_b3 (
    .clk(clk_lcd),
    .d(lcd_rdaddr[12]),
    .en(lcd_rden),
    .reset(CSI_RST_pad_neg),
    .set(1'b0),
    .q(lcd_rdaddr_piped[3]));
  reg_sr_as_w1 lcd_rdaddr_pipe_b4 (
    .clk(clk_lcd),
    .d(lcd_rdaddr[13]),
    .en(lcd_rden),
    .reset(CSI_RST_pad_neg),
    .set(1'b0),
    .q(lcd_rdaddr_piped[4]));
  reg_sr_as_w1 lcd_rdaddr_pipe_b5 (
    .clk(clk_lcd),
    .d(lcd_rdaddr[14]),
    .en(lcd_rden),
    .reset(CSI_RST_pad_neg),
    .set(1'b0),
    .q(lcd_rdaddr_piped[5]));
  reg_sr_as_w1 lcd_rdaddr_pipe_b6 (
    .clk(clk_lcd),
    .d(lcd_rdaddr[15]),
    .en(lcd_rden),
    .reset(CSI_RST_pad_neg),
    .set(1'b0),
    .q(lcd_rdaddr_piped[6]));
  reg_sr_as_w1 lcd_rdaddr_piped_pipe_b0 (
    .clk(clk_lcd),
    .d(lcd_rdaddr_piped[0]),
    .en(lcd_rden),
    .reset(CSI_RST_pad_neg),
    .set(1'b0));
  reg_sr_as_w1 lcd_rdaddr_piped_pipe_b1 (
    .clk(clk_lcd),
    .d(lcd_rdaddr_piped[1]),
    .en(lcd_rden),
    .reset(CSI_RST_pad_neg),
    .set(1'b0),
    .q(lcd_rdaddr_piped_piped[1]));
  reg_sr_as_w1 lcd_rdaddr_piped_pipe_b2 (
    .clk(clk_lcd),
    .d(lcd_rdaddr_piped[2]),
    .en(lcd_rden),
    .reset(CSI_RST_pad_neg),
    .set(1'b0),
    .q(lcd_rdaddr_piped_piped[2]));
  reg_sr_as_w1 lcd_rdaddr_piped_pipe_b3 (
    .clk(clk_lcd),
    .d(lcd_rdaddr_piped[3]),
    .en(lcd_rden),
    .reset(CSI_RST_pad_neg),
    .set(1'b0),
    .q(lcd_rdaddr_piped_piped[3]));
  reg_sr_as_w1 lcd_rdaddr_piped_pipe_b4 (
    .clk(clk_lcd),
    .d(lcd_rdaddr_piped[4]),
    .en(lcd_rden),
    .reset(CSI_RST_pad_neg),
    .set(1'b0),
    .q(lcd_rdaddr_piped_piped[4]));
  reg_sr_as_w1 lcd_rdaddr_piped_pipe_b5 (
    .clk(clk_lcd),
    .d(lcd_rdaddr_piped[5]),
    .en(lcd_rden),
    .reset(CSI_RST_pad_neg),
    .set(1'b0),
    .q(lcd_rdaddr_piped_piped[5]));
  reg_sr_as_w1 lcd_rdaddr_piped_pipe_b6 (
    .clk(clk_lcd),
    .d(lcd_rdaddr_piped[6]),
    .en(lcd_rden),
    .reset(CSI_RST_pad_neg),
    .set(1'b0),
    .q(lcd_rdaddr_piped_piped[6]));
  EG_PHY_GCLK \pll/bufg_feedback  (
    .clki(\pll/clk0_buf ),
    .clko(clk_lcd));  // al_ip/ip_pll.v(36)
  EG_PHY_PLL #(
    .CLKC0_CPHASE(19),
    .CLKC0_DIV(20),
    .CLKC0_DIV2_ENABLE("DISABLE"),
    .CLKC0_ENABLE("ENABLE"),
    .CLKC0_FPHASE(0),
    .CLKC1_CPHASE(41),
    .CLKC1_DIV(42),
    .CLKC1_DIV2_ENABLE("DISABLE"),
    .CLKC1_ENABLE("ENABLE"),
    .CLKC1_FPHASE(0),
    .CLKC2_CPHASE(125),
    .CLKC2_DIV(126),
    .CLKC2_DIV2_ENABLE("DISABLE"),
    .CLKC2_ENABLE("ENABLE"),
    .CLKC2_FPHASE(0),
    .CLKC3_CPHASE(1),
    .CLKC3_DIV(1),
    .CLKC3_DIV2_ENABLE("DISABLE"),
    .CLKC3_ENABLE("DISABLE"),
    .CLKC3_FPHASE(0),
    .CLKC4_CPHASE(1),
    .CLKC4_DIV(1),
    .CLKC4_DIV2_ENABLE("DISABLE"),
    .CLKC4_ENABLE("DISABLE"),
    .CLKC4_FPHASE(0),
    .DERIVE_PLL_CLOCKS("DISABLE"),
    .DPHASE_SOURCE("DISABLE"),
    .DYNCFG("DISABLE"),
    .FBCLK_DIV(17),
    .FEEDBK_MODE("NORMAL"),
    .FEEDBK_PATH("CLKC0_EXT"),
    .FIN("24.000"),
    .FREQ_LOCK_ACCURACY(2),
    .GEN_BASIC_CLOCK("DISABLE"),
    .GMC_GAIN(6),
    .GMC_TEST(14),
    .ICP_CURRENT(3),
    .IF_ESCLKSTSW("DISABLE"),
    .INTFB_WAKE("DISABLE"),
    .KVCO(6),
    .LPF_CAPACITOR(3),
    .LPF_RESISTOR(2),
    .NORESET("DISABLE"),
    .ODIV_MUXC0("DIV"),
    .ODIV_MUXC1("DIV"),
    .ODIV_MUXC2("DIV"),
    .ODIV_MUXC3("DIV"),
    .ODIV_MUXC4("DIV"),
    .PLLC2RST_ENA("DISABLE"),
    .PLLC34RST_ENA("DISABLE"),
    .PLLMRST_ENA("DISABLE"),
    .PLLRST_ENA("DISABLE"),
    .PLL_LOCK_MODE(0),
    .PREDIV_MUXC0("VCO"),
    .PREDIV_MUXC1("VCO"),
    .PREDIV_MUXC2("VCO"),
    .PREDIV_MUXC3("VCO"),
    .PREDIV_MUXC4("VCO"),
    .REFCLK_DIV(16),
    .REFCLK_SEL("INTERNAL"),
    .STDBY_ENABLE("DISABLE"),
    .STDBY_VCO_ENA("DISABLE"),
    .SYNC_ENABLE("DISABLE"),
    .VCO_NORESET("DISABLE"))
    \pll/pll_inst  (
    .daddr(6'b000000),
    .dclk(1'b0),
    .dcs(1'b0),
    .di(8'b00000000),
    .dwe(1'b0),
    .fbclk(clk_lcd),
    .psclk(1'b0),
    .psclksel(3'b000),
    .psdown(1'b0),
    .psstep(1'b0),
    .refclk(CLK_IN_pad),
    .reset(1'b0),
    .stdby(1'b0),
    .clkc({open_n981,open_n982,clk_sccb,clk_cam,\pll/clk0_buf }));  // al_ip/ip_pll.v(67)
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cameraReader/add0/u0  (
    .a(\u_cameraReader/pixel_counter [0]),
    .b(1'b1),
    .c(\u_cameraReader/add0/c0 ),
    .o({\u_cameraReader/add0/c1 ,\u_cameraReader/n8 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cameraReader/add0/u1  (
    .a(\u_cameraReader/pixel_counter [1]),
    .b(1'b0),
    .c(\u_cameraReader/add0/c1 ),
    .o({\u_cameraReader/add0/c2 ,\u_cameraReader/n8 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cameraReader/add0/u10  (
    .a(\u_cameraReader/pixel_counter [10]),
    .b(1'b0),
    .c(\u_cameraReader/add0/c10 ),
    .o({\u_cameraReader/add0/c11 ,\u_cameraReader/n8 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cameraReader/add0/u11  (
    .a(\u_cameraReader/pixel_counter [11]),
    .b(1'b0),
    .c(\u_cameraReader/add0/c11 ),
    .o({\u_cameraReader/add0/c12 ,\u_cameraReader/n8 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cameraReader/add0/u12  (
    .a(\u_cameraReader/pixel_counter [12]),
    .b(1'b0),
    .c(\u_cameraReader/add0/c12 ),
    .o({\u_cameraReader/add0/c13 ,\u_cameraReader/n8 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cameraReader/add0/u13  (
    .a(\u_cameraReader/pixel_counter [13]),
    .b(1'b0),
    .c(\u_cameraReader/add0/c13 ),
    .o({\u_cameraReader/add0/c14 ,\u_cameraReader/n8 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cameraReader/add0/u14  (
    .a(\u_cameraReader/pixel_counter [14]),
    .b(1'b0),
    .c(\u_cameraReader/add0/c14 ),
    .o({\u_cameraReader/add0/c15 ,\u_cameraReader/n8 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cameraReader/add0/u15  (
    .a(\u_cameraReader/pixel_counter [15]),
    .b(1'b0),
    .c(\u_cameraReader/add0/c15 ),
    .o({\u_cameraReader/add0/c16 ,\u_cameraReader/n8 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cameraReader/add0/u16  (
    .a(\u_cameraReader/pixel_counter [16]),
    .b(1'b0),
    .c(\u_cameraReader/add0/c16 ),
    .o({\u_cameraReader/add0/c17 ,\u_cameraReader/n8 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cameraReader/add0/u17  (
    .a(\u_cameraReader/pixel_counter [17]),
    .b(1'b0),
    .c(\u_cameraReader/add0/c17 ),
    .o({\u_cameraReader/add0/c18 ,\u_cameraReader/n8 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cameraReader/add0/u18  (
    .a(\u_cameraReader/pixel_counter [18]),
    .b(1'b0),
    .c(\u_cameraReader/add0/c18 ),
    .o({\u_cameraReader/add0/c19 ,\u_cameraReader/n8 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cameraReader/add0/u19  (
    .a(\u_cameraReader/pixel_counter [19]),
    .b(1'b0),
    .c(\u_cameraReader/add0/c19 ),
    .o({open_n993,\u_cameraReader/n8 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cameraReader/add0/u2  (
    .a(\u_cameraReader/pixel_counter [2]),
    .b(1'b0),
    .c(\u_cameraReader/add0/c2 ),
    .o({\u_cameraReader/add0/c3 ,\u_cameraReader/n8 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cameraReader/add0/u3  (
    .a(\u_cameraReader/pixel_counter [3]),
    .b(1'b0),
    .c(\u_cameraReader/add0/c3 ),
    .o({\u_cameraReader/add0/c4 ,\u_cameraReader/n8 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cameraReader/add0/u4  (
    .a(\u_cameraReader/pixel_counter [4]),
    .b(1'b0),
    .c(\u_cameraReader/add0/c4 ),
    .o({\u_cameraReader/add0/c5 ,\u_cameraReader/n8 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cameraReader/add0/u5  (
    .a(\u_cameraReader/pixel_counter [5]),
    .b(1'b0),
    .c(\u_cameraReader/add0/c5 ),
    .o({\u_cameraReader/add0/c6 ,\u_cameraReader/n8 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cameraReader/add0/u6  (
    .a(\u_cameraReader/pixel_counter [6]),
    .b(1'b0),
    .c(\u_cameraReader/add0/c6 ),
    .o({\u_cameraReader/add0/c7 ,\u_cameraReader/n8 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cameraReader/add0/u7  (
    .a(\u_cameraReader/pixel_counter [7]),
    .b(1'b0),
    .c(\u_cameraReader/add0/c7 ),
    .o({\u_cameraReader/add0/c8 ,\u_cameraReader/n8 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cameraReader/add0/u8  (
    .a(\u_cameraReader/pixel_counter [8]),
    .b(1'b0),
    .c(\u_cameraReader/add0/c8 ),
    .o({\u_cameraReader/add0/c9 ,\u_cameraReader/n8 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cameraReader/add0/u9  (
    .a(\u_cameraReader/pixel_counter [9]),
    .b(1'b0),
    .c(\u_cameraReader/add0/c9 ),
    .o({\u_cameraReader/add0/c10 ,\u_cameraReader/n8 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u_cameraReader/add0/ucin  (
    .a(1'b0),
    .o({\u_cameraReader/add0/c0 ,open_n996}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cameraReader/add1/u0  (
    .a(camera_addr[0]),
    .b(1'b1),
    .c(\u_cameraReader/add1/c0 ),
    .o({\u_cameraReader/add1/c1 ,\u_cameraReader/n9 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cameraReader/add1/u1  (
    .a(camera_addr[1]),
    .b(1'b0),
    .c(\u_cameraReader/add1/c1 ),
    .o({\u_cameraReader/add1/c2 ,\u_cameraReader/n9 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cameraReader/add1/u10  (
    .a(camera_addr[10]),
    .b(1'b0),
    .c(\u_cameraReader/add1/c10 ),
    .o({\u_cameraReader/add1/c11 ,\u_cameraReader/n9 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cameraReader/add1/u11  (
    .a(camera_addr[11]),
    .b(1'b0),
    .c(\u_cameraReader/add1/c11 ),
    .o({\u_cameraReader/add1/c12 ,\u_cameraReader/n9 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cameraReader/add1/u12  (
    .a(camera_addr[12]),
    .b(1'b0),
    .c(\u_cameraReader/add1/c12 ),
    .o({\u_cameraReader/add1/c13 ,\u_cameraReader/n9 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cameraReader/add1/u13  (
    .a(camera_addr[13]),
    .b(1'b0),
    .c(\u_cameraReader/add1/c13 ),
    .o({\u_cameraReader/add1/c14 ,\u_cameraReader/n9 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cameraReader/add1/u14  (
    .a(camera_addr[14]),
    .b(1'b0),
    .c(\u_cameraReader/add1/c14 ),
    .o({\u_cameraReader/add1/c15 ,\u_cameraReader/n9 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cameraReader/add1/u15  (
    .a(camera_addr[15]),
    .b(1'b0),
    .c(\u_cameraReader/add1/c15 ),
    .o({open_n997,\u_cameraReader/n9 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cameraReader/add1/u2  (
    .a(camera_addr[2]),
    .b(1'b0),
    .c(\u_cameraReader/add1/c2 ),
    .o({\u_cameraReader/add1/c3 ,\u_cameraReader/n9 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cameraReader/add1/u3  (
    .a(camera_addr[3]),
    .b(1'b0),
    .c(\u_cameraReader/add1/c3 ),
    .o({\u_cameraReader/add1/c4 ,\u_cameraReader/n9 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cameraReader/add1/u4  (
    .a(camera_addr[4]),
    .b(1'b0),
    .c(\u_cameraReader/add1/c4 ),
    .o({\u_cameraReader/add1/c5 ,\u_cameraReader/n9 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cameraReader/add1/u5  (
    .a(camera_addr[5]),
    .b(1'b0),
    .c(\u_cameraReader/add1/c5 ),
    .o({\u_cameraReader/add1/c6 ,\u_cameraReader/n9 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cameraReader/add1/u6  (
    .a(camera_addr[6]),
    .b(1'b0),
    .c(\u_cameraReader/add1/c6 ),
    .o({\u_cameraReader/add1/c7 ,\u_cameraReader/n9 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cameraReader/add1/u7  (
    .a(camera_addr[7]),
    .b(1'b0),
    .c(\u_cameraReader/add1/c7 ),
    .o({\u_cameraReader/add1/c8 ,\u_cameraReader/n9 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cameraReader/add1/u8  (
    .a(camera_addr[8]),
    .b(1'b0),
    .c(\u_cameraReader/add1/c8 ),
    .o({\u_cameraReader/add1/c9 ,\u_cameraReader/n9 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_cameraReader/add1/u9  (
    .a(camera_addr[9]),
    .b(1'b0),
    .c(\u_cameraReader/add1/c9 ),
    .o({\u_cameraReader/add1/c10 ,\u_cameraReader/n9 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u_cameraReader/add1/ucin  (
    .a(1'b0),
    .o({\u_cameraReader/add1/c0 ,open_n1000}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_cameraReader/lt0_0  (
    .a(1'b0),
    .b(\u_cameraReader/pixel_counter [0]),
    .c(\u_cameraReader/lt0_c0 ),
    .o({\u_cameraReader/lt0_c1 ,open_n1001}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_cameraReader/lt0_1  (
    .a(1'b1),
    .b(\u_cameraReader/pixel_counter [1]),
    .c(\u_cameraReader/lt0_c1 ),
    .o({\u_cameraReader/lt0_c2 ,open_n1002}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_cameraReader/lt0_10  (
    .a(1'b0),
    .b(\u_cameraReader/pixel_counter [10]),
    .c(\u_cameraReader/lt0_c10 ),
    .o({\u_cameraReader/lt0_c11 ,open_n1003}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_cameraReader/lt0_11  (
    .a(1'b0),
    .b(\u_cameraReader/pixel_counter [11]),
    .c(\u_cameraReader/lt0_c11 ),
    .o({\u_cameraReader/lt0_c12 ,open_n1004}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_cameraReader/lt0_12  (
    .a(1'b0),
    .b(\u_cameraReader/pixel_counter [12]),
    .c(\u_cameraReader/lt0_c12 ),
    .o({\u_cameraReader/lt0_c13 ,open_n1005}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_cameraReader/lt0_13  (
    .a(1'b0),
    .b(\u_cameraReader/pixel_counter [13]),
    .c(\u_cameraReader/lt0_c13 ),
    .o({\u_cameraReader/lt0_c14 ,open_n1006}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_cameraReader/lt0_14  (
    .a(1'b0),
    .b(\u_cameraReader/pixel_counter [14]),
    .c(\u_cameraReader/lt0_c14 ),
    .o({\u_cameraReader/lt0_c15 ,open_n1007}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_cameraReader/lt0_15  (
    .a(1'b0),
    .b(\u_cameraReader/pixel_counter [15]),
    .c(\u_cameraReader/lt0_c15 ),
    .o({\u_cameraReader/lt0_c16 ,open_n1008}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_cameraReader/lt0_16  (
    .a(1'b0),
    .b(\u_cameraReader/pixel_counter [16]),
    .c(\u_cameraReader/lt0_c16 ),
    .o({\u_cameraReader/lt0_c17 ,open_n1009}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_cameraReader/lt0_17  (
    .a(1'b0),
    .b(\u_cameraReader/pixel_counter [17]),
    .c(\u_cameraReader/lt0_c17 ),
    .o({\u_cameraReader/lt0_c18 ,open_n1010}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_cameraReader/lt0_18  (
    .a(1'b0),
    .b(\u_cameraReader/pixel_counter [18]),
    .c(\u_cameraReader/lt0_c18 ),
    .o({\u_cameraReader/lt0_c19 ,open_n1011}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_cameraReader/lt0_19  (
    .a(1'b0),
    .b(\u_cameraReader/pixel_counter [19]),
    .c(\u_cameraReader/lt0_c19 ),
    .o({\u_cameraReader/lt0_c20 ,open_n1012}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_cameraReader/lt0_2  (
    .a(1'b0),
    .b(\u_cameraReader/pixel_counter [2]),
    .c(\u_cameraReader/lt0_c2 ),
    .o({\u_cameraReader/lt0_c3 ,open_n1013}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_cameraReader/lt0_3  (
    .a(1'b0),
    .b(\u_cameraReader/pixel_counter [3]),
    .c(\u_cameraReader/lt0_c3 ),
    .o({\u_cameraReader/lt0_c4 ,open_n1014}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_cameraReader/lt0_4  (
    .a(1'b0),
    .b(\u_cameraReader/pixel_counter [4]),
    .c(\u_cameraReader/lt0_c4 ),
    .o({\u_cameraReader/lt0_c5 ,open_n1015}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_cameraReader/lt0_5  (
    .a(1'b0),
    .b(\u_cameraReader/pixel_counter [5]),
    .c(\u_cameraReader/lt0_c5 ),
    .o({\u_cameraReader/lt0_c6 ,open_n1016}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_cameraReader/lt0_6  (
    .a(1'b0),
    .b(\u_cameraReader/pixel_counter [6]),
    .c(\u_cameraReader/lt0_c6 ),
    .o({\u_cameraReader/lt0_c7 ,open_n1017}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_cameraReader/lt0_7  (
    .a(1'b0),
    .b(\u_cameraReader/pixel_counter [7]),
    .c(\u_cameraReader/lt0_c7 ),
    .o({\u_cameraReader/lt0_c8 ,open_n1018}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_cameraReader/lt0_8  (
    .a(1'b0),
    .b(\u_cameraReader/pixel_counter [8]),
    .c(\u_cameraReader/lt0_c8 ),
    .o({\u_cameraReader/lt0_c9 ,open_n1019}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_cameraReader/lt0_9  (
    .a(1'b0),
    .b(\u_cameraReader/pixel_counter [9]),
    .c(\u_cameraReader/lt0_c9 ),
    .o({\u_cameraReader/lt0_c10 ,open_n1020}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u_cameraReader/lt0_cin  (
    .a(1'b0),
    .o({\u_cameraReader/lt0_c0 ,open_n1023}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_cameraReader/lt0_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u_cameraReader/lt0_c20 ),
    .o({open_n1024,\u_cameraReader/n29 }));
  reg_ar_as_w1 \u_cameraReader/reg0_b0  (
    .clk(camera_wrreq),
    .d(\u_cameraReader/current_pixel [0]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(camera_wrdat[0]));  // sources/rtl/cameraReader.v(55)
  reg_ar_as_w1 \u_cameraReader/reg0_b1  (
    .clk(camera_wrreq),
    .d(\u_cameraReader/current_pixel [1]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(camera_wrdat[1]));  // sources/rtl/cameraReader.v(55)
  reg_ar_as_w1 \u_cameraReader/reg0_b10  (
    .clk(camera_wrreq),
    .d(\u_cameraReader/current_pixel [10]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(camera_wrdat[10]));  // sources/rtl/cameraReader.v(55)
  reg_ar_as_w1 \u_cameraReader/reg0_b11  (
    .clk(camera_wrreq),
    .d(\u_cameraReader/current_pixel [11]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(camera_wrdat[11]));  // sources/rtl/cameraReader.v(55)
  reg_ar_as_w1 \u_cameraReader/reg0_b12  (
    .clk(camera_wrreq),
    .d(\u_cameraReader/current_pixel [12]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(camera_wrdat[12]));  // sources/rtl/cameraReader.v(55)
  reg_ar_as_w1 \u_cameraReader/reg0_b13  (
    .clk(camera_wrreq),
    .d(\u_cameraReader/current_pixel [13]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(camera_wrdat[13]));  // sources/rtl/cameraReader.v(55)
  reg_ar_as_w1 \u_cameraReader/reg0_b14  (
    .clk(camera_wrreq),
    .d(\u_cameraReader/current_pixel [14]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(camera_wrdat[14]));  // sources/rtl/cameraReader.v(55)
  reg_ar_as_w1 \u_cameraReader/reg0_b15  (
    .clk(camera_wrreq),
    .d(\u_cameraReader/current_pixel [15]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(camera_wrdat[15]));  // sources/rtl/cameraReader.v(55)
  reg_ar_as_w1 \u_cameraReader/reg0_b2  (
    .clk(camera_wrreq),
    .d(\u_cameraReader/current_pixel [2]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(camera_wrdat[2]));  // sources/rtl/cameraReader.v(55)
  reg_ar_as_w1 \u_cameraReader/reg0_b3  (
    .clk(camera_wrreq),
    .d(\u_cameraReader/current_pixel [3]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(camera_wrdat[3]));  // sources/rtl/cameraReader.v(55)
  reg_ar_as_w1 \u_cameraReader/reg0_b4  (
    .clk(camera_wrreq),
    .d(\u_cameraReader/current_pixel [4]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(camera_wrdat[4]));  // sources/rtl/cameraReader.v(55)
  reg_ar_as_w1 \u_cameraReader/reg0_b5  (
    .clk(camera_wrreq),
    .d(\u_cameraReader/current_pixel [5]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(camera_wrdat[5]));  // sources/rtl/cameraReader.v(55)
  reg_ar_as_w1 \u_cameraReader/reg0_b6  (
    .clk(camera_wrreq),
    .d(\u_cameraReader/current_pixel [6]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(camera_wrdat[6]));  // sources/rtl/cameraReader.v(55)
  reg_ar_as_w1 \u_cameraReader/reg0_b7  (
    .clk(camera_wrreq),
    .d(\u_cameraReader/current_pixel [7]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(camera_wrdat[7]));  // sources/rtl/cameraReader.v(55)
  reg_ar_as_w1 \u_cameraReader/reg0_b8  (
    .clk(camera_wrreq),
    .d(\u_cameraReader/current_pixel [8]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(camera_wrdat[8]));  // sources/rtl/cameraReader.v(55)
  reg_ar_as_w1 \u_cameraReader/reg0_b9  (
    .clk(camera_wrreq),
    .d(\u_cameraReader/current_pixel [9]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(camera_wrdat[9]));  // sources/rtl/cameraReader.v(55)
  reg_sr_as_w1 \u_cameraReader/reg1_b0  (
    .clk(CSI_PCLK_pad),
    .d(\u_cameraReader/n8 [0]),
    .en(1'b1),
    .reset(~\u_cameraReader/mux12_b0_sel_is_2_o ),
    .set(1'b0),
    .q(\u_cameraReader/pixel_counter [0]));  // sources/rtl/cameraReader.v(95)
  reg_sr_as_w1 \u_cameraReader/reg1_b1  (
    .clk(CSI_PCLK_pad),
    .d(\u_cameraReader/n8 [1]),
    .en(1'b1),
    .reset(~\u_cameraReader/mux12_b0_sel_is_2_o ),
    .set(1'b0),
    .q(\u_cameraReader/pixel_counter [1]));  // sources/rtl/cameraReader.v(95)
  reg_sr_as_w1 \u_cameraReader/reg1_b10  (
    .clk(CSI_PCLK_pad),
    .d(\u_cameraReader/n8 [10]),
    .en(1'b1),
    .reset(~\u_cameraReader/mux12_b0_sel_is_2_o ),
    .set(1'b0),
    .q(\u_cameraReader/pixel_counter [10]));  // sources/rtl/cameraReader.v(95)
  reg_sr_as_w1 \u_cameraReader/reg1_b11  (
    .clk(CSI_PCLK_pad),
    .d(\u_cameraReader/n8 [11]),
    .en(1'b1),
    .reset(~\u_cameraReader/mux12_b0_sel_is_2_o ),
    .set(1'b0),
    .q(\u_cameraReader/pixel_counter [11]));  // sources/rtl/cameraReader.v(95)
  reg_sr_as_w1 \u_cameraReader/reg1_b12  (
    .clk(CSI_PCLK_pad),
    .d(\u_cameraReader/n8 [12]),
    .en(1'b1),
    .reset(~\u_cameraReader/mux12_b0_sel_is_2_o ),
    .set(1'b0),
    .q(\u_cameraReader/pixel_counter [12]));  // sources/rtl/cameraReader.v(95)
  reg_sr_as_w1 \u_cameraReader/reg1_b13  (
    .clk(CSI_PCLK_pad),
    .d(\u_cameraReader/n8 [13]),
    .en(1'b1),
    .reset(~\u_cameraReader/mux12_b0_sel_is_2_o ),
    .set(1'b0),
    .q(\u_cameraReader/pixel_counter [13]));  // sources/rtl/cameraReader.v(95)
  reg_sr_as_w1 \u_cameraReader/reg1_b14  (
    .clk(CSI_PCLK_pad),
    .d(\u_cameraReader/n8 [14]),
    .en(1'b1),
    .reset(~\u_cameraReader/mux12_b0_sel_is_2_o ),
    .set(1'b0),
    .q(\u_cameraReader/pixel_counter [14]));  // sources/rtl/cameraReader.v(95)
  reg_sr_as_w1 \u_cameraReader/reg1_b15  (
    .clk(CSI_PCLK_pad),
    .d(\u_cameraReader/n8 [15]),
    .en(1'b1),
    .reset(~\u_cameraReader/mux12_b0_sel_is_2_o ),
    .set(1'b0),
    .q(\u_cameraReader/pixel_counter [15]));  // sources/rtl/cameraReader.v(95)
  reg_sr_as_w1 \u_cameraReader/reg1_b16  (
    .clk(CSI_PCLK_pad),
    .d(\u_cameraReader/n8 [16]),
    .en(1'b1),
    .reset(~\u_cameraReader/mux12_b0_sel_is_2_o ),
    .set(1'b0),
    .q(\u_cameraReader/pixel_counter [16]));  // sources/rtl/cameraReader.v(95)
  reg_sr_as_w1 \u_cameraReader/reg1_b17  (
    .clk(CSI_PCLK_pad),
    .d(\u_cameraReader/n8 [17]),
    .en(1'b1),
    .reset(~\u_cameraReader/mux12_b0_sel_is_2_o ),
    .set(1'b0),
    .q(\u_cameraReader/pixel_counter [17]));  // sources/rtl/cameraReader.v(95)
  reg_sr_as_w1 \u_cameraReader/reg1_b18  (
    .clk(CSI_PCLK_pad),
    .d(\u_cameraReader/n8 [18]),
    .en(1'b1),
    .reset(~\u_cameraReader/mux12_b0_sel_is_2_o ),
    .set(1'b0),
    .q(\u_cameraReader/pixel_counter [18]));  // sources/rtl/cameraReader.v(95)
  reg_sr_as_w1 \u_cameraReader/reg1_b19  (
    .clk(CSI_PCLK_pad),
    .d(\u_cameraReader/n8 [19]),
    .en(1'b1),
    .reset(~\u_cameraReader/mux12_b0_sel_is_2_o ),
    .set(1'b0),
    .q(\u_cameraReader/pixel_counter [19]));  // sources/rtl/cameraReader.v(95)
  reg_sr_as_w1 \u_cameraReader/reg1_b2  (
    .clk(CSI_PCLK_pad),
    .d(\u_cameraReader/n8 [2]),
    .en(1'b1),
    .reset(~\u_cameraReader/mux12_b0_sel_is_2_o ),
    .set(1'b0),
    .q(\u_cameraReader/pixel_counter [2]));  // sources/rtl/cameraReader.v(95)
  reg_sr_as_w1 \u_cameraReader/reg1_b3  (
    .clk(CSI_PCLK_pad),
    .d(\u_cameraReader/n8 [3]),
    .en(1'b1),
    .reset(~\u_cameraReader/mux12_b0_sel_is_2_o ),
    .set(1'b0),
    .q(\u_cameraReader/pixel_counter [3]));  // sources/rtl/cameraReader.v(95)
  reg_sr_as_w1 \u_cameraReader/reg1_b4  (
    .clk(CSI_PCLK_pad),
    .d(\u_cameraReader/n8 [4]),
    .en(1'b1),
    .reset(~\u_cameraReader/mux12_b0_sel_is_2_o ),
    .set(1'b0),
    .q(\u_cameraReader/pixel_counter [4]));  // sources/rtl/cameraReader.v(95)
  reg_sr_as_w1 \u_cameraReader/reg1_b5  (
    .clk(CSI_PCLK_pad),
    .d(\u_cameraReader/n8 [5]),
    .en(1'b1),
    .reset(~\u_cameraReader/mux12_b0_sel_is_2_o ),
    .set(1'b0),
    .q(\u_cameraReader/pixel_counter [5]));  // sources/rtl/cameraReader.v(95)
  reg_sr_as_w1 \u_cameraReader/reg1_b6  (
    .clk(CSI_PCLK_pad),
    .d(\u_cameraReader/n8 [6]),
    .en(1'b1),
    .reset(~\u_cameraReader/mux12_b0_sel_is_2_o ),
    .set(1'b0),
    .q(\u_cameraReader/pixel_counter [6]));  // sources/rtl/cameraReader.v(95)
  reg_sr_as_w1 \u_cameraReader/reg1_b7  (
    .clk(CSI_PCLK_pad),
    .d(\u_cameraReader/n8 [7]),
    .en(1'b1),
    .reset(~\u_cameraReader/mux12_b0_sel_is_2_o ),
    .set(1'b0),
    .q(\u_cameraReader/pixel_counter [7]));  // sources/rtl/cameraReader.v(95)
  reg_sr_as_w1 \u_cameraReader/reg1_b8  (
    .clk(CSI_PCLK_pad),
    .d(\u_cameraReader/n8 [8]),
    .en(1'b1),
    .reset(~\u_cameraReader/mux12_b0_sel_is_2_o ),
    .set(1'b0),
    .q(\u_cameraReader/pixel_counter [8]));  // sources/rtl/cameraReader.v(95)
  reg_sr_as_w1 \u_cameraReader/reg1_b9  (
    .clk(CSI_PCLK_pad),
    .d(\u_cameraReader/n8 [9]),
    .en(1'b1),
    .reset(~\u_cameraReader/mux12_b0_sel_is_2_o ),
    .set(1'b0),
    .q(\u_cameraReader/pixel_counter [9]));  // sources/rtl/cameraReader.v(95)
  reg_ar_as_w1 \u_cameraReader/reg2_b0  (
    .clk(CSI_PCLK_pad),
    .d(\u_cameraReader/n21 [0]),
    .en(~CSI_RST_pad_neg),
    .reset(1'b0),
    .set(1'b0),
    .q(camera_addr[0]));  // sources/rtl/cameraReader.v(95)
  reg_ar_as_w1 \u_cameraReader/reg2_b1  (
    .clk(CSI_PCLK_pad),
    .d(\u_cameraReader/n21 [1]),
    .en(~CSI_RST_pad_neg),
    .reset(1'b0),
    .set(1'b0),
    .q(camera_addr[1]));  // sources/rtl/cameraReader.v(95)
  reg_ar_as_w1 \u_cameraReader/reg2_b10  (
    .clk(CSI_PCLK_pad),
    .d(\u_cameraReader/n21 [10]),
    .en(~CSI_RST_pad_neg),
    .reset(1'b0),
    .set(1'b0),
    .q(camera_addr[10]));  // sources/rtl/cameraReader.v(95)
  reg_ar_as_w1 \u_cameraReader/reg2_b11  (
    .clk(CSI_PCLK_pad),
    .d(\u_cameraReader/n21 [11]),
    .en(~CSI_RST_pad_neg),
    .reset(1'b0),
    .set(1'b0),
    .q(camera_addr[11]));  // sources/rtl/cameraReader.v(95)
  reg_ar_as_w1 \u_cameraReader/reg2_b12  (
    .clk(CSI_PCLK_pad),
    .d(\u_cameraReader/n21 [12]),
    .en(~CSI_RST_pad_neg),
    .reset(1'b0),
    .set(1'b0),
    .q(camera_addr[12]));  // sources/rtl/cameraReader.v(95)
  reg_ar_as_w1 \u_cameraReader/reg2_b13  (
    .clk(CSI_PCLK_pad),
    .d(\u_cameraReader/n21 [13]),
    .en(~CSI_RST_pad_neg),
    .reset(1'b0),
    .set(1'b0),
    .q(camera_addr[13]));  // sources/rtl/cameraReader.v(95)
  reg_ar_as_w1 \u_cameraReader/reg2_b14  (
    .clk(CSI_PCLK_pad),
    .d(\u_cameraReader/n21 [14]),
    .en(~CSI_RST_pad_neg),
    .reset(1'b0),
    .set(1'b0),
    .q(camera_addr[14]));  // sources/rtl/cameraReader.v(95)
  reg_ar_as_w1 \u_cameraReader/reg2_b15  (
    .clk(CSI_PCLK_pad),
    .d(\u_cameraReader/n21 [15]),
    .en(~CSI_RST_pad_neg),
    .reset(1'b0),
    .set(1'b0),
    .q(camera_addr[15]));  // sources/rtl/cameraReader.v(95)
  reg_ar_as_w1 \u_cameraReader/reg2_b2  (
    .clk(CSI_PCLK_pad),
    .d(\u_cameraReader/n21 [2]),
    .en(~CSI_RST_pad_neg),
    .reset(1'b0),
    .set(1'b0),
    .q(camera_addr[2]));  // sources/rtl/cameraReader.v(95)
  reg_ar_as_w1 \u_cameraReader/reg2_b3  (
    .clk(CSI_PCLK_pad),
    .d(\u_cameraReader/n21 [3]),
    .en(~CSI_RST_pad_neg),
    .reset(1'b0),
    .set(1'b0),
    .q(camera_addr[3]));  // sources/rtl/cameraReader.v(95)
  reg_ar_as_w1 \u_cameraReader/reg2_b4  (
    .clk(CSI_PCLK_pad),
    .d(\u_cameraReader/n21 [4]),
    .en(~CSI_RST_pad_neg),
    .reset(1'b0),
    .set(1'b0),
    .q(camera_addr[4]));  // sources/rtl/cameraReader.v(95)
  reg_ar_as_w1 \u_cameraReader/reg2_b5  (
    .clk(CSI_PCLK_pad),
    .d(\u_cameraReader/n21 [5]),
    .en(~CSI_RST_pad_neg),
    .reset(1'b0),
    .set(1'b0),
    .q(camera_addr[5]));  // sources/rtl/cameraReader.v(95)
  reg_ar_as_w1 \u_cameraReader/reg2_b6  (
    .clk(CSI_PCLK_pad),
    .d(\u_cameraReader/n21 [6]),
    .en(~CSI_RST_pad_neg),
    .reset(1'b0),
    .set(1'b0),
    .q(camera_addr[6]));  // sources/rtl/cameraReader.v(95)
  reg_ar_as_w1 \u_cameraReader/reg2_b7  (
    .clk(CSI_PCLK_pad),
    .d(\u_cameraReader/n21 [7]),
    .en(~CSI_RST_pad_neg),
    .reset(1'b0),
    .set(1'b0),
    .q(camera_addr[7]));  // sources/rtl/cameraReader.v(95)
  reg_ar_as_w1 \u_cameraReader/reg2_b8  (
    .clk(CSI_PCLK_pad),
    .d(\u_cameraReader/n21 [8]),
    .en(~CSI_RST_pad_neg),
    .reset(1'b0),
    .set(1'b0),
    .q(camera_addr[8]));  // sources/rtl/cameraReader.v(95)
  reg_ar_as_w1 \u_cameraReader/reg2_b9  (
    .clk(CSI_PCLK_pad),
    .d(\u_cameraReader/n21 [9]),
    .en(~CSI_RST_pad_neg),
    .reset(1'b0),
    .set(1'b0),
    .q(camera_addr[9]));  // sources/rtl/cameraReader.v(95)
  reg_ar_as_w1 \u_cameraReader/reg3_b0  (
    .clk(CSI_PCLK_pad),
    .d(OD_pad[7]),
    .en(\u_cameraReader/mux14_b0_sel_is_2_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cameraReader/subpixel [0]));  // sources/rtl/cameraReader.v(95)
  reg_ar_as_w1 \u_cameraReader/reg3_b1  (
    .clk(CSI_PCLK_pad),
    .d(OD_pad[6]),
    .en(\u_cameraReader/mux14_b0_sel_is_2_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cameraReader/subpixel [1]));  // sources/rtl/cameraReader.v(95)
  reg_ar_as_w1 \u_cameraReader/reg3_b2  (
    .clk(CSI_PCLK_pad),
    .d(OD_pad[5]),
    .en(\u_cameraReader/mux14_b0_sel_is_2_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cameraReader/subpixel [2]));  // sources/rtl/cameraReader.v(95)
  reg_ar_as_w1 \u_cameraReader/reg3_b3  (
    .clk(CSI_PCLK_pad),
    .d(OD_pad[4]),
    .en(\u_cameraReader/mux14_b0_sel_is_2_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cameraReader/subpixel [3]));  // sources/rtl/cameraReader.v(95)
  reg_ar_as_w1 \u_cameraReader/reg3_b4  (
    .clk(CSI_PCLK_pad),
    .d(OD_pad[3]),
    .en(\u_cameraReader/mux14_b0_sel_is_2_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cameraReader/subpixel [4]));  // sources/rtl/cameraReader.v(95)
  reg_ar_as_w1 \u_cameraReader/reg3_b5  (
    .clk(CSI_PCLK_pad),
    .d(OD_pad[2]),
    .en(\u_cameraReader/mux14_b0_sel_is_2_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cameraReader/subpixel [5]));  // sources/rtl/cameraReader.v(95)
  reg_ar_as_w1 \u_cameraReader/reg3_b6  (
    .clk(CSI_PCLK_pad),
    .d(OD_pad[1]),
    .en(\u_cameraReader/mux14_b0_sel_is_2_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cameraReader/subpixel [6]));  // sources/rtl/cameraReader.v(95)
  reg_ar_as_w1 \u_cameraReader/reg3_b7  (
    .clk(CSI_PCLK_pad),
    .d(OD_pad[0]),
    .en(\u_cameraReader/mux14_b0_sel_is_2_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cameraReader/subpixel [7]));  // sources/rtl/cameraReader.v(95)
  reg_ar_as_w1 \u_cameraReader/reg4_b0  (
    .clk(CSI_PCLK_pad),
    .d(OD_pad[7]),
    .en(\u_cameraReader/mux15_b0_sel_is_2_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cameraReader/current_pixel [0]));  // sources/rtl/cameraReader.v(95)
  reg_ar_as_w1 \u_cameraReader/reg4_b1  (
    .clk(CSI_PCLK_pad),
    .d(OD_pad[6]),
    .en(\u_cameraReader/mux15_b0_sel_is_2_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cameraReader/current_pixel [1]));  // sources/rtl/cameraReader.v(95)
  reg_ar_as_w1 \u_cameraReader/reg4_b10  (
    .clk(CSI_PCLK_pad),
    .d(\u_cameraReader/subpixel [2]),
    .en(\u_cameraReader/mux15_b0_sel_is_2_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cameraReader/current_pixel [10]));  // sources/rtl/cameraReader.v(95)
  reg_ar_as_w1 \u_cameraReader/reg4_b11  (
    .clk(CSI_PCLK_pad),
    .d(\u_cameraReader/subpixel [3]),
    .en(\u_cameraReader/mux15_b0_sel_is_2_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cameraReader/current_pixel [11]));  // sources/rtl/cameraReader.v(95)
  reg_ar_as_w1 \u_cameraReader/reg4_b12  (
    .clk(CSI_PCLK_pad),
    .d(\u_cameraReader/subpixel [4]),
    .en(\u_cameraReader/mux15_b0_sel_is_2_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cameraReader/current_pixel [12]));  // sources/rtl/cameraReader.v(95)
  reg_ar_as_w1 \u_cameraReader/reg4_b13  (
    .clk(CSI_PCLK_pad),
    .d(\u_cameraReader/subpixel [5]),
    .en(\u_cameraReader/mux15_b0_sel_is_2_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cameraReader/current_pixel [13]));  // sources/rtl/cameraReader.v(95)
  reg_ar_as_w1 \u_cameraReader/reg4_b14  (
    .clk(CSI_PCLK_pad),
    .d(\u_cameraReader/subpixel [6]),
    .en(\u_cameraReader/mux15_b0_sel_is_2_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cameraReader/current_pixel [14]));  // sources/rtl/cameraReader.v(95)
  reg_ar_as_w1 \u_cameraReader/reg4_b15  (
    .clk(CSI_PCLK_pad),
    .d(\u_cameraReader/subpixel [7]),
    .en(\u_cameraReader/mux15_b0_sel_is_2_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cameraReader/current_pixel [15]));  // sources/rtl/cameraReader.v(95)
  reg_ar_as_w1 \u_cameraReader/reg4_b2  (
    .clk(CSI_PCLK_pad),
    .d(OD_pad[5]),
    .en(\u_cameraReader/mux15_b0_sel_is_2_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cameraReader/current_pixel [2]));  // sources/rtl/cameraReader.v(95)
  reg_ar_as_w1 \u_cameraReader/reg4_b3  (
    .clk(CSI_PCLK_pad),
    .d(OD_pad[4]),
    .en(\u_cameraReader/mux15_b0_sel_is_2_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cameraReader/current_pixel [3]));  // sources/rtl/cameraReader.v(95)
  reg_ar_as_w1 \u_cameraReader/reg4_b4  (
    .clk(CSI_PCLK_pad),
    .d(OD_pad[3]),
    .en(\u_cameraReader/mux15_b0_sel_is_2_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cameraReader/current_pixel [4]));  // sources/rtl/cameraReader.v(95)
  reg_ar_as_w1 \u_cameraReader/reg4_b5  (
    .clk(CSI_PCLK_pad),
    .d(OD_pad[2]),
    .en(\u_cameraReader/mux15_b0_sel_is_2_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cameraReader/current_pixel [5]));  // sources/rtl/cameraReader.v(95)
  reg_ar_as_w1 \u_cameraReader/reg4_b6  (
    .clk(CSI_PCLK_pad),
    .d(OD_pad[1]),
    .en(\u_cameraReader/mux15_b0_sel_is_2_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cameraReader/current_pixel [6]));  // sources/rtl/cameraReader.v(95)
  reg_ar_as_w1 \u_cameraReader/reg4_b7  (
    .clk(CSI_PCLK_pad),
    .d(OD_pad[0]),
    .en(\u_cameraReader/mux15_b0_sel_is_2_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cameraReader/current_pixel [7]));  // sources/rtl/cameraReader.v(95)
  reg_ar_as_w1 \u_cameraReader/reg4_b8  (
    .clk(CSI_PCLK_pad),
    .d(\u_cameraReader/subpixel [0]),
    .en(\u_cameraReader/mux15_b0_sel_is_2_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cameraReader/current_pixel [8]));  // sources/rtl/cameraReader.v(95)
  reg_ar_as_w1 \u_cameraReader/reg4_b9  (
    .clk(CSI_PCLK_pad),
    .d(\u_cameraReader/subpixel [1]),
    .en(\u_cameraReader/mux15_b0_sel_is_2_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cameraReader/current_pixel [9]));  // sources/rtl/cameraReader.v(95)
  reg_sr_as_w1 \u_cameraReader/vsync_passed_reg  (
    .clk(CSI_PCLK_pad),
    .d(\u_cameraReader/vsync_passed_d ),
    .en(1'b1),
    .reset(CSI_RST_pad_neg),
    .set(1'b0),
    .q(\u_cameraReader/vsync_passed ));  // sources/rtl/cameraReader.v(95)
  reg_ar_as_w1 \u_cameraReader/wrclk1_reg  (
    .clk(CSI_PCLK_pad),
    .d(\u_cameraReader/n1 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cameraReader/wrclk1 ));  // sources/rtl/cameraReader.v(29)
  reg_ar_as_w1 \u_cameraReader/write_pixel_reg  (
    .clk(~\u_cameraReader/wrclk1 ),
    .d(\u_cameraReader/n2 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_cameraReader/write_pixel ));  // sources/rtl/cameraReader.v(37)
  camera_init u_camera_init (
    .clk(clk_sccb),
    .reset_n(CSI_RST_pad),
    .sda_in(TESTA_pad),
    .scl(TESTB_pad),
    .sda(sda),
    .sda_oe(sda_oe));  // sources/rtl/test_camera.v(53)
  lcd_sync u_lcd_sync (
    .clk(clk_lcd),
    .rest_n(CSI_RST_pad),
    .addr(lcd_rdaddr),
    .img_ack(lcd_rden),
    .lcd_clk(LCD_CLK_pad),
    .lcd_de(LCD_DEN_pad),
    .lcd_hsync(LCD_HSYNC_pad),
    .lcd_pwm(LCD_PWM_pad),
    .lcd_vsync(LCD_VSYNC_pad));  // sources/rtl/test_camera.v(86)
  // address_offset=0;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("INV"),
    .CSB1("INV"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \uimg/inst_32800x16_sub_000000_000  (
    .addra({camera_addr[9:0],3'b111}),
    .addrb({lcd_rdaddr[9:0],3'b111}),
    .cea(camera_wrreq),
    .ceb(lcd_rden),
    .clka(CSI_PCLK_pad),
    .clkb(clk_lcd),
    .csa({\and_Ncamera_addr[12]_o ,camera_addr[11:10]}),
    .csb({\and_Nlcd_rdaddr[12]__o ,lcd_rdaddr[11:10]}),
    .dia(camera_wrdat[8:0]),
    .rsta(CSI_RST_pad),
    .rstb(CSI_RST_pad),
    .dob({\uimg/inst_dob_i0_008 ,\uimg/inst_dob_i0_007 ,\uimg/inst_dob_i0_006 ,\uimg/inst_dob_i0_005 ,\uimg/inst_dob_i0_004 ,\uimg/inst_dob_i0_003 ,\uimg/inst_dob_i0_002 ,\uimg/inst_dob_i0_001 ,\uimg/inst_dob_i0_000 }));
  // address_offset=0;data_offset=9;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("INV"),
    .CSB1("INV"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \uimg/inst_32800x16_sub_000000_009  (
    .addra(camera_addr[12:0]),
    .addrb(lcd_rdaddr[12:0]),
    .cea(camera_wrreq),
    .ceb(lcd_rden),
    .clka(CSI_PCLK_pad),
    .clkb(clk_lcd),
    .csa(camera_addr[15:13]),
    .csb(lcd_rdaddr[15:13]),
    .dia({open_n1070,open_n1071,open_n1072,open_n1073,open_n1074,open_n1075,open_n1076,camera_wrdat[9],open_n1077}),
    .rsta(CSI_RST_pad),
    .rstb(CSI_RST_pad),
    .dob({open_n1100,open_n1101,open_n1102,open_n1103,open_n1104,open_n1105,open_n1106,open_n1107,\uimg/inst_dob_i0_009 }));
  // address_offset=0;data_offset=10;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("INV"),
    .CSB1("INV"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \uimg/inst_32800x16_sub_000000_010  (
    .addra(camera_addr[12:0]),
    .addrb(lcd_rdaddr[12:0]),
    .cea(camera_wrreq),
    .ceb(lcd_rden),
    .clka(CSI_PCLK_pad),
    .clkb(clk_lcd),
    .csa(camera_addr[15:13]),
    .csb(lcd_rdaddr[15:13]),
    .dia({open_n1108,open_n1109,open_n1110,open_n1111,open_n1112,open_n1113,open_n1114,camera_wrdat[10],open_n1115}),
    .rsta(CSI_RST_pad),
    .rstb(CSI_RST_pad),
    .dob({open_n1138,open_n1139,open_n1140,open_n1141,open_n1142,open_n1143,open_n1144,open_n1145,\uimg/inst_dob_i0_010 }));
  // address_offset=0;data_offset=11;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("INV"),
    .CSB1("INV"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \uimg/inst_32800x16_sub_000000_011  (
    .addra(camera_addr[12:0]),
    .addrb(lcd_rdaddr[12:0]),
    .cea(camera_wrreq),
    .ceb(lcd_rden),
    .clka(CSI_PCLK_pad),
    .clkb(clk_lcd),
    .csa(camera_addr[15:13]),
    .csb(lcd_rdaddr[15:13]),
    .dia({open_n1146,open_n1147,open_n1148,open_n1149,open_n1150,open_n1151,open_n1152,camera_wrdat[11],open_n1153}),
    .rsta(CSI_RST_pad),
    .rstb(CSI_RST_pad),
    .dob({open_n1176,open_n1177,open_n1178,open_n1179,open_n1180,open_n1181,open_n1182,open_n1183,\uimg/inst_dob_i0_011 }));
  // address_offset=0;data_offset=12;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("INV"),
    .CSB1("INV"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \uimg/inst_32800x16_sub_000000_012  (
    .addra(camera_addr[12:0]),
    .addrb(lcd_rdaddr[12:0]),
    .cea(camera_wrreq),
    .ceb(lcd_rden),
    .clka(CSI_PCLK_pad),
    .clkb(clk_lcd),
    .csa(camera_addr[15:13]),
    .csb(lcd_rdaddr[15:13]),
    .dia({open_n1184,open_n1185,open_n1186,open_n1187,open_n1188,open_n1189,open_n1190,camera_wrdat[12],open_n1191}),
    .rsta(CSI_RST_pad),
    .rstb(CSI_RST_pad),
    .dob({open_n1214,open_n1215,open_n1216,open_n1217,open_n1218,open_n1219,open_n1220,open_n1221,\uimg/inst_dob_i0_012 }));
  // address_offset=0;data_offset=13;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("INV"),
    .CSB1("INV"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \uimg/inst_32800x16_sub_000000_013  (
    .addra(camera_addr[12:0]),
    .addrb(lcd_rdaddr[12:0]),
    .cea(camera_wrreq),
    .ceb(lcd_rden),
    .clka(CSI_PCLK_pad),
    .clkb(clk_lcd),
    .csa(camera_addr[15:13]),
    .csb(lcd_rdaddr[15:13]),
    .dia({open_n1222,open_n1223,open_n1224,open_n1225,open_n1226,open_n1227,open_n1228,camera_wrdat[13],open_n1229}),
    .rsta(CSI_RST_pad),
    .rstb(CSI_RST_pad),
    .dob({open_n1252,open_n1253,open_n1254,open_n1255,open_n1256,open_n1257,open_n1258,open_n1259,\uimg/inst_dob_i0_013 }));
  // address_offset=0;data_offset=14;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("INV"),
    .CSB1("INV"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \uimg/inst_32800x16_sub_000000_014  (
    .addra(camera_addr[12:0]),
    .addrb(lcd_rdaddr[12:0]),
    .cea(camera_wrreq),
    .ceb(lcd_rden),
    .clka(CSI_PCLK_pad),
    .clkb(clk_lcd),
    .csa(camera_addr[15:13]),
    .csb(lcd_rdaddr[15:13]),
    .dia({open_n1260,open_n1261,open_n1262,open_n1263,open_n1264,open_n1265,open_n1266,camera_wrdat[14],open_n1267}),
    .rsta(CSI_RST_pad),
    .rstb(CSI_RST_pad),
    .dob({open_n1290,open_n1291,open_n1292,open_n1293,open_n1294,open_n1295,open_n1296,open_n1297,\uimg/inst_dob_i0_014 }));
  // address_offset=0;data_offset=15;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("INV"),
    .CSB1("INV"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \uimg/inst_32800x16_sub_000000_015  (
    .addra(camera_addr[12:0]),
    .addrb(lcd_rdaddr[12:0]),
    .cea(camera_wrreq),
    .ceb(lcd_rden),
    .clka(CSI_PCLK_pad),
    .clkb(clk_lcd),
    .csa(camera_addr[15:13]),
    .csb(lcd_rdaddr[15:13]),
    .dia({open_n1298,open_n1299,open_n1300,open_n1301,open_n1302,open_n1303,open_n1304,camera_wrdat[15],open_n1305}),
    .rsta(CSI_RST_pad),
    .rstb(CSI_RST_pad),
    .dob({open_n1328,open_n1329,open_n1330,open_n1331,open_n1332,open_n1333,open_n1334,open_n1335,\uimg/inst_dob_i0_015 }));
  // address_offset=1024;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("SIG"),
    .CSB1("INV"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \uimg/inst_32800x16_sub_001024_000  (
    .addra({camera_addr[9:0],3'b111}),
    .addrb({lcd_rdaddr[9:0],3'b111}),
    .cea(camera_wrreq),
    .ceb(lcd_rden),
    .clka(CSI_PCLK_pad),
    .clkb(clk_lcd),
    .csa({\and_Ncamera_addr[12]_o ,camera_addr[11:10]}),
    .csb({\and_Nlcd_rdaddr[12]__o ,lcd_rdaddr[11:10]}),
    .dia(camera_wrdat[8:0]),
    .rsta(CSI_RST_pad),
    .rstb(CSI_RST_pad),
    .dob({\uimg/inst_dob_i2_008 ,\uimg/inst_dob_i2_007 ,\uimg/inst_dob_i2_006 ,\uimg/inst_dob_i2_005 ,\uimg/inst_dob_i2_004 ,\uimg/inst_dob_i2_003 ,\uimg/inst_dob_i2_002 ,\uimg/inst_dob_i2_001 ,\uimg/inst_dob_i2_000 }));
  // address_offset=2048;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("INV"),
    .CSB1("SIG"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \uimg/inst_32800x16_sub_002048_000  (
    .addra({camera_addr[9:0],3'b111}),
    .addrb({lcd_rdaddr[9:0],3'b111}),
    .cea(camera_wrreq),
    .ceb(lcd_rden),
    .clka(CSI_PCLK_pad),
    .clkb(clk_lcd),
    .csa({\and_Ncamera_addr[12]_o ,camera_addr[11:10]}),
    .csb({\and_Nlcd_rdaddr[12]__o ,lcd_rdaddr[11:10]}),
    .dia(camera_wrdat[8:0]),
    .rsta(CSI_RST_pad),
    .rstb(CSI_RST_pad),
    .dob({\uimg/inst_dob_i4_008 ,\uimg/inst_dob_i4_007 ,\uimg/inst_dob_i4_006 ,\uimg/inst_dob_i4_005 ,\uimg/inst_dob_i4_004 ,\uimg/inst_dob_i4_003 ,\uimg/inst_dob_i4_002 ,\uimg/inst_dob_i4_001 ,\uimg/inst_dob_i4_000 }));
  // address_offset=3072;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("SIG"),
    .CSB1("SIG"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \uimg/inst_32800x16_sub_003072_000  (
    .addra({camera_addr[9:0],3'b111}),
    .addrb({lcd_rdaddr[9:0],3'b111}),
    .cea(camera_wrreq),
    .ceb(lcd_rden),
    .clka(CSI_PCLK_pad),
    .clkb(clk_lcd),
    .csa({\and_Ncamera_addr[12]_o ,camera_addr[11:10]}),
    .csb({\and_Nlcd_rdaddr[12]__o ,lcd_rdaddr[11:10]}),
    .dia(camera_wrdat[8:0]),
    .rsta(CSI_RST_pad),
    .rstb(CSI_RST_pad),
    .dob({\uimg/inst_dob_i6_008 ,\uimg/inst_dob_i6_007 ,\uimg/inst_dob_i6_006 ,\uimg/inst_dob_i6_005 ,\uimg/inst_dob_i6_004 ,\uimg/inst_dob_i6_003 ,\uimg/inst_dob_i6_002 ,\uimg/inst_dob_i6_001 ,\uimg/inst_dob_i6_000 }));
  // address_offset=4096;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("INV"),
    .CSB1("INV"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \uimg/inst_32800x16_sub_004096_000  (
    .addra({camera_addr[9:0],3'b111}),
    .addrb({lcd_rdaddr[9:0],3'b111}),
    .cea(camera_wrreq),
    .ceb(lcd_rden),
    .clka(CSI_PCLK_pad),
    .clkb(clk_lcd),
    .csa({\and_camera_addr[12]__o ,camera_addr[11:10]}),
    .csb({\and_lcd_rdaddr[12]_N_o ,lcd_rdaddr[11:10]}),
    .dia(camera_wrdat[8:0]),
    .rsta(CSI_RST_pad),
    .rstb(CSI_RST_pad),
    .dob({\uimg/inst_dob_i8_008 ,\uimg/inst_dob_i8_007 ,\uimg/inst_dob_i8_006 ,\uimg/inst_dob_i8_005 ,\uimg/inst_dob_i8_004 ,\uimg/inst_dob_i8_003 ,\uimg/inst_dob_i8_002 ,\uimg/inst_dob_i8_001 ,\uimg/inst_dob_i8_000 }));
  // address_offset=5120;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("SIG"),
    .CSB1("INV"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \uimg/inst_32800x16_sub_005120_000  (
    .addra({camera_addr[9:0],3'b111}),
    .addrb({lcd_rdaddr[9:0],3'b111}),
    .cea(camera_wrreq),
    .ceb(lcd_rden),
    .clka(CSI_PCLK_pad),
    .clkb(clk_lcd),
    .csa({\and_camera_addr[12]__o ,camera_addr[11:10]}),
    .csb({\and_lcd_rdaddr[12]_N_o ,lcd_rdaddr[11:10]}),
    .dia(camera_wrdat[8:0]),
    .rsta(CSI_RST_pad),
    .rstb(CSI_RST_pad),
    .dob({\uimg/inst_dob_i10_008 ,\uimg/inst_dob_i10_007 ,\uimg/inst_dob_i10_006 ,\uimg/inst_dob_i10_005 ,\uimg/inst_dob_i10_004 ,\uimg/inst_dob_i10_003 ,\uimg/inst_dob_i10_002 ,\uimg/inst_dob_i10_001 ,\uimg/inst_dob_i10_000 }));
  // address_offset=6144;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("INV"),
    .CSB1("SIG"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \uimg/inst_32800x16_sub_006144_000  (
    .addra({camera_addr[9:0],3'b111}),
    .addrb({lcd_rdaddr[9:0],3'b111}),
    .cea(camera_wrreq),
    .ceb(lcd_rden),
    .clka(CSI_PCLK_pad),
    .clkb(clk_lcd),
    .csa({\and_camera_addr[12]__o ,camera_addr[11:10]}),
    .csb({\and_lcd_rdaddr[12]_N_o ,lcd_rdaddr[11:10]}),
    .dia(camera_wrdat[8:0]),
    .rsta(CSI_RST_pad),
    .rstb(CSI_RST_pad),
    .dob({\uimg/inst_dob_i12_008 ,\uimg/inst_dob_i12_007 ,\uimg/inst_dob_i12_006 ,\uimg/inst_dob_i12_005 ,\uimg/inst_dob_i12_004 ,\uimg/inst_dob_i12_003 ,\uimg/inst_dob_i12_002 ,\uimg/inst_dob_i12_001 ,\uimg/inst_dob_i12_000 }));
  // address_offset=7168;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("SIG"),
    .CSB1("SIG"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \uimg/inst_32800x16_sub_007168_000  (
    .addra({camera_addr[9:0],3'b111}),
    .addrb({lcd_rdaddr[9:0],3'b111}),
    .cea(camera_wrreq),
    .ceb(lcd_rden),
    .clka(CSI_PCLK_pad),
    .clkb(clk_lcd),
    .csa({\and_camera_addr[12]__o ,camera_addr[11:10]}),
    .csb({\and_lcd_rdaddr[12]_N_o ,lcd_rdaddr[11:10]}),
    .dia(camera_wrdat[8:0]),
    .rsta(CSI_RST_pad),
    .rstb(CSI_RST_pad),
    .dob({\uimg/inst_dob_i14_008 ,\uimg/inst_dob_i14_007 ,\uimg/inst_dob_i14_006 ,\uimg/inst_dob_i14_005 ,\uimg/inst_dob_i14_004 ,\uimg/inst_dob_i14_003 ,\uimg/inst_dob_i14_002 ,\uimg/inst_dob_i14_001 ,\uimg/inst_dob_i14_000 }));
  // address_offset=8192;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("INV"),
    .CSB1("INV"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \uimg/inst_32800x16_sub_008192_000  (
    .addra({camera_addr[9:0],3'b111}),
    .addrb({lcd_rdaddr[9:0],3'b111}),
    .cea(camera_wrreq),
    .ceb(lcd_rden),
    .clka(CSI_PCLK_pad),
    .clkb(clk_lcd),
    .csa({\and_Ncamera_addr[12]_o_al_n197 ,camera_addr[11:10]}),
    .csb({\and_Nlcd_rdaddr[12]__o_al_n200 ,lcd_rdaddr[11:10]}),
    .dia(camera_wrdat[8:0]),
    .rsta(CSI_RST_pad),
    .rstb(CSI_RST_pad),
    .dob({\uimg/inst_dob_i16_008 ,\uimg/inst_dob_i16_007 ,\uimg/inst_dob_i16_006 ,\uimg/inst_dob_i16_005 ,\uimg/inst_dob_i16_004 ,\uimg/inst_dob_i16_003 ,\uimg/inst_dob_i16_002 ,\uimg/inst_dob_i16_001 ,\uimg/inst_dob_i16_000 }));
  // address_offset=8192;data_offset=9;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("SIG"),
    .CSB1("INV"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \uimg/inst_32800x16_sub_008192_009  (
    .addra(camera_addr[12:0]),
    .addrb(lcd_rdaddr[12:0]),
    .cea(camera_wrreq),
    .ceb(lcd_rden),
    .clka(CSI_PCLK_pad),
    .clkb(clk_lcd),
    .csa(camera_addr[15:13]),
    .csb(lcd_rdaddr[15:13]),
    .dia({open_n1512,open_n1513,open_n1514,open_n1515,open_n1516,open_n1517,open_n1518,camera_wrdat[9],open_n1519}),
    .rsta(CSI_RST_pad),
    .rstb(CSI_RST_pad),
    .dob({open_n1542,open_n1543,open_n1544,open_n1545,open_n1546,open_n1547,open_n1548,open_n1549,\uimg/inst_dob_i16_009 }));
  // address_offset=8192;data_offset=10;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("SIG"),
    .CSB1("INV"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \uimg/inst_32800x16_sub_008192_010  (
    .addra(camera_addr[12:0]),
    .addrb(lcd_rdaddr[12:0]),
    .cea(camera_wrreq),
    .ceb(lcd_rden),
    .clka(CSI_PCLK_pad),
    .clkb(clk_lcd),
    .csa(camera_addr[15:13]),
    .csb(lcd_rdaddr[15:13]),
    .dia({open_n1550,open_n1551,open_n1552,open_n1553,open_n1554,open_n1555,open_n1556,camera_wrdat[10],open_n1557}),
    .rsta(CSI_RST_pad),
    .rstb(CSI_RST_pad),
    .dob({open_n1580,open_n1581,open_n1582,open_n1583,open_n1584,open_n1585,open_n1586,open_n1587,\uimg/inst_dob_i16_010 }));
  // address_offset=8192;data_offset=11;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("SIG"),
    .CSB1("INV"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \uimg/inst_32800x16_sub_008192_011  (
    .addra(camera_addr[12:0]),
    .addrb(lcd_rdaddr[12:0]),
    .cea(camera_wrreq),
    .ceb(lcd_rden),
    .clka(CSI_PCLK_pad),
    .clkb(clk_lcd),
    .csa(camera_addr[15:13]),
    .csb(lcd_rdaddr[15:13]),
    .dia({open_n1588,open_n1589,open_n1590,open_n1591,open_n1592,open_n1593,open_n1594,camera_wrdat[11],open_n1595}),
    .rsta(CSI_RST_pad),
    .rstb(CSI_RST_pad),
    .dob({open_n1618,open_n1619,open_n1620,open_n1621,open_n1622,open_n1623,open_n1624,open_n1625,\uimg/inst_dob_i16_011 }));
  // address_offset=8192;data_offset=12;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("SIG"),
    .CSB1("INV"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \uimg/inst_32800x16_sub_008192_012  (
    .addra(camera_addr[12:0]),
    .addrb(lcd_rdaddr[12:0]),
    .cea(camera_wrreq),
    .ceb(lcd_rden),
    .clka(CSI_PCLK_pad),
    .clkb(clk_lcd),
    .csa(camera_addr[15:13]),
    .csb(lcd_rdaddr[15:13]),
    .dia({open_n1626,open_n1627,open_n1628,open_n1629,open_n1630,open_n1631,open_n1632,camera_wrdat[12],open_n1633}),
    .rsta(CSI_RST_pad),
    .rstb(CSI_RST_pad),
    .dob({open_n1656,open_n1657,open_n1658,open_n1659,open_n1660,open_n1661,open_n1662,open_n1663,\uimg/inst_dob_i16_012 }));
  // address_offset=8192;data_offset=13;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("SIG"),
    .CSB1("INV"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \uimg/inst_32800x16_sub_008192_013  (
    .addra(camera_addr[12:0]),
    .addrb(lcd_rdaddr[12:0]),
    .cea(camera_wrreq),
    .ceb(lcd_rden),
    .clka(CSI_PCLK_pad),
    .clkb(clk_lcd),
    .csa(camera_addr[15:13]),
    .csb(lcd_rdaddr[15:13]),
    .dia({open_n1664,open_n1665,open_n1666,open_n1667,open_n1668,open_n1669,open_n1670,camera_wrdat[13],open_n1671}),
    .rsta(CSI_RST_pad),
    .rstb(CSI_RST_pad),
    .dob({open_n1694,open_n1695,open_n1696,open_n1697,open_n1698,open_n1699,open_n1700,open_n1701,\uimg/inst_dob_i16_013 }));
  // address_offset=8192;data_offset=14;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("SIG"),
    .CSB1("INV"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \uimg/inst_32800x16_sub_008192_014  (
    .addra(camera_addr[12:0]),
    .addrb(lcd_rdaddr[12:0]),
    .cea(camera_wrreq),
    .ceb(lcd_rden),
    .clka(CSI_PCLK_pad),
    .clkb(clk_lcd),
    .csa(camera_addr[15:13]),
    .csb(lcd_rdaddr[15:13]),
    .dia({open_n1702,open_n1703,open_n1704,open_n1705,open_n1706,open_n1707,open_n1708,camera_wrdat[14],open_n1709}),
    .rsta(CSI_RST_pad),
    .rstb(CSI_RST_pad),
    .dob({open_n1732,open_n1733,open_n1734,open_n1735,open_n1736,open_n1737,open_n1738,open_n1739,\uimg/inst_dob_i16_014 }));
  // address_offset=8192;data_offset=15;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("SIG"),
    .CSB1("INV"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \uimg/inst_32800x16_sub_008192_015  (
    .addra(camera_addr[12:0]),
    .addrb(lcd_rdaddr[12:0]),
    .cea(camera_wrreq),
    .ceb(lcd_rden),
    .clka(CSI_PCLK_pad),
    .clkb(clk_lcd),
    .csa(camera_addr[15:13]),
    .csb(lcd_rdaddr[15:13]),
    .dia({open_n1740,open_n1741,open_n1742,open_n1743,open_n1744,open_n1745,open_n1746,camera_wrdat[15],open_n1747}),
    .rsta(CSI_RST_pad),
    .rstb(CSI_RST_pad),
    .dob({open_n1770,open_n1771,open_n1772,open_n1773,open_n1774,open_n1775,open_n1776,open_n1777,\uimg/inst_dob_i16_015 }));
  // address_offset=9216;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("SIG"),
    .CSB1("INV"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \uimg/inst_32800x16_sub_009216_000  (
    .addra({camera_addr[9:0],3'b111}),
    .addrb({lcd_rdaddr[9:0],3'b111}),
    .cea(camera_wrreq),
    .ceb(lcd_rden),
    .clka(CSI_PCLK_pad),
    .clkb(clk_lcd),
    .csa({\and_Ncamera_addr[12]_o_al_n197 ,camera_addr[11:10]}),
    .csb({\and_Nlcd_rdaddr[12]__o_al_n200 ,lcd_rdaddr[11:10]}),
    .dia(camera_wrdat[8:0]),
    .rsta(CSI_RST_pad),
    .rstb(CSI_RST_pad),
    .dob({\uimg/inst_dob_i18_008 ,\uimg/inst_dob_i18_007 ,\uimg/inst_dob_i18_006 ,\uimg/inst_dob_i18_005 ,\uimg/inst_dob_i18_004 ,\uimg/inst_dob_i18_003 ,\uimg/inst_dob_i18_002 ,\uimg/inst_dob_i18_001 ,\uimg/inst_dob_i18_000 }));
  // address_offset=10240;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("INV"),
    .CSB1("SIG"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \uimg/inst_32800x16_sub_010240_000  (
    .addra({camera_addr[9:0],3'b111}),
    .addrb({lcd_rdaddr[9:0],3'b111}),
    .cea(camera_wrreq),
    .ceb(lcd_rden),
    .clka(CSI_PCLK_pad),
    .clkb(clk_lcd),
    .csa({\and_Ncamera_addr[12]_o_al_n197 ,camera_addr[11:10]}),
    .csb({\and_Nlcd_rdaddr[12]__o_al_n200 ,lcd_rdaddr[11:10]}),
    .dia(camera_wrdat[8:0]),
    .rsta(CSI_RST_pad),
    .rstb(CSI_RST_pad),
    .dob({\uimg/inst_dob_i20_008 ,\uimg/inst_dob_i20_007 ,\uimg/inst_dob_i20_006 ,\uimg/inst_dob_i20_005 ,\uimg/inst_dob_i20_004 ,\uimg/inst_dob_i20_003 ,\uimg/inst_dob_i20_002 ,\uimg/inst_dob_i20_001 ,\uimg/inst_dob_i20_000 }));
  // address_offset=11264;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("SIG"),
    .CSB1("SIG"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \uimg/inst_32800x16_sub_011264_000  (
    .addra({camera_addr[9:0],3'b111}),
    .addrb({lcd_rdaddr[9:0],3'b111}),
    .cea(camera_wrreq),
    .ceb(lcd_rden),
    .clka(CSI_PCLK_pad),
    .clkb(clk_lcd),
    .csa({\and_Ncamera_addr[12]_o_al_n197 ,camera_addr[11:10]}),
    .csb({\and_Nlcd_rdaddr[12]__o_al_n200 ,lcd_rdaddr[11:10]}),
    .dia(camera_wrdat[8:0]),
    .rsta(CSI_RST_pad),
    .rstb(CSI_RST_pad),
    .dob({\uimg/inst_dob_i22_008 ,\uimg/inst_dob_i22_007 ,\uimg/inst_dob_i22_006 ,\uimg/inst_dob_i22_005 ,\uimg/inst_dob_i22_004 ,\uimg/inst_dob_i22_003 ,\uimg/inst_dob_i22_002 ,\uimg/inst_dob_i22_001 ,\uimg/inst_dob_i22_000 }));
  // address_offset=12288;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("INV"),
    .CSB1("INV"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \uimg/inst_32800x16_sub_012288_000  (
    .addra({camera_addr[9:0],3'b111}),
    .addrb({lcd_rdaddr[9:0],3'b111}),
    .cea(camera_wrreq),
    .ceb(lcd_rden),
    .clka(CSI_PCLK_pad),
    .clkb(clk_lcd),
    .csa({\and_camera_addr[12]__o_al_n213 ,camera_addr[11:10]}),
    .csb({\and_lcd_rdaddr[12]_l_o ,lcd_rdaddr[11:10]}),
    .dia(camera_wrdat[8:0]),
    .rsta(CSI_RST_pad),
    .rstb(CSI_RST_pad),
    .dob({\uimg/inst_dob_i24_008 ,\uimg/inst_dob_i24_007 ,\uimg/inst_dob_i24_006 ,\uimg/inst_dob_i24_005 ,\uimg/inst_dob_i24_004 ,\uimg/inst_dob_i24_003 ,\uimg/inst_dob_i24_002 ,\uimg/inst_dob_i24_001 ,\uimg/inst_dob_i24_000 }));
  // address_offset=13312;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("SIG"),
    .CSB1("INV"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \uimg/inst_32800x16_sub_013312_000  (
    .addra({camera_addr[9:0],3'b111}),
    .addrb({lcd_rdaddr[9:0],3'b111}),
    .cea(camera_wrreq),
    .ceb(lcd_rden),
    .clka(CSI_PCLK_pad),
    .clkb(clk_lcd),
    .csa({\and_camera_addr[12]__o_al_n213 ,camera_addr[11:10]}),
    .csb({\and_lcd_rdaddr[12]_l_o ,lcd_rdaddr[11:10]}),
    .dia(camera_wrdat[8:0]),
    .rsta(CSI_RST_pad),
    .rstb(CSI_RST_pad),
    .dob({\uimg/inst_dob_i26_008 ,\uimg/inst_dob_i26_007 ,\uimg/inst_dob_i26_006 ,\uimg/inst_dob_i26_005 ,\uimg/inst_dob_i26_004 ,\uimg/inst_dob_i26_003 ,\uimg/inst_dob_i26_002 ,\uimg/inst_dob_i26_001 ,\uimg/inst_dob_i26_000 }));
  // address_offset=14336;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("INV"),
    .CSB1("SIG"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \uimg/inst_32800x16_sub_014336_000  (
    .addra({camera_addr[9:0],3'b111}),
    .addrb({lcd_rdaddr[9:0],3'b111}),
    .cea(camera_wrreq),
    .ceb(lcd_rden),
    .clka(CSI_PCLK_pad),
    .clkb(clk_lcd),
    .csa({\and_camera_addr[12]__o_al_n213 ,camera_addr[11:10]}),
    .csb({\and_lcd_rdaddr[12]_l_o ,lcd_rdaddr[11:10]}),
    .dia(camera_wrdat[8:0]),
    .rsta(CSI_RST_pad),
    .rstb(CSI_RST_pad),
    .dob({\uimg/inst_dob_i28_008 ,\uimg/inst_dob_i28_007 ,\uimg/inst_dob_i28_006 ,\uimg/inst_dob_i28_005 ,\uimg/inst_dob_i28_004 ,\uimg/inst_dob_i28_003 ,\uimg/inst_dob_i28_002 ,\uimg/inst_dob_i28_001 ,\uimg/inst_dob_i28_000 }));
  // address_offset=15360;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("SIG"),
    .CSB1("SIG"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \uimg/inst_32800x16_sub_015360_000  (
    .addra({camera_addr[9:0],3'b111}),
    .addrb({lcd_rdaddr[9:0],3'b111}),
    .cea(camera_wrreq),
    .ceb(lcd_rden),
    .clka(CSI_PCLK_pad),
    .clkb(clk_lcd),
    .csa({\and_camera_addr[12]__o_al_n213 ,camera_addr[11:10]}),
    .csb({\and_lcd_rdaddr[12]_l_o ,lcd_rdaddr[11:10]}),
    .dia(camera_wrdat[8:0]),
    .rsta(CSI_RST_pad),
    .rstb(CSI_RST_pad),
    .dob({\uimg/inst_dob_i30_008 ,\uimg/inst_dob_i30_007 ,\uimg/inst_dob_i30_006 ,\uimg/inst_dob_i30_005 ,\uimg/inst_dob_i30_004 ,\uimg/inst_dob_i30_003 ,\uimg/inst_dob_i30_002 ,\uimg/inst_dob_i30_001 ,\uimg/inst_dob_i30_000 }));
  // address_offset=16384;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("INV"),
    .CSB1("INV"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \uimg/inst_32800x16_sub_016384_000  (
    .addra({camera_addr[9:0],3'b111}),
    .addrb({lcd_rdaddr[9:0],3'b111}),
    .cea(camera_wrreq),
    .ceb(lcd_rden),
    .clka(CSI_PCLK_pad),
    .clkb(clk_lcd),
    .csa({\and_Ncamera_addr[12]_o_al_n228 ,camera_addr[11:10]}),
    .csb({\and_Nlcd_rdaddr[12]__o_al_n231 ,lcd_rdaddr[11:10]}),
    .dia(camera_wrdat[8:0]),
    .rsta(CSI_RST_pad),
    .rstb(CSI_RST_pad),
    .dob({\uimg/inst_dob_i32_008 ,\uimg/inst_dob_i32_007 ,\uimg/inst_dob_i32_006 ,\uimg/inst_dob_i32_005 ,\uimg/inst_dob_i32_004 ,\uimg/inst_dob_i32_003 ,\uimg/inst_dob_i32_002 ,\uimg/inst_dob_i32_001 ,\uimg/inst_dob_i32_000 }));
  // address_offset=16384;data_offset=9;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("INV"),
    .CSB1("SIG"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \uimg/inst_32800x16_sub_016384_009  (
    .addra(camera_addr[12:0]),
    .addrb(lcd_rdaddr[12:0]),
    .cea(camera_wrreq),
    .ceb(lcd_rden),
    .clka(CSI_PCLK_pad),
    .clkb(clk_lcd),
    .csa(camera_addr[15:13]),
    .csb(lcd_rdaddr[15:13]),
    .dia({open_n1954,open_n1955,open_n1956,open_n1957,open_n1958,open_n1959,open_n1960,camera_wrdat[9],open_n1961}),
    .rsta(CSI_RST_pad),
    .rstb(CSI_RST_pad),
    .dob({open_n1984,open_n1985,open_n1986,open_n1987,open_n1988,open_n1989,open_n1990,open_n1991,\uimg/inst_dob_i32_009 }));
  // address_offset=16384;data_offset=10;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("INV"),
    .CSB1("SIG"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \uimg/inst_32800x16_sub_016384_010  (
    .addra(camera_addr[12:0]),
    .addrb(lcd_rdaddr[12:0]),
    .cea(camera_wrreq),
    .ceb(lcd_rden),
    .clka(CSI_PCLK_pad),
    .clkb(clk_lcd),
    .csa(camera_addr[15:13]),
    .csb(lcd_rdaddr[15:13]),
    .dia({open_n1992,open_n1993,open_n1994,open_n1995,open_n1996,open_n1997,open_n1998,camera_wrdat[10],open_n1999}),
    .rsta(CSI_RST_pad),
    .rstb(CSI_RST_pad),
    .dob({open_n2022,open_n2023,open_n2024,open_n2025,open_n2026,open_n2027,open_n2028,open_n2029,\uimg/inst_dob_i32_010 }));
  // address_offset=16384;data_offset=11;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("INV"),
    .CSB1("SIG"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \uimg/inst_32800x16_sub_016384_011  (
    .addra(camera_addr[12:0]),
    .addrb(lcd_rdaddr[12:0]),
    .cea(camera_wrreq),
    .ceb(lcd_rden),
    .clka(CSI_PCLK_pad),
    .clkb(clk_lcd),
    .csa(camera_addr[15:13]),
    .csb(lcd_rdaddr[15:13]),
    .dia({open_n2030,open_n2031,open_n2032,open_n2033,open_n2034,open_n2035,open_n2036,camera_wrdat[11],open_n2037}),
    .rsta(CSI_RST_pad),
    .rstb(CSI_RST_pad),
    .dob({open_n2060,open_n2061,open_n2062,open_n2063,open_n2064,open_n2065,open_n2066,open_n2067,\uimg/inst_dob_i32_011 }));
  // address_offset=16384;data_offset=12;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("INV"),
    .CSB1("SIG"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \uimg/inst_32800x16_sub_016384_012  (
    .addra(camera_addr[12:0]),
    .addrb(lcd_rdaddr[12:0]),
    .cea(camera_wrreq),
    .ceb(lcd_rden),
    .clka(CSI_PCLK_pad),
    .clkb(clk_lcd),
    .csa(camera_addr[15:13]),
    .csb(lcd_rdaddr[15:13]),
    .dia({open_n2068,open_n2069,open_n2070,open_n2071,open_n2072,open_n2073,open_n2074,camera_wrdat[12],open_n2075}),
    .rsta(CSI_RST_pad),
    .rstb(CSI_RST_pad),
    .dob({open_n2098,open_n2099,open_n2100,open_n2101,open_n2102,open_n2103,open_n2104,open_n2105,\uimg/inst_dob_i32_012 }));
  // address_offset=16384;data_offset=13;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("INV"),
    .CSB1("SIG"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \uimg/inst_32800x16_sub_016384_013  (
    .addra(camera_addr[12:0]),
    .addrb(lcd_rdaddr[12:0]),
    .cea(camera_wrreq),
    .ceb(lcd_rden),
    .clka(CSI_PCLK_pad),
    .clkb(clk_lcd),
    .csa(camera_addr[15:13]),
    .csb(lcd_rdaddr[15:13]),
    .dia({open_n2106,open_n2107,open_n2108,open_n2109,open_n2110,open_n2111,open_n2112,camera_wrdat[13],open_n2113}),
    .rsta(CSI_RST_pad),
    .rstb(CSI_RST_pad),
    .dob({open_n2136,open_n2137,open_n2138,open_n2139,open_n2140,open_n2141,open_n2142,open_n2143,\uimg/inst_dob_i32_013 }));
  // address_offset=16384;data_offset=14;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("INV"),
    .CSB1("SIG"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \uimg/inst_32800x16_sub_016384_014  (
    .addra(camera_addr[12:0]),
    .addrb(lcd_rdaddr[12:0]),
    .cea(camera_wrreq),
    .ceb(lcd_rden),
    .clka(CSI_PCLK_pad),
    .clkb(clk_lcd),
    .csa(camera_addr[15:13]),
    .csb(lcd_rdaddr[15:13]),
    .dia({open_n2144,open_n2145,open_n2146,open_n2147,open_n2148,open_n2149,open_n2150,camera_wrdat[14],open_n2151}),
    .rsta(CSI_RST_pad),
    .rstb(CSI_RST_pad),
    .dob({open_n2174,open_n2175,open_n2176,open_n2177,open_n2178,open_n2179,open_n2180,open_n2181,\uimg/inst_dob_i32_014 }));
  // address_offset=16384;data_offset=15;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("INV"),
    .CSB1("SIG"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \uimg/inst_32800x16_sub_016384_015  (
    .addra(camera_addr[12:0]),
    .addrb(lcd_rdaddr[12:0]),
    .cea(camera_wrreq),
    .ceb(lcd_rden),
    .clka(CSI_PCLK_pad),
    .clkb(clk_lcd),
    .csa(camera_addr[15:13]),
    .csb(lcd_rdaddr[15:13]),
    .dia({open_n2182,open_n2183,open_n2184,open_n2185,open_n2186,open_n2187,open_n2188,camera_wrdat[15],open_n2189}),
    .rsta(CSI_RST_pad),
    .rstb(CSI_RST_pad),
    .dob({open_n2212,open_n2213,open_n2214,open_n2215,open_n2216,open_n2217,open_n2218,open_n2219,\uimg/inst_dob_i32_015 }));
  // address_offset=17408;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("SIG"),
    .CSB1("INV"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \uimg/inst_32800x16_sub_017408_000  (
    .addra({camera_addr[9:0],3'b111}),
    .addrb({lcd_rdaddr[9:0],3'b111}),
    .cea(camera_wrreq),
    .ceb(lcd_rden),
    .clka(CSI_PCLK_pad),
    .clkb(clk_lcd),
    .csa({\and_Ncamera_addr[12]_o_al_n228 ,camera_addr[11:10]}),
    .csb({\and_Nlcd_rdaddr[12]__o_al_n231 ,lcd_rdaddr[11:10]}),
    .dia(camera_wrdat[8:0]),
    .rsta(CSI_RST_pad),
    .rstb(CSI_RST_pad),
    .dob({\uimg/inst_dob_i34_008 ,\uimg/inst_dob_i34_007 ,\uimg/inst_dob_i34_006 ,\uimg/inst_dob_i34_005 ,\uimg/inst_dob_i34_004 ,\uimg/inst_dob_i34_003 ,\uimg/inst_dob_i34_002 ,\uimg/inst_dob_i34_001 ,\uimg/inst_dob_i34_000 }));
  // address_offset=18432;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("INV"),
    .CSB1("SIG"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \uimg/inst_32800x16_sub_018432_000  (
    .addra({camera_addr[9:0],3'b111}),
    .addrb({lcd_rdaddr[9:0],3'b111}),
    .cea(camera_wrreq),
    .ceb(lcd_rden),
    .clka(CSI_PCLK_pad),
    .clkb(clk_lcd),
    .csa({\and_Ncamera_addr[12]_o_al_n228 ,camera_addr[11:10]}),
    .csb({\and_Nlcd_rdaddr[12]__o_al_n231 ,lcd_rdaddr[11:10]}),
    .dia(camera_wrdat[8:0]),
    .rsta(CSI_RST_pad),
    .rstb(CSI_RST_pad),
    .dob({\uimg/inst_dob_i36_008 ,\uimg/inst_dob_i36_007 ,\uimg/inst_dob_i36_006 ,\uimg/inst_dob_i36_005 ,\uimg/inst_dob_i36_004 ,\uimg/inst_dob_i36_003 ,\uimg/inst_dob_i36_002 ,\uimg/inst_dob_i36_001 ,\uimg/inst_dob_i36_000 }));
  // address_offset=19456;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("SIG"),
    .CSB1("SIG"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \uimg/inst_32800x16_sub_019456_000  (
    .addra({camera_addr[9:0],3'b111}),
    .addrb({lcd_rdaddr[9:0],3'b111}),
    .cea(camera_wrreq),
    .ceb(lcd_rden),
    .clka(CSI_PCLK_pad),
    .clkb(clk_lcd),
    .csa({\and_Ncamera_addr[12]_o_al_n228 ,camera_addr[11:10]}),
    .csb({\and_Nlcd_rdaddr[12]__o_al_n231 ,lcd_rdaddr[11:10]}),
    .dia(camera_wrdat[8:0]),
    .rsta(CSI_RST_pad),
    .rstb(CSI_RST_pad),
    .dob({\uimg/inst_dob_i38_008 ,\uimg/inst_dob_i38_007 ,\uimg/inst_dob_i38_006 ,\uimg/inst_dob_i38_005 ,\uimg/inst_dob_i38_004 ,\uimg/inst_dob_i38_003 ,\uimg/inst_dob_i38_002 ,\uimg/inst_dob_i38_001 ,\uimg/inst_dob_i38_000 }));
  // address_offset=20480;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("INV"),
    .CSB1("INV"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \uimg/inst_32800x16_sub_020480_000  (
    .addra({camera_addr[9:0],3'b111}),
    .addrb({lcd_rdaddr[9:0],3'b111}),
    .cea(camera_wrreq),
    .ceb(lcd_rden),
    .clka(CSI_PCLK_pad),
    .clkb(clk_lcd),
    .csa({\and_camera_addr[12]__o_al_n244 ,camera_addr[11:10]}),
    .csb({\and_lcd_rdaddr[12]_N_o_al_n247 ,lcd_rdaddr[11:10]}),
    .dia(camera_wrdat[8:0]),
    .rsta(CSI_RST_pad),
    .rstb(CSI_RST_pad),
    .dob({\uimg/inst_dob_i40_008 ,\uimg/inst_dob_i40_007 ,\uimg/inst_dob_i40_006 ,\uimg/inst_dob_i40_005 ,\uimg/inst_dob_i40_004 ,\uimg/inst_dob_i40_003 ,\uimg/inst_dob_i40_002 ,\uimg/inst_dob_i40_001 ,\uimg/inst_dob_i40_000 }));
  // address_offset=21504;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("SIG"),
    .CSB1("INV"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \uimg/inst_32800x16_sub_021504_000  (
    .addra({camera_addr[9:0],3'b111}),
    .addrb({lcd_rdaddr[9:0],3'b111}),
    .cea(camera_wrreq),
    .ceb(lcd_rden),
    .clka(CSI_PCLK_pad),
    .clkb(clk_lcd),
    .csa({\and_camera_addr[12]__o_al_n244 ,camera_addr[11:10]}),
    .csb({\and_lcd_rdaddr[12]_N_o_al_n247 ,lcd_rdaddr[11:10]}),
    .dia(camera_wrdat[8:0]),
    .rsta(CSI_RST_pad),
    .rstb(CSI_RST_pad),
    .dob({\uimg/inst_dob_i42_008 ,\uimg/inst_dob_i42_007 ,\uimg/inst_dob_i42_006 ,\uimg/inst_dob_i42_005 ,\uimg/inst_dob_i42_004 ,\uimg/inst_dob_i42_003 ,\uimg/inst_dob_i42_002 ,\uimg/inst_dob_i42_001 ,\uimg/inst_dob_i42_000 }));
  // address_offset=22528;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("INV"),
    .CSB1("SIG"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \uimg/inst_32800x16_sub_022528_000  (
    .addra({camera_addr[9:0],3'b111}),
    .addrb({lcd_rdaddr[9:0],3'b111}),
    .cea(camera_wrreq),
    .ceb(lcd_rden),
    .clka(CSI_PCLK_pad),
    .clkb(clk_lcd),
    .csa({\and_camera_addr[12]__o_al_n244 ,camera_addr[11:10]}),
    .csb({\and_lcd_rdaddr[12]_N_o_al_n247 ,lcd_rdaddr[11:10]}),
    .dia(camera_wrdat[8:0]),
    .rsta(CSI_RST_pad),
    .rstb(CSI_RST_pad),
    .dob({\uimg/inst_dob_i44_008 ,\uimg/inst_dob_i44_007 ,\uimg/inst_dob_i44_006 ,\uimg/inst_dob_i44_005 ,\uimg/inst_dob_i44_004 ,\uimg/inst_dob_i44_003 ,\uimg/inst_dob_i44_002 ,\uimg/inst_dob_i44_001 ,\uimg/inst_dob_i44_000 }));
  // address_offset=23552;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("SIG"),
    .CSB1("SIG"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \uimg/inst_32800x16_sub_023552_000  (
    .addra({camera_addr[9:0],3'b111}),
    .addrb({lcd_rdaddr[9:0],3'b111}),
    .cea(camera_wrreq),
    .ceb(lcd_rden),
    .clka(CSI_PCLK_pad),
    .clkb(clk_lcd),
    .csa({\and_camera_addr[12]__o_al_n244 ,camera_addr[11:10]}),
    .csb({\and_lcd_rdaddr[12]_N_o_al_n247 ,lcd_rdaddr[11:10]}),
    .dia(camera_wrdat[8:0]),
    .rsta(CSI_RST_pad),
    .rstb(CSI_RST_pad),
    .dob({\uimg/inst_dob_i46_008 ,\uimg/inst_dob_i46_007 ,\uimg/inst_dob_i46_006 ,\uimg/inst_dob_i46_005 ,\uimg/inst_dob_i46_004 ,\uimg/inst_dob_i46_003 ,\uimg/inst_dob_i46_002 ,\uimg/inst_dob_i46_001 ,\uimg/inst_dob_i46_000 }));
  // address_offset=24576;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("INV"),
    .CSB1("INV"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \uimg/inst_32800x16_sub_024576_000  (
    .addra({camera_addr[9:0],3'b111}),
    .addrb({lcd_rdaddr[9:0],3'b111}),
    .cea(camera_wrreq),
    .ceb(lcd_rden),
    .clka(CSI_PCLK_pad),
    .clkb(clk_lcd),
    .csa({\and_Ncamera_addr[12]_o_al_n260 ,camera_addr[11:10]}),
    .csb({\and_Nlcd_rdaddr[12]__o_al_n263 ,lcd_rdaddr[11:10]}),
    .dia(camera_wrdat[8:0]),
    .rsta(CSI_RST_pad),
    .rstb(CSI_RST_pad),
    .dob({\uimg/inst_dob_i48_008 ,\uimg/inst_dob_i48_007 ,\uimg/inst_dob_i48_006 ,\uimg/inst_dob_i48_005 ,\uimg/inst_dob_i48_004 ,\uimg/inst_dob_i48_003 ,\uimg/inst_dob_i48_002 ,\uimg/inst_dob_i48_001 ,\uimg/inst_dob_i48_000 }));
  // address_offset=24576;data_offset=9;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("SIG"),
    .CSB1("SIG"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \uimg/inst_32800x16_sub_024576_009  (
    .addra(camera_addr[12:0]),
    .addrb(lcd_rdaddr[12:0]),
    .cea(camera_wrreq),
    .ceb(lcd_rden),
    .clka(CSI_PCLK_pad),
    .clkb(clk_lcd),
    .csa(camera_addr[15:13]),
    .csb(lcd_rdaddr[15:13]),
    .dia({open_n2396,open_n2397,open_n2398,open_n2399,open_n2400,open_n2401,open_n2402,camera_wrdat[9],open_n2403}),
    .rsta(CSI_RST_pad),
    .rstb(CSI_RST_pad),
    .dob({open_n2426,open_n2427,open_n2428,open_n2429,open_n2430,open_n2431,open_n2432,open_n2433,\uimg/inst_dob_i48_009 }));
  // address_offset=24576;data_offset=10;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("SIG"),
    .CSB1("SIG"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \uimg/inst_32800x16_sub_024576_010  (
    .addra(camera_addr[12:0]),
    .addrb(lcd_rdaddr[12:0]),
    .cea(camera_wrreq),
    .ceb(lcd_rden),
    .clka(CSI_PCLK_pad),
    .clkb(clk_lcd),
    .csa(camera_addr[15:13]),
    .csb(lcd_rdaddr[15:13]),
    .dia({open_n2434,open_n2435,open_n2436,open_n2437,open_n2438,open_n2439,open_n2440,camera_wrdat[10],open_n2441}),
    .rsta(CSI_RST_pad),
    .rstb(CSI_RST_pad),
    .dob({open_n2464,open_n2465,open_n2466,open_n2467,open_n2468,open_n2469,open_n2470,open_n2471,\uimg/inst_dob_i48_010 }));
  // address_offset=24576;data_offset=11;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("SIG"),
    .CSB1("SIG"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \uimg/inst_32800x16_sub_024576_011  (
    .addra(camera_addr[12:0]),
    .addrb(lcd_rdaddr[12:0]),
    .cea(camera_wrreq),
    .ceb(lcd_rden),
    .clka(CSI_PCLK_pad),
    .clkb(clk_lcd),
    .csa(camera_addr[15:13]),
    .csb(lcd_rdaddr[15:13]),
    .dia({open_n2472,open_n2473,open_n2474,open_n2475,open_n2476,open_n2477,open_n2478,camera_wrdat[11],open_n2479}),
    .rsta(CSI_RST_pad),
    .rstb(CSI_RST_pad),
    .dob({open_n2502,open_n2503,open_n2504,open_n2505,open_n2506,open_n2507,open_n2508,open_n2509,\uimg/inst_dob_i48_011 }));
  // address_offset=24576;data_offset=12;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("SIG"),
    .CSB1("SIG"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \uimg/inst_32800x16_sub_024576_012  (
    .addra(camera_addr[12:0]),
    .addrb(lcd_rdaddr[12:0]),
    .cea(camera_wrreq),
    .ceb(lcd_rden),
    .clka(CSI_PCLK_pad),
    .clkb(clk_lcd),
    .csa(camera_addr[15:13]),
    .csb(lcd_rdaddr[15:13]),
    .dia({open_n2510,open_n2511,open_n2512,open_n2513,open_n2514,open_n2515,open_n2516,camera_wrdat[12],open_n2517}),
    .rsta(CSI_RST_pad),
    .rstb(CSI_RST_pad),
    .dob({open_n2540,open_n2541,open_n2542,open_n2543,open_n2544,open_n2545,open_n2546,open_n2547,\uimg/inst_dob_i48_012 }));
  // address_offset=24576;data_offset=13;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("SIG"),
    .CSB1("SIG"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \uimg/inst_32800x16_sub_024576_013  (
    .addra(camera_addr[12:0]),
    .addrb(lcd_rdaddr[12:0]),
    .cea(camera_wrreq),
    .ceb(lcd_rden),
    .clka(CSI_PCLK_pad),
    .clkb(clk_lcd),
    .csa(camera_addr[15:13]),
    .csb(lcd_rdaddr[15:13]),
    .dia({open_n2548,open_n2549,open_n2550,open_n2551,open_n2552,open_n2553,open_n2554,camera_wrdat[13],open_n2555}),
    .rsta(CSI_RST_pad),
    .rstb(CSI_RST_pad),
    .dob({open_n2578,open_n2579,open_n2580,open_n2581,open_n2582,open_n2583,open_n2584,open_n2585,\uimg/inst_dob_i48_013 }));
  // address_offset=24576;data_offset=14;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("SIG"),
    .CSB1("SIG"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \uimg/inst_32800x16_sub_024576_014  (
    .addra(camera_addr[12:0]),
    .addrb(lcd_rdaddr[12:0]),
    .cea(camera_wrreq),
    .ceb(lcd_rden),
    .clka(CSI_PCLK_pad),
    .clkb(clk_lcd),
    .csa(camera_addr[15:13]),
    .csb(lcd_rdaddr[15:13]),
    .dia({open_n2586,open_n2587,open_n2588,open_n2589,open_n2590,open_n2591,open_n2592,camera_wrdat[14],open_n2593}),
    .rsta(CSI_RST_pad),
    .rstb(CSI_RST_pad),
    .dob({open_n2616,open_n2617,open_n2618,open_n2619,open_n2620,open_n2621,open_n2622,open_n2623,\uimg/inst_dob_i48_014 }));
  // address_offset=24576;data_offset=15;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("SIG"),
    .CSB1("SIG"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \uimg/inst_32800x16_sub_024576_015  (
    .addra(camera_addr[12:0]),
    .addrb(lcd_rdaddr[12:0]),
    .cea(camera_wrreq),
    .ceb(lcd_rden),
    .clka(CSI_PCLK_pad),
    .clkb(clk_lcd),
    .csa(camera_addr[15:13]),
    .csb(lcd_rdaddr[15:13]),
    .dia({open_n2624,open_n2625,open_n2626,open_n2627,open_n2628,open_n2629,open_n2630,camera_wrdat[15],open_n2631}),
    .rsta(CSI_RST_pad),
    .rstb(CSI_RST_pad),
    .dob({open_n2654,open_n2655,open_n2656,open_n2657,open_n2658,open_n2659,open_n2660,open_n2661,\uimg/inst_dob_i48_015 }));
  // address_offset=25600;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("SIG"),
    .CSB1("INV"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \uimg/inst_32800x16_sub_025600_000  (
    .addra({camera_addr[9:0],3'b111}),
    .addrb({lcd_rdaddr[9:0],3'b111}),
    .cea(camera_wrreq),
    .ceb(lcd_rden),
    .clka(CSI_PCLK_pad),
    .clkb(clk_lcd),
    .csa({\and_Ncamera_addr[12]_o_al_n260 ,camera_addr[11:10]}),
    .csb({\and_Nlcd_rdaddr[12]__o_al_n263 ,lcd_rdaddr[11:10]}),
    .dia(camera_wrdat[8:0]),
    .rsta(CSI_RST_pad),
    .rstb(CSI_RST_pad),
    .dob({\uimg/inst_dob_i50_008 ,\uimg/inst_dob_i50_007 ,\uimg/inst_dob_i50_006 ,\uimg/inst_dob_i50_005 ,\uimg/inst_dob_i50_004 ,\uimg/inst_dob_i50_003 ,\uimg/inst_dob_i50_002 ,\uimg/inst_dob_i50_001 ,\uimg/inst_dob_i50_000 }));
  // address_offset=26624;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("INV"),
    .CSB1("SIG"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \uimg/inst_32800x16_sub_026624_000  (
    .addra({camera_addr[9:0],3'b111}),
    .addrb({lcd_rdaddr[9:0],3'b111}),
    .cea(camera_wrreq),
    .ceb(lcd_rden),
    .clka(CSI_PCLK_pad),
    .clkb(clk_lcd),
    .csa({\and_Ncamera_addr[12]_o_al_n260 ,camera_addr[11:10]}),
    .csb({\and_Nlcd_rdaddr[12]__o_al_n263 ,lcd_rdaddr[11:10]}),
    .dia(camera_wrdat[8:0]),
    .rsta(CSI_RST_pad),
    .rstb(CSI_RST_pad),
    .dob({\uimg/inst_dob_i52_008 ,\uimg/inst_dob_i52_007 ,\uimg/inst_dob_i52_006 ,\uimg/inst_dob_i52_005 ,\uimg/inst_dob_i52_004 ,\uimg/inst_dob_i52_003 ,\uimg/inst_dob_i52_002 ,\uimg/inst_dob_i52_001 ,\uimg/inst_dob_i52_000 }));
  // address_offset=27648;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("SIG"),
    .CSB1("SIG"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \uimg/inst_32800x16_sub_027648_000  (
    .addra({camera_addr[9:0],3'b111}),
    .addrb({lcd_rdaddr[9:0],3'b111}),
    .cea(camera_wrreq),
    .ceb(lcd_rden),
    .clka(CSI_PCLK_pad),
    .clkb(clk_lcd),
    .csa({\and_Ncamera_addr[12]_o_al_n260 ,camera_addr[11:10]}),
    .csb({\and_Nlcd_rdaddr[12]__o_al_n263 ,lcd_rdaddr[11:10]}),
    .dia(camera_wrdat[8:0]),
    .rsta(CSI_RST_pad),
    .rstb(CSI_RST_pad),
    .dob({\uimg/inst_dob_i54_008 ,\uimg/inst_dob_i54_007 ,\uimg/inst_dob_i54_006 ,\uimg/inst_dob_i54_005 ,\uimg/inst_dob_i54_004 ,\uimg/inst_dob_i54_003 ,\uimg/inst_dob_i54_002 ,\uimg/inst_dob_i54_001 ,\uimg/inst_dob_i54_000 }));
  // address_offset=28672;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("INV"),
    .CSB1("INV"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \uimg/inst_32800x16_sub_028672_000  (
    .addra({camera_addr[9:0],3'b111}),
    .addrb({lcd_rdaddr[9:0],3'b111}),
    .cea(camera_wrreq),
    .ceb(lcd_rden),
    .clka(CSI_PCLK_pad),
    .clkb(clk_lcd),
    .csa({\and_camera_addr[12]__o_al_n276 ,camera_addr[11:10]}),
    .csb({\and_lcd_rdaddr[12]_l_o_al_n279 ,lcd_rdaddr[11:10]}),
    .dia(camera_wrdat[8:0]),
    .rsta(CSI_RST_pad),
    .rstb(CSI_RST_pad),
    .dob({\uimg/inst_dob_i56_008 ,\uimg/inst_dob_i56_007 ,\uimg/inst_dob_i56_006 ,\uimg/inst_dob_i56_005 ,\uimg/inst_dob_i56_004 ,\uimg/inst_dob_i56_003 ,\uimg/inst_dob_i56_002 ,\uimg/inst_dob_i56_001 ,\uimg/inst_dob_i56_000 }));
  // address_offset=29696;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("SIG"),
    .CSB1("INV"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \uimg/inst_32800x16_sub_029696_000  (
    .addra({camera_addr[9:0],3'b111}),
    .addrb({lcd_rdaddr[9:0],3'b111}),
    .cea(camera_wrreq),
    .ceb(lcd_rden),
    .clka(CSI_PCLK_pad),
    .clkb(clk_lcd),
    .csa({\and_camera_addr[12]__o_al_n276 ,camera_addr[11:10]}),
    .csb({\and_lcd_rdaddr[12]_l_o_al_n279 ,lcd_rdaddr[11:10]}),
    .dia(camera_wrdat[8:0]),
    .rsta(CSI_RST_pad),
    .rstb(CSI_RST_pad),
    .dob({\uimg/inst_dob_i58_008 ,\uimg/inst_dob_i58_007 ,\uimg/inst_dob_i58_006 ,\uimg/inst_dob_i58_005 ,\uimg/inst_dob_i58_004 ,\uimg/inst_dob_i58_003 ,\uimg/inst_dob_i58_002 ,\uimg/inst_dob_i58_001 ,\uimg/inst_dob_i58_000 }));
  // address_offset=30720;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("INV"),
    .CSB1("SIG"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \uimg/inst_32800x16_sub_030720_000  (
    .addra({camera_addr[9:0],3'b111}),
    .addrb({lcd_rdaddr[9:0],3'b111}),
    .cea(camera_wrreq),
    .ceb(lcd_rden),
    .clka(CSI_PCLK_pad),
    .clkb(clk_lcd),
    .csa({\and_camera_addr[12]__o_al_n276 ,camera_addr[11:10]}),
    .csb({\and_lcd_rdaddr[12]_l_o_al_n279 ,lcd_rdaddr[11:10]}),
    .dia(camera_wrdat[8:0]),
    .rsta(CSI_RST_pad),
    .rstb(CSI_RST_pad),
    .dob({\uimg/inst_dob_i60_008 ,\uimg/inst_dob_i60_007 ,\uimg/inst_dob_i60_006 ,\uimg/inst_dob_i60_005 ,\uimg/inst_dob_i60_004 ,\uimg/inst_dob_i60_003 ,\uimg/inst_dob_i60_002 ,\uimg/inst_dob_i60_001 ,\uimg/inst_dob_i60_000 }));
  // address_offset=31744;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("SIG"),
    .CSB1("SIG"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("1"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \uimg/inst_32800x16_sub_031744_000  (
    .addra({camera_addr[9:0],3'b111}),
    .addrb({lcd_rdaddr[9:0],3'b111}),
    .cea(camera_wrreq),
    .ceb(lcd_rden),
    .clka(CSI_PCLK_pad),
    .clkb(clk_lcd),
    .csa({\and_camera_addr[12]__o_al_n276 ,camera_addr[11:10]}),
    .csb({\and_lcd_rdaddr[12]_l_o_al_n279 ,lcd_rdaddr[11:10]}),
    .dia(camera_wrdat[8:0]),
    .rsta(CSI_RST_pad),
    .rstb(CSI_RST_pad),
    .dob({\uimg/inst_dob_i62_008 ,\uimg/inst_dob_i62_007 ,\uimg/inst_dob_i62_006 ,\uimg/inst_dob_i62_005 ,\uimg/inst_dob_i62_004 ,\uimg/inst_dob_i62_003 ,\uimg/inst_dob_i62_002 ,\uimg/inst_dob_i62_001 ,\uimg/inst_dob_i62_000 }));
  // address_offset=32768;data_offset=0;depth=32;width=16;num_section=1;width_per_section=16;section_size=16;working_depth=512;working_width=18;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("1"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("INV"),
    .CSB1("INV"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("18"),
    .DATA_WIDTH_B("18"),
    .MODE("PDPW8K"),
    .OCEAMUX("1"),
    .OCEBMUX("1"),
    .REGMODE_A("OUTREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("INV"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \uimg/inst_32800x16_sub_032768_000  (
    .addra({camera_addr[8:0],4'b1111}),
    .addrb({lcd_rdaddr[8:0],4'b1111}),
    .clka(CSI_PCLK_pad),
    .clkb(clk_lcd),
    .csa({\and_Ncamera_addr[11]_o_and_camera_wrreq ,camera_addr[10:9]}),
    .csb({\and_Nlcd_rdaddr[11]__o_and_lcd_rden ,lcd_rdaddr[10:9]}),
    .dia(camera_wrdat[8:0]),
    .dib({open_n2818,open_n2819,camera_wrdat[15:9]}),
    .rsta(CSI_RST_pad),
    .rstb(CSI_RST_pad),
    .doa({\uimg/inst_dob_i64_008 ,\uimg/inst_dob_i64_007 ,\uimg/inst_dob_i64_006 ,\uimg/inst_dob_i64_005 ,\uimg/inst_dob_i64_004 ,\uimg/inst_dob_i64_003 ,\uimg/inst_dob_i64_002 ,\uimg/inst_dob_i64_001 ,\uimg/inst_dob_i64_000 }),
    .dob({open_n2824,open_n2825,\uimg/inst_dob_i64_015 ,\uimg/inst_dob_i64_014 ,\uimg/inst_dob_i64_013 ,\uimg/inst_dob_i64_012 ,\uimg/inst_dob_i64_011 ,\uimg/inst_dob_i64_010 ,\uimg/inst_dob_i64_009 }));

endmodule 

module reg_sr_as_w1
  (
  clk,
  d,
  en,
  reset,
  set,
  q
  );

  input clk;
  input d;
  input en;
  input reset;
  input set;
  output q;

  parameter REGSET = "RESET";
  wire enout;
  wire resetout;

  AL_MUX u_en0 (
    .i0(q),
    .i1(d),
    .sel(en),
    .o(enout));
  AL_MUX u_reset0 (
    .i0(enout),
    .i1(1'b0),
    .sel(reset),
    .o(resetout));
  AL_DFF #(
    .INI((REGSET == "SET") ? 1'b1 : 1'b0))
    u_seq0 (
    .clk(clk),
    .d(resetout),
    .reset(1'b0),
    .set(set),
    .q(q));

endmodule 

module reg_ar_as_w1
  (
  clk,
  d,
  en,
  reset,
  set,
  q
  );

  input clk;
  input d;
  input en;
  input reset;
  input set;
  output q;

  parameter REGSET = "RESET";
  wire enout;

  AL_MUX u_en0 (
    .i0(q),
    .i1(d),
    .sel(en),
    .o(enout));
  AL_DFF #(
    .INI((REGSET == "SET") ? 1'b1 : 1'b0))
    u_seq0 (
    .clk(clk),
    .d(enout),
    .reset(reset),
    .set(set),
    .q(q));

endmodule 

module camera_init  // sources/rtl/camera_init.v(1)
  (
  clk,
  reset_n,
  sda_in,
  ready,
  scl,
  sda,
  sda_oe
  );

  input clk;  // sources/rtl/camera_init.v(3)
  input reset_n;  // sources/rtl/camera_init.v(4)
  input sda_in;  // sources/rtl/camera_init.v(10)
  output ready;  // sources/rtl/camera_init.v(6)
  output scl;  // sources/rtl/camera_init.v(11)
  output sda;  // sources/rtl/camera_init.v(9)
  output sda_oe;  // sources/rtl/camera_init.v(8)

  parameter REGS_TO_INIT = 178;
  // localparam CAMERA_IDLE = 18;
  // localparam CAMERA_INIT_1 = 11;
  // localparam CAMERA_INIT_2 = 12;
  // localparam CAMERA_INIT_3 = 13;
  // localparam CAMERA_INIT_4 = 14;
  // localparam CAMERA_INIT_5 = 15;
  // localparam CAMERA_INIT_6 = 16;
  // localparam CAMERA_INIT_7 = 17;
  // localparam CONTROL_REG = 3'b000;
  // localparam SLAVE_ADDRESS = 3'b001;
  // localparam SLAVE_DATA_1 = 3'b011;
  // localparam SLAVE_DATA_2 = 3'b100;
  // localparam SLAVE_REG_ADDRESS = 3'b010;
  wire [7:0] cnt;  // sources/rtl/camera_init.v(47)
  wire [7:0] counter;  // sources/rtl/camera_init.v(46)
  wire [7:0] data_in_bus;  // sources/rtl/camera_init.v(32)
  wire [8:0] divider2;  // sources/rtl/camera_init.v(52)
  wire [8:0] n0;
  wire [15:0] n186;
  wire [15:0] n187;
  wire [15:0] n189;
  wire [15:0] n190;
  wire [15:0] n193;
  wire [15:0] n197;
  wire [15:0] n198;
  wire [15:0] n200;
  wire [15:0] n202;
  wire [15:0] n203;
  wire [15:0] n205;
  wire [15:0] n206;
  wire [15:0] n208;
  wire [15:0] n210;
  wire [15:0] n213;
  wire [15:0] n214;
  wire [15:0] n215;
  wire [15:0] n216;
  wire [15:0] n217;
  wire [15:0] n221;
  wire [15:0] n225;
  wire [15:0] n227;
  wire [15:0] n246;
  wire [15:0] n247;
  wire [15:0] n258;
  wire [15:0] n275;
  wire [7:0] n369;
  wire [7:0] n372;
  wire [7:0] n373;
  wire [7:0] n375;
  wire [2:0] n385;
  wire [2:0] reg_address;  // sources/rtl/camera_init.v(33)
  wire  \sel0_b0/B4 ;
  wire  \sel0_b3/B3 ;
  wire [7:0] state_next;  // sources/rtl/camera_init.v(50)
  wire _al_u2838_o;
  wire _al_u2839_o;
  wire _al_u2842_o;
  wire _al_u2843_o;
  wire _al_u2844_o;
  wire _al_u2853_o;
  wire _al_u2854_o;
  wire _al_u2858_o;
  wire _al_u2860_o;
  wire _al_u2863_o;
  wire _al_u2865_o;
  wire _al_u2867_o;
  wire _al_u2869_o;
  wire _al_u2871_o;
  wire _al_u2872_o;
  wire _al_u2873_o;
  wire _al_u2874_o;
  wire _al_u2875_o;
  wire _al_u2877_o;
  wire _al_u2879_o;
  wire _al_u2882_o;
  wire _al_u2884_o;
  wire _al_u2885_o;
  wire _al_u2886_o;
  wire _al_u2887_o;
  wire _al_u2888_o;
  wire _al_u2889_o;
  wire _al_u2890_o;
  wire _al_u2891_o;
  wire _al_u2892_o;
  wire _al_u2894_o;
  wire _al_u2895_o;
  wire _al_u2897_o;
  wire _al_u2898_o;
  wire _al_u2899_o;
  wire _al_u2900_o;
  wire _al_u2902_o;
  wire _al_u2903_o;
  wire _al_u2904_o;
  wire _al_u2905_o;
  wire _al_u2906_o;
  wire _al_u2907_o;
  wire _al_u2908_o;
  wire _al_u2909_o;
  wire _al_u2911_o;
  wire _al_u2912_o;
  wire _al_u2913_o;
  wire _al_u2914_o;
  wire _al_u2915_o;
  wire _al_u2916_o;
  wire _al_u2917_o;
  wire _al_u2918_o;
  wire _al_u2919_o;
  wire _al_u2920_o;
  wire _al_u2921_o;
  wire _al_u2922_o;
  wire _al_u2923_o;
  wire _al_u2924_o;
  wire _al_u2925_o;
  wire _al_u2926_o;
  wire _al_u2927_o;
  wire _al_u2928_o;
  wire _al_u2929_o;
  wire _al_u2930_o;
  wire _al_u2932_o;
  wire _al_u2933_o;
  wire _al_u2935_o;
  wire _al_u2936_o;
  wire _al_u2937_o;
  wire _al_u2938_o;
  wire _al_u2939_o;
  wire _al_u2940_o;
  wire _al_u2941_o;
  wire _al_u2943_o;
  wire _al_u2945_o;
  wire _al_u2946_o;
  wire _al_u2947_o;
  wire _al_u2949_o;
  wire _al_u2950_o;
  wire _al_u2951_o;
  wire _al_u2952_o;
  wire _al_u2953_o;
  wire _al_u2955_o;
  wire _al_u2956_o;
  wire _al_u2958_o;
  wire _al_u2959_o;
  wire _al_u2963_o;
  wire _al_u2964_o;
  wire _al_u2965_o;
  wire _al_u2966_o;
  wire _al_u2968_o;
  wire _al_u2969_o;
  wire _al_u2970_o;
  wire _al_u2972_o;
  wire _al_u2974_o;
  wire _al_u2975_o;
  wire _al_u2976_o;
  wire _al_u2977_o;
  wire _al_u2979_o;
  wire _al_u2980_o;
  wire _al_u2982_o;
  wire _al_u2984_o;
  wire _al_u2985_o;
  wire _al_u2986_o;
  wire _al_u2987_o;
  wire _al_u2989_o;
  wire _al_u2990_o;
  wire _al_u2991_o;
  wire _al_u2993_o;
  wire _al_u2994_o;
  wire _al_u2995_o;
  wire _al_u2996_o;
  wire _al_u2997_o;
  wire _al_u2998_o;
  wire _al_u2999_o;
  wire _al_u3000_o;
  wire _al_u3001_o;
  wire _al_u3002_o;
  wire _al_u3003_o;
  wire _al_u3004_o;
  wire _al_u3005_o;
  wire _al_u3006_o;
  wire _al_u3007_o;
  wire _al_u3008_o;
  wire _al_u3010_o;
  wire _al_u3011_o;
  wire _al_u3012_o;
  wire _al_u3013_o;
  wire _al_u3014_o;
  wire _al_u3015_o;
  wire _al_u3016_o;
  wire _al_u3017_o;
  wire _al_u3019_o;
  wire _al_u3020_o;
  wire _al_u3021_o;
  wire _al_u3022_o;
  wire _al_u3023_o;
  wire _al_u3024_o;
  wire _al_u3025_o;
  wire _al_u3026_o;
  wire _al_u3027_o;
  wire _al_u3028_o;
  wire _al_u3030_o;
  wire _al_u3031_o;
  wire _al_u3032_o;
  wire _al_u3033_o;
  wire _al_u3034_o;
  wire _al_u3035_o;
  wire _al_u3036_o;
  wire _al_u3037_o;
  wire _al_u3038_o;
  wire _al_u3039_o;
  wire _al_u3040_o;
  wire _al_u3041_o;
  wire _al_u3042_o;
  wire _al_u3043_o;
  wire _al_u3044_o;
  wire _al_u3045_o;
  wire _al_u3046_o;
  wire _al_u3047_o;
  wire _al_u3048_o;
  wire _al_u3049_o;
  wire _al_u3050_o;
  wire _al_u3052_o;
  wire _al_u3054_o;
  wire _al_u3055_o;
  wire _al_u3056_o;
  wire _al_u3057_o;
  wire _al_u3058_o;
  wire _al_u3059_o;
  wire _al_u3061_o;
  wire _al_u3064_o;
  wire _al_u3065_o;
  wire _al_u3066_o;
  wire _al_u3067_o;
  wire _al_u3068_o;
  wire _al_u3069_o;
  wire _al_u3070_o;
  wire _al_u3071_o;
  wire _al_u3072_o;
  wire _al_u3073_o;
  wire _al_u3074_o;
  wire _al_u3075_o;
  wire _al_u3076_o;
  wire _al_u3077_o;
  wire _al_u3078_o;
  wire _al_u3079_o;
  wire _al_u3080_o;
  wire _al_u3081_o;
  wire _al_u3083_o;
  wire _al_u3084_o;
  wire _al_u3085_o;
  wire _al_u3086_o;
  wire _al_u3087_o;
  wire _al_u3088_o;
  wire _al_u3089_o;
  wire _al_u3090_o;
  wire _al_u3091_o;
  wire _al_u3092_o;
  wire _al_u3093_o;
  wire _al_u3094_o;
  wire _al_u3095_o;
  wire _al_u3096_o;
  wire _al_u3097_o;
  wire _al_u3098_o;
  wire _al_u3099_o;
  wire _al_u3101_o;
  wire _al_u3102_o;
  wire _al_u3103_o;
  wire _al_u3104_o;
  wire _al_u3105_o;
  wire _al_u3106_o;
  wire _al_u3107_o;
  wire _al_u3108_o;
  wire _al_u3109_o;
  wire _al_u3110_o;
  wire _al_u3111_o;
  wire _al_u3112_o;
  wire _al_u3113_o;
  wire _al_u3114_o;
  wire _al_u3115_o;
  wire _al_u3117_o;
  wire _al_u3118_o;
  wire _al_u3120_o;
  wire _al_u3121_o;
  wire _al_u3122_o;
  wire _al_u3124_o;
  wire _al_u3129_o;
  wire _al_u3132_o;
  wire _al_u3134_o;
  wire _al_u3135_o;
  wire _al_u3136_o;
  wire _al_u3137_o;
  wire _al_u3138_o;
  wire _al_u3139_o;
  wire _al_u3141_o;
  wire _al_u3142_o;
  wire _al_u3143_o;
  wire _al_u3144_o;
  wire _al_u3145_o;
  wire _al_u3146_o;
  wire _al_u3147_o;
  wire _al_u3148_o;
  wire _al_u3150_o;
  wire _al_u3151_o;
  wire _al_u3152_o;
  wire _al_u3153_o;
  wire _al_u3155_o;
  wire _al_u3156_o;
  wire _al_u3158_o;
  wire _al_u3160_o;
  wire _al_u3162_o;
  wire _al_u3163_o;
  wire _al_u3164_o;
  wire _al_u3165_o;
  wire _al_u3167_o;
  wire _al_u3168_o;
  wire _al_u3169_o;
  wire _al_u3171_o;
  wire _al_u3174_o;
  wire _al_u3176_o;
  wire _al_u3177_o;
  wire _al_u3180_o;
  wire _al_u3181_o;
  wire _al_u3182_o;
  wire _al_u3183_o;
  wire _al_u3184_o;
  wire _al_u3185_o;
  wire _al_u3186_o;
  wire _al_u3187_o;
  wire _al_u3188_o;
  wire _al_u3189_o;
  wire _al_u3191_o;
  wire _al_u3193_o;
  wire _al_u3194_o;
  wire _al_u3195_o;
  wire _al_u3196_o;
  wire _al_u3197_o;
  wire _al_u3198_o;
  wire _al_u3199_o;
  wire _al_u3200_o;
  wire _al_u3201_o;
  wire _al_u3202_o;
  wire _al_u3203_o;
  wire _al_u3204_o;
  wire _al_u3205_o;
  wire _al_u3206_o;
  wire _al_u3207_o;
  wire _al_u3208_o;
  wire _al_u3209_o;
  wire _al_u3210_o;
  wire _al_u3211_o;
  wire _al_u3213_o;
  wire _al_u3214_o;
  wire _al_u3215_o;
  wire _al_u3216_o;
  wire _al_u3217_o;
  wire _al_u3218_o;
  wire _al_u3219_o;
  wire _al_u3220_o;
  wire _al_u3221_o;
  wire _al_u3222_o;
  wire _al_u3223_o;
  wire _al_u3224_o;
  wire _al_u3225_o;
  wire _al_u3226_o;
  wire _al_u3227_o;
  wire _al_u3228_o;
  wire _al_u3229_o;
  wire _al_u3230_o;
  wire _al_u3231_o;
  wire _al_u3232_o;
  wire _al_u3233_o;
  wire _al_u3234_o;
  wire _al_u3235_o;
  wire _al_u3236_o;
  wire _al_u3237_o;
  wire _al_u3239_o;
  wire _al_u3240_o;
  wire _al_u3241_o;
  wire _al_u3244_o;
  wire _al_u3245_o;
  wire _al_u3249_o;
  wire _al_u3250_o;
  wire _al_u3252_o;
  wire _al_u3253_o;
  wire _al_u3256_o;
  wire _al_u3257_o;
  wire _al_u3258_o;
  wire _al_u3262_o;
  wire _al_u3263_o;
  wire _al_u3264_o;
  wire _al_u3265_o;
  wire _al_u3266_o;
  wire _al_u3267_o;
  wire _al_u3268_o;
  wire _al_u3269_o;
  wire _al_u3270_o;
  wire _al_u3271_o;
  wire _al_u3272_o;
  wire _al_u3273_o;
  wire _al_u3274_o;
  wire _al_u3275_o;
  wire _al_u3276_o;
  wire _al_u3277_o;
  wire _al_u3278_o;
  wire _al_u3279_o;
  wire _al_u3280_o;
  wire _al_u3281_o;
  wire _al_u3282_o;
  wire _al_u3283_o;
  wire _al_u3284_o;
  wire _al_u3286_o;
  wire _al_u3287_o;
  wire _al_u3289_o;
  wire _al_u3290_o;
  wire _al_u3291_o;
  wire _al_u3292_o;
  wire _al_u3293_o;
  wire _al_u3294_o;
  wire _al_u3295_o;
  wire _al_u3296_o;
  wire _al_u3297_o;
  wire _al_u3298_o;
  wire _al_u3299_o;
  wire _al_u3300_o;
  wire _al_u3301_o;
  wire _al_u3302_o;
  wire _al_u3304_o;
  wire _al_u3308_o;
  wire _al_u3311_o;
  wire _al_u3314_o;
  wire _al_u3315_o;
  wire _al_u3316_o;
  wire _al_u3317_o;
  wire _al_u3318_o;
  wire _al_u3319_o;
  wire _al_u3320_o;
  wire _al_u3321_o;
  wire _al_u3322_o;
  wire _al_u3323_o;
  wire _al_u3325_o;
  wire _al_u3326_o;
  wire _al_u3327_o;
  wire _al_u3330_o;
  wire _al_u3331_o;
  wire _al_u3332_o;
  wire _al_u3333_o;
  wire _al_u3334_o;
  wire _al_u3335_o;
  wire _al_u3336_o;
  wire _al_u3337_o;
  wire _al_u3338_o;
  wire _al_u3339_o;
  wire _al_u3340_o;
  wire _al_u3341_o;
  wire _al_u3342_o;
  wire _al_u3343_o;
  wire _al_u3344_o;
  wire _al_u3345_o;
  wire _al_u3348_o;
  wire _al_u3349_o;
  wire _al_u3352_o;
  wire _al_u3353_o;
  wire _al_u3354_o;
  wire _al_u3355_o;
  wire _al_u3357_o;
  wire _al_u3359_o;
  wire _al_u3360_o;
  wire _al_u3361_o;
  wire _al_u3362_o;
  wire _al_u3363_o;
  wire _al_u3364_o;
  wire _al_u3365_o;
  wire _al_u3366_o;
  wire _al_u3367_o;
  wire _al_u3368_o;
  wire _al_u3369_o;
  wire _al_u3370_o;
  wire _al_u3371_o;
  wire _al_u3372_o;
  wire _al_u3373_o;
  wire _al_u3374_o;
  wire _al_u3375_o;
  wire _al_u3376_o;
  wire _al_u3377_o;
  wire _al_u3378_o;
  wire _al_u3379_o;
  wire _al_u3380_o;
  wire _al_u3381_o;
  wire _al_u3382_o;
  wire _al_u3383_o;
  wire _al_u3384_o;
  wire _al_u3385_o;
  wire _al_u3386_o;
  wire _al_u3387_o;
  wire _al_u3388_o;
  wire _al_u3391_o;
  wire _al_u3393_o;
  wire _al_u3396_o;
  wire _al_u3397_o;
  wire _al_u3398_o;
  wire _al_u3400_o;
  wire _al_u3401_o;
  wire _al_u3402_o;
  wire _al_u3403_o;
  wire _al_u3406_o;
  wire _al_u3407_o;
  wire _al_u3408_o;
  wire _al_u3409_o;
  wire _al_u3410_o;
  wire _al_u3411_o;
  wire _al_u3412_o;
  wire _al_u3413_o;
  wire _al_u3414_o;
  wire _al_u3415_o;
  wire _al_u3416_o;
  wire _al_u3417_o;
  wire _al_u3418_o;
  wire _al_u3419_o;
  wire _al_u3420_o;
  wire _al_u3421_o;
  wire _al_u3422_o;
  wire _al_u3423_o;
  wire _al_u3425_o;
  wire _al_u3426_o;
  wire _al_u3427_o;
  wire _al_u3428_o;
  wire _al_u3429_o;
  wire _al_u3430_o;
  wire _al_u3431_o;
  wire _al_u3432_o;
  wire _al_u3433_o;
  wire _al_u3434_o;
  wire _al_u3435_o;
  wire _al_u3436_o;
  wire _al_u3437_o;
  wire _al_u3438_o;
  wire _al_u3439_o;
  wire _al_u3440_o;
  wire _al_u3441_o;
  wire _al_u3442_o;
  wire _al_u3443_o;
  wire _al_u3444_o;
  wire _al_u3445_o;
  wire _al_u3449_o;
  wire _al_u3453_o;
  wire _al_u3454_o;
  wire _al_u3455_o;
  wire _al_u3456_o;
  wire _al_u3457_o;
  wire _al_u3458_o;
  wire _al_u3459_o;
  wire _al_u3460_o;
  wire _al_u3462_o;
  wire _al_u3463_o;
  wire _al_u3464_o;
  wire _al_u3465_o;
  wire _al_u3467_o;
  wire _al_u3468_o;
  wire _al_u3471_o;
  wire _al_u3473_o;
  wire _al_u3474_o;
  wire _al_u3475_o;
  wire _al_u3476_o;
  wire _al_u3477_o;
  wire _al_u3478_o;
  wire _al_u3479_o;
  wire _al_u3480_o;
  wire _al_u3481_o;
  wire _al_u3482_o;
  wire _al_u3483_o;
  wire _al_u3484_o;
  wire _al_u3485_o;
  wire _al_u3486_o;
  wire _al_u3487_o;
  wire _al_u3488_o;
  wire _al_u3489_o;
  wire _al_u3490_o;
  wire _al_u3491_o;
  wire _al_u3492_o;
  wire _al_u3493_o;
  wire _al_u3494_o;
  wire _al_u3495_o;
  wire _al_u3496_o;
  wire _al_u3497_o;
  wire _al_u3499_o;
  wire _al_u3500_o;
  wire _al_u3501_o;
  wire _al_u3502_o;
  wire _al_u3503_o;
  wire _al_u3504_o;
  wire _al_u3505_o;
  wire _al_u3507_o;
  wire _al_u3508_o;
  wire _al_u3509_o;
  wire _al_u3510_o;
  wire _al_u3511_o;
  wire _al_u3512_o;
  wire _al_u3513_o;
  wire _al_u3514_o;
  wire _al_u3515_o;
  wire _al_u3516_o;
  wire _al_u3517_o;
  wire _al_u3518_o;
  wire _al_u3519_o;
  wire _al_u3520_o;
  wire _al_u3521_o;
  wire _al_u3522_o;
  wire _al_u3523_o;
  wire _al_u3524_o;
  wire _al_u3525_o;
  wire _al_u3530_o;
  wire _al_u3532_o;
  wire _al_u3533_o;
  wire _al_u3534_o;
  wire _al_u3535_o;
  wire _al_u3536_o;
  wire _al_u3537_o;
  wire _al_u3538_o;
  wire _al_u3539_o;
  wire _al_u3540_o;
  wire _al_u3541_o;
  wire _al_u3542_o;
  wire _al_u3545_o;
  wire _al_u3546_o;
  wire _al_u3547_o;
  wire _al_u3548_o;
  wire _al_u3549_o;
  wire _al_u3550_o;
  wire _al_u3551_o;
  wire _al_u3552_o;
  wire _al_u3553_o;
  wire _al_u3554_o;
  wire _al_u3555_o;
  wire _al_u3556_o;
  wire _al_u3557_o;
  wire _al_u3558_o;
  wire _al_u3559_o;
  wire _al_u3560_o;
  wire _al_u3562_o;
  wire _al_u3563_o;
  wire _al_u3564_o;
  wire _al_u3565_o;
  wire _al_u3566_o;
  wire _al_u3570_o;
  wire _al_u3574_o;
  wire _al_u3575_o;
  wire _al_u3576_o;
  wire _al_u3577_o;
  wire _al_u3578_o;
  wire _al_u3579_o;
  wire _al_u3580_o;
  wire _al_u3581_o;
  wire _al_u3582_o;
  wire _al_u3583_o;
  wire _al_u3584_o;
  wire _al_u3585_o;
  wire _al_u3586_o;
  wire _al_u3588_o;
  wire _al_u3589_o;
  wire _al_u3590_o;
  wire _al_u3591_o;
  wire _al_u3592_o;
  wire _al_u3593_o;
  wire _al_u3594_o;
  wire _al_u3595_o;
  wire _al_u3596_o;
  wire _al_u3598_o;
  wire _al_u3599_o;
  wire _al_u3600_o;
  wire _al_u3601_o;
  wire _al_u3602_o;
  wire _al_u3603_o;
  wire _al_u3604_o;
  wire _al_u3606_o;
  wire _al_u3607_o;
  wire _al_u3608_o;
  wire _al_u3609_o;
  wire _al_u3610_o;
  wire _al_u3611_o;
  wire _al_u3612_o;
  wire _al_u3613_o;
  wire _al_u3614_o;
  wire _al_u3615_o;
  wire _al_u3616_o;
  wire _al_u3617_o;
  wire _al_u3618_o;
  wire _al_u3619_o;
  wire _al_u3620_o;
  wire _al_u3621_o;
  wire \add0/c0 ;
  wire \add0/c1 ;
  wire \add0/c2 ;
  wire \add0/c3 ;
  wire \add0/c4 ;
  wire \add0/c5 ;
  wire \add0/c6 ;
  wire \add0/c7 ;
  wire \add0/c8 ;
  wire \add1/c0 ;
  wire \add1/c1 ;
  wire \add1/c2 ;
  wire \add1/c3 ;
  wire \add1/c4 ;
  wire \add1/c5 ;
  wire \add1/c6 ;
  wire \add1/c7 ;
  wire \add2/c0 ;
  wire \add2/c1 ;
  wire \add2/c2 ;
  wire \add2/c3 ;
  wire \add2/c4 ;
  wire \add2/c5 ;
  wire \add2/c6 ;
  wire \add2/c7 ;
  wire bus_write;  // sources/rtl/camera_init.v(34)
  wire mux103_b1_sel_is_2_o;
  wire mux104_b11_sel_is_2_o;
  wire mux107_b0_sel_is_2_o;
  wire mux111_b0_sel_is_2_o;
  wire mux115_b2_sel_is_2_o;
  wire mux117_b5_sel_is_2_o;
  wire mux119_b3_sel_is_0_o;
  wire mux120_b3_sel_is_2_o;
  wire mux120_b7_sel_is_2_o;
  wire mux121_b7_sel_is_2_o;
  wire mux124_b0_sel_is_0_o;
  wire mux124_b11_sel_is_2_o;
  wire mux127_b5_sel_is_2_o;
  wire mux129_b0_sel_is_2_o;
  wire mux129_b8_sel_is_2_o;
  wire mux12_b9_sel_is_2_o_neg_lutinv;
  wire mux130_b1_sel_is_2_o;
  wire mux132_b0_sel_is_0_o;
  wire mux132_b3_sel_is_2_o;
  wire mux134_b0_sel_is_2_o;
  wire mux135_b11_sel_is_0_o;
  wire mux136_b0_sel_is_2_o;
  wire mux136_b1_sel_is_0_o;
  wire mux136_b7_sel_is_2_o;
  wire mux137_b2_sel_is_2_o;
  wire mux137_b5_sel_is_2_o;
  wire mux139_b0_sel_is_2_o;
  wire mux13_b2_sel_is_2_o;
  wire mux140_b11_sel_is_2_o;
  wire mux141_b1_sel_is_2_o;
  wire mux146_b12_sel_is_2_o;
  wire mux147_b12_sel_is_2_o;
  wire mux147_b3_sel_is_2_o;
  wire mux14_b0_sel_is_2_o;
  wire mux14_b11_sel_is_2_o;
  wire mux150_b0_sel_is_2_o;
  wire mux152_b0_sel_is_2_o;
  wire mux159_b3_sel_is_2_o;
  wire mux168_b4_sel_is_2_o;
  wire mux169_b0_sel_is_2_o;
  wire mux16_b11_sel_is_2_o;
  wire mux16_b1_sel_is_0_o;
  wire mux170_b10_sel_is_0_o;
  wire mux170_b2_sel_is_2_o;
  wire mux174_b0_sel_is_0_o;
  wire mux182_b0_sel_is_2_o;
  wire mux182_b1_sel_is_2_o;
  wire mux185_b0_sel_is_2_o;
  wire mux18_b6_sel_is_2_o;
  wire mux19_b2_sel_is_0_o;
  wire mux22_b11_sel_is_2_o;
  wire mux30_b12_sel_is_2_o;
  wire mux30_b1_sel_is_2_o;
  wire mux33_b0_sel_is_2_o;
  wire mux38_b12_sel_is_2_o;
  wire mux38_b1_sel_is_2_o;
  wire mux47_b0_sel_is_2_o;
  wire mux47_b1_sel_is_2_o;
  wire mux48_b1_sel_is_2_o;
  wire mux49_b0_sel_is_2_o;
  wire mux52_b1_sel_is_2_o;
  wire mux57_b3_sel_is_2_o;
  wire mux5_b5_sel_is_2_o;
  wire mux60_b10_sel_is_2_o;
  wire mux60_b1_sel_is_2_o;
  wire mux61_b0_sel_is_2_o;
  wire mux61_b3_sel_is_2_o;
  wire mux63_b12_sel_is_2_o;
  wire mux63_b1_sel_is_2_o;
  wire mux67_b0_sel_is_2_o;
  wire mux68_b1_sel_is_2_o;
  wire mux70_b2_sel_is_0_o;
  wire mux75_b5_sel_is_2_o;
  wire mux75_b6_sel_is_2_o;
  wire mux77_b8_sel_is_2_o;
  wire mux84_b4_sel_is_2_o;
  wire mux85_b0_sel_is_2_o;
  wire mux87_b0_sel_is_2_o;
  wire mux89_b1_sel_is_2_o;
  wire mux92_b0_sel_is_0_o;
  wire mux92_b7_sel_is_2_o;
  wire mux93_b3_sel_is_2_o;
  wire mux94_b0_sel_is_2_o;
  wire mux96_b0_sel_is_2_o;
  wire mux97_b15_sel_is_2_o;
  wire mux97_b5_sel_is_2_o;
  wire mux9_b12_sel_is_2_o;
  wire n366;
  wire n376_lutinv;
  wire n377_lutinv;
  wire n378_lutinv;
  wire n380_lutinv;
  wire n381;
  wire n383;
  wire ready_out;  // sources/rtl/camera_init.v(35)
  wire \sel2_b0/or_or_B4_B5_o_or_B6__o ;
  wire \sel2_b1/or_B6_or_B7_B8_o_o ;
  wire \sel2_b2/or_B6_or_B7_B8_o_o ;
  wire \sel2_b3/or_B6_or_B7_B8_o_o ;
  wire \sel2_b4/or_B6_or_B7_B8_o_o ;
  wire \sel2_b5/or_B6_or_B7_B8_o_o ;
  wire \sel2_b6/or_B6_or_B7_B8_o_o ;
  wire \sel2_b7/or_B6_or_B7_B8_o_o ;
  wire success_out;  // sources/rtl/camera_init.v(36)

  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u2838 (
    .a(state_next[2]),
    .b(n369[6]),
    .c(n369[7]),
    .o(_al_u2838_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*~B*A)"),
    .INIT(16'h0020))
    _al_u2839 (
    .a(_al_u2838_o),
    .b(state_next[3]),
    .c(state_next[4]),
    .d(n369[5]),
    .o(_al_u2839_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u2840 (
    .a(_al_u2839_o),
    .b(state_next[0]),
    .c(state_next[1]),
    .o(n381));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u2841 (
    .a(_al_u2839_o),
    .b(state_next[0]),
    .c(state_next[1]),
    .o(n383));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u2842 (
    .a(counter[1]),
    .b(counter[2]),
    .c(counter[3]),
    .o(_al_u2842_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*B*A)"),
    .INIT(16'h0800))
    _al_u2843 (
    .a(counter[4]),
    .b(counter[5]),
    .c(counter[6]),
    .d(counter[7]),
    .o(_al_u2843_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u2844 (
    .a(_al_u2842_o),
    .b(_al_u2843_o),
    .c(counter[0]),
    .o(_al_u2844_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2845 (
    .a(_al_u2844_o),
    .b(n373[7]),
    .o(n375[7]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2846 (
    .a(_al_u2844_o),
    .b(n373[6]),
    .o(n375[6]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2847 (
    .a(_al_u2844_o),
    .b(n373[5]),
    .o(n375[5]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2848 (
    .a(_al_u2844_o),
    .b(n373[4]),
    .o(n375[4]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2849 (
    .a(_al_u2844_o),
    .b(n373[3]),
    .o(n375[3]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2850 (
    .a(_al_u2844_o),
    .b(n373[2]),
    .o(n375[2]));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    _al_u2851 (
    .a(_al_u2844_o),
    .b(n373[1]),
    .o(n375[1]));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    _al_u2852 (
    .a(_al_u2844_o),
    .b(n373[0]),
    .o(n375[0]));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u2853 (
    .a(state_next[3]),
    .b(state_next[4]),
    .c(n369[5]),
    .o(_al_u2853_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    _al_u2854 (
    .a(_al_u2853_o),
    .b(state_next[2]),
    .c(n369[6]),
    .d(n369[7]),
    .o(_al_u2854_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u2855 (
    .a(_al_u2854_o),
    .b(reset_n),
    .c(state_next[1]),
    .o(mux182_b1_sel_is_2_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u2856 (
    .a(_al_u2854_o),
    .b(state_next[0]),
    .c(state_next[1]),
    .o(n378_lutinv));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u2857 (
    .a(_al_u2838_o),
    .b(_al_u2853_o),
    .c(state_next[0]),
    .d(state_next[1]),
    .o(n376_lutinv));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u2858 (
    .a(n378_lutinv),
    .b(n376_lutinv),
    .o(_al_u2858_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2859 (
    .a(_al_u2858_o),
    .b(reset_n),
    .o(mux182_b0_sel_is_2_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u2860 (
    .a(_al_u2854_o),
    .b(state_next[0]),
    .o(_al_u2860_o));
  AL_MAP_LUT2 #(
    .EQN("~(~B*A)"),
    .INIT(4'hd))
    _al_u2861 (
    .a(_al_u2858_o),
    .b(_al_u2860_o),
    .o(n366));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u2862 (
    .a(n381),
    .b(_al_u2844_o),
    .c(reset_n),
    .o(mux185_b0_sel_is_2_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u2863 (
    .a(_al_u2854_o),
    .b(n376_lutinv),
    .o(_al_u2863_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u2864 (
    .a(_al_u2854_o),
    .b(state_next[0]),
    .c(state_next[1]),
    .o(n380_lutinv));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u2865 (
    .a(_al_u2863_o),
    .b(n380_lutinv),
    .c(ready_out),
    .o(_al_u2865_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u2866 (
    .a(_al_u2860_o),
    .b(state_next[1]),
    .o(n377_lutinv));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u2867 (
    .a(_al_u2858_o),
    .b(n377_lutinv),
    .c(n381),
    .o(_al_u2867_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u2868 (
    .a(_al_u2839_o),
    .b(state_next[0]),
    .c(state_next[1]),
    .o(\sel0_b0/B4 ));
  AL_MAP_LUT4 #(
    .EQN("~(A*~((~D*B))*~(C)+A*(~D*B)*~(C)+~(A)*(~D*B)*C+A*(~D*B)*C)"),
    .INIT(16'hf535))
    _al_u2869 (
    .a(\sel0_b0/B4 ),
    .b(n380_lutinv),
    .c(ready_out),
    .d(success_out),
    .o(_al_u2869_o));
  AL_MAP_LUT4 #(
    .EQN("~(C*B*~(D*~A))"),
    .INIT(16'h7f3f))
    _al_u2870 (
    .a(_al_u2865_o),
    .b(_al_u2867_o),
    .c(_al_u2869_o),
    .d(state_next[2]),
    .o(n369[2]));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u2871 (
    .a(n380_lutinv),
    .b(_al_u2844_o),
    .c(success_out),
    .o(_al_u2871_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u2872 (
    .a(cnt[4]),
    .b(cnt[5]),
    .c(cnt[6]),
    .d(cnt[7]),
    .o(_al_u2872_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*~B*~A)"),
    .INIT(16'h0010))
    _al_u2873 (
    .a(cnt[0]),
    .b(cnt[1]),
    .c(cnt[2]),
    .d(cnt[3]),
    .o(_al_u2873_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2874 (
    .a(_al_u2872_o),
    .b(_al_u2873_o),
    .o(_al_u2874_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u2875 (
    .a(_al_u2871_o),
    .b(_al_u2860_o),
    .c(_al_u2874_o),
    .o(_al_u2875_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C*~A))"),
    .INIT(8'h73))
    _al_u2876 (
    .a(_al_u2865_o),
    .b(_al_u2875_o),
    .c(state_next[0]),
    .o(n369[0]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~(~B*A))"),
    .INIT(16'hd000))
    _al_u2877 (
    .a(_al_u2844_o),
    .b(_al_u2874_o),
    .c(ready_out),
    .d(success_out),
    .o(_al_u2877_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u2878 (
    .a(n380_lutinv),
    .b(_al_u2877_o),
    .o(\sel0_b3/B3 ));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u2879 (
    .a(_al_u2863_o),
    .b(\sel0_b3/B3 ),
    .c(state_next[3]),
    .o(_al_u2879_o));
  AL_MAP_LUT4 #(
    .EQN("~(B*A*~(~D*C))"),
    .INIT(16'h77f7))
    _al_u2880 (
    .a(_al_u2867_o),
    .b(_al_u2879_o),
    .c(\sel0_b0/B4 ),
    .d(ready_out),
    .o(n369[3]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+~(A)*~(B)*C+A*~(B)*C+A*B*C)"),
    .INIT(8'hb2))
    _al_u2881 (
    .a(state_next[4]),
    .b(n369[3]),
    .c(state_next[3]),
    .o(n369[4]));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D)*~((~B*~A))+~C*D*~((~B*~A))+~(~C)*D*(~B*~A)+~C*D*(~B*~A))"),
    .INIT(16'h1f0e))
    _al_u2882 (
    .a(\sel0_b0/B4 ),
    .b(n380_lutinv),
    .c(ready_out),
    .d(n378_lutinv),
    .o(_al_u2882_o));
  AL_MAP_LUT4 #(
    .EQN("~(~C*~A*~(D*B))"),
    .INIT(16'hfefa))
    _al_u2883 (
    .a(_al_u2882_o),
    .b(_al_u2863_o),
    .c(_al_u2871_o),
    .d(state_next[1]),
    .o(n369[1]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u2884 (
    .a(counter[0]),
    .b(counter[1]),
    .c(counter[2]),
    .d(counter[3]),
    .o(_al_u2884_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*A)"),
    .INIT(16'h0002))
    _al_u2885 (
    .a(counter[4]),
    .b(counter[5]),
    .c(counter[6]),
    .d(counter[7]),
    .o(_al_u2885_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2886 (
    .a(counter[2]),
    .b(counter[3]),
    .o(_al_u2886_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u2887 (
    .a(_al_u2886_o),
    .b(counter[0]),
    .c(counter[1]),
    .o(_al_u2887_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*B*~A)"),
    .INIT(16'h0400))
    _al_u2888 (
    .a(counter[4]),
    .b(counter[5]),
    .c(counter[6]),
    .d(counter[7]),
    .o(_al_u2888_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2889 (
    .a(_al_u2887_o),
    .b(_al_u2888_o),
    .o(_al_u2889_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2890 (
    .a(_al_u2884_o),
    .b(_al_u2888_o),
    .o(_al_u2890_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*B*A)"),
    .INIT(16'h0800))
    _al_u2891 (
    .a(counter[0]),
    .b(counter[1]),
    .c(counter[2]),
    .d(counter[3]),
    .o(_al_u2891_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2892 (
    .a(_al_u2891_o),
    .b(_al_u2888_o),
    .o(_al_u2892_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u2893 (
    .a(_al_u2889_o),
    .b(_al_u2890_o),
    .c(_al_u2892_o),
    .o(mux5_b5_sel_is_2_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u2894 (
    .a(counter[0]),
    .b(counter[1]),
    .c(counter[2]),
    .d(counter[3]),
    .o(_al_u2894_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2895 (
    .a(_al_u2894_o),
    .b(_al_u2888_o),
    .o(_al_u2895_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u2896 (
    .a(_al_u2844_o),
    .b(_al_u2895_o),
    .o(n186[0]));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u2897 (
    .a(counter[0]),
    .b(counter[1]),
    .o(_al_u2897_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2898 (
    .a(_al_u2897_o),
    .b(_al_u2886_o),
    .o(_al_u2898_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u2899 (
    .a(counter[1]),
    .b(counter[2]),
    .c(counter[3]),
    .o(_al_u2899_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2900 (
    .a(_al_u2899_o),
    .b(_al_u2888_o),
    .o(_al_u2900_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u2901 (
    .a(_al_u2898_o),
    .b(_al_u2900_o),
    .c(_al_u2888_o),
    .o(mux9_b12_sel_is_2_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u2902 (
    .a(mux5_b5_sel_is_2_o),
    .b(n186[0]),
    .c(mux9_b12_sel_is_2_o),
    .o(_al_u2902_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u2903 (
    .a(counter[2]),
    .b(counter[3]),
    .o(_al_u2903_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u2904 (
    .a(_al_u2903_o),
    .b(counter[0]),
    .c(counter[1]),
    .o(_al_u2904_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u2905 (
    .a(counter[2]),
    .b(counter[3]),
    .o(_al_u2905_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*(D@C))"),
    .INIT(16'h0880))
    _al_u2906 (
    .a(_al_u2905_o),
    .b(_al_u2888_o),
    .c(counter[0]),
    .d(counter[1]),
    .o(_al_u2906_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    _al_u2907 (
    .a(counter[0]),
    .b(counter[1]),
    .c(counter[2]),
    .d(counter[3]),
    .o(_al_u2907_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*~A)"),
    .INIT(8'h04))
    _al_u2908 (
    .a(counter[1]),
    .b(counter[2]),
    .c(counter[3]),
    .o(_al_u2908_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(~A*~(~D*B)))"),
    .INIT(16'ha0e0))
    _al_u2909 (
    .a(_al_u2907_o),
    .b(_al_u2908_o),
    .c(_al_u2888_o),
    .d(counter[0]),
    .o(_al_u2909_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~B*~(D*A))"),
    .INIT(16'h0103))
    _al_u2910 (
    .a(_al_u2904_o),
    .b(_al_u2906_o),
    .c(_al_u2909_o),
    .d(_al_u2888_o),
    .o(mux13_b2_sel_is_2_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2911 (
    .a(_al_u2842_o),
    .b(_al_u2888_o),
    .o(_al_u2911_o));
  AL_MAP_LUT4 #(
    .EQN("(~(B*A)*~(D)*~(C)+~(B*A)*D*~(C)+~(~(B*A))*D*C+~(B*A)*D*C)"),
    .INIT(16'hf707))
    _al_u2912 (
    .a(_al_u2902_o),
    .b(mux13_b2_sel_is_2_o),
    .c(_al_u2911_o),
    .d(counter[0]),
    .o(_al_u2912_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2913 (
    .a(counter[2]),
    .b(counter[3]),
    .o(_al_u2913_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2914 (
    .a(_al_u2897_o),
    .b(_al_u2913_o),
    .o(_al_u2914_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*A)"),
    .INIT(16'h0200))
    _al_u2915 (
    .a(counter[4]),
    .b(counter[5]),
    .c(counter[6]),
    .d(counter[7]),
    .o(_al_u2915_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2916 (
    .a(_al_u2914_o),
    .b(_al_u2915_o),
    .o(_al_u2916_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(~B*~A))"),
    .INIT(8'he0))
    _al_u2917 (
    .a(_al_u2887_o),
    .b(_al_u2891_o),
    .c(_al_u2915_o),
    .o(_al_u2917_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u2918 (
    .a(_al_u2916_o),
    .b(_al_u2917_o),
    .o(_al_u2918_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    _al_u2919 (
    .a(_al_u2912_o),
    .b(_al_u2918_o),
    .c(_al_u2915_o),
    .o(_al_u2919_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2920 (
    .a(_al_u2904_o),
    .b(_al_u2915_o),
    .o(_al_u2920_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2921 (
    .a(_al_u2907_o),
    .b(_al_u2915_o),
    .o(_al_u2921_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u2922 (
    .a(_al_u2920_o),
    .b(_al_u2921_o),
    .o(_al_u2922_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2923 (
    .a(_al_u2905_o),
    .b(_al_u2915_o),
    .o(_al_u2923_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u2924 (
    .a(_al_u2919_o),
    .b(_al_u2922_o),
    .c(_al_u2923_o),
    .d(counter[1]),
    .o(_al_u2924_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*~A)"),
    .INIT(16'h4000))
    _al_u2925 (
    .a(counter[0]),
    .b(counter[1]),
    .c(counter[2]),
    .d(counter[3]),
    .o(_al_u2925_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*~A)"),
    .INIT(16'h0100))
    _al_u2926 (
    .a(counter[4]),
    .b(counter[5]),
    .c(counter[6]),
    .d(counter[7]),
    .o(_al_u2926_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2927 (
    .a(_al_u2925_o),
    .b(_al_u2926_o),
    .o(_al_u2927_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2928 (
    .a(_al_u2894_o),
    .b(_al_u2926_o),
    .o(_al_u2928_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u2929 (
    .a(_al_u2927_o),
    .b(_al_u2928_o),
    .o(_al_u2929_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2930 (
    .a(_al_u2842_o),
    .b(_al_u2915_o),
    .o(_al_u2930_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(A*~(D)*~(C)+A*D*~(C)+~(A)*D*C+A*D*C))"),
    .INIT(16'h04c4))
    _al_u2931 (
    .a(_al_u2924_o),
    .b(_al_u2929_o),
    .c(_al_u2930_o),
    .d(counter[0]),
    .o(n217[6]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(~B*~A))"),
    .INIT(8'he0))
    _al_u2932 (
    .a(_al_u2887_o),
    .b(_al_u2891_o),
    .c(_al_u2926_o),
    .o(_al_u2932_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2933 (
    .a(_al_u2914_o),
    .b(_al_u2926_o),
    .o(_al_u2933_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u2934 (
    .a(n217[6]),
    .b(_al_u2932_o),
    .c(_al_u2933_o),
    .o(n221[6]));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u2935 (
    .a(_al_u2898_o),
    .b(_al_u2899_o),
    .c(counter[0]),
    .o(_al_u2935_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2936 (
    .a(_al_u2908_o),
    .b(_al_u2899_o),
    .c(counter[0]),
    .o(_al_u2936_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u2937 (
    .a(_al_u2935_o),
    .b(_al_u2936_o),
    .o(_al_u2937_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u2938 (
    .a(_al_u2908_o),
    .b(counter[0]),
    .o(_al_u2938_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(~B*A))"),
    .INIT(8'hd0))
    _al_u2939 (
    .a(_al_u2937_o),
    .b(_al_u2938_o),
    .c(_al_u2926_o),
    .o(_al_u2939_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2940 (
    .a(_al_u2904_o),
    .b(_al_u2926_o),
    .o(_al_u2940_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2941 (
    .a(_al_u2842_o),
    .b(_al_u2926_o),
    .o(_al_u2941_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u2942 (
    .a(_al_u2940_o),
    .b(_al_u2941_o),
    .o(mux47_b1_sel_is_2_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2943 (
    .a(_al_u2907_o),
    .b(_al_u2926_o),
    .o(_al_u2943_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*~A)"),
    .INIT(8'h04))
    _al_u2944 (
    .a(_al_u2939_o),
    .b(mux47_b1_sel_is_2_o),
    .c(_al_u2943_o),
    .o(mux47_b0_sel_is_2_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*A)"),
    .INIT(16'h0080))
    _al_u2945 (
    .a(counter[4]),
    .b(counter[5]),
    .c(counter[6]),
    .d(counter[7]),
    .o(_al_u2945_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2946 (
    .a(_al_u2925_o),
    .b(_al_u2945_o),
    .o(_al_u2946_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2947 (
    .a(_al_u2894_o),
    .b(_al_u2945_o),
    .o(_al_u2947_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u2948 (
    .a(mux47_b0_sel_is_2_o),
    .b(_al_u2946_o),
    .c(_al_u2947_o),
    .o(mux49_b0_sel_is_2_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u2949 (
    .a(_al_u2886_o),
    .b(counter[0]),
    .c(counter[1]),
    .o(_al_u2949_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u2950 (
    .a(_al_u2949_o),
    .b(_al_u2887_o),
    .o(_al_u2950_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u2951 (
    .a(_al_u2898_o),
    .b(_al_u2899_o),
    .o(_al_u2951_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B*A))"),
    .INIT(8'h70))
    _al_u2952 (
    .a(_al_u2950_o),
    .b(_al_u2951_o),
    .c(_al_u2945_o),
    .o(_al_u2952_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u2953 (
    .a(_al_u2907_o),
    .b(_al_u2908_o),
    .o(_al_u2953_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u2954 (
    .a(_al_u2952_o),
    .b(_al_u2953_o),
    .c(_al_u2945_o),
    .o(mux60_b10_sel_is_2_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(~B*~A))"),
    .INIT(8'he0))
    _al_u2955 (
    .a(_al_u2914_o),
    .b(_al_u2884_o),
    .c(_al_u2945_o),
    .o(_al_u2955_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2956 (
    .a(_al_u2891_o),
    .b(_al_u2945_o),
    .o(_al_u2956_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u2957 (
    .a(_al_u2955_o),
    .b(_al_u2956_o),
    .o(mux52_b1_sel_is_2_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2958 (
    .a(_al_u2904_o),
    .b(_al_u2945_o),
    .o(_al_u2958_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2959 (
    .a(_al_u2842_o),
    .b(_al_u2945_o),
    .o(_al_u2959_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    _al_u2960 (
    .a(mux60_b10_sel_is_2_o),
    .b(mux52_b1_sel_is_2_o),
    .c(_al_u2958_o),
    .d(_al_u2959_o),
    .o(mux63_b1_sel_is_2_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2961 (
    .a(mux49_b0_sel_is_2_o),
    .b(mux63_b1_sel_is_2_o),
    .o(mux63_b12_sel_is_2_o));
  AL_MAP_LUT2 #(
    .EQN("~(B@A)"),
    .INIT(4'h9))
    _al_u2962 (
    .a(n221[6]),
    .b(mux63_b12_sel_is_2_o),
    .o(n246[6]));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*~A)"),
    .INIT(16'h0040))
    _al_u2963 (
    .a(counter[4]),
    .b(counter[5]),
    .c(counter[6]),
    .d(counter[7]),
    .o(_al_u2963_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2964 (
    .a(_al_u2899_o),
    .b(_al_u2963_o),
    .o(_al_u2964_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u2965 (
    .a(_al_u2964_o),
    .b(counter[0]),
    .o(_al_u2965_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2966 (
    .a(_al_u2908_o),
    .b(_al_u2963_o),
    .o(_al_u2966_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u2967 (
    .a(_al_u2965_o),
    .b(_al_u2966_o),
    .o(mux75_b5_sel_is_2_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2968 (
    .a(_al_u2898_o),
    .b(_al_u2963_o),
    .o(_al_u2968_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u2969 (
    .a(_al_u2899_o),
    .b(_al_u2963_o),
    .c(counter[0]),
    .o(_al_u2969_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u2970 (
    .a(_al_u2968_o),
    .b(_al_u2969_o),
    .o(_al_u2970_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2971 (
    .a(mux75_b5_sel_is_2_o),
    .b(_al_u2970_o),
    .o(mux75_b6_sel_is_2_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(~B*~A))"),
    .INIT(8'he0))
    _al_u2972 (
    .a(_al_u2884_o),
    .b(_al_u2925_o),
    .c(_al_u2963_o),
    .o(_al_u2972_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u2973 (
    .a(_al_u2914_o),
    .b(_al_u2972_o),
    .c(_al_u2963_o),
    .o(mux67_b0_sel_is_2_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u2974 (
    .a(n246[6]),
    .b(mux75_b6_sel_is_2_o),
    .c(mux67_b0_sel_is_2_o),
    .o(_al_u2974_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*~B*A)"),
    .INIT(16'h0020))
    _al_u2975 (
    .a(counter[4]),
    .b(counter[5]),
    .c(counter[6]),
    .d(counter[7]),
    .o(_al_u2975_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(~B*~A))"),
    .INIT(8'he0))
    _al_u2976 (
    .a(_al_u2914_o),
    .b(_al_u2884_o),
    .c(_al_u2975_o),
    .o(_al_u2976_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2977 (
    .a(_al_u2891_o),
    .b(_al_u2975_o),
    .o(_al_u2977_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u2978 (
    .a(_al_u2976_o),
    .b(_al_u2977_o),
    .o(mux84_b4_sel_is_2_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2979 (
    .a(_al_u2887_o),
    .b(_al_u2975_o),
    .o(_al_u2979_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2980 (
    .a(_al_u2925_o),
    .b(_al_u2975_o),
    .o(_al_u2980_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u2981 (
    .a(mux84_b4_sel_is_2_o),
    .b(_al_u2979_o),
    .c(_al_u2980_o),
    .o(mux85_b0_sel_is_2_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(~B*~A))"),
    .INIT(8'he0))
    _al_u2982 (
    .a(_al_u2898_o),
    .b(_al_u2949_o),
    .c(_al_u2975_o),
    .o(_al_u2982_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u2983 (
    .a(mux85_b0_sel_is_2_o),
    .b(_al_u2982_o),
    .o(mux87_b0_sel_is_2_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2984 (
    .a(_al_u2894_o),
    .b(_al_u2975_o),
    .o(_al_u2984_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u2985 (
    .a(_al_u2974_o),
    .b(mux87_b0_sel_is_2_o),
    .c(_al_u2984_o),
    .o(_al_u2985_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2986 (
    .a(_al_u2938_o),
    .b(_al_u2975_o),
    .o(_al_u2986_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2987 (
    .a(_al_u2907_o),
    .b(_al_u2975_o),
    .o(_al_u2987_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u2988 (
    .a(_al_u2986_o),
    .b(_al_u2987_o),
    .o(mux92_b0_sel_is_0_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2989 (
    .a(_al_u2908_o),
    .b(counter[0]),
    .o(_al_u2989_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2990 (
    .a(_al_u2989_o),
    .b(_al_u2975_o),
    .o(_al_u2990_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2991 (
    .a(_al_u2904_o),
    .b(_al_u2975_o),
    .o(_al_u2991_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u2992 (
    .a(mux92_b0_sel_is_0_o),
    .b(_al_u2990_o),
    .c(_al_u2991_o),
    .o(mux93_b3_sel_is_2_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*~B*~A)"),
    .INIT(16'h0010))
    _al_u2993 (
    .a(counter[4]),
    .b(counter[5]),
    .c(counter[6]),
    .d(counter[7]),
    .o(_al_u2993_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2994 (
    .a(_al_u2914_o),
    .b(_al_u2993_o),
    .o(_al_u2994_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2995 (
    .a(_al_u2884_o),
    .b(_al_u2993_o),
    .o(_al_u2995_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u2996 (
    .a(_al_u2994_o),
    .b(_al_u2995_o),
    .o(_al_u2996_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2997 (
    .a(_al_u2925_o),
    .b(_al_u2993_o),
    .o(_al_u2997_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2998 (
    .a(_al_u2894_o),
    .b(_al_u2993_o),
    .o(_al_u2998_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u2999 (
    .a(_al_u2842_o),
    .b(_al_u2975_o),
    .c(counter[0]),
    .o(_al_u2999_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u3000 (
    .a(_al_u2997_o),
    .b(_al_u2998_o),
    .c(_al_u2999_o),
    .o(_al_u3000_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3001 (
    .a(_al_u2842_o),
    .b(_al_u2975_o),
    .c(counter[0]),
    .o(_al_u3001_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*A)"),
    .INIT(16'h0080))
    _al_u3002 (
    .a(mux93_b3_sel_is_2_o),
    .b(_al_u2996_o),
    .c(_al_u3000_o),
    .d(_al_u3001_o),
    .o(_al_u3002_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u3003 (
    .a(_al_u2985_o),
    .b(_al_u3002_o),
    .c(_al_u2994_o),
    .o(_al_u3003_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3004 (
    .a(_al_u2936_o),
    .b(_al_u2993_o),
    .o(_al_u3004_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3005 (
    .a(_al_u2886_o),
    .b(_al_u2993_o),
    .o(_al_u3005_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u3006 (
    .a(_al_u3003_o),
    .b(_al_u3004_o),
    .c(_al_u3005_o),
    .o(_al_u3006_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3007 (
    .a(_al_u2904_o),
    .b(_al_u2993_o),
    .o(_al_u3007_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3008 (
    .a(_al_u2842_o),
    .b(_al_u2993_o),
    .o(_al_u3008_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3009 (
    .a(_al_u3007_o),
    .b(_al_u3008_o),
    .o(mux111_b0_sel_is_2_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    _al_u3010 (
    .a(counter[4]),
    .b(counter[5]),
    .c(counter[6]),
    .d(counter[7]),
    .o(_al_u3010_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3011 (
    .a(_al_u2894_o),
    .b(_al_u3010_o),
    .o(_al_u3011_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3012 (
    .a(mux111_b0_sel_is_2_o),
    .b(_al_u3011_o),
    .o(_al_u3012_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3013 (
    .a(_al_u2914_o),
    .b(_al_u3010_o),
    .o(_al_u3013_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3014 (
    .a(_al_u2884_o),
    .b(_al_u3010_o),
    .o(_al_u3014_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3015 (
    .a(_al_u2925_o),
    .b(_al_u3010_o),
    .o(_al_u3015_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3016 (
    .a(_al_u3014_o),
    .b(_al_u3015_o),
    .o(_al_u3016_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u3017 (
    .a(_al_u3013_o),
    .b(_al_u3016_o),
    .o(_al_u3017_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3018 (
    .a(_al_u3012_o),
    .b(_al_u3017_o),
    .o(mux115_b2_sel_is_2_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3019 (
    .a(_al_u3006_o),
    .b(mux115_b2_sel_is_2_o),
    .o(_al_u3019_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3020 (
    .a(_al_u3013_o),
    .b(_al_u3014_o),
    .o(_al_u3020_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*A))"),
    .INIT(8'hc4))
    _al_u3021 (
    .a(_al_u3019_o),
    .b(_al_u3020_o),
    .c(_al_u3010_o),
    .o(_al_u3021_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3022 (
    .a(_al_u2887_o),
    .b(_al_u3010_o),
    .o(_al_u3022_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3023 (
    .a(_al_u3021_o),
    .b(_al_u3022_o),
    .o(_al_u3023_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3024 (
    .a(_al_u2898_o),
    .b(_al_u3010_o),
    .o(_al_u3024_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3025 (
    .a(_al_u3023_o),
    .b(_al_u3024_o),
    .o(_al_u3025_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*~A)"),
    .INIT(16'h0004))
    _al_u3026 (
    .a(counter[4]),
    .b(counter[5]),
    .c(counter[6]),
    .d(counter[7]),
    .o(_al_u3026_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3027 (
    .a(_al_u2914_o),
    .b(_al_u3026_o),
    .o(_al_u3027_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3028 (
    .a(_al_u2891_o),
    .b(_al_u3026_o),
    .o(_al_u3028_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3029 (
    .a(_al_u3027_o),
    .b(_al_u3028_o),
    .o(mux132_b0_sel_is_0_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3030 (
    .a(_al_u2884_o),
    .b(_al_u3026_o),
    .o(_al_u3030_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3031 (
    .a(mux132_b0_sel_is_0_o),
    .b(_al_u3030_o),
    .o(_al_u3031_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3032 (
    .a(_al_u2936_o),
    .b(_al_u3010_o),
    .o(_al_u3032_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*A))"),
    .INIT(8'hc4))
    _al_u3033 (
    .a(_al_u3025_o),
    .b(_al_u3031_o),
    .c(_al_u3032_o),
    .o(_al_u3033_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3034 (
    .a(_al_u2938_o),
    .b(_al_u3026_o),
    .o(_al_u3034_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*(~C*~(D)*~(A)+~C*D*~(A)+~(~C)*D*A+~C*D*A))"),
    .INIT(16'h2301))
    _al_u3035 (
    .a(_al_u3033_o),
    .b(_al_u3034_o),
    .c(_al_u3028_o),
    .d(_al_u3026_o),
    .o(_al_u3035_o));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    _al_u3036 (
    .a(_al_u2884_o),
    .b(_al_u2885_o),
    .c(_al_u3035_o),
    .o(_al_u3036_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3037 (
    .a(_al_u2891_o),
    .b(_al_u2885_o),
    .o(_al_u3037_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3038 (
    .a(_al_u3036_o),
    .b(_al_u3037_o),
    .o(_al_u3038_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3039 (
    .a(_al_u2908_o),
    .b(_al_u2885_o),
    .o(_al_u3039_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3040 (
    .a(_al_u2899_o),
    .b(_al_u2885_o),
    .o(_al_u3040_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3041 (
    .a(_al_u3039_o),
    .b(_al_u3040_o),
    .o(_al_u3041_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3042 (
    .a(_al_u2898_o),
    .b(_al_u2885_o),
    .o(_al_u3042_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3043 (
    .a(_al_u3038_o),
    .b(_al_u3041_o),
    .c(_al_u3042_o),
    .o(_al_u3043_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u3044 (
    .a(_al_u3041_o),
    .b(counter[0]),
    .o(_al_u3044_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3045 (
    .a(_al_u3043_o),
    .b(_al_u3044_o),
    .o(_al_u3045_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u3046 (
    .a(counter[4]),
    .b(counter[5]),
    .c(counter[6]),
    .d(counter[7]),
    .o(_al_u3046_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3047 (
    .a(_al_u3046_o),
    .b(_al_u2925_o),
    .o(_al_u3047_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3048 (
    .a(_al_u3045_o),
    .b(_al_u3047_o),
    .o(_al_u3048_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(~B*~A))"),
    .INIT(8'he0))
    _al_u3049 (
    .a(_al_u2898_o),
    .b(_al_u2949_o),
    .c(_al_u3046_o),
    .o(_al_u3049_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3050 (
    .a(_al_u3046_o),
    .b(_al_u2899_o),
    .o(_al_u3050_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3051 (
    .a(_al_u3049_o),
    .b(_al_u3050_o),
    .o(mux169_b0_sel_is_2_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3052 (
    .a(_al_u2989_o),
    .b(_al_u3046_o),
    .o(_al_u3052_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3053 (
    .a(mux169_b0_sel_is_2_o),
    .b(_al_u3052_o),
    .o(mux170_b2_sel_is_2_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3054 (
    .a(_al_u2914_o),
    .b(_al_u3046_o),
    .o(_al_u3054_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3055 (
    .a(_al_u3048_o),
    .b(mux170_b2_sel_is_2_o),
    .c(_al_u3054_o),
    .o(_al_u3055_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3056 (
    .a(_al_u2989_o),
    .b(_al_u2888_o),
    .o(_al_u3056_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3057 (
    .a(_al_u2899_o),
    .b(_al_u2888_o),
    .o(_al_u3057_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3058 (
    .a(_al_u3056_o),
    .b(_al_u3057_o),
    .o(_al_u3058_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3059 (
    .a(_al_u2894_o),
    .b(_al_u2915_o),
    .o(_al_u3059_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u3060 (
    .a(_al_u3059_o),
    .b(_al_u2911_o),
    .c(counter[0]),
    .o(mux16_b1_sel_is_0_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3061 (
    .a(_al_u2842_o),
    .b(_al_u2888_o),
    .c(counter[0]),
    .o(_al_u3061_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~B*~(D*A))"),
    .INIT(16'h0103))
    _al_u3062 (
    .a(_al_u2904_o),
    .b(_al_u2909_o),
    .c(_al_u3061_o),
    .d(_al_u2888_o),
    .o(mux14_b11_sel_is_2_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3063 (
    .a(mux16_b1_sel_is_0_o),
    .b(mux14_b11_sel_is_2_o),
    .o(mux16_b11_sel_is_2_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3064 (
    .a(_al_u3058_o),
    .b(mux16_b11_sel_is_2_o),
    .o(_al_u3064_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3065 (
    .a(_al_u2842_o),
    .b(_al_u2843_o),
    .o(_al_u3065_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(~D*~C))"),
    .INIT(16'h8880))
    _al_u3066 (
    .a(_al_u2913_o),
    .b(_al_u2888_o),
    .c(counter[0]),
    .d(counter[1]),
    .o(_al_u3066_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~B*~(~D*A))"),
    .INIT(16'h0301))
    _al_u3067 (
    .a(_al_u3065_o),
    .b(_al_u2892_o),
    .c(_al_u3066_o),
    .d(counter[0]),
    .o(_al_u3067_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u3068 (
    .a(_al_u2886_o),
    .b(_al_u2888_o),
    .c(counter[0]),
    .d(counter[1]),
    .o(_al_u3068_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3069 (
    .a(_al_u3064_o),
    .b(_al_u3067_o),
    .c(_al_u3068_o),
    .o(_al_u3069_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3070 (
    .a(_al_u3069_o),
    .b(_al_u2918_o),
    .c(_al_u2928_o),
    .o(_al_u3070_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3071 (
    .a(_al_u2884_o),
    .b(_al_u2926_o),
    .o(_al_u3071_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3072 (
    .a(_al_u2933_o),
    .b(_al_u3071_o),
    .o(_al_u3072_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3073 (
    .a(_al_u3070_o),
    .b(_al_u3072_o),
    .o(_al_u3073_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3074 (
    .a(_al_u2949_o),
    .b(_al_u2926_o),
    .o(_al_u3074_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3075 (
    .a(_al_u3073_o),
    .b(_al_u3074_o),
    .o(_al_u3075_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(~B*~A))"),
    .INIT(8'he0))
    _al_u3076 (
    .a(_al_u2949_o),
    .b(_al_u2887_o),
    .c(_al_u2975_o),
    .o(_al_u3076_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3077 (
    .a(_al_u3076_o),
    .b(_al_u2977_o),
    .o(_al_u3077_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3078 (
    .a(_al_u2898_o),
    .b(_al_u2975_o),
    .o(_al_u3078_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3079 (
    .a(_al_u2899_o),
    .b(_al_u2975_o),
    .o(_al_u3079_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3080 (
    .a(_al_u3078_o),
    .b(_al_u3079_o),
    .o(_al_u3080_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*A)"),
    .INIT(16'h0080))
    _al_u3081 (
    .a(mux92_b0_sel_is_0_o),
    .b(_al_u3077_o),
    .c(_al_u3080_o),
    .d(_al_u2990_o),
    .o(_al_u3081_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*~A)"),
    .INIT(8'h04))
    _al_u3082 (
    .a(_al_u2991_o),
    .b(_al_u3000_o),
    .c(_al_u3001_o),
    .o(mux97_b15_sel_is_2_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3083 (
    .a(_al_u3075_o),
    .b(_al_u3081_o),
    .c(mux97_b15_sel_is_2_o),
    .o(_al_u3083_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u3084 (
    .a(_al_u3083_o),
    .b(_al_u3005_o),
    .c(_al_u2897_o),
    .o(_al_u3084_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3085 (
    .a(_al_u3011_o),
    .b(_al_u3015_o),
    .o(_al_u3085_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3086 (
    .a(_al_u3085_o),
    .b(_al_u3014_o),
    .o(_al_u3086_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*B))"),
    .INIT(8'ha2))
    _al_u3087 (
    .a(_al_u3086_o),
    .b(_al_u3008_o),
    .c(counter[0]),
    .o(_al_u3087_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3088 (
    .a(_al_u2938_o),
    .b(_al_u2993_o),
    .o(_al_u3088_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3089 (
    .a(_al_u2907_o),
    .b(_al_u2993_o),
    .o(_al_u3089_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u3090 (
    .a(_al_u3088_o),
    .b(_al_u3007_o),
    .c(_al_u3089_o),
    .o(_al_u3090_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(~B*~A))"),
    .INIT(8'he0))
    _al_u3091 (
    .a(_al_u2989_o),
    .b(_al_u2899_o),
    .c(_al_u2993_o),
    .o(_al_u3091_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3092 (
    .a(_al_u3090_o),
    .b(_al_u3091_o),
    .o(_al_u3092_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3093 (
    .a(_al_u3084_o),
    .b(_al_u3087_o),
    .c(_al_u3092_o),
    .o(_al_u3093_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(~B*~A))"),
    .INIT(8'he0))
    _al_u3094 (
    .a(_al_u2904_o),
    .b(_al_u2842_o),
    .c(_al_u3010_o),
    .o(_al_u3094_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u3095 (
    .a(_al_u3094_o),
    .b(_al_u2953_o),
    .c(_al_u3010_o),
    .o(_al_u3095_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3096 (
    .a(_al_u3093_o),
    .b(_al_u3095_o),
    .o(_al_u3096_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3097 (
    .a(_al_u3096_o),
    .b(_al_u3031_o),
    .o(_al_u3097_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3098 (
    .a(_al_u2898_o),
    .b(_al_u3026_o),
    .o(_al_u3098_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3099 (
    .a(_al_u2949_o),
    .b(_al_u3026_o),
    .o(_al_u3099_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3100 (
    .a(_al_u3098_o),
    .b(_al_u3099_o),
    .o(mux135_b11_sel_is_0_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3101 (
    .a(_al_u2899_o),
    .b(_al_u3026_o),
    .o(_al_u3101_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3102 (
    .a(_al_u3101_o),
    .b(counter[0]),
    .o(_al_u3102_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3103 (
    .a(_al_u3097_o),
    .b(mux135_b11_sel_is_0_o),
    .c(_al_u3102_o),
    .o(_al_u3103_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    _al_u3104 (
    .a(_al_u2904_o),
    .b(_al_u3026_o),
    .c(_al_u2842_o),
    .o(_al_u3104_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(~B*~A))"),
    .INIT(8'he0))
    _al_u3105 (
    .a(_al_u2925_o),
    .b(_al_u2894_o),
    .c(_al_u2885_o),
    .o(_al_u3105_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u3106 (
    .a(_al_u3103_o),
    .b(_al_u3104_o),
    .c(_al_u3105_o),
    .o(_al_u3106_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3107 (
    .a(_al_u2842_o),
    .b(_al_u2885_o),
    .o(_al_u3107_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3108 (
    .a(_al_u3107_o),
    .b(counter[0]),
    .o(_al_u3108_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3109 (
    .a(_al_u3106_o),
    .b(_al_u3108_o),
    .o(_al_u3109_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3110 (
    .a(_al_u3109_o),
    .b(_al_u3052_o),
    .o(_al_u3110_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3111 (
    .a(_al_u2904_o),
    .b(_al_u3046_o),
    .o(_al_u3111_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3112 (
    .a(_al_u3110_o),
    .b(_al_u3111_o),
    .o(_al_u3112_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3113 (
    .a(_al_u2842_o),
    .b(_al_u3046_o),
    .c(counter[0]),
    .o(_al_u3113_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(B*~(~D*A)))"),
    .INIT(16'h030b))
    _al_u3114 (
    .a(_al_u3112_o),
    .b(n377_lutinv),
    .c(n376_lutinv),
    .d(_al_u3113_o),
    .o(_al_u3114_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3115 (
    .a(_al_u2842_o),
    .b(_al_u3046_o),
    .c(counter[0]),
    .o(_al_u3115_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3116 (
    .a(_al_u3111_o),
    .b(_al_u3115_o),
    .o(mux174_b0_sel_is_0_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3117 (
    .a(mux174_b0_sel_is_0_o),
    .b(_al_u3113_o),
    .o(_al_u3117_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3118 (
    .a(_al_u3117_o),
    .b(n378_lutinv),
    .o(_al_u3118_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C*A))"),
    .INIT(8'hb3))
    _al_u3119 (
    .a(_al_u3055_o),
    .b(_al_u3114_o),
    .c(_al_u3118_o),
    .o(\sel2_b6/or_B6_or_B7_B8_o_o ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3120 (
    .a(_al_u2886_o),
    .b(_al_u2888_o),
    .o(_al_u3120_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3121 (
    .a(n186[0]),
    .b(_al_u3120_o),
    .o(_al_u3121_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(~B*~A))"),
    .INIT(8'he0))
    _al_u3122 (
    .a(_al_u3121_o),
    .b(_al_u2949_o),
    .c(mux9_b12_sel_is_2_o),
    .o(_al_u3122_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3123 (
    .a(_al_u3122_o),
    .b(mux13_b2_sel_is_2_o),
    .o(n197[2]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3124 (
    .a(_al_u2884_o),
    .b(_al_u2915_o),
    .o(_al_u3124_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3125 (
    .a(_al_u2916_o),
    .b(_al_u3124_o),
    .o(mux19_b2_sel_is_0_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3126 (
    .a(n197[2]),
    .b(mux19_b2_sel_is_0_o),
    .c(mux16_b1_sel_is_0_o),
    .o(n214[2]));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u3127 (
    .a(_al_u3072_o),
    .b(_al_u3074_o),
    .c(_al_u2932_o),
    .o(mux38_b12_sel_is_2_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3128 (
    .a(mux38_b12_sel_is_2_o),
    .b(_al_u2929_o),
    .o(mux38_b1_sel_is_2_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3129 (
    .a(n214[2]),
    .b(mux38_b1_sel_is_2_o),
    .o(_al_u3129_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*~A))"),
    .INIT(8'h32))
    _al_u3130 (
    .a(_al_u3129_o),
    .b(_al_u2939_o),
    .c(_al_u3074_o),
    .o(n227[2]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3131 (
    .a(mux60_b10_sel_is_2_o),
    .b(mux52_b1_sel_is_2_o),
    .o(mux60_b1_sel_is_2_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3132 (
    .a(mux60_b1_sel_is_2_o),
    .b(_al_u2946_o),
    .o(_al_u3132_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3133 (
    .a(mux47_b1_sel_is_2_o),
    .b(_al_u2947_o),
    .o(mux48_b1_sel_is_2_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u3134 (
    .a(_al_u2947_o),
    .b(_al_u2941_o),
    .c(counter[0]),
    .o(_al_u3134_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(D*~(C*A)))"),
    .INIT(16'h80cc))
    _al_u3135 (
    .a(n227[2]),
    .b(_al_u3132_o),
    .c(mux48_b1_sel_is_2_o),
    .d(_al_u3134_o),
    .o(_al_u3135_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B)*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+A*~(B)*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h32aa))
    _al_u3136 (
    .a(_al_u3135_o),
    .b(_al_u2904_o),
    .c(_al_u2907_o),
    .d(_al_u2945_o),
    .o(_al_u3136_o));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'h47))
    _al_u3137 (
    .a(_al_u2925_o),
    .b(_al_u2963_o),
    .c(_al_u3136_o),
    .o(_al_u3137_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3138 (
    .a(_al_u2887_o),
    .b(_al_u2963_o),
    .o(_al_u3138_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3139 (
    .a(_al_u2949_o),
    .b(_al_u2963_o),
    .o(_al_u3139_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3140 (
    .a(_al_u3138_o),
    .b(_al_u3139_o),
    .o(mux70_b2_sel_is_0_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3141 (
    .a(mux70_b2_sel_is_0_o),
    .b(_al_u2968_o),
    .o(_al_u3141_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3142 (
    .a(_al_u3137_o),
    .b(_al_u3141_o),
    .c(mux75_b5_sel_is_2_o),
    .o(_al_u3142_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3143 (
    .a(_al_u2904_o),
    .b(_al_u2963_o),
    .o(_al_u3143_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3144 (
    .a(_al_u2907_o),
    .b(_al_u2963_o),
    .o(_al_u3144_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3145 (
    .a(_al_u3143_o),
    .b(_al_u3144_o),
    .o(_al_u3145_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3146 (
    .a(_al_u2938_o),
    .b(_al_u2963_o),
    .o(_al_u3146_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    _al_u3147 (
    .a(_al_u3142_o),
    .b(_al_u3145_o),
    .c(_al_u3146_o),
    .o(_al_u3147_o));
  AL_MAP_LUT3 #(
    .EQN("~(~A*~(B)*~(C)+~A*B*~(C)+~(~A)*B*C+~A*B*C)"),
    .INIT(8'h3a))
    _al_u3148 (
    .a(_al_u3147_o),
    .b(_al_u2884_o),
    .c(_al_u2975_o),
    .o(_al_u3148_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*A)"),
    .INIT(16'h0080))
    _al_u3149 (
    .a(mux92_b0_sel_is_0_o),
    .b(_al_u3080_o),
    .c(mux97_b15_sel_is_2_o),
    .d(_al_u2990_o),
    .o(mux97_b5_sel_is_2_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*A))"),
    .INIT(8'hc4))
    _al_u3150 (
    .a(_al_u3148_o),
    .b(mux97_b5_sel_is_2_o),
    .c(_al_u2977_o),
    .o(_al_u3150_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3151 (
    .a(_al_u3150_o),
    .b(_al_u3005_o),
    .o(_al_u3151_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3152 (
    .a(_al_u3151_o),
    .b(_al_u3088_o),
    .o(_al_u3152_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3153 (
    .a(_al_u2949_o),
    .b(_al_u3010_o),
    .o(_al_u3153_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3154 (
    .a(_al_u3024_o),
    .b(_al_u3153_o),
    .o(mux119_b3_sel_is_0_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3155 (
    .a(_al_u2905_o),
    .b(_al_u3010_o),
    .o(_al_u3155_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3156 (
    .a(_al_u3155_o),
    .b(counter[0]),
    .c(counter[1]),
    .o(_al_u3156_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3157 (
    .a(mux119_b3_sel_is_0_o),
    .b(_al_u3156_o),
    .o(mux120_b3_sel_is_2_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(~B*~A))"),
    .INIT(8'he0))
    _al_u3158 (
    .a(_al_u2887_o),
    .b(_al_u2891_o),
    .c(_al_u3010_o),
    .o(_al_u3158_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3159 (
    .a(mux120_b3_sel_is_2_o),
    .b(_al_u3158_o),
    .o(mux120_b7_sel_is_2_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u3160 (
    .a(_al_u3155_o),
    .b(counter[0]),
    .c(counter[1]),
    .o(_al_u3160_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3161 (
    .a(mux120_b7_sel_is_2_o),
    .b(_al_u3160_o),
    .o(mux121_b7_sel_is_2_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3162 (
    .a(_al_u3155_o),
    .b(counter[1]),
    .o(_al_u3162_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*A)"),
    .INIT(16'h0080))
    _al_u3163 (
    .a(_al_u3152_o),
    .b(mux121_b7_sel_is_2_o),
    .c(mux115_b2_sel_is_2_o),
    .d(_al_u3162_o),
    .o(_al_u3163_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3164 (
    .a(_al_u3162_o),
    .b(counter[0]),
    .o(_al_u3164_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(~B*~A))"),
    .INIT(8'he0))
    _al_u3165 (
    .a(_al_u2925_o),
    .b(_al_u2894_o),
    .c(_al_u3026_o),
    .o(_al_u3165_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(~D*C*B))"),
    .INIT(16'h5515))
    _al_u3166 (
    .a(_al_u3165_o),
    .b(_al_u2842_o),
    .c(_al_u3010_o),
    .d(counter[0]),
    .o(mux129_b8_sel_is_2_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(~D*~C))"),
    .INIT(16'h8880))
    _al_u3167 (
    .a(_al_u2903_o),
    .b(_al_u3010_o),
    .c(counter[0]),
    .d(counter[1]),
    .o(_al_u3167_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*~(~B*~A))"),
    .INIT(16'h00e0))
    _al_u3168 (
    .a(_al_u3163_o),
    .b(_al_u3164_o),
    .c(mux129_b8_sel_is_2_o),
    .d(_al_u3167_o),
    .o(_al_u3168_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3169 (
    .a(_al_u3168_o),
    .b(mux132_b0_sel_is_0_o),
    .o(_al_u3169_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3170 (
    .a(_al_u3102_o),
    .b(_al_u3098_o),
    .o(mux136_b1_sel_is_0_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3171 (
    .a(_al_u3101_o),
    .b(counter[0]),
    .o(_al_u3171_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3172 (
    .a(mux136_b1_sel_is_0_o),
    .b(_al_u3171_o),
    .o(mux137_b5_sel_is_2_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3173 (
    .a(mux137_b5_sel_is_2_o),
    .b(_al_u3099_o),
    .o(mux137_b2_sel_is_2_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(~B*~A))"),
    .INIT(8'he0))
    _al_u3174 (
    .a(_al_u2907_o),
    .b(_al_u2908_o),
    .c(_al_u3026_o),
    .o(_al_u3174_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u3175 (
    .a(_al_u2904_o),
    .b(_al_u3174_o),
    .c(_al_u3026_o),
    .o(mux141_b1_sel_is_2_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3176 (
    .a(_al_u2914_o),
    .b(_al_u2885_o),
    .o(_al_u3176_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(~B*~A))"),
    .INIT(8'he0))
    _al_u3177 (
    .a(_al_u2884_o),
    .b(_al_u2925_o),
    .c(_al_u2885_o),
    .o(_al_u3177_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u3178 (
    .a(_al_u3177_o),
    .b(_al_u2894_o),
    .c(_al_u2885_o),
    .o(mux146_b12_sel_is_2_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u3179 (
    .a(_al_u3176_o),
    .b(mux146_b12_sel_is_2_o),
    .o(mux147_b12_sel_is_2_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*A)"),
    .INIT(16'h0080))
    _al_u3180 (
    .a(mux137_b2_sel_is_2_o),
    .b(mux141_b1_sel_is_2_o),
    .c(mux147_b12_sel_is_2_o),
    .d(_al_u3104_o),
    .o(_al_u3180_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u3181 (
    .a(_al_u3169_o),
    .b(_al_u3180_o),
    .c(_al_u3176_o),
    .o(_al_u3181_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3182 (
    .a(_al_u3046_o),
    .b(_al_u2894_o),
    .o(_al_u3182_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3183 (
    .a(_al_u3047_o),
    .b(_al_u3182_o),
    .o(_al_u3183_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3184 (
    .a(_al_u3046_o),
    .b(_al_u2884_o),
    .o(_al_u3184_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3185 (
    .a(_al_u3183_o),
    .b(_al_u3184_o),
    .o(_al_u3185_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3186 (
    .a(_al_u3107_o),
    .b(counter[0]),
    .o(_al_u3186_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3187 (
    .a(_al_u3185_o),
    .b(_al_u3186_o),
    .o(_al_u3187_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3188 (
    .a(_al_u2949_o),
    .b(_al_u2885_o),
    .o(_al_u3188_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(~B*~A))"),
    .INIT(8'he0))
    _al_u3189 (
    .a(_al_u2887_o),
    .b(_al_u2891_o),
    .c(_al_u2885_o),
    .o(_al_u3189_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3190 (
    .a(_al_u3188_o),
    .b(_al_u3189_o),
    .o(mux150_b0_sel_is_2_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u3191 (
    .a(_al_u2935_o),
    .b(_al_u2885_o),
    .o(_al_u3191_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3192 (
    .a(mux150_b0_sel_is_2_o),
    .b(_al_u3191_o),
    .o(mux152_b0_sel_is_2_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3193 (
    .a(_al_u2907_o),
    .b(_al_u3026_o),
    .o(_al_u3193_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u3194 (
    .a(_al_u3034_o),
    .b(_al_u3193_o),
    .c(_al_u3107_o),
    .o(_al_u3194_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(~A*~(~D*B)))"),
    .INIT(16'ha0e0))
    _al_u3195 (
    .a(_al_u2907_o),
    .b(_al_u2908_o),
    .c(_al_u2885_o),
    .d(counter[0]),
    .o(_al_u3195_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u3196 (
    .a(_al_u2904_o),
    .b(_al_u3195_o),
    .c(_al_u2885_o),
    .o(_al_u3196_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u3197 (
    .a(mux152_b0_sel_is_2_o),
    .b(_al_u3194_o),
    .c(_al_u3196_o),
    .d(_al_u3041_o),
    .o(_al_u3197_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3198 (
    .a(_al_u3181_o),
    .b(_al_u3187_o),
    .c(_al_u3197_o),
    .o(_al_u3198_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u3199 (
    .a(_al_u3198_o),
    .b(_al_u3046_o),
    .c(_al_u2891_o),
    .o(_al_u3199_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3200 (
    .a(_al_u3199_o),
    .b(_al_u3118_o),
    .c(mux170_b2_sel_is_2_o),
    .o(_al_u3200_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3201 (
    .a(_al_u3065_o),
    .b(_al_u2890_o),
    .o(_al_u3201_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u3202 (
    .a(_al_u2889_o),
    .b(_al_u3201_o),
    .o(_al_u3202_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(~B*A))"),
    .INIT(8'h0d))
    _al_u3203 (
    .a(_al_u3202_o),
    .b(_al_u2900_o),
    .c(_al_u2906_o),
    .o(_al_u3203_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3204 (
    .a(_al_u2925_o),
    .b(_al_u2915_o),
    .o(_al_u3204_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3205 (
    .a(_al_u3204_o),
    .b(_al_u3124_o),
    .o(_al_u3205_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*~A)"),
    .INIT(8'h04))
    _al_u3206 (
    .a(_al_u3203_o),
    .b(_al_u3205_o),
    .c(_al_u2909_o),
    .o(_al_u3206_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3207 (
    .a(_al_u2887_o),
    .b(_al_u2915_o),
    .o(_al_u3207_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3208 (
    .a(_al_u3206_o),
    .b(_al_u3207_o),
    .o(_al_u3208_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3209 (
    .a(_al_u2936_o),
    .b(_al_u2915_o),
    .o(_al_u3209_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u3210 (
    .a(_al_u3208_o),
    .b(_al_u2920_o),
    .c(_al_u3209_o),
    .o(_al_u3210_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3211 (
    .a(_al_u2930_o),
    .b(counter[0]),
    .o(_al_u3211_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u3212 (
    .a(_al_u3211_o),
    .b(_al_u2929_o),
    .o(mux33_b0_sel_is_2_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3213 (
    .a(_al_u3210_o),
    .b(mux33_b0_sel_is_2_o),
    .o(_al_u3213_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*~B))"),
    .INIT(8'h8a))
    _al_u3214 (
    .a(_al_u3213_o),
    .b(_al_u2891_o),
    .c(_al_u2926_o),
    .o(_al_u3214_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*~(~D*~A))"),
    .INIT(16'hc080))
    _al_u3215 (
    .a(_al_u3214_o),
    .b(mux49_b0_sel_is_2_o),
    .c(mux52_b1_sel_is_2_o),
    .d(_al_u3074_o),
    .o(_al_u3215_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3216 (
    .a(_al_u3215_o),
    .b(_al_u3081_o),
    .o(_al_u3216_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3217 (
    .a(_al_u3216_o),
    .b(_al_u2997_o),
    .o(_al_u3217_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3218 (
    .a(_al_u3005_o),
    .b(counter[0]),
    .c(counter[1]),
    .o(_al_u3218_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3219 (
    .a(_al_u2994_o),
    .b(_al_u3218_o),
    .o(_al_u3219_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3220 (
    .a(_al_u2899_o),
    .b(_al_u2993_o),
    .o(_al_u3220_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3221 (
    .a(_al_u3220_o),
    .b(counter[0]),
    .o(_al_u3221_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3222 (
    .a(_al_u3217_o),
    .b(_al_u3219_o),
    .c(_al_u3221_o),
    .o(_al_u3222_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u3223 (
    .a(_al_u3222_o),
    .b(_al_u2903_o),
    .c(_al_u2993_o),
    .o(_al_u3223_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3224 (
    .a(_al_u3223_o),
    .b(_al_u3020_o),
    .o(_al_u3224_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3225 (
    .a(_al_u3224_o),
    .b(_al_u3156_o),
    .o(_al_u3225_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u3226 (
    .a(_al_u3225_o),
    .b(_al_u3094_o),
    .c(_al_u3030_o),
    .o(_al_u3226_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3227 (
    .a(_al_u2887_o),
    .b(_al_u3026_o),
    .o(_al_u3227_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3228 (
    .a(_al_u3099_o),
    .b(_al_u3227_o),
    .o(_al_u3228_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3229 (
    .a(_al_u3226_o),
    .b(_al_u3228_o),
    .o(_al_u3229_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u3230 (
    .a(_al_u3229_o),
    .b(_al_u2905_o),
    .c(_al_u3026_o),
    .o(_al_u3230_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*B))"),
    .INIT(8'ha2))
    _al_u3231 (
    .a(_al_u3230_o),
    .b(_al_u2885_o),
    .c(_al_u2894_o),
    .o(_al_u3231_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~A*~(D*C))"),
    .INIT(16'h0111))
    _al_u3232 (
    .a(_al_u3231_o),
    .b(_al_u3044_o),
    .c(_al_u2907_o),
    .d(_al_u2885_o),
    .o(_al_u3232_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3233 (
    .a(_al_u3232_o),
    .b(_al_u3108_o),
    .o(_al_u3233_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3234 (
    .a(_al_u2949_o),
    .b(_al_u3046_o),
    .o(_al_u3234_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    _al_u3235 (
    .a(_al_u2914_o),
    .b(_al_u3046_o),
    .c(_al_u2891_o),
    .o(_al_u3235_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u3236 (
    .a(_al_u3233_o),
    .b(_al_u3234_o),
    .c(_al_u3235_o),
    .o(_al_u3236_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3237 (
    .a(_al_u3050_o),
    .b(counter[0]),
    .o(_al_u3237_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3238 (
    .a(_al_u3052_o),
    .b(_al_u3237_o),
    .o(mux170_b10_sel_is_0_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    _al_u3239 (
    .a(_al_u2938_o),
    .b(_al_u3046_o),
    .c(_al_u2907_o),
    .o(_al_u3239_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u3240 (
    .a(mux170_b10_sel_is_0_o),
    .b(_al_u3239_o),
    .c(_al_u3111_o),
    .o(_al_u3240_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3241 (
    .a(_al_u3236_o),
    .b(_al_u3240_o),
    .o(_al_u3241_o));
  AL_MAP_LUT4 #(
    .EQN("~(~A*~(C*~(~D*B)))"),
    .INIT(16'hfaba))
    _al_u3242 (
    .a(_al_u3200_o),
    .b(_al_u3241_o),
    .c(n377_lutinv),
    .d(_al_u3113_o),
    .o(\sel2_b2/or_B6_or_B7_B8_o_o ));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*~A)"),
    .INIT(8'h04))
    _al_u3243 (
    .a(_al_u2889_o),
    .b(_al_u3067_o),
    .c(_al_u2844_o),
    .o(n190[7]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(C*B*A))"),
    .INIT(16'h007f))
    _al_u3244 (
    .a(_al_u3058_o),
    .b(n190[7]),
    .c(mux14_b11_sel_is_2_o),
    .d(_al_u2911_o),
    .o(_al_u3244_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3245 (
    .a(_al_u2949_o),
    .b(_al_u2915_o),
    .o(_al_u3245_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3246 (
    .a(_al_u2918_o),
    .b(_al_u3245_o),
    .o(mux22_b11_sel_is_2_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3247 (
    .a(_al_u3205_o),
    .b(_al_u3059_o),
    .o(mux18_b6_sel_is_2_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    _al_u3248 (
    .a(_al_u3244_o),
    .b(mux22_b11_sel_is_2_o),
    .c(mux18_b6_sel_is_2_o),
    .o(n210[7]));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3249 (
    .a(n210[7]),
    .b(_al_u2922_o),
    .c(mux33_b0_sel_is_2_o),
    .o(_al_u3249_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(B*~(~D*~A)))"),
    .INIT(16'h0307))
    _al_u3250 (
    .a(_al_u3249_o),
    .b(mux38_b12_sel_is_2_o),
    .c(_al_u3074_o),
    .d(_al_u2927_o),
    .o(_al_u3250_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u3251 (
    .a(_al_u3250_o),
    .b(_al_u2935_o),
    .c(_al_u2926_o),
    .o(n225[7]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3252 (
    .a(mux63_b1_sel_is_2_o),
    .b(mux48_b1_sel_is_2_o),
    .o(_al_u3252_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(~B*~A))"),
    .INIT(8'he0))
    _al_u3253 (
    .a(_al_u2938_o),
    .b(_al_u2907_o),
    .c(_al_u2926_o),
    .o(_al_u3253_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    _al_u3254 (
    .a(n225[7]),
    .b(_al_u3252_o),
    .c(_al_u3253_o),
    .d(_al_u2946_o),
    .o(n247[7]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3255 (
    .a(n247[7]),
    .b(mux67_b0_sel_is_2_o),
    .o(n258[7]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3256 (
    .a(_al_u2842_o),
    .b(_al_u2963_o),
    .o(_al_u3256_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3257 (
    .a(_al_u3145_o),
    .b(_al_u3256_o),
    .o(_al_u3257_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*A)"),
    .INIT(16'h0002))
    _al_u3258 (
    .a(mux92_b0_sel_is_0_o),
    .b(_al_u2990_o),
    .c(_al_u2984_o),
    .d(_al_u2980_o),
    .o(_al_u3258_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3259 (
    .a(_al_u3080_o),
    .b(_al_u3076_o),
    .o(mux89_b1_sel_is_2_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u3260 (
    .a(_al_u3257_o),
    .b(_al_u3258_o),
    .c(mux89_b1_sel_is_2_o),
    .d(mux84_b4_sel_is_2_o),
    .o(mux92_b7_sel_is_2_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3261 (
    .a(n258[7]),
    .b(mux92_b7_sel_is_2_o),
    .o(n275[7]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3262 (
    .a(n275[7]),
    .b(_al_u3001_o),
    .o(_al_u3262_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*~B))"),
    .INIT(8'h8a))
    _al_u3263 (
    .a(_al_u3262_o),
    .b(_al_u2897_o),
    .c(_al_u2993_o),
    .o(_al_u3263_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u3264 (
    .a(_al_u3221_o),
    .b(_al_u3005_o),
    .c(_al_u2897_o),
    .o(_al_u3264_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u3265 (
    .a(_al_u3263_o),
    .b(_al_u3264_o),
    .o(_al_u3265_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u3266 (
    .a(_al_u3265_o),
    .b(_al_u3012_o),
    .o(_al_u3266_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3267 (
    .a(_al_u3266_o),
    .b(mux121_b7_sel_is_2_o),
    .o(_al_u3267_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3268 (
    .a(_al_u2842_o),
    .b(_al_u3010_o),
    .c(counter[0]),
    .o(_al_u3268_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~C*~(~D*A)))"),
    .INIT(16'hc0c8))
    _al_u3269 (
    .a(_al_u3267_o),
    .b(mux129_b8_sel_is_2_o),
    .c(_al_u3268_o),
    .d(_al_u3167_o),
    .o(_al_u3269_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u3270 (
    .a(_al_u3269_o),
    .b(_al_u2925_o),
    .c(_al_u3026_o),
    .o(_al_u3270_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3271 (
    .a(_al_u3270_o),
    .b(_al_u3027_o),
    .o(_al_u3271_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(~B*~A))"),
    .INIT(8'he0))
    _al_u3272 (
    .a(_al_u2904_o),
    .b(_al_u2907_o),
    .c(_al_u3026_o),
    .o(_al_u3272_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u3273 (
    .a(_al_u3271_o),
    .b(_al_u3171_o),
    .c(_al_u3272_o),
    .o(_al_u3273_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u3274 (
    .a(_al_u3273_o),
    .b(mux146_b12_sel_is_2_o),
    .o(_al_u3274_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3275 (
    .a(_al_u3274_o),
    .b(_al_u3188_o),
    .o(_al_u3275_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u3276 (
    .a(_al_u2953_o),
    .b(_al_u2885_o),
    .o(_al_u3276_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(~A*~(D)*~(C)+~A*D*~(C)+~(~A)*D*C+~A*D*C))"),
    .INIT(16'h0232))
    _al_u3277 (
    .a(_al_u3275_o),
    .b(_al_u3276_o),
    .c(_al_u3040_o),
    .d(counter[0]),
    .o(_al_u3277_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(~B*~A))"),
    .INIT(8'he0))
    _al_u3278 (
    .a(_al_u2904_o),
    .b(_al_u2842_o),
    .c(_al_u2885_o),
    .o(_al_u3278_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*~A))"),
    .INIT(8'h32))
    _al_u3279 (
    .a(_al_u3277_o),
    .b(_al_u3278_o),
    .c(_al_u3195_o),
    .o(_al_u3279_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3280 (
    .a(_al_u3235_o),
    .b(_al_u3184_o),
    .o(_al_u3280_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3281 (
    .a(_al_u3279_o),
    .b(_al_u3280_o),
    .c(_al_u3047_o),
    .o(_al_u3281_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3282 (
    .a(_al_u3281_o),
    .b(mux170_b2_sel_is_2_o),
    .c(_al_u3111_o),
    .o(_al_u3282_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3283 (
    .a(_al_u3282_o),
    .b(n378_lutinv),
    .c(_al_u3113_o),
    .o(_al_u3283_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3284 (
    .a(_al_u2930_o),
    .b(counter[0]),
    .o(_al_u3284_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3285 (
    .a(_al_u2922_o),
    .b(_al_u3284_o),
    .o(mux30_b1_sel_is_2_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(~B*A))"),
    .INIT(8'hd0))
    _al_u3286 (
    .a(_al_u2935_o),
    .b(_al_u2949_o),
    .c(_al_u2915_o),
    .o(_al_u3286_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u3287 (
    .a(_al_u2923_o),
    .b(counter[0]),
    .c(counter[1]),
    .o(_al_u3287_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u3288 (
    .a(mux30_b1_sel_is_2_o),
    .b(_al_u3286_o),
    .c(_al_u3287_o),
    .o(mux30_b12_sel_is_2_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    _al_u3289 (
    .a(mux30_b12_sel_is_2_o),
    .b(mux33_b0_sel_is_2_o),
    .c(_al_u2976_o),
    .d(_al_u2945_o),
    .o(_al_u3289_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(~B*~A))"),
    .INIT(8'he0))
    _al_u3290 (
    .a(_al_u2898_o),
    .b(_al_u2949_o),
    .c(_al_u2888_o),
    .o(_al_u3290_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u3291 (
    .a(_al_u3290_o),
    .b(_al_u3067_o),
    .o(_al_u3291_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3292 (
    .a(_al_u3256_o),
    .b(counter[0]),
    .o(_al_u3292_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u3293 (
    .a(_al_u3292_o),
    .b(_al_u2984_o),
    .c(_al_u2980_o),
    .o(_al_u3293_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3294 (
    .a(_al_u3289_o),
    .b(_al_u3291_o),
    .c(_al_u3293_o),
    .o(_al_u3294_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u3295 (
    .a(_al_u2916_o),
    .b(_al_u2917_o),
    .c(_al_u3124_o),
    .o(_al_u3295_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3296 (
    .a(mux38_b12_sel_is_2_o),
    .b(_al_u3295_o),
    .c(_al_u3204_o),
    .o(_al_u3296_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*A)"),
    .INIT(16'h0080))
    _al_u3297 (
    .a(_al_u3294_o),
    .b(mux47_b0_sel_is_2_o),
    .c(_al_u3296_o),
    .d(_al_u2963_o),
    .o(_al_u3297_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3298 (
    .a(_al_u3297_o),
    .b(_al_u2996_o),
    .c(mux97_b15_sel_is_2_o),
    .o(_al_u3298_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*B))"),
    .INIT(8'ha2))
    _al_u3299 (
    .a(_al_u3298_o),
    .b(_al_u3220_o),
    .c(counter[0]),
    .o(_al_u3299_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3300 (
    .a(_al_u3299_o),
    .b(_al_u3090_o),
    .o(_al_u3300_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3301 (
    .a(_al_u3300_o),
    .b(_al_u3052_o),
    .o(_al_u3301_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3302 (
    .a(_al_u3301_o),
    .b(_al_u3111_o),
    .o(_al_u3302_o));
  AL_MAP_LUT4 #(
    .EQN("~(~A*~(C*~(~D*B)))"),
    .INIT(16'hfaba))
    _al_u3303 (
    .a(_al_u3283_o),
    .b(_al_u3302_o),
    .c(n377_lutinv),
    .d(_al_u3113_o),
    .o(\sel2_b7/or_B6_or_B7_B8_o_o ));
  AL_MAP_LUT3 #(
    .EQN("(C*~(~B*~A))"),
    .INIT(8'he0))
    _al_u3304 (
    .a(_al_u2884_o),
    .b(_al_u2925_o),
    .c(_al_u2888_o),
    .o(_al_u3304_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~A*~(D*~C))"),
    .INIT(16'h1011))
    _al_u3305 (
    .a(_al_u2844_o),
    .b(_al_u2895_o),
    .c(_al_u2890_o),
    .d(_al_u3304_o),
    .o(n187[3]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u3306 (
    .a(_al_u2889_o),
    .b(n187[3]),
    .o(n189[3]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u3307 (
    .a(_al_u3056_o),
    .b(mux14_b11_sel_is_2_o),
    .o(mux14_b0_sel_is_2_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3308 (
    .a(_al_u2899_o),
    .b(_al_u2888_o),
    .c(counter[0]),
    .o(_al_u3308_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~D*~(C*A)))"),
    .INIT(16'hcc80))
    _al_u3309 (
    .a(n189[3]),
    .b(mux14_b0_sel_is_2_o),
    .c(mux9_b12_sel_is_2_o),
    .d(_al_u3308_o),
    .o(n198[3]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3310 (
    .a(n198[3]),
    .b(_al_u3059_o),
    .o(n200[3]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3311 (
    .a(_al_u2891_o),
    .b(_al_u2915_o),
    .o(_al_u3311_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u3312 (
    .a(n200[3]),
    .b(_al_u3311_o),
    .c(_al_u3124_o),
    .o(n205[3]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*~B))"),
    .INIT(8'h8a))
    _al_u3313 (
    .a(n205[3]),
    .b(_al_u2935_o),
    .c(_al_u2915_o),
    .o(n208[3]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*B))"),
    .INIT(8'ha2))
    _al_u3314 (
    .a(n208[3]),
    .b(_al_u2923_o),
    .c(counter[1]),
    .o(_al_u3314_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u3315 (
    .a(mux38_b1_sel_is_2_o),
    .b(_al_u2920_o),
    .c(_al_u2930_o),
    .o(_al_u3315_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3316 (
    .a(_al_u2923_o),
    .b(_al_u2897_o),
    .o(_al_u3316_o));
  AL_MAP_LUT4 #(
    .EQN("~(~C*~((~D*~A))*~(B)+~C*(~D*~A)*~(B)+~(~C)*(~D*~A)*B+~C*(~D*~A)*B)"),
    .INIT(16'hfcb8))
    _al_u3317 (
    .a(_al_u3314_o),
    .b(_al_u3315_o),
    .c(_al_u3074_o),
    .d(_al_u3316_o),
    .o(_al_u3317_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u3318 (
    .a(_al_u2937_o),
    .b(_al_u2926_o),
    .o(_al_u3318_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3319 (
    .a(_al_u2989_o),
    .b(_al_u2926_o),
    .o(_al_u3319_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(~D*~(~B*A)))"),
    .INIT(16'h0f02))
    _al_u3320 (
    .a(_al_u3317_o),
    .b(_al_u3318_o),
    .c(_al_u3253_o),
    .d(_al_u3319_o),
    .o(_al_u3320_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3321 (
    .a(_al_u3320_o),
    .b(_al_u2941_o),
    .o(_al_u3321_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(~B*~A))"),
    .INIT(8'he0))
    _al_u3322 (
    .a(_al_u2914_o),
    .b(_al_u2891_o),
    .c(_al_u2963_o),
    .o(_al_u3322_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3323 (
    .a(_al_u2884_o),
    .b(_al_u2963_o),
    .o(_al_u3323_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3324 (
    .a(_al_u3322_o),
    .b(_al_u3323_o),
    .o(mux68_b1_sel_is_2_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(~B*~A))"),
    .INIT(8'he0))
    _al_u3325 (
    .a(_al_u2925_o),
    .b(_al_u2894_o),
    .c(_al_u2963_o),
    .o(_al_u3325_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3326 (
    .a(mux68_b1_sel_is_2_o),
    .b(_al_u3325_o),
    .o(_al_u3326_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3327 (
    .a(_al_u3326_o),
    .b(_al_u2959_o),
    .o(_al_u3327_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3328 (
    .a(_al_u2952_o),
    .b(_al_u2956_o),
    .o(mux57_b3_sel_is_2_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D*~(C*~B)))"),
    .INIT(16'h20aa))
    _al_u3329 (
    .a(mux57_b3_sel_is_2_o),
    .b(_al_u2904_o),
    .c(_al_u2953_o),
    .d(_al_u2945_o),
    .o(mux61_b3_sel_is_2_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3330 (
    .a(_al_u3327_o),
    .b(mux61_b3_sel_is_2_o),
    .o(_al_u3330_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3331 (
    .a(_al_u3321_o),
    .b(_al_u3330_o),
    .c(_al_u2946_o),
    .o(_al_u3331_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3332 (
    .a(_al_u2891_o),
    .b(_al_u2963_o),
    .o(_al_u3332_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    _al_u3333 (
    .a(_al_u3331_o),
    .b(mux70_b2_sel_is_0_o),
    .c(_al_u3332_o),
    .o(_al_u3333_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u3334 (
    .a(_al_u3333_o),
    .b(_al_u3143_o),
    .c(_al_u2964_o),
    .o(_al_u3334_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3335 (
    .a(_al_u3334_o),
    .b(_al_u2984_o),
    .o(_al_u3335_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3336 (
    .a(_al_u2914_o),
    .b(_al_u2975_o),
    .o(_al_u3336_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u3337 (
    .a(_al_u3335_o),
    .b(_al_u3336_o),
    .c(_al_u3076_o),
    .o(_al_u3337_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3338 (
    .a(_al_u3337_o),
    .b(mux93_b3_sel_is_2_o),
    .o(_al_u3338_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*~C))"),
    .INIT(16'h8088))
    _al_u3339 (
    .a(_al_u3338_o),
    .b(_al_u3000_o),
    .c(_al_u2995_o),
    .d(_al_u2993_o),
    .o(_al_u3339_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u3340 (
    .a(_al_u3005_o),
    .b(counter[0]),
    .c(counter[1]),
    .o(_al_u3340_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3341 (
    .a(_al_u3221_o),
    .b(_al_u3340_o),
    .o(_al_u3341_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*~A)"),
    .INIT(8'h04))
    _al_u3342 (
    .a(_al_u3339_o),
    .b(_al_u3341_o),
    .c(_al_u3089_o),
    .o(_al_u3342_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*A))"),
    .INIT(8'hc4))
    _al_u3343 (
    .a(_al_u3342_o),
    .b(_al_u3087_o),
    .c(_al_u3008_o),
    .o(_al_u3343_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*~A))"),
    .INIT(8'h23))
    _al_u3344 (
    .a(_al_u3343_o),
    .b(_al_u3013_o),
    .c(_al_u3016_o),
    .o(_al_u3344_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3345 (
    .a(_al_u2907_o),
    .b(_al_u3010_o),
    .o(_al_u3345_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3346 (
    .a(_al_u3164_o),
    .b(_al_u3345_o),
    .o(mux124_b0_sel_is_0_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3347 (
    .a(mux124_b0_sel_is_0_o),
    .b(_al_u3155_o),
    .o(mux124_b11_sel_is_2_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3348 (
    .a(_al_u2894_o),
    .b(_al_u3026_o),
    .o(_al_u3348_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3349 (
    .a(_al_u3094_o),
    .b(_al_u3348_o),
    .o(_al_u3349_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D*~(~C*~B)))"),
    .INIT(16'h02aa))
    _al_u3350 (
    .a(_al_u3349_o),
    .b(_al_u2884_o),
    .c(_al_u2925_o),
    .d(_al_u3026_o),
    .o(mux130_b1_sel_is_2_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u3351 (
    .a(mux124_b11_sel_is_2_o),
    .b(mux130_b1_sel_is_2_o),
    .c(mux132_b0_sel_is_0_o),
    .d(mux119_b3_sel_is_0_o),
    .o(mux132_b3_sel_is_2_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3352 (
    .a(_al_u3344_o),
    .b(mux132_b3_sel_is_2_o),
    .c(mux137_b2_sel_is_2_o),
    .o(_al_u3352_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3353 (
    .a(_al_u3352_o),
    .b(_al_u3034_o),
    .o(_al_u3353_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3354 (
    .a(_al_u2842_o),
    .b(_al_u3026_o),
    .c(counter[0]),
    .o(_al_u3354_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3355 (
    .a(mux147_b12_sel_is_2_o),
    .b(_al_u3354_o),
    .o(_al_u3355_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3356 (
    .a(_al_u3355_o),
    .b(_al_u3104_o),
    .o(mux147_b3_sel_is_2_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3357 (
    .a(_al_u3353_o),
    .b(mux147_b3_sel_is_2_o),
    .c(_al_u3037_o),
    .o(_al_u3357_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u3358 (
    .a(_al_u3278_o),
    .b(_al_u2907_o),
    .c(_al_u2885_o),
    .o(mux159_b3_sel_is_2_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u3359 (
    .a(_al_u2951_o),
    .b(_al_u2885_o),
    .o(_al_u3359_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3360 (
    .a(_al_u3357_o),
    .b(mux159_b3_sel_is_2_o),
    .c(_al_u3359_o),
    .o(_al_u3360_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3361 (
    .a(_al_u3360_o),
    .b(_al_u3047_o),
    .o(_al_u3361_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3362 (
    .a(_al_u2887_o),
    .b(_al_u3046_o),
    .o(_al_u3362_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D*~C*A))"),
    .INIT(16'h3133))
    _al_u3363 (
    .a(_al_u3361_o),
    .b(_al_u3234_o),
    .c(_al_u3362_o),
    .d(mux170_b2_sel_is_2_o),
    .o(_al_u3363_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u3364 (
    .a(_al_u3081_o),
    .b(_al_u2991_o),
    .c(_al_u3001_o),
    .o(_al_u3364_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3365 (
    .a(_al_u3065_o),
    .b(counter[0]),
    .o(_al_u3365_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u3366 (
    .a(_al_u2889_o),
    .b(_al_u3365_o),
    .c(_al_u2892_o),
    .o(_al_u3366_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3367 (
    .a(_al_u3058_o),
    .b(_al_u3366_o),
    .o(_al_u3367_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3368 (
    .a(_al_u3367_o),
    .b(_al_u3124_o),
    .o(_al_u3368_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u3369 (
    .a(_al_u2921_o),
    .b(_al_u3368_o),
    .o(_al_u3369_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(B*~(~C*A)))"),
    .INIT(16'h003b))
    _al_u3370 (
    .a(_al_u3369_o),
    .b(mux33_b0_sel_is_2_o),
    .c(_al_u2930_o),
    .d(_al_u2927_o),
    .o(_al_u3370_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u3371 (
    .a(_al_u3370_o),
    .b(_al_u2891_o),
    .c(_al_u2926_o),
    .o(_al_u3371_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u3372 (
    .a(_al_u3364_o),
    .b(_al_u2998_o),
    .c(_al_u3371_o),
    .o(_al_u3372_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3373 (
    .a(_al_u3372_o),
    .b(_al_u2995_o),
    .o(_al_u3373_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3374 (
    .a(_al_u3373_o),
    .b(_al_u3218_o),
    .o(_al_u3374_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3375 (
    .a(_al_u3374_o),
    .b(_al_u3012_o),
    .c(_al_u3088_o),
    .o(_al_u3375_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3376 (
    .a(_al_u3375_o),
    .b(_al_u3014_o),
    .o(_al_u3376_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3377 (
    .a(mux119_b3_sel_is_0_o),
    .b(_al_u3022_o),
    .o(_al_u3377_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3378 (
    .a(_al_u3376_o),
    .b(_al_u3377_o),
    .o(_al_u3378_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3379 (
    .a(_al_u3378_o),
    .b(_al_u3349_o),
    .o(_al_u3379_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u3380 (
    .a(_al_u3379_o),
    .b(_al_u3227_o),
    .c(_al_u3030_o),
    .o(_al_u3380_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3381 (
    .a(_al_u3380_o),
    .b(_al_u3102_o),
    .o(_al_u3381_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u3382 (
    .a(_al_u3381_o),
    .b(_al_u2904_o),
    .c(_al_u3026_o),
    .o(_al_u3382_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(D*C))"),
    .INIT(16'h0444))
    _al_u3383 (
    .a(_al_u3186_o),
    .b(_al_u3183_o),
    .c(_al_u2907_o),
    .d(_al_u2885_o),
    .o(_al_u3383_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3384 (
    .a(_al_u3382_o),
    .b(_al_u3355_o),
    .c(_al_u3383_o),
    .o(_al_u3384_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3385 (
    .a(_al_u3384_o),
    .b(_al_u3054_o),
    .o(_al_u3385_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u3386 (
    .a(_al_u3385_o),
    .b(_al_u2898_o),
    .c(_al_u3046_o),
    .o(_al_u3386_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3387 (
    .a(_al_u3386_o),
    .b(_al_u3240_o),
    .o(_al_u3387_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*A))"),
    .INIT(8'hc4))
    _al_u3388 (
    .a(_al_u3387_o),
    .b(n377_lutinv),
    .c(_al_u3113_o),
    .o(_al_u3388_o));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*~A))"),
    .INIT(8'hdc))
    _al_u3389 (
    .a(_al_u3363_o),
    .b(_al_u3388_o),
    .c(_al_u3118_o),
    .o(\sel2_b3/or_B6_or_B7_B8_o_o ));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u3390 (
    .a(n187[3]),
    .b(_al_u3057_o),
    .c(_al_u3120_o),
    .o(n193[4]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~D*~(C*A)))"),
    .INIT(16'hcc80))
    _al_u3391 (
    .a(mux16_b11_sel_is_2_o),
    .b(_al_u3295_o),
    .c(n193[4]),
    .d(_al_u3061_o),
    .o(_al_u3391_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(~B*~A))"),
    .INIT(8'h0e))
    _al_u3392 (
    .a(_al_u3391_o),
    .b(_al_u3207_o),
    .c(_al_u3245_o),
    .o(n206[4]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u3393 (
    .a(n206[4]),
    .b(_al_u3209_o),
    .c(_al_u2923_o),
    .o(_al_u3393_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u3394 (
    .a(_al_u3393_o),
    .b(_al_u2920_o),
    .c(_al_u2930_o),
    .o(n215[4]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3395 (
    .a(n215[4]),
    .b(_al_u2927_o),
    .o(n216[4]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*A)"),
    .INIT(16'h0002))
    _al_u3396 (
    .a(n216[4]),
    .b(_al_u3318_o),
    .c(_al_u3074_o),
    .d(_al_u2932_o),
    .o(_al_u3396_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~B*~(~D*~A))"),
    .INIT(16'h0302))
    _al_u3397 (
    .a(_al_u3396_o),
    .b(_al_u2940_o),
    .c(_al_u3253_o),
    .d(_al_u3319_o),
    .o(_al_u3397_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u3398 (
    .a(_al_u3134_o),
    .b(_al_u2946_o),
    .c(_al_u3397_o),
    .o(_al_u3398_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u3399 (
    .a(mux61_b3_sel_is_2_o),
    .b(_al_u2914_o),
    .c(_al_u2945_o),
    .o(mux61_b0_sel_is_2_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3400 (
    .a(_al_u3398_o),
    .b(mux61_b0_sel_is_2_o),
    .c(_al_u3327_o),
    .o(_al_u3400_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3401 (
    .a(_al_u3400_o),
    .b(_al_u2970_o),
    .c(_al_u3139_o),
    .o(_al_u3401_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u3402 (
    .a(_al_u3401_o),
    .b(_al_u3256_o),
    .c(_al_u2966_o),
    .o(_al_u3402_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*~A))"),
    .INIT(8'h8c))
    _al_u3403 (
    .a(_al_u3402_o),
    .b(mux84_b4_sel_is_2_o),
    .c(_al_u3293_o),
    .o(_al_u3403_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u3404 (
    .a(mux92_b0_sel_is_0_o),
    .b(_al_u2991_o),
    .c(_al_u3001_o),
    .o(mux94_b0_sel_is_2_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u3405 (
    .a(mux94_b0_sel_is_2_o),
    .b(_al_u2998_o),
    .c(_al_u2999_o),
    .o(mux96_b0_sel_is_2_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3406 (
    .a(mux96_b0_sel_is_2_o),
    .b(_al_u3079_o),
    .o(_al_u3406_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u3407 (
    .a(_al_u3406_o),
    .b(_al_u2982_o),
    .c(_al_u2990_o),
    .o(_al_u3407_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(B*A))"),
    .INIT(8'h07))
    _al_u3408 (
    .a(_al_u3403_o),
    .b(_al_u3407_o),
    .c(_al_u2998_o),
    .o(_al_u3408_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u3409 (
    .a(_al_u3408_o),
    .b(_al_u3005_o),
    .c(_al_u2997_o),
    .o(_al_u3409_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3410 (
    .a(_al_u2908_o),
    .b(_al_u2993_o),
    .o(_al_u3410_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u3411 (
    .a(_al_u3409_o),
    .b(_al_u3340_o),
    .c(_al_u3410_o),
    .o(_al_u3411_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3412 (
    .a(_al_u3411_o),
    .b(_al_u3007_o),
    .o(_al_u3412_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3413 (
    .a(mux120_b7_sel_is_2_o),
    .b(_al_u3087_o),
    .c(_al_u3013_o),
    .o(_al_u3413_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(~D*~(B*A)))"),
    .INIT(16'h0f08))
    _al_u3414 (
    .a(_al_u3412_o),
    .b(_al_u3413_o),
    .c(_al_u3032_o),
    .d(_al_u3156_o),
    .o(_al_u3414_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3415 (
    .a(_al_u2903_o),
    .b(_al_u3010_o),
    .o(_al_u3415_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3416 (
    .a(_al_u3414_o),
    .b(_al_u3415_o),
    .o(_al_u3416_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u3417 (
    .a(_al_u2913_o),
    .b(_al_u3026_o),
    .c(counter[0]),
    .d(counter[1]),
    .o(_al_u3417_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3418 (
    .a(_al_u3416_o),
    .b(mux137_b2_sel_is_2_o),
    .c(_al_u3417_o),
    .o(_al_u3418_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3419 (
    .a(_al_u3418_o),
    .b(_al_u3034_o),
    .o(_al_u3419_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3420 (
    .a(mux147_b3_sel_is_2_o),
    .b(mux150_b0_sel_is_2_o),
    .o(_al_u3420_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(~D*~(B*A)))"),
    .INIT(16'h0f08))
    _al_u3421 (
    .a(_al_u3419_o),
    .b(_al_u3420_o),
    .c(_al_u3359_o),
    .d(_al_u3188_o),
    .o(_al_u3421_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3422 (
    .a(_al_u3421_o),
    .b(_al_u3186_o),
    .o(_al_u3422_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~A*~(D*C)))"),
    .INIT(16'hc888))
    _al_u3423 (
    .a(_al_u2898_o),
    .b(_al_u3046_o),
    .c(_al_u2899_o),
    .d(counter[0]),
    .o(_al_u3423_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~B*~(D*~A))"),
    .INIT(16'h0203))
    _al_u3424 (
    .a(_al_u2950_o),
    .b(_al_u3235_o),
    .c(_al_u3423_o),
    .d(_al_u3046_o),
    .o(mux168_b4_sel_is_2_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3425 (
    .a(_al_u3422_o),
    .b(mux168_b4_sel_is_2_o),
    .c(_al_u3052_o),
    .o(_al_u3425_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u3426 (
    .a(mux63_b12_sel_is_2_o),
    .b(_al_u2963_o),
    .c(mux92_b7_sel_is_2_o),
    .o(_al_u3426_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3427 (
    .a(mux30_b12_sel_is_2_o),
    .b(_al_u3211_o),
    .o(_al_u3427_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D*~(~C*~B)))"),
    .INIT(16'h02aa))
    _al_u3428 (
    .a(_al_u3366_o),
    .b(_al_u2898_o),
    .c(_al_u2899_o),
    .d(_al_u2888_o),
    .o(_al_u3428_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3429 (
    .a(_al_u3428_o),
    .b(mux16_b11_sel_is_2_o),
    .c(_al_u3056_o),
    .o(_al_u3429_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3430 (
    .a(_al_u3427_o),
    .b(_al_u3429_o),
    .o(_al_u3430_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3431 (
    .a(_al_u3430_o),
    .b(_al_u2927_o),
    .o(_al_u3431_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3432 (
    .a(_al_u3426_o),
    .b(_al_u3431_o),
    .o(_al_u3432_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3433 (
    .a(_al_u3432_o),
    .b(_al_u3264_o),
    .c(_al_u3000_o),
    .o(_al_u3433_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3434 (
    .a(_al_u3433_o),
    .b(_al_u3088_o),
    .o(_al_u3434_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~B*A)*~(D)*~(C)+~(~B*A)*D*~(C)+~(~(~B*A))*D*C+~(~B*A)*D*C)"),
    .INIT(16'hfd0d))
    _al_u3435 (
    .a(_al_u3434_o),
    .b(_al_u3007_o),
    .c(_al_u3008_o),
    .d(counter[0]),
    .o(_al_u3435_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u3436 (
    .a(_al_u3435_o),
    .b(_al_u3014_o),
    .c(_al_u3010_o),
    .o(_al_u3436_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(B*~A))"),
    .INIT(8'h0b))
    _al_u3437 (
    .a(_al_u3436_o),
    .b(mux130_b1_sel_is_2_o),
    .c(_al_u3030_o),
    .o(_al_u3437_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u3438 (
    .a(_al_u3437_o),
    .b(_al_u3102_o),
    .c(_al_u3354_o),
    .o(_al_u3438_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u3439 (
    .a(_al_u3188_o),
    .b(_al_u3042_o),
    .c(_al_u3040_o),
    .o(_al_u3439_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3440 (
    .a(_al_u3438_o),
    .b(_al_u3439_o),
    .o(_al_u3440_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(~B*~A))"),
    .INIT(8'he0))
    _al_u3441 (
    .a(_al_u3440_o),
    .b(_al_u3044_o),
    .c(_al_u3196_o),
    .o(_al_u3441_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    _al_u3442 (
    .a(_al_u2887_o),
    .b(_al_u3046_o),
    .c(_al_u2891_o),
    .o(_al_u3442_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3443 (
    .a(_al_u3441_o),
    .b(_al_u3187_o),
    .c(_al_u3442_o),
    .o(_al_u3443_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u3444 (
    .a(_al_u3443_o),
    .b(_al_u3052_o),
    .c(_al_u3050_o),
    .o(_al_u3444_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B*A))"),
    .INIT(8'h70))
    _al_u3445 (
    .a(_al_u3444_o),
    .b(_al_u3117_o),
    .c(n377_lutinv),
    .o(_al_u3445_o));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    _al_u3446 (
    .a(_al_u3425_o),
    .b(_al_u3445_o),
    .c(_al_u3118_o),
    .o(\sel2_b4/or_B6_or_B7_B8_o_o ));
  AL_MAP_LUT4 #(
    .EQN("(~C*B*~(~D*~A))"),
    .INIT(16'h0c08))
    _al_u3447 (
    .a(_al_u3122_o),
    .b(mux16_b11_sel_is_2_o),
    .c(_al_u3056_o),
    .d(_al_u3308_o),
    .o(n200[0]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3448 (
    .a(n200[0]),
    .b(_al_u3124_o),
    .o(n202[0]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3449 (
    .a(_al_u2898_o),
    .b(_al_u2915_o),
    .o(_al_u3449_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u3450 (
    .a(n202[0]),
    .b(_al_u2917_o),
    .c(_al_u3449_o),
    .o(n210[0]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3451 (
    .a(n210[0]),
    .b(_al_u2922_o),
    .o(n213[0]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3452 (
    .a(n213[0]),
    .b(mux33_b0_sel_is_2_o),
    .o(n216[0]));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3453 (
    .a(n216[0]),
    .b(mux49_b0_sel_is_2_o),
    .c(_al_u2932_o),
    .o(_al_u3453_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3454 (
    .a(_al_u3453_o),
    .b(mux61_b0_sel_is_2_o),
    .o(_al_u3454_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u3455 (
    .a(_al_u3454_o),
    .b(_al_u3322_o),
    .c(_al_u2972_o),
    .o(_al_u3455_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3456 (
    .a(_al_u3455_o),
    .b(_al_u3139_o),
    .o(_al_u3456_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3457 (
    .a(_al_u3456_o),
    .b(_al_u2965_o),
    .o(_al_u3457_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u3458 (
    .a(_al_u3457_o),
    .b(_al_u3146_o),
    .c(_al_u3144_o),
    .o(_al_u3458_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3459 (
    .a(_al_u3458_o),
    .b(_al_u3292_o),
    .o(_al_u3459_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3460 (
    .a(_al_u3459_o),
    .b(_al_u3406_o),
    .c(mux87_b0_sel_is_2_o),
    .o(_al_u3460_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3461 (
    .a(_al_u3088_o),
    .b(_al_u3004_o),
    .o(mux107_b0_sel_is_2_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3462 (
    .a(_al_u3460_o),
    .b(mux107_b0_sel_is_2_o),
    .c(_al_u3005_o),
    .o(_al_u3462_o));
  AL_MAP_LUT2 #(
    .EQN("~(B@A)"),
    .INIT(4'h9))
    _al_u3463 (
    .a(_al_u3462_o),
    .b(mux111_b0_sel_is_2_o),
    .o(_al_u3463_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3464 (
    .a(_al_u3463_o),
    .b(mux120_b3_sel_is_2_o),
    .c(_al_u3017_o),
    .o(_al_u3464_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(~A*~(D*~B)))"),
    .INIT(16'h0b0a))
    _al_u3465 (
    .a(_al_u3464_o),
    .b(_al_u2935_o),
    .c(_al_u3160_o),
    .d(_al_u3010_o),
    .o(_al_u3465_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*~A)"),
    .INIT(8'h04))
    _al_u3466 (
    .a(_al_u3164_o),
    .b(mux129_b8_sel_is_2_o),
    .c(_al_u3167_o),
    .o(mux129_b0_sel_is_2_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3467 (
    .a(_al_u3465_o),
    .b(mux129_b0_sel_is_2_o),
    .o(_al_u3467_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3468 (
    .a(_al_u3227_o),
    .b(_al_u3028_o),
    .o(_al_u3468_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3469 (
    .a(mux135_b11_sel_is_0_o),
    .b(_al_u3468_o),
    .c(_al_u3102_o),
    .o(mux136_b7_sel_is_2_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3470 (
    .a(mux136_b7_sel_is_2_o),
    .b(_al_u3027_o),
    .o(mux136_b0_sel_is_2_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3471 (
    .a(_al_u2908_o),
    .b(_al_u3026_o),
    .o(_al_u3471_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u3472 (
    .a(mux136_b0_sel_is_2_o),
    .b(_al_u3171_o),
    .c(_al_u3471_o),
    .o(mux139_b0_sel_is_2_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3473 (
    .a(_al_u3467_o),
    .b(mux139_b0_sel_is_2_o),
    .c(_al_u3355_o),
    .o(_al_u3473_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(~B*~A))"),
    .INIT(8'he0))
    _al_u3474 (
    .a(_al_u2914_o),
    .b(_al_u2884_o),
    .c(_al_u2885_o),
    .o(_al_u3474_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    _al_u3475 (
    .a(_al_u3473_o),
    .b(mux152_b0_sel_is_2_o),
    .c(_al_u3474_o),
    .o(_al_u3475_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3476 (
    .a(_al_u3276_o),
    .b(_al_u3278_o),
    .o(_al_u3476_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~C*~(D*A)))"),
    .INIT(16'hc8c0))
    _al_u3477 (
    .a(_al_u3475_o),
    .b(_al_u3280_o),
    .c(_al_u3108_o),
    .d(_al_u3476_o),
    .o(_al_u3477_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3478 (
    .a(_al_u3477_o),
    .b(mux169_b0_sel_is_2_o),
    .o(_al_u3478_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3479 (
    .a(_al_u3478_o),
    .b(mux174_b0_sel_is_0_o),
    .c(n378_lutinv),
    .o(_al_u3479_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3480 (
    .a(_al_u3065_o),
    .b(_al_u3304_o),
    .o(_al_u3480_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u3481 (
    .a(_al_u3480_o),
    .b(_al_u3308_o),
    .c(_al_u3068_o),
    .o(_al_u3481_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3482 (
    .a(_al_u2938_o),
    .b(_al_u2888_o),
    .o(_al_u3482_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3483 (
    .a(_al_u3481_o),
    .b(_al_u3482_o),
    .o(_al_u3483_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(~B*~A))"),
    .INIT(8'he0))
    _al_u3484 (
    .a(_al_u2904_o),
    .b(_al_u2842_o),
    .c(_al_u2888_o),
    .o(_al_u3484_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*A*~(~D*C))"),
    .INIT(16'h2202))
    _al_u3485 (
    .a(_al_u3483_o),
    .b(_al_u2916_o),
    .c(_al_u3484_o),
    .d(counter[0]),
    .o(_al_u3485_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3486 (
    .a(_al_u3449_o),
    .b(_al_u2923_o),
    .o(_al_u3486_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*~B))"),
    .INIT(8'ha8))
    _al_u3487 (
    .a(_al_u3485_o),
    .b(_al_u3486_o),
    .c(counter[0]),
    .o(_al_u3487_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3488 (
    .a(_al_u3487_o),
    .b(_al_u2929_o),
    .c(_al_u2922_o),
    .o(_al_u3488_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3489 (
    .a(_al_u3488_o),
    .b(_al_u2933_o),
    .o(_al_u3489_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(~C*~B*A))"),
    .INIT(16'hfd00))
    _al_u3490 (
    .a(_al_u2937_o),
    .b(_al_u2938_o),
    .c(_al_u2949_o),
    .d(_al_u2926_o),
    .o(_al_u3490_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3491 (
    .a(_al_u2959_o),
    .b(_al_u3325_o),
    .o(_al_u3491_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*~A)"),
    .INIT(16'h0004))
    _al_u3492 (
    .a(_al_u2958_o),
    .b(_al_u3491_o),
    .c(_al_u2972_o),
    .d(_al_u2943_o),
    .o(_al_u3492_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    _al_u3493 (
    .a(mux47_b1_sel_is_2_o),
    .b(_al_u3492_o),
    .c(_al_u2946_o),
    .d(_al_u2947_o),
    .o(_al_u3493_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u3494 (
    .a(mux60_b1_sel_is_2_o),
    .b(_al_u3490_o),
    .c(_al_u3493_o),
    .o(_al_u3494_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*~B))"),
    .INIT(8'ha8))
    _al_u3495 (
    .a(_al_u3489_o),
    .b(_al_u2956_o),
    .c(_al_u3494_o),
    .o(_al_u3495_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u3496 (
    .a(_al_u2953_o),
    .b(_al_u2963_o),
    .o(_al_u3496_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3497 (
    .a(_al_u3496_o),
    .b(_al_u2964_o),
    .o(_al_u3497_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    _al_u3498 (
    .a(_al_u3141_o),
    .b(_al_u3497_o),
    .c(_al_u3143_o),
    .d(_al_u3322_o),
    .o(mux77_b8_sel_is_2_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(~B*~A))"),
    .INIT(8'he0))
    _al_u3499 (
    .a(_al_u2884_o),
    .b(_al_u2925_o),
    .c(_al_u2975_o),
    .o(_al_u3499_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u3500 (
    .a(_al_u3256_o),
    .b(_al_u2984_o),
    .c(_al_u3499_o),
    .o(_al_u3500_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3501 (
    .a(mux77_b8_sel_is_2_o),
    .b(_al_u3500_o),
    .o(_al_u3501_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    _al_u3502 (
    .a(_al_u3495_o),
    .b(_al_u3501_o),
    .c(_al_u3323_o),
    .o(_al_u3502_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3503 (
    .a(_al_u3502_o),
    .b(_al_u3077_o),
    .c(_al_u3079_o),
    .o(_al_u3503_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3504 (
    .a(_al_u3503_o),
    .b(_al_u2986_o),
    .o(_al_u3504_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u3505 (
    .a(_al_u3504_o),
    .b(_al_u2991_o),
    .c(_al_u3000_o),
    .o(_al_u3505_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3506 (
    .a(_al_u2994_o),
    .b(_al_u3005_o),
    .o(mux103_b1_sel_is_2_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u3507 (
    .a(_al_u3505_o),
    .b(mux103_b1_sel_is_2_o),
    .c(counter[0]),
    .o(_al_u3507_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D*~(~C*~B)))"),
    .INIT(16'h02aa))
    _al_u3508 (
    .a(_al_u3090_o),
    .b(_al_u2989_o),
    .c(_al_u2842_o),
    .d(_al_u2993_o),
    .o(_al_u3508_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3509 (
    .a(_al_u3507_o),
    .b(_al_u3508_o),
    .c(_al_u3020_o),
    .o(_al_u3509_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3510 (
    .a(_al_u3509_o),
    .b(_al_u3153_o),
    .o(_al_u3510_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3511 (
    .a(_al_u3162_o),
    .b(_al_u3156_o),
    .o(_al_u3511_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3512 (
    .a(_al_u3510_o),
    .b(_al_u3511_o),
    .c(_al_u3268_o),
    .o(_al_u3512_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3513 (
    .a(_al_u3512_o),
    .b(_al_u3028_o),
    .o(_al_u3513_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3514 (
    .a(_al_u3513_o),
    .b(_al_u3098_o),
    .o(_al_u3514_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(~B*~(~C*A)))"),
    .INIT(16'h00ce))
    _al_u3515 (
    .a(_al_u3514_o),
    .b(_al_u3034_o),
    .c(_al_u3471_o),
    .d(_al_u3193_o),
    .o(_al_u3515_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3516 (
    .a(_al_u3515_o),
    .b(_al_u3354_o),
    .o(_al_u3516_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3517 (
    .a(_al_u3176_o),
    .b(_al_u3037_o),
    .o(_al_u3517_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3518 (
    .a(_al_u3516_o),
    .b(_al_u3517_o),
    .c(_al_u3040_o),
    .o(_al_u3518_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3519 (
    .a(_al_u3108_o),
    .b(_al_u3195_o),
    .o(_al_u3519_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3520 (
    .a(_al_u3518_o),
    .b(_al_u3519_o),
    .o(_al_u3520_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u3521 (
    .a(_al_u3520_o),
    .b(_al_u3184_o),
    .c(_al_u3182_o),
    .o(_al_u3521_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3522 (
    .a(_al_u3521_o),
    .b(_al_u3362_o),
    .o(_al_u3522_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u3523 (
    .a(_al_u3522_o),
    .b(_al_u3052_o),
    .c(_al_u3423_o),
    .o(_al_u3523_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3524 (
    .a(_al_u3523_o),
    .b(_al_u3111_o),
    .o(_al_u3524_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3525 (
    .a(_al_u3113_o),
    .b(state_next[1]),
    .o(_al_u3525_o));
  AL_MAP_LUT4 #(
    .EQN("~(~A*~(C*~(D*B)))"),
    .INIT(16'hbafa))
    _al_u3526 (
    .a(_al_u3479_o),
    .b(_al_u3524_o),
    .c(_al_u2860_o),
    .d(_al_u3525_o),
    .o(\sel2_b0/or_or_B4_B5_o_or_B6__o ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    _al_u3527 (
    .a(_al_u2902_o),
    .b(mux16_b11_sel_is_2_o),
    .c(_al_u2906_o),
    .o(n200[5]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3528 (
    .a(n200[5]),
    .b(mux19_b2_sel_is_0_o),
    .o(n203[5]));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u3529 (
    .a(n203[5]),
    .b(_al_u3286_o),
    .c(_al_u3207_o),
    .o(n208[5]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*B))"),
    .INIT(8'ha2))
    _al_u3530 (
    .a(n208[5]),
    .b(_al_u2923_o),
    .c(counter[1]),
    .o(_al_u3530_o));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~((~C*~A))*~(B)+~D*(~C*~A)*~(B)+~(~D)*(~C*~A)*B+~D*(~C*~A)*B)"),
    .INIT(16'hfbc8))
    _al_u3531 (
    .a(_al_u3530_o),
    .b(mux38_b1_sel_is_2_o),
    .c(_al_u3316_o),
    .d(_al_u2949_o),
    .o(n221[5]));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u3532 (
    .a(n221[5]),
    .b(_al_u2939_o),
    .c(_al_u2945_o),
    .o(_al_u3532_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3533 (
    .a(_al_u3532_o),
    .b(_al_u2972_o),
    .o(_al_u3533_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3534 (
    .a(_al_u3533_o),
    .b(mux70_b2_sel_is_0_o),
    .c(mux75_b5_sel_is_2_o),
    .o(_al_u3534_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3535 (
    .a(_al_u3534_o),
    .b(_al_u3292_o),
    .o(_al_u3535_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3536 (
    .a(_al_u3535_o),
    .b(mux85_b0_sel_is_2_o),
    .o(_al_u3536_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3537 (
    .a(_al_u3536_o),
    .b(mux97_b5_sel_is_2_o),
    .o(_al_u3537_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3538 (
    .a(_al_u3537_o),
    .b(_al_u3219_o),
    .c(_al_u3340_o),
    .o(_al_u3538_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*B))"),
    .INIT(8'ha2))
    _al_u3539 (
    .a(_al_u3538_o),
    .b(_al_u3220_o),
    .c(counter[0]),
    .o(_al_u3539_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3540 (
    .a(_al_u3539_o),
    .b(mux111_b0_sel_is_2_o),
    .c(_al_u3088_o),
    .o(_al_u3540_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3541 (
    .a(_al_u3008_o),
    .b(counter[0]),
    .o(_al_u3541_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3542 (
    .a(_al_u3540_o),
    .b(_al_u3541_o),
    .o(_al_u3542_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3543 (
    .a(_al_u3020_o),
    .b(_al_u3158_o),
    .o(mux117_b5_sel_is_2_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    _al_u3544 (
    .a(mux117_b5_sel_is_2_o),
    .b(mux119_b3_sel_is_0_o),
    .c(_al_u3155_o),
    .d(_al_u3415_o),
    .o(mux127_b5_sel_is_2_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u3545 (
    .a(_al_u3542_o),
    .b(mux127_b5_sel_is_2_o),
    .o(_al_u3545_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3546 (
    .a(_al_u3545_o),
    .b(_al_u3417_o),
    .o(_al_u3546_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3547 (
    .a(_al_u3546_o),
    .b(mux137_b5_sel_is_2_o),
    .o(_al_u3547_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3548 (
    .a(_al_u3547_o),
    .b(mux147_b3_sel_is_2_o),
    .c(_al_u3197_o),
    .o(_al_u3548_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u3549 (
    .a(_al_u3548_o),
    .b(_al_u3235_o),
    .c(_al_u3423_o),
    .o(_al_u3549_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u3550 (
    .a(_al_u3549_o),
    .b(_al_u3046_o),
    .c(_al_u2908_o),
    .o(_al_u3550_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3551 (
    .a(_al_u2889_o),
    .b(_al_u3066_o),
    .o(_al_u3551_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3552 (
    .a(_al_u3427_o),
    .b(_al_u3551_o),
    .o(_al_u3552_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u3553 (
    .a(_al_u3552_o),
    .b(_al_u2932_o),
    .c(_al_u2927_o),
    .o(_al_u3553_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3554 (
    .a(_al_u3553_o),
    .b(_al_u3081_o),
    .o(_al_u3554_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*~B))"),
    .INIT(8'h8a))
    _al_u3555 (
    .a(_al_u3554_o),
    .b(_al_u2951_o),
    .c(_al_u2993_o),
    .o(_al_u3555_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3556 (
    .a(_al_u3555_o),
    .b(_al_u3090_o),
    .c(_al_u3008_o),
    .o(_al_u3556_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(~B*~A))"),
    .INIT(8'he0))
    _al_u3557 (
    .a(_al_u2914_o),
    .b(_al_u2891_o),
    .c(_al_u3010_o),
    .o(_al_u3557_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3558 (
    .a(_al_u3556_o),
    .b(_al_u3557_o),
    .o(_al_u3558_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*A)"),
    .INIT(16'h0080))
    _al_u3559 (
    .a(_al_u3558_o),
    .b(_al_u3031_o),
    .c(_al_u3095_o),
    .d(_al_u3165_o),
    .o(_al_u3559_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3560 (
    .a(_al_u3559_o),
    .b(_al_u3098_o),
    .o(_al_u3560_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3561 (
    .a(_al_u3171_o),
    .b(_al_u3174_o),
    .o(mux140_b11_sel_is_2_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3562 (
    .a(_al_u3560_o),
    .b(mux140_b11_sel_is_2_o),
    .o(_al_u3562_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3563 (
    .a(_al_u3562_o),
    .b(_al_u3439_o),
    .c(_al_u3276_o),
    .o(_al_u3563_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3564 (
    .a(_al_u3563_o),
    .b(_al_u3187_o),
    .c(_al_u3054_o),
    .o(_al_u3564_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3565 (
    .a(_al_u3564_o),
    .b(_al_u3240_o),
    .o(_al_u3565_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*A))"),
    .INIT(8'hc4))
    _al_u3566 (
    .a(_al_u3565_o),
    .b(n377_lutinv),
    .c(_al_u3113_o),
    .o(_al_u3566_o));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~B*~(C*A))"),
    .INIT(16'hffec))
    _al_u3567 (
    .a(_al_u3550_o),
    .b(_al_u3566_o),
    .c(_al_u3118_o),
    .d(n376_lutinv),
    .o(\sel2_b5/or_B6_or_B7_B8_o_o ));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B)*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0eaa))
    _al_u3568 (
    .a(_al_u3121_o),
    .b(_al_u2898_o),
    .c(_al_u2899_o),
    .d(_al_u2888_o),
    .o(n193[1]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u3569 (
    .a(n193[1]),
    .b(mux14_b11_sel_is_2_o),
    .c(_al_u3061_o),
    .o(n197[1]));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*A)"),
    .INIT(16'h0080))
    _al_u3570 (
    .a(n197[1]),
    .b(mux19_b2_sel_is_0_o),
    .c(mux16_b1_sel_is_0_o),
    .d(_al_u3204_o),
    .o(_al_u3570_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(~B*~A))"),
    .INIT(8'h0e))
    _al_u3571 (
    .a(_al_u3570_o),
    .b(_al_u2916_o),
    .c(_al_u2917_o),
    .o(n205[1]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~C*~(D*A)))"),
    .INIT(16'hc8c0))
    _al_u3572 (
    .a(n205[1]),
    .b(mux30_b1_sel_is_2_o),
    .c(_al_u3287_o),
    .d(_al_u3486_o),
    .o(n214[1]));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3573 (
    .a(n214[1]),
    .b(mux38_b1_sel_is_2_o),
    .c(_al_u3318_o),
    .o(n225[1]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3574 (
    .a(n225[1]),
    .b(_al_u3252_o),
    .o(_al_u3574_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3575 (
    .a(_al_u3574_o),
    .b(mux68_b1_sel_is_2_o),
    .o(_al_u3575_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u3576 (
    .a(_al_u3575_o),
    .b(_al_u2949_o),
    .c(_al_u2963_o),
    .o(_al_u3576_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u3577 (
    .a(_al_u3143_o),
    .b(_al_u3256_o),
    .c(counter[0]),
    .o(_al_u3577_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3578 (
    .a(_al_u3576_o),
    .b(_al_u3577_o),
    .c(_al_u3146_o),
    .o(_al_u3578_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3579 (
    .a(_al_u3578_o),
    .b(_al_u2984_o),
    .o(_al_u3579_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3580 (
    .a(_al_u3579_o),
    .b(mux89_b1_sel_is_2_o),
    .c(_al_u3336_o),
    .o(_al_u3580_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3581 (
    .a(_al_u3580_o),
    .b(mux94_b0_sel_is_2_o),
    .o(_al_u3581_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3582 (
    .a(_al_u3581_o),
    .b(mux103_b1_sel_is_2_o),
    .c(_al_u2998_o),
    .o(_al_u3582_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3583 (
    .a(_al_u3582_o),
    .b(mux107_b0_sel_is_2_o),
    .o(_al_u3583_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3584 (
    .a(_al_u3583_o),
    .b(mux111_b0_sel_is_2_o),
    .c(_al_u3015_o),
    .o(_al_u3584_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3585 (
    .a(_al_u3584_o),
    .b(_al_u3557_o),
    .o(_al_u3585_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3586 (
    .a(_al_u3585_o),
    .b(mux124_b11_sel_is_2_o),
    .c(_al_u3153_o),
    .o(_al_u3586_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u3587 (
    .a(_al_u3468_o),
    .b(_al_u3027_o),
    .c(_al_u3099_o),
    .o(mux134_b0_sel_is_2_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3588 (
    .a(mux134_b0_sel_is_2_o),
    .b(mux130_b1_sel_is_2_o),
    .o(_al_u3588_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(B*~(~D*~A)))"),
    .INIT(16'h0307))
    _al_u3589 (
    .a(_al_u3586_o),
    .b(_al_u3588_o),
    .c(_al_u3099_o),
    .d(_al_u3345_o),
    .o(_al_u3589_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    _al_u3590 (
    .a(_al_u3589_o),
    .b(mux136_b1_sel_is_0_o),
    .c(mux141_b1_sel_is_2_o),
    .o(_al_u3590_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u3591 (
    .a(_al_u3590_o),
    .b(_al_u3355_o),
    .c(_al_u3176_o),
    .o(_al_u3591_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u3592 (
    .a(_al_u3591_o),
    .b(_al_u3191_o),
    .c(_al_u3189_o),
    .o(_al_u3592_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3593 (
    .a(_al_u3592_o),
    .b(_al_u3278_o),
    .o(_al_u3593_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u3594 (
    .a(_al_u3280_o),
    .b(_al_u3049_o),
    .c(_al_u3362_o),
    .o(_al_u3594_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u3595 (
    .a(_al_u3052_o),
    .b(_al_u3050_o),
    .c(counter[0]),
    .o(_al_u3595_o));
  AL_MAP_LUT4 #(
    .EQN("~(D*~((C*A))*~(B)+D*(C*A)*~(B)+~(D)*(C*A)*B+D*(C*A)*B)"),
    .INIT(16'h4c7f))
    _al_u3596 (
    .a(_al_u3593_o),
    .b(_al_u3594_o),
    .c(_al_u3595_o),
    .d(_al_u2898_o),
    .o(_al_u3596_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3597 (
    .a(_al_u2906_o),
    .b(_al_u3120_o),
    .o(mux12_b9_sel_is_2_o_neg_lutinv));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*B))"),
    .INIT(8'ha2))
    _al_u3598 (
    .a(mux16_b1_sel_is_0_o),
    .b(mux12_b9_sel_is_2_o_neg_lutinv),
    .c(_al_u3484_o),
    .o(_al_u3598_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u3599 (
    .a(_al_u3598_o),
    .b(_al_u3245_o),
    .c(_al_u3204_o),
    .o(_al_u3599_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    _al_u3600 (
    .a(_al_u2920_o),
    .b(_al_u3316_o),
    .c(_al_u3599_o),
    .o(_al_u3600_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3601 (
    .a(_al_u3600_o),
    .b(mux33_b0_sel_is_2_o),
    .c(_al_u3071_o),
    .o(_al_u3601_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3602 (
    .a(_al_u3601_o),
    .b(_al_u3494_o),
    .o(_al_u3602_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    _al_u3603 (
    .a(_al_u2997_o),
    .b(_al_u2999_o),
    .c(_al_u3602_o),
    .o(_al_u3603_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3604 (
    .a(_al_u3603_o),
    .b(_al_u2994_o),
    .o(_al_u3604_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*~B))"),
    .INIT(8'h8a))
    _al_u3605 (
    .a(_al_u3264_o),
    .b(_al_u2950_o),
    .c(_al_u2993_o),
    .o(mux104_b11_sel_is_2_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3606 (
    .a(_al_u3604_o),
    .b(mux104_b11_sel_is_2_o),
    .o(_al_u3606_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3607 (
    .a(_al_u3606_o),
    .b(_al_u3007_o),
    .o(_al_u3607_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3608 (
    .a(_al_u3607_o),
    .b(mux117_b5_sel_is_2_o),
    .c(_al_u3011_o),
    .o(_al_u3608_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3609 (
    .a(_al_u3608_o),
    .b(_al_u3155_o),
    .o(_al_u3609_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*C)*~(B*~A))"),
    .INIT(16'h0bbb))
    _al_u3610 (
    .a(_al_u3609_o),
    .b(mux124_b0_sel_is_0_o),
    .c(_al_u2904_o),
    .d(_al_u3010_o),
    .o(_al_u3610_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u3611 (
    .a(_al_u3027_o),
    .b(_al_u3610_o),
    .o(_al_u3611_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3612 (
    .a(_al_u3611_o),
    .b(mux135_b11_sel_is_0_o),
    .c(_al_u3101_o),
    .o(_al_u3612_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*~A))"),
    .INIT(8'h32))
    _al_u3613 (
    .a(_al_u3612_o),
    .b(_al_u3104_o),
    .c(_al_u3102_o),
    .o(_al_u3613_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u3614 (
    .a(_al_u3613_o),
    .b(_al_u2884_o),
    .c(_al_u2885_o),
    .o(_al_u3614_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3615 (
    .a(_al_u3614_o),
    .b(mux150_b0_sel_is_2_o),
    .o(_al_u3615_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u3616 (
    .a(_al_u3615_o),
    .b(_al_u3040_o),
    .c(_al_u3044_o),
    .o(_al_u3616_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3617 (
    .a(_al_u3185_o),
    .b(_al_u3278_o),
    .o(_al_u3617_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3618 (
    .a(_al_u3616_o),
    .b(_al_u3617_o),
    .o(_al_u3618_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3619 (
    .a(_al_u3618_o),
    .b(_al_u3362_o),
    .o(_al_u3619_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u3620 (
    .a(_al_u3619_o),
    .b(_al_u3046_o),
    .c(_al_u2908_o),
    .o(_al_u3620_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B*A))"),
    .INIT(8'h70))
    _al_u3621 (
    .a(_al_u3620_o),
    .b(_al_u3117_o),
    .c(n377_lutinv),
    .o(_al_u3621_o));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*~A))"),
    .INIT(8'hdc))
    _al_u3622 (
    .a(_al_u3596_o),
    .b(_al_u3621_o),
    .c(_al_u3118_o),
    .o(\sel2_b1/or_B6_or_B7_B8_o_o ));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add0/u0  (
    .a(divider2[0]),
    .b(1'b1),
    .c(\add0/c0 ),
    .o({\add0/c1 ,n0[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add0/u1  (
    .a(divider2[1]),
    .b(1'b0),
    .c(\add0/c1 ),
    .o({\add0/c2 ,n0[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add0/u2  (
    .a(divider2[2]),
    .b(1'b0),
    .c(\add0/c2 ),
    .o({\add0/c3 ,n0[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add0/u3  (
    .a(divider2[3]),
    .b(1'b0),
    .c(\add0/c3 ),
    .o({\add0/c4 ,n0[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add0/u4  (
    .a(divider2[4]),
    .b(1'b0),
    .c(\add0/c4 ),
    .o({\add0/c5 ,n0[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add0/u5  (
    .a(divider2[5]),
    .b(1'b0),
    .c(\add0/c5 ),
    .o({\add0/c6 ,n0[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add0/u6  (
    .a(divider2[6]),
    .b(1'b0),
    .c(\add0/c6 ),
    .o({\add0/c7 ,n0[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add0/u7  (
    .a(divider2[7]),
    .b(1'b0),
    .c(\add0/c7 ),
    .o({\add0/c8 ,n0[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add0/u8  (
    .a(divider2[8]),
    .b(1'b0),
    .c(\add0/c8 ),
    .o({open_n0,n0[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \add0/ucin  (
    .a(1'b0),
    .o({\add0/c0 ,open_n3}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add1/u0  (
    .a(cnt[0]),
    .b(1'b1),
    .c(\add1/c0 ),
    .o({\add1/c1 ,n372[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add1/u1  (
    .a(cnt[1]),
    .b(1'b0),
    .c(\add1/c1 ),
    .o({\add1/c2 ,n372[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add1/u2  (
    .a(cnt[2]),
    .b(1'b0),
    .c(\add1/c2 ),
    .o({\add1/c3 ,n372[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add1/u3  (
    .a(cnt[3]),
    .b(1'b0),
    .c(\add1/c3 ),
    .o({\add1/c4 ,n372[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add1/u4  (
    .a(cnt[4]),
    .b(1'b0),
    .c(\add1/c4 ),
    .o({\add1/c5 ,n372[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add1/u5  (
    .a(cnt[5]),
    .b(1'b0),
    .c(\add1/c5 ),
    .o({\add1/c6 ,n372[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add1/u6  (
    .a(cnt[6]),
    .b(1'b0),
    .c(\add1/c6 ),
    .o({\add1/c7 ,n372[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add1/u7  (
    .a(cnt[7]),
    .b(1'b0),
    .c(\add1/c7 ),
    .o({open_n4,n372[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \add1/ucin  (
    .a(1'b0),
    .o({\add1/c0 ,open_n7}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add2/u0  (
    .a(counter[0]),
    .b(1'b1),
    .c(\add2/c0 ),
    .o({\add2/c1 ,n373[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add2/u1  (
    .a(counter[1]),
    .b(1'b0),
    .c(\add2/c1 ),
    .o({\add2/c2 ,n373[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add2/u2  (
    .a(counter[2]),
    .b(1'b0),
    .c(\add2/c2 ),
    .o({\add2/c3 ,n373[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add2/u3  (
    .a(counter[3]),
    .b(1'b0),
    .c(\add2/c3 ),
    .o({\add2/c4 ,n373[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add2/u4  (
    .a(counter[4]),
    .b(1'b0),
    .c(\add2/c4 ),
    .o({\add2/c5 ,n373[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add2/u5  (
    .a(counter[5]),
    .b(1'b0),
    .c(\add2/c5 ),
    .o({\add2/c6 ,n373[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add2/u6  (
    .a(counter[6]),
    .b(1'b0),
    .c(\add2/c6 ),
    .o({\add2/c7 ,n373[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add2/u7  (
    .a(counter[7]),
    .b(1'b0),
    .c(\add2/c7 ),
    .o({open_n8,n373[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \add2/ucin  (
    .a(1'b0),
    .o({\add2/c0 ,open_n11}));
  reg_sr_as_w1 bus_write_reg (
    .clk(divider2[8]),
    .d(n366),
    .en(1'b1),
    .reset(~reset_n),
    .set(1'b0),
    .q(bus_write));  // sources/rtl/camera_init.v(434)
  i2c_module i2c_write_module (
    .address({1'b0,reg_address[1:0]}),
    .clk(clk),
    .reset_n(reset_n),
    .sda_in(sda_in),
    .write(bus_write),
    .writedata(data_in_bus),
    .ready(ready_out),
    .scl_out(scl),
    .sda(sda),
    .sda_oe(sda_oe),
    .success_out(success_out));  // sources/rtl/camera_init.v(38)
  reg_ar_as_w1 ready_reg (
    .clk(clk),
    .d(n383),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(ready));  // sources/rtl/camera_init.v(271)
  reg_ar_ss_w1 reg0_b0 (
    .clk(divider2[8]),
    .d(n369[0]),
    .en(1'b1),
    .reset(1'b0),
    .set(~reset_n),
    .q(state_next[0]));  // sources/rtl/camera_init.v(347)
  reg_ar_ss_w1 reg0_b1 (
    .clk(divider2[8]),
    .d(n369[1]),
    .en(1'b1),
    .reset(1'b0),
    .set(~reset_n),
    .q(state_next[1]));  // sources/rtl/camera_init.v(347)
  reg_sr_as_w1 reg0_b2 (
    .clk(divider2[8]),
    .d(n369[2]),
    .en(1'b1),
    .reset(~reset_n),
    .set(1'b0),
    .q(state_next[2]));  // sources/rtl/camera_init.v(347)
  reg_ar_ss_w1 reg0_b3 (
    .clk(divider2[8]),
    .d(n369[3]),
    .en(1'b1),
    .reset(1'b0),
    .set(~reset_n),
    .q(state_next[3]));  // sources/rtl/camera_init.v(347)
  reg_sr_as_w1 reg0_b4 (
    .clk(divider2[8]),
    .d(n369[4]),
    .en(1'b1),
    .reset(~reset_n),
    .set(1'b0),
    .q(state_next[4]));  // sources/rtl/camera_init.v(347)
  reg_sr_as_w1 reg0_b5 (
    .clk(divider2[8]),
    .d(n369[5]),
    .en(1'b1),
    .reset(~reset_n),
    .set(1'b0),
    .q(n369[5]));  // sources/rtl/camera_init.v(347)
  reg_sr_as_w1 reg0_b6 (
    .clk(divider2[8]),
    .d(n369[6]),
    .en(1'b1),
    .reset(~reset_n),
    .set(1'b0),
    .q(n369[6]));  // sources/rtl/camera_init.v(347)
  reg_sr_as_w1 reg0_b7 (
    .clk(divider2[8]),
    .d(n369[7]),
    .en(1'b1),
    .reset(~reset_n),
    .set(1'b0),
    .q(n369[7]));  // sources/rtl/camera_init.v(347)
  reg_sr_as_w1 reg1_b0 (
    .clk(divider2[8]),
    .d(1'b1),
    .en(1'b1),
    .reset(~mux182_b0_sel_is_2_o),
    .set(1'b0),
    .q(reg_address[0]));  // sources/rtl/camera_init.v(434)
  reg_sr_as_w1 reg1_b1 (
    .clk(divider2[8]),
    .d(1'b1),
    .en(1'b1),
    .reset(~mux182_b1_sel_is_2_o),
    .set(1'b0),
    .q(reg_address[1]));  // sources/rtl/camera_init.v(434)
  reg_sr_as_w1 reg2_b0 (
    .clk(divider2[8]),
    .d(\sel2_b0/or_or_B4_B5_o_or_B6__o ),
    .en(1'b1),
    .reset(~reset_n),
    .set(1'b0),
    .q(data_in_bus[0]));  // sources/rtl/camera_init.v(434)
  reg_sr_as_w1 reg2_b1 (
    .clk(divider2[8]),
    .d(\sel2_b1/or_B6_or_B7_B8_o_o ),
    .en(1'b1),
    .reset(~reset_n),
    .set(1'b0),
    .q(data_in_bus[1]));  // sources/rtl/camera_init.v(434)
  reg_sr_as_w1 reg2_b2 (
    .clk(divider2[8]),
    .d(\sel2_b2/or_B6_or_B7_B8_o_o ),
    .en(1'b1),
    .reset(~reset_n),
    .set(1'b0),
    .q(data_in_bus[2]));  // sources/rtl/camera_init.v(434)
  reg_sr_as_w1 reg2_b3 (
    .clk(divider2[8]),
    .d(\sel2_b3/or_B6_or_B7_B8_o_o ),
    .en(1'b1),
    .reset(~reset_n),
    .set(1'b0),
    .q(data_in_bus[3]));  // sources/rtl/camera_init.v(434)
  reg_sr_as_w1 reg2_b4 (
    .clk(divider2[8]),
    .d(\sel2_b4/or_B6_or_B7_B8_o_o ),
    .en(1'b1),
    .reset(~reset_n),
    .set(1'b0),
    .q(data_in_bus[4]));  // sources/rtl/camera_init.v(434)
  reg_sr_as_w1 reg2_b5 (
    .clk(divider2[8]),
    .d(\sel2_b5/or_B6_or_B7_B8_o_o ),
    .en(1'b1),
    .reset(~reset_n),
    .set(1'b0),
    .q(data_in_bus[5]));  // sources/rtl/camera_init.v(434)
  reg_sr_as_w1 reg2_b6 (
    .clk(divider2[8]),
    .d(\sel2_b6/or_B6_or_B7_B8_o_o ),
    .en(1'b1),
    .reset(~reset_n),
    .set(1'b0),
    .q(data_in_bus[6]));  // sources/rtl/camera_init.v(434)
  reg_sr_as_w1 reg2_b7 (
    .clk(divider2[8]),
    .d(\sel2_b7/or_B6_or_B7_B8_o_o ),
    .en(1'b1),
    .reset(~reset_n),
    .set(1'b0),
    .q(data_in_bus[7]));  // sources/rtl/camera_init.v(434)
  reg_sr_as_w1 reg3_b0 (
    .clk(divider2[8]),
    .d(n375[0]),
    .en(n381),
    .reset(~reset_n),
    .set(1'b0),
    .q(counter[0]));  // sources/rtl/camera_init.v(434)
  reg_sr_as_w1 reg3_b1 (
    .clk(divider2[8]),
    .d(n375[1]),
    .en(n381),
    .reset(~reset_n),
    .set(1'b0),
    .q(counter[1]));  // sources/rtl/camera_init.v(434)
  reg_sr_as_w1 reg3_b2 (
    .clk(divider2[8]),
    .d(n375[2]),
    .en(n381),
    .reset(~reset_n),
    .set(1'b0),
    .q(counter[2]));  // sources/rtl/camera_init.v(434)
  reg_sr_as_w1 reg3_b3 (
    .clk(divider2[8]),
    .d(n375[3]),
    .en(n381),
    .reset(~reset_n),
    .set(1'b0),
    .q(counter[3]));  // sources/rtl/camera_init.v(434)
  reg_sr_as_w1 reg3_b4 (
    .clk(divider2[8]),
    .d(n375[4]),
    .en(n381),
    .reset(~reset_n),
    .set(1'b0),
    .q(counter[4]));  // sources/rtl/camera_init.v(434)
  reg_sr_as_w1 reg3_b5 (
    .clk(divider2[8]),
    .d(n375[5]),
    .en(n381),
    .reset(~reset_n),
    .set(1'b0),
    .q(counter[5]));  // sources/rtl/camera_init.v(434)
  reg_sr_as_w1 reg3_b6 (
    .clk(divider2[8]),
    .d(n375[6]),
    .en(n381),
    .reset(~reset_n),
    .set(1'b0),
    .q(counter[6]));  // sources/rtl/camera_init.v(434)
  reg_sr_as_w1 reg3_b7 (
    .clk(divider2[8]),
    .d(n375[7]),
    .en(n381),
    .reset(~reset_n),
    .set(1'b0),
    .q(counter[7]));  // sources/rtl/camera_init.v(434)
  reg_ar_as_w1 reg4_b0 (
    .clk(divider2[8]),
    .d(n372[0]),
    .en(mux185_b0_sel_is_2_o),
    .reset(1'b0),
    .set(1'b0),
    .q(cnt[0]));  // sources/rtl/camera_init.v(434)
  reg_ar_as_w1 reg4_b1 (
    .clk(divider2[8]),
    .d(n372[1]),
    .en(mux185_b0_sel_is_2_o),
    .reset(1'b0),
    .set(1'b0),
    .q(cnt[1]));  // sources/rtl/camera_init.v(434)
  reg_ar_as_w1 reg4_b2 (
    .clk(divider2[8]),
    .d(n372[2]),
    .en(mux185_b0_sel_is_2_o),
    .reset(1'b0),
    .set(1'b0),
    .q(cnt[2]));  // sources/rtl/camera_init.v(434)
  reg_ar_as_w1 reg4_b3 (
    .clk(divider2[8]),
    .d(n372[3]),
    .en(mux185_b0_sel_is_2_o),
    .reset(1'b0),
    .set(1'b0),
    .q(cnt[3]));  // sources/rtl/camera_init.v(434)
  reg_ar_as_w1 reg4_b4 (
    .clk(divider2[8]),
    .d(n372[4]),
    .en(mux185_b0_sel_is_2_o),
    .reset(1'b0),
    .set(1'b0),
    .q(cnt[4]));  // sources/rtl/camera_init.v(434)
  reg_ar_as_w1 reg4_b5 (
    .clk(divider2[8]),
    .d(n372[5]),
    .en(mux185_b0_sel_is_2_o),
    .reset(1'b0),
    .set(1'b0),
    .q(cnt[5]));  // sources/rtl/camera_init.v(434)
  reg_ar_as_w1 reg4_b6 (
    .clk(divider2[8]),
    .d(n372[6]),
    .en(mux185_b0_sel_is_2_o),
    .reset(1'b0),
    .set(1'b0),
    .q(cnt[6]));  // sources/rtl/camera_init.v(434)
  reg_ar_as_w1 reg4_b7 (
    .clk(divider2[8]),
    .d(n372[7]),
    .en(mux185_b0_sel_is_2_o),
    .reset(1'b0),
    .set(1'b0),
    .q(cnt[7]));  // sources/rtl/camera_init.v(434)
  reg_ar_as_w1 reg5_b0 (
    .clk(clk),
    .d(n0[0]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(divider2[0]));  // sources/rtl/camera_init.v(57)
  reg_ar_as_w1 reg5_b1 (
    .clk(clk),
    .d(n0[1]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(divider2[1]));  // sources/rtl/camera_init.v(57)
  reg_ar_as_w1 reg5_b2 (
    .clk(clk),
    .d(n0[2]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(divider2[2]));  // sources/rtl/camera_init.v(57)
  reg_ar_as_w1 reg5_b3 (
    .clk(clk),
    .d(n0[3]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(divider2[3]));  // sources/rtl/camera_init.v(57)
  reg_ar_as_w1 reg5_b4 (
    .clk(clk),
    .d(n0[4]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(divider2[4]));  // sources/rtl/camera_init.v(57)
  reg_ar_as_w1 reg5_b5 (
    .clk(clk),
    .d(n0[5]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(divider2[5]));  // sources/rtl/camera_init.v(57)
  reg_ar_as_w1 reg5_b6 (
    .clk(clk),
    .d(n0[6]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(divider2[6]));  // sources/rtl/camera_init.v(57)
  reg_ar_as_w1 reg5_b7 (
    .clk(clk),
    .d(n0[7]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(divider2[7]));  // sources/rtl/camera_init.v(57)
  reg_ar_as_w1 reg5_b8 (
    .clk(clk),
    .d(n0[8]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(divider2[8]));  // sources/rtl/camera_init.v(57)

endmodule 

module lcd_sync  // sources/rtl/lcd_sync.v(2)
  (
  clk,
  rest_n,
  addr,
  hsync_cnt,
  img_ack,
  lcd_clk,
  lcd_de,
  lcd_hsync,
  lcd_pwm,
  lcd_vsync,
  vsync_cnt
  );

  input clk;  // sources/rtl/lcd_sync.v(11)
  input rest_n;  // sources/rtl/lcd_sync.v(12)
  output [15:0] addr;  // sources/rtl/lcd_sync.v(21)
  output [10:0] hsync_cnt;  // sources/rtl/lcd_sync.v(18)
  output img_ack;  // sources/rtl/lcd_sync.v(20)
  output lcd_clk;  // sources/rtl/lcd_sync.v(13)
  output lcd_de;  // sources/rtl/lcd_sync.v(17)
  output lcd_hsync;  // sources/rtl/lcd_sync.v(15)
  output lcd_pwm;  // sources/rtl/lcd_sync.v(14)
  output lcd_vsync;  // sources/rtl/lcd_sync.v(16)
  output [10:0] vsync_cnt;  // sources/rtl/lcd_sync.v(19)

  parameter IMG_H = 164;
  parameter IMG_W = 200;
  parameter IMG_X = 0;
  parameter IMG_Y = 0;
  // localparam TH = 800;
  // localparam THB = 160;
  // localparam TV = 525;
  // localparam TVB = 45;
  // localparam VGA_H = 640;
  // localparam VGA_V = 480;
  wire [10:0] n2;
  wire [11:0] n22;
  wire [39:0] n29;
  wire [10:0] n3;
  wire [15:0] n31;
  wire [10:0] n4;
  wire [12:0] n6;
  wire [6:0] n7;
  wire _al_u41_o;
  wire _al_u42_o;
  wire _al_u43_o;
  wire _al_u45_o;
  wire _al_u46_o;
  wire _al_u47_o;
  wire \add0/c0 ;
  wire \add0/c1 ;
  wire \add0/c10 ;
  wire \add0/c2 ;
  wire \add0/c3 ;
  wire \add0/c4 ;
  wire \add0/c5 ;
  wire \add0/c6 ;
  wire \add0/c7 ;
  wire \add0/c8 ;
  wire \add0/c9 ;
  wire \add1/c0 ;
  wire \add1/c1 ;
  wire \add1/c10 ;
  wire \add1/c2 ;
  wire \add1/c3 ;
  wire \add1/c4 ;
  wire \add1/c5 ;
  wire \add1/c6 ;
  wire \add1/c7 ;
  wire \add1/c8 ;
  wire \add1/c9 ;
  wire lt0_c0;
  wire lt0_c1;
  wire lt0_c10;
  wire lt0_c11;
  wire lt0_c2;
  wire lt0_c3;
  wire lt0_c4;
  wire lt0_c5;
  wire lt0_c6;
  wire lt0_c7;
  wire lt0_c8;
  wire lt0_c9;
  wire lt1_c0;
  wire lt1_c1;
  wire lt1_c10;
  wire lt1_c11;
  wire lt1_c2;
  wire lt1_c3;
  wire lt1_c4;
  wire lt1_c5;
  wire lt1_c6;
  wire lt1_c7;
  wire lt1_c8;
  wire lt1_c9;
  wire lt2_c0;
  wire lt2_c1;
  wire lt2_c10;
  wire lt2_c11;
  wire lt2_c2;
  wire lt2_c3;
  wire lt2_c4;
  wire lt2_c5;
  wire lt2_c6;
  wire lt2_c7;
  wire lt2_c8;
  wire lt2_c9;
  wire lt3_c0;
  wire lt3_c1;
  wire lt3_c10;
  wire lt3_c11;
  wire lt3_c2;
  wire lt3_c3;
  wire lt3_c4;
  wire lt3_c5;
  wire lt3_c6;
  wire lt3_c7;
  wire lt3_c8;
  wire lt3_c9;
  wire lt4_c0;
  wire lt4_c1;
  wire lt4_c10;
  wire lt4_c11;
  wire lt4_c2;
  wire lt4_c3;
  wire lt4_c4;
  wire lt4_c5;
  wire lt4_c6;
  wire lt4_c7;
  wire lt4_c8;
  wire lt4_c9;
  wire lt5_c0;
  wire lt5_c1;
  wire lt5_c10;
  wire lt5_c11;
  wire lt5_c2;
  wire lt5_c3;
  wire lt5_c4;
  wire lt5_c5;
  wire lt5_c6;
  wire lt5_c7;
  wire lt5_c8;
  wire lt5_c9;
  wire lt6_c0;
  wire lt6_c1;
  wire lt6_c10;
  wire lt6_c11;
  wire lt6_c2;
  wire lt6_c3;
  wire lt6_c4;
  wire lt6_c5;
  wire lt6_c6;
  wire lt6_c7;
  wire lt6_c8;
  wire lt6_c9;
  wire lt7_c0;
  wire lt7_c1;
  wire lt7_c10;
  wire lt7_c11;
  wire lt7_c2;
  wire lt7_c3;
  wire lt7_c4;
  wire lt7_c5;
  wire lt7_c6;
  wire lt7_c7;
  wire lt7_c8;
  wire lt7_c9;
  wire lt8_2_c0;
  wire lt8_2_c1;
  wire lt8_2_c10;
  wire lt8_2_c11;
  wire lt8_2_c12;
  wire lt8_2_c2;
  wire lt8_2_c3;
  wire lt8_2_c4;
  wire lt8_2_c5;
  wire lt8_2_c6;
  wire lt8_2_c7;
  wire lt8_2_c8;
  wire lt8_2_c9;
  wire lt9_2_c0;
  wire lt9_2_c1;
  wire lt9_2_c10;
  wire lt9_2_c11;
  wire lt9_2_c12;
  wire lt9_2_c2;
  wire lt9_2_c3;
  wire lt9_2_c4;
  wire lt9_2_c5;
  wire lt9_2_c6;
  wire lt9_2_c7;
  wire lt9_2_c8;
  wire lt9_2_c9;
  wire mux3_b0_sel_is_0_o;
  wire n0;
  wire n10;
  wire n11;
  wire n12;
  wire n13;
  wire n14;
  wire n16;
  wire n18;
  wire n20;
  wire n23;
  wire n9;
  wire \sub0/c0 ;
  wire \sub0/c1 ;
  wire \sub0/c2 ;
  wire \sub0/c3 ;
  wire \sub0/c4 ;
  wire \sub0/c5 ;
  wire \sub0/c6 ;
  wire \sub1/c0 ;
  wire \sub1/c1 ;
  wire \sub1/c10 ;
  wire \sub1/c11 ;
  wire \sub1/c2 ;
  wire \sub1/c3 ;
  wire \sub1/c4 ;
  wire \sub1/c5 ;
  wire \sub1/c6 ;
  wire \sub1/c7 ;
  wire \sub1/c8 ;
  wire \sub1/c9 ;
  wire \u2/c0 ;
  wire \u2/c1 ;
  wire \u2/c10 ;
  wire \u2/c11 ;
  wire \u2/c12 ;
  wire \u2/c2 ;
  wire \u2/c3 ;
  wire \u2/c4 ;
  wire \u2/c5 ;
  wire \u2/c6 ;
  wire \u2/c7 ;
  wire \u2/c8 ;
  wire \u2/c9 ;

  assign lcd_pwm = rest_n;
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u20 (
    .a(n9),
    .b(n10),
    .o(lcd_hsync));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u21 (
    .a(n11),
    .b(n12),
    .o(lcd_vsync));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u22 (
    .a(clk),
    .b(lcd_pwm),
    .o(lcd_clk));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u23 (
    .a(n13),
    .b(n14),
    .c(n16),
    .d(n18),
    .o(lcd_de));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u24 (
    .a(lcd_de),
    .b(n20),
    .c(n23),
    .o(img_ack));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u25 (
    .a(lcd_de),
    .b(n20),
    .c(n23),
    .d(n6[6]),
    .o(n31[9]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u26 (
    .a(lcd_de),
    .b(n20),
    .c(n23),
    .d(n6[5]),
    .o(n31[8]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u27 (
    .a(lcd_de),
    .b(n20),
    .c(n23),
    .d(n6[4]),
    .o(n31[7]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u28 (
    .a(lcd_de),
    .b(n20),
    .c(n23),
    .d(n6[3]),
    .o(n31[6]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u29 (
    .a(lcd_de),
    .b(n20),
    .c(n23),
    .d(n6[2]),
    .o(n31[5]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u30 (
    .a(lcd_de),
    .b(n20),
    .c(n23),
    .d(n6[1]),
    .o(n31[4]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u31 (
    .a(lcd_de),
    .b(n20),
    .c(n23),
    .d(n6[0]),
    .o(n31[3]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u32 (
    .a(lcd_de),
    .b(n20),
    .c(n23),
    .d(hsync_cnt[2]),
    .o(n31[2]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u33 (
    .a(lcd_de),
    .b(n20),
    .c(n23),
    .d(n6[12]),
    .o(n31[15]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u34 (
    .a(lcd_de),
    .b(n20),
    .c(n23),
    .d(n6[11]),
    .o(n31[14]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u35 (
    .a(lcd_de),
    .b(n20),
    .c(n23),
    .d(n6[10]),
    .o(n31[13]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u36 (
    .a(lcd_de),
    .b(n20),
    .c(n23),
    .d(n6[9]),
    .o(n31[12]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u37 (
    .a(lcd_de),
    .b(n20),
    .c(n23),
    .d(n6[8]),
    .o(n31[11]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u38 (
    .a(lcd_de),
    .b(n20),
    .c(n23),
    .d(n6[7]),
    .o(n31[10]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u39 (
    .a(lcd_de),
    .b(n20),
    .c(n23),
    .d(hsync_cnt[1]),
    .o(n31[1]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u40 (
    .a(lcd_de),
    .b(n20),
    .c(n23),
    .d(hsync_cnt[0]),
    .o(n31[0]));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    _al_u41 (
    .a(hsync_cnt[7]),
    .b(hsync_cnt[8]),
    .c(hsync_cnt[9]),
    .o(_al_u41_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*~B*~A)"),
    .INIT(16'h0010))
    _al_u42 (
    .a(hsync_cnt[3]),
    .b(hsync_cnt[4]),
    .c(hsync_cnt[5]),
    .d(hsync_cnt[6]),
    .o(_al_u42_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u43 (
    .a(hsync_cnt[0]),
    .b(hsync_cnt[1]),
    .c(hsync_cnt[10]),
    .d(hsync_cnt[2]),
    .o(_al_u43_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u44 (
    .a(_al_u41_o),
    .b(_al_u42_o),
    .c(_al_u43_o),
    .o(n0));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    _al_u45 (
    .a(vsync_cnt[7]),
    .b(vsync_cnt[8]),
    .c(vsync_cnt[9]),
    .o(_al_u45_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*A)"),
    .INIT(16'h0002))
    _al_u46 (
    .a(vsync_cnt[3]),
    .b(vsync_cnt[4]),
    .c(vsync_cnt[5]),
    .d(vsync_cnt[6]),
    .o(_al_u46_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*A)"),
    .INIT(16'h0200))
    _al_u47 (
    .a(vsync_cnt[0]),
    .b(vsync_cnt[1]),
    .c(vsync_cnt[10]),
    .d(vsync_cnt[2]),
    .o(_al_u47_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C*B*A))"),
    .INIT(16'h7f00))
    _al_u48 (
    .a(_al_u45_o),
    .b(_al_u46_o),
    .c(_al_u47_o),
    .d(n2[9]),
    .o(n3[9]));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C*B*A))"),
    .INIT(16'h7f00))
    _al_u49 (
    .a(_al_u45_o),
    .b(_al_u46_o),
    .c(_al_u47_o),
    .d(n2[8]),
    .o(n3[8]));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C*B*A))"),
    .INIT(16'h7f00))
    _al_u50 (
    .a(_al_u45_o),
    .b(_al_u46_o),
    .c(_al_u47_o),
    .d(n2[7]),
    .o(n3[7]));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C*B*A))"),
    .INIT(16'h7f00))
    _al_u51 (
    .a(_al_u45_o),
    .b(_al_u46_o),
    .c(_al_u47_o),
    .d(n2[6]),
    .o(n3[6]));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C*B*A))"),
    .INIT(16'h7f00))
    _al_u52 (
    .a(_al_u45_o),
    .b(_al_u46_o),
    .c(_al_u47_o),
    .d(n2[5]),
    .o(n3[5]));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C*B*A))"),
    .INIT(16'h7f00))
    _al_u53 (
    .a(_al_u45_o),
    .b(_al_u46_o),
    .c(_al_u47_o),
    .d(n2[4]),
    .o(n3[4]));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C*B*A))"),
    .INIT(16'h7f00))
    _al_u54 (
    .a(_al_u45_o),
    .b(_al_u46_o),
    .c(_al_u47_o),
    .d(n2[3]),
    .o(n3[3]));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C*B*A))"),
    .INIT(16'h7f00))
    _al_u55 (
    .a(_al_u45_o),
    .b(_al_u46_o),
    .c(_al_u47_o),
    .d(n2[2]),
    .o(n3[2]));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C*B*A))"),
    .INIT(16'h7f00))
    _al_u56 (
    .a(_al_u45_o),
    .b(_al_u46_o),
    .c(_al_u47_o),
    .d(n2[10]),
    .o(n3[10]));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C*B*A))"),
    .INIT(16'h7f00))
    _al_u57 (
    .a(_al_u45_o),
    .b(_al_u46_o),
    .c(_al_u47_o),
    .d(n2[1]),
    .o(n3[1]));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C*B*A))"),
    .INIT(16'h7f00))
    _al_u58 (
    .a(_al_u45_o),
    .b(_al_u46_o),
    .c(_al_u47_o),
    .d(n2[0]),
    .o(n3[0]));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C*B*A))"),
    .INIT(16'h7f00))
    _al_u59 (
    .a(_al_u41_o),
    .b(_al_u42_o),
    .c(_al_u43_o),
    .d(lcd_pwm),
    .o(mux3_b0_sel_is_0_o));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add0/u0  (
    .a(vsync_cnt[0]),
    .b(1'b1),
    .c(\add0/c0 ),
    .o({\add0/c1 ,n2[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add0/u1  (
    .a(vsync_cnt[1]),
    .b(1'b0),
    .c(\add0/c1 ),
    .o({\add0/c2 ,n2[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add0/u10  (
    .a(vsync_cnt[10]),
    .b(1'b0),
    .c(\add0/c10 ),
    .o({open_n0,n2[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add0/u2  (
    .a(vsync_cnt[2]),
    .b(1'b0),
    .c(\add0/c2 ),
    .o({\add0/c3 ,n2[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add0/u3  (
    .a(vsync_cnt[3]),
    .b(1'b0),
    .c(\add0/c3 ),
    .o({\add0/c4 ,n2[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add0/u4  (
    .a(vsync_cnt[4]),
    .b(1'b0),
    .c(\add0/c4 ),
    .o({\add0/c5 ,n2[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add0/u5  (
    .a(vsync_cnt[5]),
    .b(1'b0),
    .c(\add0/c5 ),
    .o({\add0/c6 ,n2[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add0/u6  (
    .a(vsync_cnt[6]),
    .b(1'b0),
    .c(\add0/c6 ),
    .o({\add0/c7 ,n2[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add0/u7  (
    .a(vsync_cnt[7]),
    .b(1'b0),
    .c(\add0/c7 ),
    .o({\add0/c8 ,n2[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add0/u8  (
    .a(vsync_cnt[8]),
    .b(1'b0),
    .c(\add0/c8 ),
    .o({\add0/c9 ,n2[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add0/u9  (
    .a(vsync_cnt[9]),
    .b(1'b0),
    .c(\add0/c9 ),
    .o({\add0/c10 ,n2[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \add0/ucin  (
    .a(1'b0),
    .o({\add0/c0 ,open_n3}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add1/u0  (
    .a(hsync_cnt[0]),
    .b(1'b1),
    .c(\add1/c0 ),
    .o({\add1/c1 ,n4[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add1/u1  (
    .a(hsync_cnt[1]),
    .b(1'b0),
    .c(\add1/c1 ),
    .o({\add1/c2 ,n4[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add1/u10  (
    .a(hsync_cnt[10]),
    .b(1'b0),
    .c(\add1/c10 ),
    .o({open_n4,n4[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add1/u2  (
    .a(hsync_cnt[2]),
    .b(1'b0),
    .c(\add1/c2 ),
    .o({\add1/c3 ,n4[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add1/u3  (
    .a(hsync_cnt[3]),
    .b(1'b0),
    .c(\add1/c3 ),
    .o({\add1/c4 ,n4[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add1/u4  (
    .a(hsync_cnt[4]),
    .b(1'b0),
    .c(\add1/c4 ),
    .o({\add1/c5 ,n4[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add1/u5  (
    .a(hsync_cnt[5]),
    .b(1'b0),
    .c(\add1/c5 ),
    .o({\add1/c6 ,n4[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add1/u6  (
    .a(hsync_cnt[6]),
    .b(1'b0),
    .c(\add1/c6 ),
    .o({\add1/c7 ,n4[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add1/u7  (
    .a(hsync_cnt[7]),
    .b(1'b0),
    .c(\add1/c7 ),
    .o({\add1/c8 ,n4[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add1/u8  (
    .a(hsync_cnt[8]),
    .b(1'b0),
    .c(\add1/c8 ),
    .o({\add1/c9 ,n4[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add1/u9  (
    .a(hsync_cnt[9]),
    .b(1'b0),
    .c(\add1/c9 ),
    .o({\add1/c10 ,n4[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \add1/ucin  (
    .a(1'b0),
    .o({\add1/c0 ,open_n7}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt0_0 (
    .a(1'b0),
    .b(hsync_cnt[0]),
    .c(lt0_c0),
    .o({lt0_c1,open_n8}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt0_1 (
    .a(1'b0),
    .b(hsync_cnt[1]),
    .c(lt0_c1),
    .o({lt0_c2,open_n9}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt0_10 (
    .a(1'b0),
    .b(hsync_cnt[10]),
    .c(lt0_c10),
    .o({lt0_c11,open_n10}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt0_2 (
    .a(1'b0),
    .b(hsync_cnt[2]),
    .c(lt0_c2),
    .o({lt0_c3,open_n11}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt0_3 (
    .a(1'b0),
    .b(hsync_cnt[3]),
    .c(lt0_c3),
    .o({lt0_c4,open_n12}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt0_4 (
    .a(1'b1),
    .b(hsync_cnt[4]),
    .c(lt0_c4),
    .o({lt0_c5,open_n13}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt0_5 (
    .a(1'b0),
    .b(hsync_cnt[5]),
    .c(lt0_c5),
    .o({lt0_c6,open_n14}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt0_6 (
    .a(1'b0),
    .b(hsync_cnt[6]),
    .c(lt0_c6),
    .o({lt0_c7,open_n15}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt0_7 (
    .a(1'b0),
    .b(hsync_cnt[7]),
    .c(lt0_c7),
    .o({lt0_c8,open_n16}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt0_8 (
    .a(1'b0),
    .b(hsync_cnt[8]),
    .c(lt0_c8),
    .o({lt0_c9,open_n17}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt0_9 (
    .a(1'b0),
    .b(hsync_cnt[9]),
    .c(lt0_c9),
    .o({lt0_c10,open_n18}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    lt0_cin (
    .a(1'b1),
    .o({lt0_c0,open_n21}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt0_cout (
    .a(1'b0),
    .b(1'b1),
    .c(lt0_c11),
    .o({open_n22,n9}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt1_0 (
    .a(hsync_cnt[0]),
    .b(1'b0),
    .c(lt1_c0),
    .o({lt1_c1,open_n23}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt1_1 (
    .a(hsync_cnt[1]),
    .b(1'b0),
    .c(lt1_c1),
    .o({lt1_c2,open_n24}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt1_10 (
    .a(hsync_cnt[10]),
    .b(1'b0),
    .c(lt1_c10),
    .o({lt1_c11,open_n25}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt1_2 (
    .a(hsync_cnt[2]),
    .b(1'b0),
    .c(lt1_c2),
    .o({lt1_c3,open_n26}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt1_3 (
    .a(hsync_cnt[3]),
    .b(1'b0),
    .c(lt1_c3),
    .o({lt1_c4,open_n27}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt1_4 (
    .a(hsync_cnt[4]),
    .b(1'b1),
    .c(lt1_c4),
    .o({lt1_c5,open_n28}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt1_5 (
    .a(hsync_cnt[5]),
    .b(1'b1),
    .c(lt1_c5),
    .o({lt1_c6,open_n29}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt1_6 (
    .a(hsync_cnt[6]),
    .b(1'b1),
    .c(lt1_c6),
    .o({lt1_c7,open_n30}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt1_7 (
    .a(hsync_cnt[7]),
    .b(1'b0),
    .c(lt1_c7),
    .o({lt1_c8,open_n31}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt1_8 (
    .a(hsync_cnt[8]),
    .b(1'b0),
    .c(lt1_c8),
    .o({lt1_c9,open_n32}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt1_9 (
    .a(hsync_cnt[9]),
    .b(1'b0),
    .c(lt1_c9),
    .o({lt1_c10,open_n33}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    lt1_cin (
    .a(1'b0),
    .o({lt1_c0,open_n36}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt1_cout (
    .a(1'b0),
    .b(1'b1),
    .c(lt1_c11),
    .o({open_n37,n10}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt2_0 (
    .a(1'b0),
    .b(vsync_cnt[0]),
    .c(lt2_c0),
    .o({lt2_c1,open_n38}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt2_1 (
    .a(1'b1),
    .b(vsync_cnt[1]),
    .c(lt2_c1),
    .o({lt2_c2,open_n39}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt2_10 (
    .a(1'b0),
    .b(vsync_cnt[10]),
    .c(lt2_c10),
    .o({lt2_c11,open_n40}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt2_2 (
    .a(1'b0),
    .b(vsync_cnt[2]),
    .c(lt2_c2),
    .o({lt2_c3,open_n41}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt2_3 (
    .a(1'b1),
    .b(vsync_cnt[3]),
    .c(lt2_c3),
    .o({lt2_c4,open_n42}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt2_4 (
    .a(1'b0),
    .b(vsync_cnt[4]),
    .c(lt2_c4),
    .o({lt2_c5,open_n43}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt2_5 (
    .a(1'b0),
    .b(vsync_cnt[5]),
    .c(lt2_c5),
    .o({lt2_c6,open_n44}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt2_6 (
    .a(1'b0),
    .b(vsync_cnt[6]),
    .c(lt2_c6),
    .o({lt2_c7,open_n45}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt2_7 (
    .a(1'b0),
    .b(vsync_cnt[7]),
    .c(lt2_c7),
    .o({lt2_c8,open_n46}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt2_8 (
    .a(1'b0),
    .b(vsync_cnt[8]),
    .c(lt2_c8),
    .o({lt2_c9,open_n47}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt2_9 (
    .a(1'b0),
    .b(vsync_cnt[9]),
    .c(lt2_c9),
    .o({lt2_c10,open_n48}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    lt2_cin (
    .a(1'b1),
    .o({lt2_c0,open_n51}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt2_cout (
    .a(1'b0),
    .b(1'b1),
    .c(lt2_c11),
    .o({open_n52,n11}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt3_0 (
    .a(vsync_cnt[0]),
    .b(1'b0),
    .c(lt3_c0),
    .o({lt3_c1,open_n53}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt3_1 (
    .a(vsync_cnt[1]),
    .b(1'b0),
    .c(lt3_c1),
    .o({lt3_c2,open_n54}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt3_10 (
    .a(vsync_cnt[10]),
    .b(1'b0),
    .c(lt3_c10),
    .o({lt3_c11,open_n55}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt3_2 (
    .a(vsync_cnt[2]),
    .b(1'b1),
    .c(lt3_c2),
    .o({lt3_c3,open_n56}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt3_3 (
    .a(vsync_cnt[3]),
    .b(1'b1),
    .c(lt3_c3),
    .o({lt3_c4,open_n57}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt3_4 (
    .a(vsync_cnt[4]),
    .b(1'b0),
    .c(lt3_c4),
    .o({lt3_c5,open_n58}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt3_5 (
    .a(vsync_cnt[5]),
    .b(1'b0),
    .c(lt3_c5),
    .o({lt3_c6,open_n59}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt3_6 (
    .a(vsync_cnt[6]),
    .b(1'b0),
    .c(lt3_c6),
    .o({lt3_c7,open_n60}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt3_7 (
    .a(vsync_cnt[7]),
    .b(1'b0),
    .c(lt3_c7),
    .o({lt3_c8,open_n61}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt3_8 (
    .a(vsync_cnt[8]),
    .b(1'b0),
    .c(lt3_c8),
    .o({lt3_c9,open_n62}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt3_9 (
    .a(vsync_cnt[9]),
    .b(1'b0),
    .c(lt3_c9),
    .o({lt3_c10,open_n63}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    lt3_cin (
    .a(1'b0),
    .o({lt3_c0,open_n66}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt3_cout (
    .a(1'b0),
    .b(1'b1),
    .c(lt3_c11),
    .o({open_n67,n12}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt4_0 (
    .a(1'b0),
    .b(hsync_cnt[0]),
    .c(lt4_c0),
    .o({lt4_c1,open_n68}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt4_1 (
    .a(1'b0),
    .b(hsync_cnt[1]),
    .c(lt4_c1),
    .o({lt4_c2,open_n69}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt4_10 (
    .a(1'b0),
    .b(hsync_cnt[10]),
    .c(lt4_c10),
    .o({lt4_c11,open_n70}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt4_2 (
    .a(1'b0),
    .b(hsync_cnt[2]),
    .c(lt4_c2),
    .o({lt4_c3,open_n71}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt4_3 (
    .a(1'b0),
    .b(hsync_cnt[3]),
    .c(lt4_c3),
    .o({lt4_c4,open_n72}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt4_4 (
    .a(1'b0),
    .b(hsync_cnt[4]),
    .c(lt4_c4),
    .o({lt4_c5,open_n73}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt4_5 (
    .a(1'b1),
    .b(hsync_cnt[5]),
    .c(lt4_c5),
    .o({lt4_c6,open_n74}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt4_6 (
    .a(1'b0),
    .b(hsync_cnt[6]),
    .c(lt4_c6),
    .o({lt4_c7,open_n75}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt4_7 (
    .a(1'b1),
    .b(hsync_cnt[7]),
    .c(lt4_c7),
    .o({lt4_c8,open_n76}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt4_8 (
    .a(1'b0),
    .b(hsync_cnt[8]),
    .c(lt4_c8),
    .o({lt4_c9,open_n77}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt4_9 (
    .a(1'b0),
    .b(hsync_cnt[9]),
    .c(lt4_c9),
    .o({lt4_c10,open_n78}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    lt4_cin (
    .a(1'b1),
    .o({lt4_c0,open_n81}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt4_cout (
    .a(1'b0),
    .b(1'b1),
    .c(lt4_c11),
    .o({open_n82,n13}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt5_0 (
    .a(hsync_cnt[0]),
    .b(1'b0),
    .c(lt5_c0),
    .o({lt5_c1,open_n83}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt5_1 (
    .a(hsync_cnt[1]),
    .b(1'b0),
    .c(lt5_c1),
    .o({lt5_c2,open_n84}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt5_10 (
    .a(hsync_cnt[10]),
    .b(1'b0),
    .c(lt5_c10),
    .o({lt5_c11,open_n85}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt5_2 (
    .a(hsync_cnt[2]),
    .b(1'b0),
    .c(lt5_c2),
    .o({lt5_c3,open_n86}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt5_3 (
    .a(hsync_cnt[3]),
    .b(1'b0),
    .c(lt5_c3),
    .o({lt5_c4,open_n87}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt5_4 (
    .a(hsync_cnt[4]),
    .b(1'b0),
    .c(lt5_c4),
    .o({lt5_c5,open_n88}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt5_5 (
    .a(hsync_cnt[5]),
    .b(1'b1),
    .c(lt5_c5),
    .o({lt5_c6,open_n89}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt5_6 (
    .a(hsync_cnt[6]),
    .b(1'b0),
    .c(lt5_c6),
    .o({lt5_c7,open_n90}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt5_7 (
    .a(hsync_cnt[7]),
    .b(1'b0),
    .c(lt5_c7),
    .o({lt5_c8,open_n91}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt5_8 (
    .a(hsync_cnt[8]),
    .b(1'b1),
    .c(lt5_c8),
    .o({lt5_c9,open_n92}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt5_9 (
    .a(hsync_cnt[9]),
    .b(1'b1),
    .c(lt5_c9),
    .o({lt5_c10,open_n93}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    lt5_cin (
    .a(1'b1),
    .o({lt5_c0,open_n96}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt5_cout (
    .a(1'b0),
    .b(1'b1),
    .c(lt5_c11),
    .o({open_n97,n14}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt6_0 (
    .a(1'b1),
    .b(vsync_cnt[0]),
    .c(lt6_c0),
    .o({lt6_c1,open_n98}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt6_1 (
    .a(1'b0),
    .b(vsync_cnt[1]),
    .c(lt6_c1),
    .o({lt6_c2,open_n99}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt6_10 (
    .a(1'b0),
    .b(vsync_cnt[10]),
    .c(lt6_c10),
    .o({lt6_c11,open_n100}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt6_2 (
    .a(1'b1),
    .b(vsync_cnt[2]),
    .c(lt6_c2),
    .o({lt6_c3,open_n101}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt6_3 (
    .a(1'b1),
    .b(vsync_cnt[3]),
    .c(lt6_c3),
    .o({lt6_c4,open_n102}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt6_4 (
    .a(1'b0),
    .b(vsync_cnt[4]),
    .c(lt6_c4),
    .o({lt6_c5,open_n103}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt6_5 (
    .a(1'b1),
    .b(vsync_cnt[5]),
    .c(lt6_c5),
    .o({lt6_c6,open_n104}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt6_6 (
    .a(1'b0),
    .b(vsync_cnt[6]),
    .c(lt6_c6),
    .o({lt6_c7,open_n105}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt6_7 (
    .a(1'b0),
    .b(vsync_cnt[7]),
    .c(lt6_c7),
    .o({lt6_c8,open_n106}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt6_8 (
    .a(1'b0),
    .b(vsync_cnt[8]),
    .c(lt6_c8),
    .o({lt6_c9,open_n107}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt6_9 (
    .a(1'b0),
    .b(vsync_cnt[9]),
    .c(lt6_c9),
    .o({lt6_c10,open_n108}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    lt6_cin (
    .a(1'b1),
    .o({lt6_c0,open_n111}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt6_cout (
    .a(1'b0),
    .b(1'b1),
    .c(lt6_c11),
    .o({open_n112,n16}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt7_0 (
    .a(vsync_cnt[0]),
    .b(1'b1),
    .c(lt7_c0),
    .o({lt7_c1,open_n113}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt7_1 (
    .a(vsync_cnt[1]),
    .b(1'b0),
    .c(lt7_c1),
    .o({lt7_c2,open_n114}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt7_10 (
    .a(vsync_cnt[10]),
    .b(1'b0),
    .c(lt7_c10),
    .o({lt7_c11,open_n115}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt7_2 (
    .a(vsync_cnt[2]),
    .b(1'b1),
    .c(lt7_c2),
    .o({lt7_c3,open_n116}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt7_3 (
    .a(vsync_cnt[3]),
    .b(1'b1),
    .c(lt7_c3),
    .o({lt7_c4,open_n117}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt7_4 (
    .a(vsync_cnt[4]),
    .b(1'b0),
    .c(lt7_c4),
    .o({lt7_c5,open_n118}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt7_5 (
    .a(vsync_cnt[5]),
    .b(1'b0),
    .c(lt7_c5),
    .o({lt7_c6,open_n119}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt7_6 (
    .a(vsync_cnt[6]),
    .b(1'b0),
    .c(lt7_c6),
    .o({lt7_c7,open_n120}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt7_7 (
    .a(vsync_cnt[7]),
    .b(1'b0),
    .c(lt7_c7),
    .o({lt7_c8,open_n121}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt7_8 (
    .a(vsync_cnt[8]),
    .b(1'b0),
    .c(lt7_c8),
    .o({lt7_c9,open_n122}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt7_9 (
    .a(vsync_cnt[9]),
    .b(1'b1),
    .c(lt7_c9),
    .o({lt7_c10,open_n123}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    lt7_cin (
    .a(1'b0),
    .o({lt7_c0,open_n126}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt7_cout (
    .a(1'b0),
    .b(1'b1),
    .c(lt7_c11),
    .o({open_n127,n18}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt8_2_0 (
    .a(hsync_cnt[0]),
    .b(1'b0),
    .c(lt8_2_c0),
    .o({lt8_2_c1,open_n128}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt8_2_1 (
    .a(hsync_cnt[1]),
    .b(1'b0),
    .c(lt8_2_c1),
    .o({lt8_2_c2,open_n129}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt8_2_10 (
    .a(n7[5]),
    .b(1'b0),
    .c(lt8_2_c10),
    .o({lt8_2_c11,open_n130}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt8_2_11 (
    .a(n7[6]),
    .b(1'b0),
    .c(lt8_2_c11),
    .o({lt8_2_c12,open_n131}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt8_2_2 (
    .a(hsync_cnt[2]),
    .b(1'b0),
    .c(lt8_2_c2),
    .o({lt8_2_c3,open_n132}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt8_2_3 (
    .a(hsync_cnt[3]),
    .b(1'b1),
    .c(lt8_2_c3),
    .o({lt8_2_c4,open_n133}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt8_2_4 (
    .a(hsync_cnt[4]),
    .b(1'b0),
    .c(lt8_2_c4),
    .o({lt8_2_c5,open_n134}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt8_2_5 (
    .a(n7[0]),
    .b(1'b0),
    .c(lt8_2_c5),
    .o({lt8_2_c6,open_n135}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt8_2_6 (
    .a(n7[1]),
    .b(1'b1),
    .c(lt8_2_c6),
    .o({lt8_2_c7,open_n136}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt8_2_7 (
    .a(n7[2]),
    .b(1'b1),
    .c(lt8_2_c7),
    .o({lt8_2_c8,open_n137}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt8_2_8 (
    .a(n7[3]),
    .b(1'b0),
    .c(lt8_2_c8),
    .o({lt8_2_c9,open_n138}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt8_2_9 (
    .a(n7[4]),
    .b(1'b0),
    .c(lt8_2_c9),
    .o({lt8_2_c10,open_n139}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    lt8_2_cin (
    .a(1'b0),
    .o({lt8_2_c0,open_n142}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt8_2_cout (
    .a(1'b0),
    .b(1'b1),
    .c(lt8_2_c12),
    .o({open_n143,n20}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt9_2_0 (
    .a(n22[0]),
    .b(1'b0),
    .c(lt9_2_c0),
    .o({lt9_2_c1,open_n144}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt9_2_1 (
    .a(n22[1]),
    .b(1'b0),
    .c(lt9_2_c1),
    .o({lt9_2_c2,open_n145}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt9_2_10 (
    .a(n22[10]),
    .b(1'b0),
    .c(lt9_2_c10),
    .o({lt9_2_c11,open_n146}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt9_2_11 (
    .a(n22[11]),
    .b(1'b0),
    .c(lt9_2_c11),
    .o({lt9_2_c12,open_n147}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt9_2_2 (
    .a(n22[2]),
    .b(1'b1),
    .c(lt9_2_c2),
    .o({lt9_2_c3,open_n148}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt9_2_3 (
    .a(n22[3]),
    .b(1'b0),
    .c(lt9_2_c3),
    .o({lt9_2_c4,open_n149}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt9_2_4 (
    .a(n22[4]),
    .b(1'b0),
    .c(lt9_2_c4),
    .o({lt9_2_c5,open_n150}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt9_2_5 (
    .a(n22[5]),
    .b(1'b1),
    .c(lt9_2_c5),
    .o({lt9_2_c6,open_n151}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt9_2_6 (
    .a(n22[6]),
    .b(1'b0),
    .c(lt9_2_c6),
    .o({lt9_2_c7,open_n152}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt9_2_7 (
    .a(n22[7]),
    .b(1'b1),
    .c(lt9_2_c7),
    .o({lt9_2_c8,open_n153}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt9_2_8 (
    .a(n22[8]),
    .b(1'b0),
    .c(lt9_2_c8),
    .o({lt9_2_c9,open_n154}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt9_2_9 (
    .a(n22[9]),
    .b(1'b0),
    .c(lt9_2_c9),
    .o({lt9_2_c10,open_n155}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    lt9_2_cin (
    .a(1'b0),
    .o({lt9_2_c0,open_n158}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    lt9_2_cout (
    .a(1'b0),
    .b(1'b1),
    .c(lt9_2_c12),
    .o({open_n159,n23}));
  EG_PHY_MULT18 #(
    .INPUTREGA("DISABLE"),
    .INPUTREGB("DISABLE"),
    .MODE("MULT18X18C"),
    .OUTPUTREG("DISABLE"),
    .SIGNEDAMUX("0"),
    .SIGNEDBMUX("0"))
    mult0_ (
    .a({5'b00000,n22[11],n22}),
    .b(18'b000000000000011001),
    .p({open_n243,open_n244,open_n245,open_n246,open_n247,open_n248,open_n249,open_n250,open_n251,open_n252,open_n253,open_n254,open_n255,open_n256,open_n257,open_n258,open_n259,open_n260,open_n261,open_n262,open_n263,open_n264,open_n265,n29[15:3]}));
  reg_sr_as_w1 reg0_b0 (
    .clk(clk),
    .d(n3[0]),
    .en(n0),
    .reset(~lcd_pwm),
    .set(1'b0),
    .q(vsync_cnt[0]));  // sources/rtl/lcd_sync.v(56)
  reg_sr_as_w1 reg0_b1 (
    .clk(clk),
    .d(n3[1]),
    .en(n0),
    .reset(~lcd_pwm),
    .set(1'b0),
    .q(vsync_cnt[1]));  // sources/rtl/lcd_sync.v(56)
  reg_sr_as_w1 reg0_b10 (
    .clk(clk),
    .d(n3[10]),
    .en(n0),
    .reset(~lcd_pwm),
    .set(1'b0),
    .q(vsync_cnt[10]));  // sources/rtl/lcd_sync.v(56)
  reg_sr_as_w1 reg0_b2 (
    .clk(clk),
    .d(n3[2]),
    .en(n0),
    .reset(~lcd_pwm),
    .set(1'b0),
    .q(vsync_cnt[2]));  // sources/rtl/lcd_sync.v(56)
  reg_sr_as_w1 reg0_b3 (
    .clk(clk),
    .d(n3[3]),
    .en(n0),
    .reset(~lcd_pwm),
    .set(1'b0),
    .q(vsync_cnt[3]));  // sources/rtl/lcd_sync.v(56)
  reg_sr_as_w1 reg0_b4 (
    .clk(clk),
    .d(n3[4]),
    .en(n0),
    .reset(~lcd_pwm),
    .set(1'b0),
    .q(vsync_cnt[4]));  // sources/rtl/lcd_sync.v(56)
  reg_sr_as_w1 reg0_b5 (
    .clk(clk),
    .d(n3[5]),
    .en(n0),
    .reset(~lcd_pwm),
    .set(1'b0),
    .q(vsync_cnt[5]));  // sources/rtl/lcd_sync.v(56)
  reg_sr_as_w1 reg0_b6 (
    .clk(clk),
    .d(n3[6]),
    .en(n0),
    .reset(~lcd_pwm),
    .set(1'b0),
    .q(vsync_cnt[6]));  // sources/rtl/lcd_sync.v(56)
  reg_sr_as_w1 reg0_b7 (
    .clk(clk),
    .d(n3[7]),
    .en(n0),
    .reset(~lcd_pwm),
    .set(1'b0),
    .q(vsync_cnt[7]));  // sources/rtl/lcd_sync.v(56)
  reg_sr_as_w1 reg0_b8 (
    .clk(clk),
    .d(n3[8]),
    .en(n0),
    .reset(~lcd_pwm),
    .set(1'b0),
    .q(vsync_cnt[8]));  // sources/rtl/lcd_sync.v(56)
  reg_sr_as_w1 reg0_b9 (
    .clk(clk),
    .d(n3[9]),
    .en(n0),
    .reset(~lcd_pwm),
    .set(1'b0),
    .q(vsync_cnt[9]));  // sources/rtl/lcd_sync.v(56)
  reg_ar_as_w1 reg1_b0 (
    .clk(clk),
    .d(n31[0]),
    .en(1'b1),
    .reset(~lcd_pwm),
    .set(1'b0),
    .q(addr[0]));  // sources/rtl/lcd_sync.v(81)
  reg_ar_as_w1 reg1_b1 (
    .clk(clk),
    .d(n31[1]),
    .en(1'b1),
    .reset(~lcd_pwm),
    .set(1'b0),
    .q(addr[1]));  // sources/rtl/lcd_sync.v(81)
  reg_ar_as_w1 reg1_b10 (
    .clk(clk),
    .d(n31[10]),
    .en(1'b1),
    .reset(~lcd_pwm),
    .set(1'b0),
    .q(addr[10]));  // sources/rtl/lcd_sync.v(81)
  reg_ar_as_w1 reg1_b11 (
    .clk(clk),
    .d(n31[11]),
    .en(1'b1),
    .reset(~lcd_pwm),
    .set(1'b0),
    .q(addr[11]));  // sources/rtl/lcd_sync.v(81)
  reg_ar_as_w1 reg1_b12 (
    .clk(clk),
    .d(n31[12]),
    .en(1'b1),
    .reset(~lcd_pwm),
    .set(1'b0),
    .q(addr[12]));  // sources/rtl/lcd_sync.v(81)
  reg_ar_as_w1 reg1_b13 (
    .clk(clk),
    .d(n31[13]),
    .en(1'b1),
    .reset(~lcd_pwm),
    .set(1'b0),
    .q(addr[13]));  // sources/rtl/lcd_sync.v(81)
  reg_ar_as_w1 reg1_b14 (
    .clk(clk),
    .d(n31[14]),
    .en(1'b1),
    .reset(~lcd_pwm),
    .set(1'b0),
    .q(addr[14]));  // sources/rtl/lcd_sync.v(81)
  reg_ar_as_w1 reg1_b15 (
    .clk(clk),
    .d(n31[15]),
    .en(1'b1),
    .reset(~lcd_pwm),
    .set(1'b0),
    .q(addr[15]));  // sources/rtl/lcd_sync.v(81)
  reg_ar_as_w1 reg1_b2 (
    .clk(clk),
    .d(n31[2]),
    .en(1'b1),
    .reset(~lcd_pwm),
    .set(1'b0),
    .q(addr[2]));  // sources/rtl/lcd_sync.v(81)
  reg_ar_as_w1 reg1_b3 (
    .clk(clk),
    .d(n31[3]),
    .en(1'b1),
    .reset(~lcd_pwm),
    .set(1'b0),
    .q(addr[3]));  // sources/rtl/lcd_sync.v(81)
  reg_ar_as_w1 reg1_b4 (
    .clk(clk),
    .d(n31[4]),
    .en(1'b1),
    .reset(~lcd_pwm),
    .set(1'b0),
    .q(addr[4]));  // sources/rtl/lcd_sync.v(81)
  reg_ar_as_w1 reg1_b5 (
    .clk(clk),
    .d(n31[5]),
    .en(1'b1),
    .reset(~lcd_pwm),
    .set(1'b0),
    .q(addr[5]));  // sources/rtl/lcd_sync.v(81)
  reg_ar_as_w1 reg1_b6 (
    .clk(clk),
    .d(n31[6]),
    .en(1'b1),
    .reset(~lcd_pwm),
    .set(1'b0),
    .q(addr[6]));  // sources/rtl/lcd_sync.v(81)
  reg_ar_as_w1 reg1_b7 (
    .clk(clk),
    .d(n31[7]),
    .en(1'b1),
    .reset(~lcd_pwm),
    .set(1'b0),
    .q(addr[7]));  // sources/rtl/lcd_sync.v(81)
  reg_ar_as_w1 reg1_b8 (
    .clk(clk),
    .d(n31[8]),
    .en(1'b1),
    .reset(~lcd_pwm),
    .set(1'b0),
    .q(addr[8]));  // sources/rtl/lcd_sync.v(81)
  reg_ar_as_w1 reg1_b9 (
    .clk(clk),
    .d(n31[9]),
    .en(1'b1),
    .reset(~lcd_pwm),
    .set(1'b0),
    .q(addr[9]));  // sources/rtl/lcd_sync.v(81)
  reg_sr_as_w1 reg2_b0 (
    .clk(clk),
    .d(n4[0]),
    .en(1'b1),
    .reset(~mux3_b0_sel_is_0_o),
    .set(1'b0),
    .q(hsync_cnt[0]));  // sources/rtl/lcd_sync.v(56)
  reg_sr_as_w1 reg2_b1 (
    .clk(clk),
    .d(n4[1]),
    .en(1'b1),
    .reset(~mux3_b0_sel_is_0_o),
    .set(1'b0),
    .q(hsync_cnt[1]));  // sources/rtl/lcd_sync.v(56)
  reg_sr_as_w1 reg2_b10 (
    .clk(clk),
    .d(n4[10]),
    .en(1'b1),
    .reset(~mux3_b0_sel_is_0_o),
    .set(1'b0),
    .q(hsync_cnt[10]));  // sources/rtl/lcd_sync.v(56)
  reg_sr_as_w1 reg2_b2 (
    .clk(clk),
    .d(n4[2]),
    .en(1'b1),
    .reset(~mux3_b0_sel_is_0_o),
    .set(1'b0),
    .q(hsync_cnt[2]));  // sources/rtl/lcd_sync.v(56)
  reg_sr_as_w1 reg2_b3 (
    .clk(clk),
    .d(n4[3]),
    .en(1'b1),
    .reset(~mux3_b0_sel_is_0_o),
    .set(1'b0),
    .q(hsync_cnt[3]));  // sources/rtl/lcd_sync.v(56)
  reg_sr_as_w1 reg2_b4 (
    .clk(clk),
    .d(n4[4]),
    .en(1'b1),
    .reset(~mux3_b0_sel_is_0_o),
    .set(1'b0),
    .q(hsync_cnt[4]));  // sources/rtl/lcd_sync.v(56)
  reg_sr_as_w1 reg2_b5 (
    .clk(clk),
    .d(n4[5]),
    .en(1'b1),
    .reset(~mux3_b0_sel_is_0_o),
    .set(1'b0),
    .q(hsync_cnt[5]));  // sources/rtl/lcd_sync.v(56)
  reg_sr_as_w1 reg2_b6 (
    .clk(clk),
    .d(n4[6]),
    .en(1'b1),
    .reset(~mux3_b0_sel_is_0_o),
    .set(1'b0),
    .q(hsync_cnt[6]));  // sources/rtl/lcd_sync.v(56)
  reg_sr_as_w1 reg2_b7 (
    .clk(clk),
    .d(n4[7]),
    .en(1'b1),
    .reset(~mux3_b0_sel_is_0_o),
    .set(1'b0),
    .q(hsync_cnt[7]));  // sources/rtl/lcd_sync.v(56)
  reg_sr_as_w1 reg2_b8 (
    .clk(clk),
    .d(n4[8]),
    .en(1'b1),
    .reset(~mux3_b0_sel_is_0_o),
    .set(1'b0),
    .q(hsync_cnt[8]));  // sources/rtl/lcd_sync.v(56)
  reg_sr_as_w1 reg2_b9 (
    .clk(clk),
    .d(n4[9]),
    .en(1'b1),
    .reset(~mux3_b0_sel_is_0_o),
    .set(1'b0),
    .q(hsync_cnt[9]));  // sources/rtl/lcd_sync.v(56)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \sub0/u0  (
    .a(hsync_cnt[5]),
    .b(1'b1),
    .c(\sub0/c0 ),
    .o({\sub0/c1 ,n7[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \sub0/u1  (
    .a(hsync_cnt[6]),
    .b(1'b0),
    .c(\sub0/c1 ),
    .o({\sub0/c2 ,n7[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \sub0/u2  (
    .a(hsync_cnt[7]),
    .b(1'b1),
    .c(\sub0/c2 ),
    .o({\sub0/c3 ,n7[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \sub0/u3  (
    .a(hsync_cnt[8]),
    .b(1'b0),
    .c(\sub0/c3 ),
    .o({\sub0/c4 ,n7[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \sub0/u4  (
    .a(hsync_cnt[9]),
    .b(1'b0),
    .c(\sub0/c4 ),
    .o({\sub0/c5 ,n7[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \sub0/u5  (
    .a(hsync_cnt[10]),
    .b(1'b0),
    .c(\sub0/c5 ),
    .o({\sub0/c6 ,n7[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    \sub0/ucin  (
    .a(1'b0),
    .o({\sub0/c0 ,open_n268}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \sub0/ucout  (
    .c(\sub0/c6 ),
    .o({open_n271,n7[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \sub1/u0  (
    .a(vsync_cnt[0]),
    .b(1'b1),
    .c(\sub1/c0 ),
    .o({\sub1/c1 ,n22[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \sub1/u1  (
    .a(vsync_cnt[1]),
    .b(1'b0),
    .c(\sub1/c1 ),
    .o({\sub1/c2 ,n22[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \sub1/u10  (
    .a(vsync_cnt[10]),
    .b(1'b0),
    .c(\sub1/c10 ),
    .o({\sub1/c11 ,n22[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \sub1/u2  (
    .a(vsync_cnt[2]),
    .b(1'b1),
    .c(\sub1/c2 ),
    .o({\sub1/c3 ,n22[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \sub1/u3  (
    .a(vsync_cnt[3]),
    .b(1'b1),
    .c(\sub1/c3 ),
    .o({\sub1/c4 ,n22[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \sub1/u4  (
    .a(vsync_cnt[4]),
    .b(1'b0),
    .c(\sub1/c4 ),
    .o({\sub1/c5 ,n22[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \sub1/u5  (
    .a(vsync_cnt[5]),
    .b(1'b1),
    .c(\sub1/c5 ),
    .o({\sub1/c6 ,n22[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \sub1/u6  (
    .a(vsync_cnt[6]),
    .b(1'b0),
    .c(\sub1/c6 ),
    .o({\sub1/c7 ,n22[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \sub1/u7  (
    .a(vsync_cnt[7]),
    .b(1'b0),
    .c(\sub1/c7 ),
    .o({\sub1/c8 ,n22[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \sub1/u8  (
    .a(vsync_cnt[8]),
    .b(1'b0),
    .c(\sub1/c8 ),
    .o({\sub1/c9 ,n22[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \sub1/u9  (
    .a(vsync_cnt[9]),
    .b(1'b0),
    .c(\sub1/c9 ),
    .o({\sub1/c10 ,n22[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    \sub1/ucin  (
    .a(1'b0),
    .o({\sub1/c0 ,open_n274}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \sub1/ucout  (
    .c(\sub1/c11 ),
    .o({open_n277,n22[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2/u0  (
    .a(hsync_cnt[3]),
    .b(n29[3]),
    .c(\u2/c0 ),
    .o({\u2/c1 ,n6[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2/u1  (
    .a(hsync_cnt[4]),
    .b(n29[4]),
    .c(\u2/c1 ),
    .o({\u2/c2 ,n6[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2/u10  (
    .a(n7[6]),
    .b(n29[13]),
    .c(\u2/c10 ),
    .o({\u2/c11 ,n6[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2/u11  (
    .a(n7[6]),
    .b(n29[14]),
    .c(\u2/c11 ),
    .o({\u2/c12 ,n6[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2/u12  (
    .a(n7[6]),
    .b(n29[15]),
    .c(\u2/c12 ),
    .o({open_n278,n6[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2/u2  (
    .a(n7[0]),
    .b(n29[5]),
    .c(\u2/c2 ),
    .o({\u2/c3 ,n6[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2/u3  (
    .a(n7[1]),
    .b(n29[6]),
    .c(\u2/c3 ),
    .o({\u2/c4 ,n6[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2/u4  (
    .a(n7[2]),
    .b(n29[7]),
    .c(\u2/c4 ),
    .o({\u2/c5 ,n6[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2/u5  (
    .a(n7[3]),
    .b(n29[8]),
    .c(\u2/c5 ),
    .o({\u2/c6 ,n6[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2/u6  (
    .a(n7[4]),
    .b(n29[9]),
    .c(\u2/c6 ),
    .o({\u2/c7 ,n6[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2/u7  (
    .a(n7[5]),
    .b(n29[10]),
    .c(\u2/c7 ),
    .o({\u2/c8 ,n6[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2/u8  (
    .a(n7[6]),
    .b(n29[11]),
    .c(\u2/c8 ),
    .o({\u2/c9 ,n6[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2/u9  (
    .a(n7[6]),
    .b(n29[12]),
    .c(\u2/c9 ),
    .o({\u2/c10 ,n6[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2/ucin  (
    .a(1'b0),
    .o({\u2/c0 ,open_n281}));

endmodule 

module i2c_module  // sources/rtl/i2c_module.v(2)
  (
  address,
  clk,
  reset_n,
  sda_in,
  write,
  writedata,
  ready,
  scl_out,
  sda,
  sda_oe,
  success_out
  );

  input [2:0] address;  // sources/rtl/i2c_module.v(14)
  input clk;  // sources/rtl/i2c_module.v(3)
  input reset_n;  // sources/rtl/i2c_module.v(4)
  input sda_in;  // sources/rtl/i2c_module.v(7)
  input write;  // sources/rtl/i2c_module.v(13)
  input [7:0] writedata;  // sources/rtl/i2c_module.v(12)
  output ready;  // sources/rtl/i2c_module.v(16)
  output scl_out;  // sources/rtl/i2c_module.v(10)
  output sda;  // sources/rtl/i2c_module.v(8)
  output sda_oe;  // sources/rtl/i2c_module.v(6)
  output success_out;  // sources/rtl/i2c_module.v(17)

  // localparam STATE_ADDRESS_ACK = 10;
  // localparam STATE_ADDRESS_BIT_1 = 2;
  // localparam STATE_ADDRESS_BIT_2 = 3;
  // localparam STATE_ADDRESS_BIT_3 = 4;
  // localparam STATE_ADDRESS_BIT_4 = 5;
  // localparam STATE_ADDRESS_BIT_5 = 6;
  // localparam STATE_ADDRESS_BIT_6 = 7;
  // localparam STATE_ADDRESS_BIT_7 = 8;
  // localparam STATE_ADDRESS_BIT_8 = 9;
  // localparam STATE_ADDRESS_START = 1;
  // localparam STATE_ADDRESS_START_2 = 111;
  // localparam STATE_ADDRESS_START_3 = 112;
  // localparam STATE_DATA_ACK = 28;
  // localparam STATE_DATA_BIT_1 = 20;
  // localparam STATE_DATA_BIT_2 = 21;
  // localparam STATE_DATA_BIT_3 = 22;
  // localparam STATE_DATA_BIT_4 = 23;
  // localparam STATE_DATA_BIT_5 = 24;
  // localparam STATE_DATA_BIT_6 = 25;
  // localparam STATE_DATA_BIT_7 = 26;
  // localparam STATE_DATA_BIT_8 = 27;
  // localparam STATE_IDLE = 0;
  // localparam STATE_REG_ACK = 19;
  // localparam STATE_REG_BIT_1 = 11;
  // localparam STATE_REG_BIT_2 = 12;
  // localparam STATE_REG_BIT_3 = 13;
  // localparam STATE_REG_BIT_4 = 14;
  // localparam STATE_REG_BIT_5 = 15;
  // localparam STATE_REG_BIT_6 = 16;
  // localparam STATE_REG_BIT_7 = 17;
  // localparam STATE_REG_BIT_8 = 18;
  // localparam STATE_STOP = 29;
  // localparam STATE_STOP_1 = 30;
  // localparam STATE_STOP_2 = 31;
  // localparam STATE_TRANSIT_1 = 102;
  // localparam STATE_TRANSIT_2 = 192;
  wire [7:0] control_reg;  // sources/rtl/i2c_module.v(85)
  wire [7:0] divider2;  // sources/rtl/i2c_module.v(71)
  wire [7:0] n1;
  wire [7:0] n99;
  wire  \sel0_b0/B1 ;
  wire  \sel0_b0/B35 ;
  wire  \sel0_b1/B10 ;
  wire  \sel0_b1/B23 ;
  wire  \sel0_b2/B11 ;
  wire  \sel0_b2/B12 ;
  wire  \sel0_b2/B20 ;
  wire  \sel0_b2/B21 ;
  wire  \sel0_b2/B29 ;
  wire  \sel0_b2/B3 ;
  wire  \sel0_b2/B4 ;
  wire  \sel0_b3/B22 ;
  wire  \sel0_b3/B26 ;
  wire  \sel0_b3/B8 ;
  wire  \sel0_b4/B16 ;
  wire  \sel0_b4/B17 ;
  wire  \sel0_b4/B9 ;
  wire  \sel0_b5/B34 ;
  wire  \sel1/B33 ;
  wire  \sel5/B3 ;
  wire [7:0] slave_address;  // sources/rtl/i2c_module.v(86)
  wire [7:0] slave_data_1;  // sources/rtl/i2c_module.v(88)
  wire [7:0] slave_reg_address;  // sources/rtl/i2c_module.v(87)
  wire [7:0] state_next;  // sources/rtl/i2c_module.v(21)
  wire _al_u107_o;
  wire _al_u108_o;
  wire _al_u112_o;
  wire _al_u113_o;
  wire _al_u114_o;
  wire _al_u116_o;
  wire _al_u120_o;
  wire _al_u121_o;
  wire _al_u122_o;
  wire _al_u125_o;
  wire _al_u126_o;
  wire _al_u128_o;
  wire _al_u130_o;
  wire _al_u131_o;
  wire _al_u132_o;
  wire _al_u133_o;
  wire _al_u134_o;
  wire _al_u135_o;
  wire _al_u137_o;
  wire _al_u138_o;
  wire _al_u140_o;
  wire _al_u141_o;
  wire _al_u142_o;
  wire _al_u143_o;
  wire _al_u144_o;
  wire _al_u145_o;
  wire _al_u146_o;
  wire _al_u148_o;
  wire _al_u149_o;
  wire _al_u150_o;
  wire _al_u152_o;
  wire _al_u153_o;
  wire _al_u154_o;
  wire _al_u155_o;
  wire _al_u156_o;
  wire _al_u157_o;
  wire _al_u159_o;
  wire _al_u160_o;
  wire _al_u163_o;
  wire _al_u164_o;
  wire _al_u165_o;
  wire _al_u167_o;
  wire _al_u169_o;
  wire _al_u170_o;
  wire _al_u171_o;
  wire _al_u174_o;
  wire _al_u175_o;
  wire _al_u176_o;
  wire _al_u179_o;
  wire _al_u180_o;
  wire _al_u182_o;
  wire _al_u184_o;
  wire _al_u185_o;
  wire _al_u186_o;
  wire _al_u188_o;
  wire _al_u192_o;
  wire _al_u193_o;
  wire _al_u194_o;
  wire _al_u195_o;
  wire _al_u196_o;
  wire _al_u197_o;
  wire _al_u199_o;
  wire _al_u201_o;
  wire _al_u202_o;
  wire _al_u204_o;
  wire _al_u205_o;
  wire _al_u206_o;
  wire _al_u207_o;
  wire _al_u208_o;
  wire _al_u209_o;
  wire _al_u210_o;
  wire _al_u211_o;
  wire _al_u212_o;
  wire _al_u213_o;
  wire _al_u214_o;
  wire _al_u215_o;
  wire _al_u216_o;
  wire _al_u218_o;
  wire _al_u220_o;
  wire _al_u221_o;
  wire _al_u222_o;
  wire _al_u223_o;
  wire _al_u225_o;
  wire _al_u226_o;
  wire _al_u227_o;
  wire _al_u228_o;
  wire _al_u230_o;
  wire _al_u231_o;
  wire _al_u232_o;
  wire _al_u233_o;
  wire _al_u234_o;
  wire _al_u235_o;
  wire _al_u237_o;
  wire _al_u238_o;
  wire _al_u240_o;
  wire _al_u242_o;
  wire _al_u243_o;
  wire _al_u244_o;
  wire _al_u245_o;
  wire _al_u246_o;
  wire _al_u247_o;
  wire _al_u248_o;
  wire _al_u249_o;
  wire _al_u250_o;
  wire _al_u252_o;
  wire _al_u254_o;
  wire _al_u257_o;
  wire _al_u258_o;
  wire _al_u259_o;
  wire _al_u260_o;
  wire _al_u262_o;
  wire _al_u263_o;
  wire _al_u264_o;
  wire _al_u265_o;
  wire _al_u267_o;
  wire _al_u268_o;
  wire _al_u271_o;
  wire _al_u272_o;
  wire _al_u273_o;
  wire _al_u275_o;
  wire _al_u276_o;
  wire _al_u277_o;
  wire _al_u279_o;
  wire _al_u280_o;
  wire _al_u281_o;
  wire _al_u282_o;
  wire _al_u283_o;
  wire _al_u284_o;
  wire _al_u285_o;
  wire _al_u286_o;
  wire _al_u287_o;
  wire _al_u288_o;
  wire _al_u289_o;
  wire _al_u290_o;
  wire _al_u291_o;
  wire _al_u293_o;
  wire _al_u294_o;
  wire _al_u295_o;
  wire _al_u296_o;
  wire _al_u297_o;
  wire _al_u298_o;
  wire _al_u299_o;
  wire _al_u300_o;
  wire _al_u301_o;
  wire _al_u302_o;
  wire _al_u303_o;
  wire _al_u304_o;
  wire _al_u307_o;
  wire _al_u308_o;
  wire _al_u310_o;
  wire _al_u311_o;
  wire ack_ok;  // sources/rtl/i2c_module.v(143)
  wire \add0/c0 ;
  wire \add0/c1 ;
  wire \add0/c2 ;
  wire \add0/c3 ;
  wire \add0/c4 ;
  wire \add0/c5 ;
  wire \add0/c6 ;
  wire \add0/c7 ;
  wire clk_div_neg;
  wire mux4_b0_sel_is_3_o;
  wire mux5_b0_sel_is_3_o;
  wire mux6_b0_sel_is_3_o;
  wire mux7_b0_sel_is_3_o;
  wire mux9_b0_sel_is_0_o;
  wire n106_lutinv;
  wire n107_lutinv;
  wire n146_lutinv;
  wire n155_lutinv;
  wire n158_lutinv;
  wire n164_lutinv;
  wire n168_lutinv;
  wire n169_lutinv;
  wire n180_lutinv;
  wire n181_lutinv;
  wire n183_lutinv;
  wire n184;
  wire n186;
  wire n188;
  wire n190;
  wire n191_lutinv;
  wire n192;
  wire n194;
  wire n2;
  wire n20;
  wire n28;
  wire n29;
  wire n33;
  wire n80_lutinv;
  wire n81_lutinv;
  wire n88_lutinv;
  wire n94_lutinv;
  wire scl_output_enable;  // sources/rtl/i2c_module.v(120)
  wire scl_output_zero;  // sources/rtl/i2c_module.v(121)
  wire \sel0_b3/or_or_B13_B14_o_or_B_o_lutinv ;
  wire success;  // sources/rtl/i2c_module.v(141)

  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u103 (
    .a(address[1]),
    .b(address[0]),
    .c(write),
    .o(mux4_b0_sel_is_3_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    _al_u104 (
    .a(address[1]),
    .b(address[0]),
    .c(write),
    .o(mux6_b0_sel_is_3_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    _al_u105 (
    .a(address[1]),
    .b(address[0]),
    .c(write),
    .o(mux7_b0_sel_is_3_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u106 (
    .a(address[1]),
    .b(address[0]),
    .c(write),
    .o(mux5_b0_sel_is_3_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u107 (
    .a(state_next[4]),
    .b(state_next[5]),
    .c(state_next[6]),
    .d(state_next[7]),
    .o(_al_u107_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u108 (
    .a(state_next[0]),
    .b(state_next[1]),
    .c(state_next[2]),
    .d(state_next[3]),
    .o(_al_u108_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u109 (
    .a(_al_u107_o),
    .b(_al_u108_o),
    .o(n146_lutinv));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u110 (
    .a(n146_lutinv),
    .b(reset_n),
    .o(mux9_b0_sel_is_0_o));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'h47))
    _al_u111 (
    .a(scl_out),
    .b(scl_output_enable),
    .c(scl_output_zero),
    .o(n20));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*A)"),
    .INIT(16'h0002))
    _al_u112 (
    .a(state_next[4]),
    .b(state_next[5]),
    .c(state_next[6]),
    .d(state_next[7]),
    .o(_al_u112_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u113 (
    .a(state_next[0]),
    .b(state_next[1]),
    .o(_al_u113_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u114 (
    .a(state_next[2]),
    .b(state_next[3]),
    .o(_al_u114_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u115 (
    .a(_al_u112_o),
    .b(_al_u113_o),
    .c(_al_u114_o),
    .o(\sel0_b2/B3 ));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*A)"),
    .INIT(16'h0002))
    _al_u116 (
    .a(state_next[0]),
    .b(state_next[1]),
    .c(state_next[2]),
    .d(state_next[3]),
    .o(_al_u116_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u117 (
    .a(_al_u107_o),
    .b(_al_u116_o),
    .o(\sel0_b0/B35 ));
  AL_MAP_LUT4 #(
    .EQN("~(~(C*~B)*~(D*A))"),
    .INIT(16'hba30))
    _al_u118 (
    .a(\sel0_b2/B3 ),
    .b(\sel0_b0/B35 ),
    .c(success_out),
    .d(success),
    .o(n33));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    _al_u119 (
    .a(_al_u112_o),
    .b(_al_u114_o),
    .c(state_next[0]),
    .d(state_next[1]),
    .o(\sel0_b2/B4 ));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*B*~A)"),
    .INIT(16'h0400))
    _al_u120 (
    .a(state_next[0]),
    .b(state_next[1]),
    .c(state_next[2]),
    .d(state_next[3]),
    .o(_al_u120_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    _al_u121 (
    .a(state_next[0]),
    .b(state_next[1]),
    .c(state_next[2]),
    .d(state_next[3]),
    .o(_al_u121_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u122 (
    .a(_al_u107_o),
    .b(_al_u112_o),
    .c(_al_u120_o),
    .d(_al_u121_o),
    .o(_al_u122_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~(B*~A))"),
    .INIT(16'h0b00))
    _al_u123 (
    .a(\sel0_b2/B4 ),
    .b(_al_u122_o),
    .c(sda_in),
    .d(n28),
    .o(n29));
  AL_MAP_LUT4 #(
    .EQN("(B*A*(D@C))"),
    .INIT(16'h0880))
    _al_u124 (
    .a(_al_u107_o),
    .b(_al_u114_o),
    .c(state_next[0]),
    .d(state_next[1]),
    .o(n88_lutinv));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u125 (
    .a(state_next[2]),
    .b(state_next[3]),
    .o(_al_u125_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u126 (
    .a(state_next[0]),
    .b(state_next[1]),
    .o(_al_u126_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u127 (
    .a(_al_u107_o),
    .b(_al_u125_o),
    .c(_al_u126_o),
    .o(\sel0_b3/B22 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u128 (
    .a(state_next[0]),
    .b(state_next[1]),
    .o(_al_u128_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u129 (
    .a(_al_u128_o),
    .b(_al_u107_o),
    .c(_al_u114_o),
    .o(\sel0_b2/B21 ));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u130 (
    .a(n88_lutinv),
    .b(\sel0_b3/B22 ),
    .c(\sel0_b2/B21 ),
    .o(_al_u130_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*~A)"),
    .INIT(16'h0100))
    _al_u131 (
    .a(state_next[0]),
    .b(state_next[1]),
    .c(state_next[2]),
    .d(state_next[3]),
    .o(_al_u131_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*A)"),
    .INIT(16'h0080))
    _al_u132 (
    .a(state_next[0]),
    .b(state_next[1]),
    .c(state_next[2]),
    .d(state_next[3]),
    .o(_al_u132_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u133 (
    .a(state_next[0]),
    .b(state_next[1]),
    .c(state_next[3]),
    .o(_al_u133_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(~D*~C*~B))"),
    .INIT(16'haaa8))
    _al_u134 (
    .a(_al_u107_o),
    .b(_al_u131_o),
    .c(_al_u132_o),
    .d(_al_u133_o),
    .o(_al_u134_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*~B*~A)"),
    .INIT(16'h0010))
    _al_u135 (
    .a(state_next[0]),
    .b(state_next[1]),
    .c(state_next[2]),
    .d(state_next[3]),
    .o(_al_u135_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*~B))"),
    .INIT(8'ha8))
    _al_u136 (
    .a(_al_u107_o),
    .b(_al_u121_o),
    .c(_al_u135_o),
    .o(n80_lutinv));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*~A)"),
    .INIT(16'h0040))
    _al_u137 (
    .a(state_next[0]),
    .b(state_next[1]),
    .c(state_next[2]),
    .d(state_next[3]),
    .o(_al_u137_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*~B*A)"),
    .INIT(16'h0020))
    _al_u138 (
    .a(state_next[0]),
    .b(state_next[1]),
    .c(state_next[2]),
    .d(state_next[3]),
    .o(_al_u138_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*~B))"),
    .INIT(8'ha8))
    _al_u139 (
    .a(_al_u107_o),
    .b(_al_u137_o),
    .c(_al_u138_o),
    .o(n81_lutinv));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*~A)"),
    .INIT(16'h0004))
    _al_u140 (
    .a(state_next[0]),
    .b(state_next[1]),
    .c(state_next[2]),
    .d(state_next[3]),
    .o(_al_u140_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*A)"),
    .INIT(16'h0080))
    _al_u141 (
    .a(state_next[4]),
    .b(state_next[5]),
    .c(state_next[6]),
    .d(state_next[7]),
    .o(_al_u141_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*C)*~(B*A))"),
    .INIT(16'h0777))
    _al_u142 (
    .a(_al_u107_o),
    .b(_al_u140_o),
    .c(_al_u108_o),
    .d(_al_u141_o),
    .o(_al_u142_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*~A)"),
    .INIT(16'h0100))
    _al_u143 (
    .a(_al_u134_o),
    .b(n80_lutinv),
    .c(n81_lutinv),
    .d(_al_u142_o),
    .o(_al_u143_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*~A)"),
    .INIT(16'h1000))
    _al_u144 (
    .a(state_next[4]),
    .b(state_next[5]),
    .c(state_next[6]),
    .d(state_next[7]),
    .o(_al_u144_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*C)*~(B*A))"),
    .INIT(16'h0777))
    _al_u145 (
    .a(_al_u112_o),
    .b(_al_u138_o),
    .c(_al_u108_o),
    .d(_al_u144_o),
    .o(_al_u145_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*~B))"),
    .INIT(8'ha8))
    _al_u146 (
    .a(_al_u112_o),
    .b(_al_u135_o),
    .c(_al_u137_o),
    .o(_al_u146_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u147 (
    .a(_al_u112_o),
    .b(_al_u116_o),
    .o(\sel0_b4/B16 ));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u148 (
    .a(state_next[0]),
    .b(state_next[1]),
    .c(state_next[2]),
    .d(state_next[3]),
    .o(_al_u148_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u149 (
    .a(_al_u107_o),
    .b(_al_u112_o),
    .c(_al_u108_o),
    .d(_al_u148_o),
    .o(_al_u149_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*A)"),
    .INIT(16'h0200))
    _al_u150 (
    .a(_al_u145_o),
    .b(_al_u146_o),
    .c(\sel0_b4/B16 ),
    .d(_al_u149_o),
    .o(_al_u150_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u151 (
    .a(_al_u112_o),
    .b(_al_u132_o),
    .o(\sel0_b4/B9 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u152 (
    .a(_al_u112_o),
    .b(_al_u125_o),
    .o(_al_u152_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*~A)"),
    .INIT(16'h0040))
    _al_u153 (
    .a(state_next[4]),
    .b(state_next[5]),
    .c(state_next[6]),
    .d(state_next[7]),
    .o(_al_u153_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u154 (
    .a(_al_u112_o),
    .b(_al_u137_o),
    .c(_al_u140_o),
    .d(_al_u153_o),
    .o(_al_u154_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    _al_u155 (
    .a(\sel0_b4/B9 ),
    .b(_al_u152_o),
    .c(_al_u154_o),
    .o(_al_u155_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u156 (
    .a(_al_u130_o),
    .b(_al_u143_o),
    .c(_al_u150_o),
    .d(_al_u155_o),
    .o(_al_u156_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*~A)"),
    .INIT(16'h4000))
    _al_u157 (
    .a(state_next[0]),
    .b(state_next[1]),
    .c(state_next[2]),
    .d(state_next[3]),
    .o(_al_u157_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u158 (
    .a(_al_u112_o),
    .b(_al_u157_o),
    .o(n180_lutinv));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u159 (
    .a(\sel0_b0/B35 ),
    .b(n180_lutinv),
    .o(_al_u159_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~(B*A))"),
    .INIT(16'h7000))
    _al_u160 (
    .a(_al_u156_o),
    .b(_al_u159_o),
    .c(n28),
    .d(scl_output_zero),
    .o(_al_u160_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u161 (
    .a(_al_u112_o),
    .b(_al_u148_o),
    .o(n181_lutinv));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u162 (
    .a(_al_u148_o),
    .b(_al_u153_o),
    .o(\sel0_b5/B34 ));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(~D*~(~C*~A)))"),
    .INIT(16'h3301))
    _al_u163 (
    .a(\sel0_b2/B3 ),
    .b(n181_lutinv),
    .c(\sel0_b5/B34 ),
    .d(n28),
    .o(_al_u163_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u164 (
    .a(_al_u163_o),
    .b(\sel0_b5/B34 ),
    .c(scl_output_zero),
    .o(_al_u164_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*C)*~(B*~A))"),
    .INIT(16'hbb0b))
    _al_u165 (
    .a(\sel0_b2/B4 ),
    .b(_al_u122_o),
    .c(n28),
    .d(scl_output_zero),
    .o(_al_u165_o));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~B*~A)"),
    .INIT(8'hfe))
    _al_u166 (
    .a(_al_u160_o),
    .b(_al_u164_o),
    .c(_al_u165_o),
    .o(n194));
  AL_MAP_LUT4 #(
    .EQN("(~(D*C)*~(B*A))"),
    .INIT(16'h0777))
    _al_u167 (
    .a(_al_u107_o),
    .b(_al_u120_o),
    .c(_al_u137_o),
    .d(_al_u153_o),
    .o(_al_u167_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*~B))"),
    .INIT(8'ha8))
    _al_u168 (
    .a(_al_u112_o),
    .b(_al_u121_o),
    .c(_al_u140_o),
    .o(n94_lutinv));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*~B*~A)"),
    .INIT(16'h0010))
    _al_u169 (
    .a(\sel0_b4/B9 ),
    .b(_al_u152_o),
    .c(_al_u167_o),
    .d(n94_lutinv),
    .o(_al_u169_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u170 (
    .a(_al_u130_o),
    .b(_al_u143_o),
    .c(_al_u150_o),
    .d(_al_u169_o),
    .o(_al_u170_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~(B*A))"),
    .INIT(16'h7000))
    _al_u171 (
    .a(_al_u170_o),
    .b(_al_u159_o),
    .c(n28),
    .d(success),
    .o(_al_u171_o));
  AL_MAP_LUT4 #(
    .EQN("(A*(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C))"),
    .INIT(16'ha808))
    _al_u172 (
    .a(\sel0_b2/B4 ),
    .b(ack_ok),
    .c(n28),
    .d(success),
    .o(\sel5/B3 ));
  AL_MAP_LUT4 #(
    .EQN("~(~C*~A*~(D*~B))"),
    .INIT(16'hfbfa))
    _al_u173 (
    .a(_al_u171_o),
    .b(_al_u163_o),
    .c(\sel5/B3 ),
    .d(success),
    .o(n192));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*~A)"),
    .INIT(8'h04))
    _al_u174 (
    .a(\sel0_b0/B35 ),
    .b(_al_u122_o),
    .c(n180_lutinv),
    .o(_al_u174_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(A*~(C*~B)))"),
    .INIT(16'h7500))
    _al_u175 (
    .a(_al_u163_o),
    .b(_al_u174_o),
    .c(n28),
    .d(scl_output_enable),
    .o(_al_u175_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(B*~(~D*~C)))"),
    .INIT(16'h1115))
    _al_u176 (
    .a(_al_u175_o),
    .b(\sel0_b2/B4 ),
    .c(ack_ok),
    .d(n28),
    .o(_al_u176_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*C)*~(B*A))"),
    .INIT(16'h7707))
    _al_u177 (
    .a(_al_u176_o),
    .b(_al_u156_o),
    .c(n28),
    .d(scl_output_enable),
    .o(n188));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u178 (
    .a(_al_u112_o),
    .b(_al_u114_o),
    .o(n191_lutinv));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u179 (
    .a(n191_lutinv),
    .b(\sel0_b5/B34 ),
    .o(_al_u179_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u180 (
    .a(_al_u170_o),
    .b(_al_u179_o),
    .o(_al_u180_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u181 (
    .a(_al_u112_o),
    .b(_al_u121_o),
    .o(n168_lutinv));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u182 (
    .a(n168_lutinv),
    .b(ack_ok),
    .o(_al_u182_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((~B*~A))+C*D*~((~B*~A))+~(C)*D*(~B*~A)+C*D*(~B*~A))"),
    .INIT(16'hf1e0))
    _al_u183 (
    .a(_al_u180_o),
    .b(n28),
    .c(state_next[7]),
    .d(_al_u182_o),
    .o(n99[7]));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*~A)"),
    .INIT(8'h04))
    _al_u184 (
    .a(_al_u122_o),
    .b(ack_ok),
    .c(n28),
    .o(_al_u184_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(B)*~(A)+~C*B*~(A)+~(~C)*B*A+~C*B*A)"),
    .INIT(8'h8d))
    _al_u185 (
    .a(\sel0_b0/B35 ),
    .b(n28),
    .c(_al_u184_o),
    .o(_al_u185_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u186 (
    .a(\sel0_b5/B34 ),
    .b(_al_u185_o),
    .o(_al_u186_o));
  AL_MAP_LUT4 #(
    .EQN("~(D*~(B*~(~C*~A)))"),
    .INIT(16'hc8ff))
    _al_u187 (
    .a(_al_u180_o),
    .b(state_next[6]),
    .c(n28),
    .d(_al_u186_o),
    .o(n99[6]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u188 (
    .a(_al_u185_o),
    .b(state_next[5]),
    .o(_al_u188_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(~D*~C*~A))"),
    .INIT(16'h3332))
    _al_u189 (
    .a(_al_u180_o),
    .b(_al_u188_o),
    .c(n28),
    .d(state_next[3]),
    .o(n99[5]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u190 (
    .a(_al_u108_o),
    .b(_al_u144_o),
    .o(n169_lutinv));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u191 (
    .a(_al_u112_o),
    .b(_al_u108_o),
    .o(\sel0_b4/B17 ));
  AL_MAP_LUT4 #(
    .EQN("(A*~(~D*~C*~B))"),
    .INIT(16'haaa8))
    _al_u192 (
    .a(_al_u112_o),
    .b(_al_u116_o),
    .c(_al_u138_o),
    .d(_al_u140_o),
    .o(_al_u192_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u193 (
    .a(n169_lutinv),
    .b(_al_u146_o),
    .c(\sel0_b4/B17 ),
    .d(_al_u192_o),
    .o(_al_u193_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*A)"),
    .INIT(16'h0002))
    _al_u194 (
    .a(_al_u193_o),
    .b(\sel0_b2/B4 ),
    .c(\sel0_b4/B9 ),
    .d(_al_u152_o),
    .o(_al_u194_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u195 (
    .a(\sel0_b2/B3 ),
    .b(\sel0_b5/B34 ),
    .o(_al_u195_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h7735))
    _al_u196 (
    .a(_al_u194_o),
    .b(_al_u195_o),
    .c(n28),
    .d(state_next[4]),
    .o(_al_u196_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u197 (
    .a(_al_u122_o),
    .b(ack_ok),
    .c(n28),
    .o(_al_u197_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u198 (
    .a(_al_u107_o),
    .b(_al_u148_o),
    .o(n164_lutinv));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u199 (
    .a(n180_lutinv),
    .b(n164_lutinv),
    .c(n28),
    .o(_al_u199_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u200 (
    .a(_al_u112_o),
    .b(_al_u148_o),
    .c(n28),
    .o(\sel0_b0/B1 ));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*~A)"),
    .INIT(8'h04))
    _al_u201 (
    .a(_al_u197_o),
    .b(_al_u199_o),
    .c(\sel0_b0/B1 ),
    .o(_al_u201_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hd151))
    _al_u202 (
    .a(_al_u201_o),
    .b(n28),
    .c(state_next[4]),
    .d(state_next[5]),
    .o(_al_u202_o));
  AL_MAP_LUT4 #(
    .EQN("~(~C*~B*~(D*A))"),
    .INIT(16'hfefc))
    _al_u203 (
    .a(_al_u180_o),
    .b(_al_u196_o),
    .c(_al_u202_o),
    .d(state_next[4]),
    .o(n99[4]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*C)*~(B*A))"),
    .INIT(16'h0777))
    _al_u204 (
    .a(_al_u107_o),
    .b(_al_u133_o),
    .c(_al_u137_o),
    .d(_al_u153_o),
    .o(_al_u204_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*~B))"),
    .INIT(8'h8a))
    _al_u205 (
    .a(_al_u125_o),
    .b(state_next[0]),
    .c(state_next[1]),
    .o(_al_u205_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*~B*~A)"),
    .INIT(16'h0010))
    _al_u206 (
    .a(n88_lutinv),
    .b(\sel0_b2/B21 ),
    .c(_al_u204_o),
    .d(_al_u205_o),
    .o(_al_u206_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u207 (
    .a(_al_u206_o),
    .b(\sel0_b2/B4 ),
    .c(_al_u152_o),
    .o(_al_u207_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u208 (
    .a(_al_u207_o),
    .b(n28),
    .c(state_next[3]),
    .o(_al_u208_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(~B*~A))"),
    .INIT(8'he0))
    _al_u209 (
    .a(n180_lutinv),
    .b(n164_lutinv),
    .c(n28),
    .o(_al_u209_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*B))"),
    .INIT(8'ha2))
    _al_u210 (
    .a(_al_u197_o),
    .b(n28),
    .c(state_next[3]),
    .o(_al_u210_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u211 (
    .a(\sel0_b2/B3 ),
    .b(\sel0_b4/B9 ),
    .c(n28),
    .o(_al_u211_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*~B))"),
    .INIT(8'ha8))
    _al_u212 (
    .a(_al_u107_o),
    .b(_al_u116_o),
    .c(_al_u132_o),
    .o(_al_u212_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u213 (
    .a(_al_u212_o),
    .b(n28),
    .o(_al_u213_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(~B*~A))"),
    .INIT(8'h0e))
    _al_u214 (
    .a(n181_lutinv),
    .b(\sel0_b5/B34 ),
    .c(n28),
    .o(_al_u214_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u215 (
    .a(_al_u211_o),
    .b(_al_u213_o),
    .c(_al_u214_o),
    .o(_al_u215_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    _al_u216 (
    .a(_al_u209_o),
    .b(_al_u210_o),
    .c(_al_u215_o),
    .o(_al_u216_o));
  AL_MAP_LUT4 #(
    .EQN("~(C*~B*~(D*A))"),
    .INIT(16'hefcf))
    _al_u217 (
    .a(_al_u180_o),
    .b(_al_u208_o),
    .c(_al_u216_o),
    .d(state_next[3]),
    .o(n99[3]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u218 (
    .a(_al_u145_o),
    .b(_al_u146_o),
    .o(_al_u218_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u219 (
    .a(_al_u107_o),
    .b(_al_u120_o),
    .o(n158_lutinv));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u220 (
    .a(\sel0_b0/B35 ),
    .b(n158_lutinv),
    .c(n80_lutinv),
    .d(n81_lutinv),
    .o(_al_u220_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u221 (
    .a(_al_u125_o),
    .b(_al_u126_o),
    .o(_al_u221_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u222 (
    .a(\sel0_b2/B4 ),
    .b(_al_u221_o),
    .c(_al_u112_o),
    .o(_al_u222_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u223 (
    .a(_al_u130_o),
    .b(_al_u218_o),
    .c(_al_u220_o),
    .d(_al_u222_o),
    .o(_al_u223_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u224 (
    .a(n168_lutinv),
    .b(ack_ok),
    .c(n28),
    .o(\sel0_b3/or_or_B13_B14_o_or_B_o_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(~D*C*B))"),
    .INIT(16'h5515))
    _al_u225 (
    .a(\sel0_b2/B3 ),
    .b(n28),
    .c(state_next[2]),
    .d(state_next[0]),
    .o(_al_u225_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    _al_u226 (
    .a(\sel0_b3/or_or_B13_B14_o_or_B_o_lutinv ),
    .b(_al_u214_o),
    .c(_al_u225_o),
    .o(_al_u226_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    _al_u227 (
    .a(_al_u223_o),
    .b(_al_u226_o),
    .c(n28),
    .o(_al_u227_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u228 (
    .a(n28),
    .b(_al_u179_o),
    .o(_al_u228_o));
  AL_MAP_LUT4 #(
    .EQN("~(B*~(D*~(~C*~A)))"),
    .INIT(16'hfb33))
    _al_u229 (
    .a(_al_u180_o),
    .b(_al_u227_o),
    .c(_al_u228_o),
    .d(state_next[2]),
    .o(n99[2]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u230 (
    .a(n81_lutinv),
    .b(_al_u142_o),
    .o(_al_u230_o));
  AL_MAP_LUT3 #(
    .EQN("(A*(C@B))"),
    .INIT(8'h28))
    _al_u231 (
    .a(_al_u152_o),
    .b(state_next[0]),
    .c(state_next[1]),
    .o(_al_u231_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(~C*~B*A))"),
    .INIT(16'h00fd))
    _al_u232 (
    .a(_al_u230_o),
    .b(_al_u231_o),
    .c(\sel0_b0/B35 ),
    .d(n28),
    .o(_al_u232_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u233 (
    .a(\sel0_b2/B3 ),
    .b(n180_lutinv),
    .o(_al_u233_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*C)*~(B*~A))"),
    .INIT(16'h0bbb))
    _al_u234 (
    .a(_al_u233_o),
    .b(n28),
    .c(_al_u107_o),
    .d(_al_u184_o),
    .o(_al_u234_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u235 (
    .a(n88_lutinv),
    .b(_al_u204_o),
    .o(_al_u235_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u236 (
    .a(_al_u112_o),
    .b(_al_u137_o),
    .o(\sel0_b1/B10 ));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(~C*~B*A))"),
    .INIT(16'h00fd))
    _al_u237 (
    .a(_al_u235_o),
    .b(\sel0_b1/B10 ),
    .c(_al_u192_o),
    .d(n28),
    .o(_al_u237_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*~A)"),
    .INIT(16'h0004))
    _al_u238 (
    .a(_al_u232_o),
    .b(_al_u234_o),
    .c(_al_u237_o),
    .d(_al_u214_o),
    .o(_al_u238_o));
  AL_MAP_LUT4 #(
    .EQN("~(B*~(C*~(~D*~A)))"),
    .INIT(16'hf3b3))
    _al_u239 (
    .a(_al_u180_o),
    .b(_al_u238_o),
    .c(state_next[1]),
    .d(_al_u228_o),
    .o(n99[1]));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u240 (
    .a(\sel0_b2/B4 ),
    .b(_al_u152_o),
    .c(state_next[0]),
    .o(_al_u240_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u241 (
    .a(_al_u107_o),
    .b(_al_u131_o),
    .o(\sel0_b3/B26 ));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u242 (
    .a(\sel0_b2/B21 ),
    .b(\sel0_b3/B26 ),
    .c(_al_u146_o),
    .o(_al_u242_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*~B))"),
    .INIT(8'ha8))
    _al_u243 (
    .a(_al_u107_o),
    .b(_al_u135_o),
    .c(_al_u137_o),
    .o(_al_u243_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*~B))"),
    .INIT(8'ha8))
    _al_u244 (
    .a(_al_u107_o),
    .b(_al_u157_o),
    .c(_al_u140_o),
    .o(_al_u244_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*~A)"),
    .INIT(16'h0004))
    _al_u245 (
    .a(\sel0_b4/B17 ),
    .b(_al_u154_o),
    .c(_al_u243_o),
    .d(_al_u244_o),
    .o(_al_u245_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*~A)"),
    .INIT(16'h4000))
    _al_u246 (
    .a(_al_u197_o),
    .b(_al_u240_o),
    .c(_al_u242_o),
    .d(_al_u245_o),
    .o(_al_u246_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~(~B*~A))"),
    .INIT(16'h0e00))
    _al_u247 (
    .a(n191_lutinv),
    .b(\sel0_b5/B34 ),
    .c(n28),
    .d(state_next[0]),
    .o(_al_u247_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u248 (
    .a(_al_u247_o),
    .b(n146_lutinv),
    .c(control_reg[0]),
    .o(_al_u248_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u249 (
    .a(n28),
    .b(state_next[0]),
    .o(_al_u249_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~C*~(~D*A)))"),
    .INIT(16'hc0c8))
    _al_u250 (
    .a(_al_u246_o),
    .b(_al_u248_o),
    .c(_al_u249_o),
    .d(_al_u228_o),
    .o(_al_u250_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C*A))"),
    .INIT(8'hb3))
    _al_u251 (
    .a(_al_u180_o),
    .b(_al_u250_o),
    .c(state_next[0]),
    .o(n99[0]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u252 (
    .a(_al_u114_o),
    .b(state_next[0]),
    .o(_al_u252_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u253 (
    .a(n28),
    .b(ready),
    .o(n107_lutinv));
  AL_MAP_LUT4 #(
    .EQN("(D*~(~C*~B*A))"),
    .INIT(16'hfd00))
    _al_u254 (
    .a(_al_u170_o),
    .b(\sel0_b0/B35 ),
    .c(_al_u252_o),
    .d(n107_lutinv),
    .o(_al_u254_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u255 (
    .a(_al_u170_o),
    .b(_al_u179_o),
    .c(\sel0_b0/B35 ),
    .o(n183_lutinv));
  AL_MAP_LUT4 #(
    .EQN("~(~B*~A*~(D*~C))"),
    .INIT(16'hefee))
    _al_u256 (
    .a(_al_u254_o),
    .b(n183_lutinv),
    .c(_al_u163_o),
    .d(ready),
    .o(n190));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u257 (
    .a(n80_lutinv),
    .b(_al_u149_o),
    .o(_al_u257_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u258 (
    .a(_al_u218_o),
    .b(_al_u231_o),
    .c(_al_u257_o),
    .o(_al_u258_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u259 (
    .a(_al_u116_o),
    .b(_al_u132_o),
    .o(_al_u259_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    _al_u260 (
    .a(_al_u252_o),
    .b(_al_u167_o),
    .c(_al_u259_o),
    .o(_al_u260_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u261 (
    .a(_al_u112_o),
    .b(_al_u131_o),
    .o(\sel0_b3/B8 ));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u262 (
    .a(n168_lutinv),
    .b(\sel0_b3/B26 ),
    .c(\sel0_b3/B8 ),
    .o(_al_u262_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u263 (
    .a(_al_u130_o),
    .b(_al_u230_o),
    .c(_al_u260_o),
    .d(_al_u262_o),
    .o(_al_u263_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(B*A))"),
    .INIT(8'h07))
    _al_u264 (
    .a(_al_u258_o),
    .b(_al_u263_o),
    .c(n28),
    .o(_al_u264_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf5d0))
    _al_u265 (
    .a(_al_u195_o),
    .b(n181_lutinv),
    .c(sda_oe),
    .d(n28),
    .o(_al_u265_o));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~B*~A)"),
    .INIT(8'hfe))
    _al_u266 (
    .a(n183_lutinv),
    .b(_al_u264_o),
    .c(_al_u265_o),
    .o(n186));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u267 (
    .a(n28),
    .b(slave_address[7]),
    .o(_al_u267_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u268 (
    .a(_al_u267_o),
    .b(_al_u141_o),
    .o(_al_u268_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u269 (
    .a(_al_u107_o),
    .b(_al_u113_o),
    .c(_al_u114_o),
    .o(\sel0_b2/B20 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u270 (
    .a(_al_u107_o),
    .b(_al_u138_o),
    .o(\sel0_b2/B29 ));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u271 (
    .a(n28),
    .b(slave_address[3]),
    .o(_al_u271_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u272 (
    .a(n28),
    .b(slave_reg_address[4]),
    .o(_al_u272_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u273 (
    .a(\sel0_b2/B20 ),
    .b(\sel0_b2/B29 ),
    .c(_al_u271_o),
    .d(_al_u272_o),
    .o(_al_u273_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u274 (
    .a(_al_u137_o),
    .b(_al_u153_o),
    .o(\sel0_b1/B23 ));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u275 (
    .a(n28),
    .b(slave_address[2]),
    .o(_al_u275_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u276 (
    .a(_al_u107_o),
    .b(_al_u137_o),
    .c(_al_u275_o),
    .o(_al_u276_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D*~C*A))"),
    .INIT(16'h3133))
    _al_u277 (
    .a(\sel0_b1/B23 ),
    .b(_al_u276_o),
    .c(n28),
    .d(slave_reg_address[7]),
    .o(_al_u277_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u278 (
    .a(_al_u112_o),
    .b(_al_u138_o),
    .o(\sel0_b2/B11 ));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u279 (
    .a(n28),
    .b(slave_data_1[5]),
    .o(_al_u279_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u280 (
    .a(n28),
    .b(slave_data_1[4]),
    .o(_al_u280_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u281 (
    .a(\sel0_b2/B11 ),
    .b(\sel0_b1/B10 ),
    .c(_al_u279_o),
    .d(_al_u280_o),
    .o(_al_u281_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*~A)"),
    .INIT(16'h4000))
    _al_u282 (
    .a(_al_u268_o),
    .b(_al_u273_o),
    .c(_al_u277_o),
    .d(_al_u281_o),
    .o(_al_u282_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u283 (
    .a(n28),
    .b(slave_address[0]),
    .o(_al_u283_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u284 (
    .a(\sel0_b3/B26 ),
    .b(_al_u283_o),
    .o(_al_u284_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u285 (
    .a(n28),
    .b(slave_reg_address[3]),
    .o(_al_u285_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u286 (
    .a(n28),
    .b(slave_address[6]),
    .o(_al_u286_o));
  AL_MAP_LUT4 #(
    .EQN("~((D*B)*~(A)*~(C)+(D*B)*A*~(C)+~((D*B))*A*C+(D*B)*A*C)"),
    .INIT(16'h535f))
    _al_u287 (
    .a(_al_u285_o),
    .b(_al_u286_o),
    .c(_al_u157_o),
    .d(_al_u244_o),
    .o(_al_u287_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u288 (
    .a(_al_u113_o),
    .b(n28),
    .c(slave_data_1[1]),
    .o(_al_u288_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u289 (
    .a(n28),
    .b(slave_data_1[2]),
    .o(_al_u289_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u290 (
    .a(_al_u152_o),
    .b(\sel0_b3/B8 ),
    .c(_al_u288_o),
    .d(_al_u289_o),
    .o(_al_u290_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    _al_u291 (
    .a(_al_u284_o),
    .b(_al_u287_o),
    .c(_al_u290_o),
    .o(_al_u291_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u292 (
    .a(\sel0_b5/B34 ),
    .b(n28),
    .c(sda),
    .o(\sel1/B33 ));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u293 (
    .a(_al_u282_o),
    .b(_al_u291_o),
    .c(\sel1/B33 ),
    .o(_al_u293_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u294 (
    .a(_al_u107_o),
    .b(_al_u121_o),
    .c(slave_address[5]),
    .o(_al_u294_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u295 (
    .a(_al_u107_o),
    .b(_al_u135_o),
    .c(slave_address[4]),
    .o(_al_u295_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~B*~(D*A))"),
    .INIT(16'h0103))
    _al_u296 (
    .a(\sel0_b3/B22 ),
    .b(_al_u294_o),
    .c(_al_u295_o),
    .d(slave_reg_address[6]),
    .o(_al_u296_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(A*~(D*B)))"),
    .INIT(16'h0d05))
    _al_u297 (
    .a(_al_u296_o),
    .b(\sel0_b2/B21 ),
    .c(n28),
    .d(slave_reg_address[5]),
    .o(_al_u297_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u298 (
    .a(\sel0_b4/B16 ),
    .b(\sel0_b4/B9 ),
    .c(slave_reg_address[0]),
    .d(slave_data_1[3]),
    .o(_al_u298_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(~B*~(~C*A)))"),
    .INIT(16'hce00))
    _al_u299 (
    .a(\sel0_b2/B3 ),
    .b(n181_lutinv),
    .c(n28),
    .d(sda),
    .o(_al_u299_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u300 (
    .a(_al_u120_o),
    .b(n28),
    .c(slave_data_1[0]),
    .o(_al_u300_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u301 (
    .a(_al_u152_o),
    .b(_al_u300_o),
    .o(_al_u301_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~B*~(~D*~A))"),
    .INIT(16'h0302))
    _al_u302 (
    .a(_al_u298_o),
    .b(_al_u299_o),
    .c(_al_u301_o),
    .d(n28),
    .o(_al_u302_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u303 (
    .a(n180_lutinv),
    .b(\sel0_b4/B17 ),
    .c(slave_reg_address[1]),
    .o(_al_u303_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u304 (
    .a(n169_lutinv),
    .b(n164_lutinv),
    .c(slave_reg_address[2]),
    .d(slave_data_1[7]),
    .o(_al_u304_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u305 (
    .a(_al_u107_o),
    .b(_al_u132_o),
    .o(n155_lutinv));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u306 (
    .a(_al_u112_o),
    .b(_al_u135_o),
    .o(\sel0_b2/B12 ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u307 (
    .a(n155_lutinv),
    .b(\sel0_b2/B12 ),
    .c(slave_address[1]),
    .d(slave_data_1[6]),
    .o(_al_u307_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(C*B*A))"),
    .INIT(16'h007f))
    _al_u308 (
    .a(_al_u303_o),
    .b(_al_u304_o),
    .c(_al_u307_o),
    .d(n28),
    .o(_al_u308_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u309 (
    .a(n28),
    .b(sda),
    .o(n106_lutinv));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u310 (
    .a(n106_lutinv),
    .b(_al_u195_o),
    .o(_al_u310_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*~A)"),
    .INIT(16'h0004))
    _al_u311 (
    .a(_al_u297_o),
    .b(_al_u302_o),
    .c(_al_u308_o),
    .d(_al_u310_o),
    .o(_al_u311_o));
  AL_MAP_LUT3 #(
    .EQN("~(C*B*~A)"),
    .INIT(8'hbf))
    _al_u312 (
    .a(n183_lutinv),
    .b(_al_u293_o),
    .c(_al_u311_o),
    .o(n184));
  AL_MAP_LUT1 #(
    .EQN("(~A)"),
    .INIT(2'h1))
    _al_u313 (
    .a(reset_n),
    .o(n2));
  AL_MAP_LUT1 #(
    .EQN("(~A)"),
    .INIT(2'h1))
    _al_u314 (
    .a(n28),
    .o(clk_div_neg));
  reg_ar_as_w1 ack_ok_reg (
    .clk(divider2[7]),
    .d(n29),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(ack_ok));  // sources/rtl/i2c_module.v(153)
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add0/u0  (
    .a(divider2[0]),
    .b(1'b1),
    .c(\add0/c0 ),
    .o({\add0/c1 ,n1[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add0/u1  (
    .a(divider2[1]),
    .b(1'b0),
    .c(\add0/c1 ),
    .o({\add0/c2 ,n1[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add0/u2  (
    .a(divider2[2]),
    .b(1'b0),
    .c(\add0/c2 ),
    .o({\add0/c3 ,n1[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add0/u3  (
    .a(divider2[3]),
    .b(1'b0),
    .c(\add0/c3 ),
    .o({\add0/c4 ,n1[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add0/u4  (
    .a(divider2[4]),
    .b(1'b0),
    .c(\add0/c4 ),
    .o({\add0/c5 ,n1[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add0/u5  (
    .a(divider2[5]),
    .b(1'b0),
    .c(\add0/c5 ),
    .o({\add0/c6 ,n1[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add0/u6  (
    .a(divider2[6]),
    .b(1'b0),
    .c(\add0/c6 ),
    .o({\add0/c7 ,n1[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add0/u7  (
    .a(divider2[7]),
    .b(1'b0),
    .c(\add0/c7 ),
    .o({open_n0,n1[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \add0/ucin  (
    .a(1'b0),
    .o({\add0/c0 ,open_n3}));
  reg_ar_as_w1 clk_div_reg (
    .clk(divider2[7]),
    .d(clk_div_neg),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(n28));  // sources/rtl/i2c_module.v(76)
  reg_ar_ss_w1 ready_reg (
    .clk(~divider2[7]),
    .d(n190),
    .en(1'b1),
    .reset(1'b0),
    .set(~reset_n),
    .q(ready));  // sources/rtl/i2c_module.v(1066)
  reg_ar_as_w1 reg0_b0 (
    .clk(clk),
    .d(n1[0]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(divider2[0]));  // sources/rtl/i2c_module.v(81)
  reg_ar_as_w1 reg0_b1 (
    .clk(clk),
    .d(n1[1]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(divider2[1]));  // sources/rtl/i2c_module.v(81)
  reg_ar_as_w1 reg0_b2 (
    .clk(clk),
    .d(n1[2]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(divider2[2]));  // sources/rtl/i2c_module.v(81)
  reg_ar_as_w1 reg0_b3 (
    .clk(clk),
    .d(n1[3]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(divider2[3]));  // sources/rtl/i2c_module.v(81)
  reg_ar_as_w1 reg0_b4 (
    .clk(clk),
    .d(n1[4]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(divider2[4]));  // sources/rtl/i2c_module.v(81)
  reg_ar_as_w1 reg0_b5 (
    .clk(clk),
    .d(n1[5]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(divider2[5]));  // sources/rtl/i2c_module.v(81)
  reg_ar_as_w1 reg0_b6 (
    .clk(clk),
    .d(n1[6]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(divider2[6]));  // sources/rtl/i2c_module.v(81)
  reg_ar_as_w1 reg0_b7 (
    .clk(clk),
    .d(n1[7]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(divider2[7]));  // sources/rtl/i2c_module.v(81)
  reg_sr_as_w1 reg1_b0 (
    .clk(clk),
    .d(writedata[0]),
    .en(mux7_b0_sel_is_3_o),
    .reset(~mux9_b0_sel_is_0_o),
    .set(1'b0),
    .q(control_reg[0]));  // sources/rtl/i2c_module.v(117)
  reg_sr_as_w1 reg2_b0 (
    .clk(clk),
    .d(writedata[0]),
    .en(mux6_b0_sel_is_3_o),
    .reset(n2),
    .set(1'b0),
    .q(slave_address[0]));  // sources/rtl/i2c_module.v(117)
  reg_sr_as_w1 reg2_b1 (
    .clk(clk),
    .d(writedata[1]),
    .en(mux6_b0_sel_is_3_o),
    .reset(n2),
    .set(1'b0),
    .q(slave_address[1]));  // sources/rtl/i2c_module.v(117)
  reg_sr_as_w1 reg2_b2 (
    .clk(clk),
    .d(writedata[2]),
    .en(mux6_b0_sel_is_3_o),
    .reset(n2),
    .set(1'b0),
    .q(slave_address[2]));  // sources/rtl/i2c_module.v(117)
  reg_sr_as_w1 reg2_b3 (
    .clk(clk),
    .d(writedata[3]),
    .en(mux6_b0_sel_is_3_o),
    .reset(n2),
    .set(1'b0),
    .q(slave_address[3]));  // sources/rtl/i2c_module.v(117)
  reg_sr_as_w1 reg2_b4 (
    .clk(clk),
    .d(writedata[4]),
    .en(mux6_b0_sel_is_3_o),
    .reset(n2),
    .set(1'b0),
    .q(slave_address[4]));  // sources/rtl/i2c_module.v(117)
  reg_sr_as_w1 reg2_b5 (
    .clk(clk),
    .d(writedata[5]),
    .en(mux6_b0_sel_is_3_o),
    .reset(n2),
    .set(1'b0),
    .q(slave_address[5]));  // sources/rtl/i2c_module.v(117)
  reg_sr_as_w1 reg2_b6 (
    .clk(clk),
    .d(writedata[6]),
    .en(mux6_b0_sel_is_3_o),
    .reset(n2),
    .set(1'b0),
    .q(slave_address[6]));  // sources/rtl/i2c_module.v(117)
  reg_sr_as_w1 reg2_b7 (
    .clk(clk),
    .d(writedata[7]),
    .en(mux6_b0_sel_is_3_o),
    .reset(n2),
    .set(1'b0),
    .q(slave_address[7]));  // sources/rtl/i2c_module.v(117)
  reg_sr_as_w1 reg3_b0 (
    .clk(clk),
    .d(writedata[0]),
    .en(mux5_b0_sel_is_3_o),
    .reset(n2),
    .set(1'b0),
    .q(slave_reg_address[0]));  // sources/rtl/i2c_module.v(117)
  reg_sr_as_w1 reg3_b1 (
    .clk(clk),
    .d(writedata[1]),
    .en(mux5_b0_sel_is_3_o),
    .reset(n2),
    .set(1'b0),
    .q(slave_reg_address[1]));  // sources/rtl/i2c_module.v(117)
  reg_sr_as_w1 reg3_b2 (
    .clk(clk),
    .d(writedata[2]),
    .en(mux5_b0_sel_is_3_o),
    .reset(n2),
    .set(1'b0),
    .q(slave_reg_address[2]));  // sources/rtl/i2c_module.v(117)
  reg_sr_as_w1 reg3_b3 (
    .clk(clk),
    .d(writedata[3]),
    .en(mux5_b0_sel_is_3_o),
    .reset(n2),
    .set(1'b0),
    .q(slave_reg_address[3]));  // sources/rtl/i2c_module.v(117)
  reg_sr_as_w1 reg3_b4 (
    .clk(clk),
    .d(writedata[4]),
    .en(mux5_b0_sel_is_3_o),
    .reset(n2),
    .set(1'b0),
    .q(slave_reg_address[4]));  // sources/rtl/i2c_module.v(117)
  reg_sr_as_w1 reg3_b5 (
    .clk(clk),
    .d(writedata[5]),
    .en(mux5_b0_sel_is_3_o),
    .reset(n2),
    .set(1'b0),
    .q(slave_reg_address[5]));  // sources/rtl/i2c_module.v(117)
  reg_sr_as_w1 reg3_b6 (
    .clk(clk),
    .d(writedata[6]),
    .en(mux5_b0_sel_is_3_o),
    .reset(n2),
    .set(1'b0),
    .q(slave_reg_address[6]));  // sources/rtl/i2c_module.v(117)
  reg_sr_as_w1 reg3_b7 (
    .clk(clk),
    .d(writedata[7]),
    .en(mux5_b0_sel_is_3_o),
    .reset(n2),
    .set(1'b0),
    .q(slave_reg_address[7]));  // sources/rtl/i2c_module.v(117)
  reg_sr_as_w1 reg4_b0 (
    .clk(clk),
    .d(writedata[0]),
    .en(mux4_b0_sel_is_3_o),
    .reset(n2),
    .set(1'b0),
    .q(slave_data_1[0]));  // sources/rtl/i2c_module.v(117)
  reg_sr_as_w1 reg4_b1 (
    .clk(clk),
    .d(writedata[1]),
    .en(mux4_b0_sel_is_3_o),
    .reset(n2),
    .set(1'b0),
    .q(slave_data_1[1]));  // sources/rtl/i2c_module.v(117)
  reg_sr_as_w1 reg4_b2 (
    .clk(clk),
    .d(writedata[2]),
    .en(mux4_b0_sel_is_3_o),
    .reset(n2),
    .set(1'b0),
    .q(slave_data_1[2]));  // sources/rtl/i2c_module.v(117)
  reg_sr_as_w1 reg4_b3 (
    .clk(clk),
    .d(writedata[3]),
    .en(mux4_b0_sel_is_3_o),
    .reset(n2),
    .set(1'b0),
    .q(slave_data_1[3]));  // sources/rtl/i2c_module.v(117)
  reg_sr_as_w1 reg4_b4 (
    .clk(clk),
    .d(writedata[4]),
    .en(mux4_b0_sel_is_3_o),
    .reset(n2),
    .set(1'b0),
    .q(slave_data_1[4]));  // sources/rtl/i2c_module.v(117)
  reg_sr_as_w1 reg4_b5 (
    .clk(clk),
    .d(writedata[5]),
    .en(mux4_b0_sel_is_3_o),
    .reset(n2),
    .set(1'b0),
    .q(slave_data_1[5]));  // sources/rtl/i2c_module.v(117)
  reg_sr_as_w1 reg4_b6 (
    .clk(clk),
    .d(writedata[6]),
    .en(mux4_b0_sel_is_3_o),
    .reset(n2),
    .set(1'b0),
    .q(slave_data_1[6]));  // sources/rtl/i2c_module.v(117)
  reg_sr_as_w1 reg4_b7 (
    .clk(clk),
    .d(writedata[7]),
    .en(mux4_b0_sel_is_3_o),
    .reset(n2),
    .set(1'b0),
    .q(slave_data_1[7]));  // sources/rtl/i2c_module.v(117)
  reg_sr_as_w1 reg5_b0 (
    .clk(~divider2[7]),
    .d(n99[0]),
    .en(1'b1),
    .reset(n2),
    .set(1'b0),
    .q(state_next[0]));  // sources/rtl/i2c_module.v(510)
  reg_sr_as_w1 reg5_b1 (
    .clk(~divider2[7]),
    .d(n99[1]),
    .en(1'b1),
    .reset(n2),
    .set(1'b0),
    .q(state_next[1]));  // sources/rtl/i2c_module.v(510)
  reg_sr_as_w1 reg5_b2 (
    .clk(~divider2[7]),
    .d(n99[2]),
    .en(1'b1),
    .reset(n2),
    .set(1'b0),
    .q(state_next[2]));  // sources/rtl/i2c_module.v(510)
  reg_sr_as_w1 reg5_b3 (
    .clk(~divider2[7]),
    .d(n99[3]),
    .en(1'b1),
    .reset(n2),
    .set(1'b0),
    .q(state_next[3]));  // sources/rtl/i2c_module.v(510)
  reg_sr_as_w1 reg5_b4 (
    .clk(~divider2[7]),
    .d(n99[4]),
    .en(1'b1),
    .reset(n2),
    .set(1'b0),
    .q(state_next[4]));  // sources/rtl/i2c_module.v(510)
  reg_sr_as_w1 reg5_b5 (
    .clk(~divider2[7]),
    .d(n99[5]),
    .en(1'b1),
    .reset(n2),
    .set(1'b0),
    .q(state_next[5]));  // sources/rtl/i2c_module.v(510)
  reg_sr_as_w1 reg5_b6 (
    .clk(~divider2[7]),
    .d(n99[6]),
    .en(1'b1),
    .reset(n2),
    .set(1'b0),
    .q(state_next[6]));  // sources/rtl/i2c_module.v(510)
  reg_sr_as_w1 reg5_b7 (
    .clk(~divider2[7]),
    .d(n99[7]),
    .en(1'b1),
    .reset(n2),
    .set(1'b0),
    .q(state_next[7]));  // sources/rtl/i2c_module.v(510)
  reg_ar_as_w1 scl_out_reg (
    .clk(divider2[7]),
    .d(n20),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(scl_out));  // sources/rtl/i2c_module.v(137)
  reg_sr_as_w1 scl_output_enable_reg (
    .clk(~divider2[7]),
    .d(n188),
    .en(1'b1),
    .reset(~reset_n),
    .set(1'b0),
    .q(scl_output_enable));  // sources/rtl/i2c_module.v(1066)
  reg_ar_as_w1 scl_output_zero_reg (
    .clk(~divider2[7]),
    .d(n194),
    .en(~n2),
    .reset(1'b0),
    .set(1'b0),
    .q(scl_output_zero));  // sources/rtl/i2c_module.v(1066)
  reg_ar_ss_w1 sda_oe_reg (
    .clk(~divider2[7]),
    .d(n186),
    .en(1'b1),
    .reset(1'b0),
    .set(~reset_n),
    .q(sda_oe));  // sources/rtl/i2c_module.v(1066)
  reg_ar_ss_w1 sda_reg (
    .clk(~divider2[7]),
    .d(n184),
    .en(1'b1),
    .reset(1'b0),
    .set(~reset_n),
    .q(sda));  // sources/rtl/i2c_module.v(1066)
  reg_ar_as_w1 success_out_reg (
    .clk(~divider2[7]),
    .d(n33),
    .en(n28),
    .reset(1'b0),
    .set(1'b0),
    .q(success_out));  // sources/rtl/i2c_module.v(167)
  reg_sr_as_w1 success_reg (
    .clk(~divider2[7]),
    .d(n192),
    .en(1'b1),
    .reset(~reset_n),
    .set(1'b0),
    .q(success));  // sources/rtl/i2c_module.v(1066)

endmodule 

module reg_ar_ss_w1
  (
  clk,
  d,
  en,
  reset,
  set,
  q
  );

  input clk;
  input d;
  input en;
  input reset;
  input set;
  output q;

  parameter REGSET = "RESET";
  wire enout;
  wire setout;

  AL_MUX u_en0 (
    .i0(q),
    .i1(d),
    .sel(en),
    .o(enout));
  AL_DFF #(
    .INI((REGSET == "SET") ? 1'b1 : 1'b0))
    u_seq0 (
    .clk(clk),
    .d(setout),
    .reset(reset),
    .set(1'b0),
    .q(q));
  AL_MUX u_set0 (
    .i0(enout),
    .i1(1'b1),
    .sel(set),
    .o(setout));

endmodule 

module AL_MUX
  (
  input i0,
  input i1,
  input sel,
  output o
  );

  wire not_sel, sel_i0, sel_i1;
  not u0 (not_sel, sel);
  and u1 (sel_i1, sel, i1);
  and u2 (sel_i0, not_sel, i0);
  or u3 (o, sel_i1, sel_i0);

endmodule

module AL_DFF
  (
  input reset,
  input set,
  input clk,
  input d,
  output reg q
  );

  parameter INI = 1'b0;

  always @(posedge reset or posedge set or posedge clk)
  begin
    if (reset)
      q <= 1'b0;
    else if (set)
      q <= 1'b1;
    else
      q <= d;
  end

endmodule

