// Verilog netlist created by TD v4.6.12906
// Tue Jul 30 09:10:03 2019

`timescale 1ns / 1ps
module test_camera  // sources/rtl/test_camera.v(14)
  (
  cam_data,
  cam_href,
  cam_pclk,
  cam_vsync,
  clk_24m,
  rst_n,
  cam_pwdn,
  cam_rst,
  cam_soic,
  cam_xclk,
  vga_b,
  vga_clk,
  vga_g,
  vga_hsync,
  vga_r,
  vga_vsync,
  cam_soid
  );

  input [7:0] cam_data;  // sources/rtl/test_camera.v(27)
  input cam_href;  // sources/rtl/test_camera.v(21)
  input cam_pclk;  // sources/rtl/test_camera.v(19)
  input cam_vsync;  // sources/rtl/test_camera.v(22)
  input clk_24m;  // sources/rtl/test_camera.v(16)
  input rst_n;  // sources/rtl/test_camera.v(17)
  output cam_pwdn;  // sources/rtl/test_camera.v(23)
  output cam_rst;  // sources/rtl/test_camera.v(24)
  output cam_soic;  // sources/rtl/test_camera.v(25)
  output cam_xclk;  // sources/rtl/test_camera.v(20)
  output [7:0] vga_b;  // sources/rtl/test_camera.v(31)
  output vga_clk;  // sources/rtl/test_camera.v(32)
  output [7:0] vga_g;  // sources/rtl/test_camera.v(30)
  output vga_hsync;  // sources/rtl/test_camera.v(33)
  output [7:0] vga_r;  // sources/rtl/test_camera.v(29)
  output vga_vsync;  // sources/rtl/test_camera.v(34)
  inout cam_soid;  // sources/rtl/test_camera.v(26)

  wire [19:0] camera_addr;  // sources/rtl/test_camera.v(45)
  wire [15:0] camera_wrdat;  // sources/rtl/test_camera.v(44)
  wire [15:0] \u_camera_reader/current_pixel ;  // sources/rtl/camera_reader.v(37)
  wire [19:0] \u_camera_reader/n18 ;
  wire [19:0] \u_camera_reader/n19 ;
  wire [19:0] \u_camera_reader/n21 ;
  wire [19:0] \u_camera_reader/n8 ;
  wire [19:0] \u_camera_reader/n9 ;
  wire [19:0] \u_camera_reader/pixel_counter ;  // sources/rtl/camera_reader.v(32)
  wire [7:0] \u_camera_reader/subpixel ;  // sources/rtl/camera_reader.v(36)
  wire [15:0] vga_rdaddr;  // sources/rtl/test_camera.v(59)
  wire [15:0] vga_rddat;  // sources/rtl/test_camera.v(58)
  wire camera_wrreq;  // sources/rtl/test_camera.v(42)
  wire clk_cam;  // sources/rtl/test_camera.v(39)
  wire clk_lcd;  // sources/rtl/test_camera.v(38)
  wire clk_sccb;  // sources/rtl/test_camera.v(40)
  wire n0;
  wire n1;
  wire sda;  // sources/rtl/test_camera.v(50)
  wire sda_oe;  // sources/rtl/test_camera.v(49)
  wire \u_camera_reader/mux10_b0_sel_is_2_o ;
  wire \u_camera_reader/mux11_b0_sel_is_2_o ;
  wire \u_camera_reader/mux13_b0_sel_is_2_o ;
  wire \u_camera_reader/mux14_b0_sel_is_2_o ;
  wire \u_camera_reader/mux4_b0_sel_is_0_o ;
  wire \u_camera_reader/mux4_b0_sel_is_0_o_neg ;
  wire \u_camera_reader/mux5_b0_sel_is_3_o ;
  wire \u_camera_reader/mux6_b0_sel_is_1_o ;
  wire \u_camera_reader/mux8_b0_sel_is_0_o ;
  wire \u_camera_reader/n0 ;
  wire \u_camera_reader/n1 ;
  wire \u_camera_reader/n13 ;
  wire \u_camera_reader/n13_neg ;
  wire \u_camera_reader/n2 ;
  wire \u_camera_reader/n27 ;
  wire \u_camera_reader/n28 ;
  wire \u_camera_reader/n3 ;
  wire \u_camera_reader/n3_neg ;
  wire \u_camera_reader/n4 ;
  wire \u_camera_reader/n4_neg ;
  wire \u_camera_reader/n5 ;
  wire \u_camera_reader/n6 ;
  wire \u_camera_reader/n6_neg ;
  wire \u_camera_reader/n7 ;
  wire \u_camera_reader/n7_neg ;
  wire \u_camera_reader/vsync_passed ;  // sources/rtl/camera_reader.v(34)
  wire \u_camera_reader/wrclk1 ;  // sources/rtl/camera_reader.v(38)
  wire \u_camera_reader/write_pixel ;  // sources/rtl/camera_reader.v(35)
  wire \u_pll/clk0_buf ;  // al_ip/ip_pll.v(34)
  wire vga_rden;  // sources/rtl/test_camera.v(57)

  assign cam_rst = rst_n;
  assign cam_pwdn = 1'b0;
  assign vga_b[2] = 1'b0;
  assign vga_b[1] = 1'b0;
  assign vga_b[0] = 1'b0;
  assign vga_g[1] = 1'b0;
  assign vga_g[0] = 1'b0;
  assign vga_r[2] = 1'b0;
  assign vga_r[1] = 1'b0;
  assign vga_r[0] = 1'b0;
  binary_mux_s1_w1 mux0_b0 (
    .i0(1'b0),
    .i1(vga_rddat[11]),
    .sel(vga_rden),
    .o(vga_r[3]));  // sources/rtl/test_camera.v(67)
  binary_mux_s1_w1 mux0_b1 (
    .i0(1'b0),
    .i1(vga_rddat[12]),
    .sel(vga_rden),
    .o(vga_r[4]));  // sources/rtl/test_camera.v(67)
  binary_mux_s1_w1 mux0_b2 (
    .i0(1'b0),
    .i1(vga_rddat[13]),
    .sel(vga_rden),
    .o(vga_r[5]));  // sources/rtl/test_camera.v(67)
  binary_mux_s1_w1 mux0_b3 (
    .i0(1'b0),
    .i1(vga_rddat[14]),
    .sel(vga_rden),
    .o(vga_r[6]));  // sources/rtl/test_camera.v(67)
  binary_mux_s1_w1 mux0_b4 (
    .i0(1'b0),
    .i1(vga_rddat[15]),
    .sel(vga_rden),
    .o(vga_r[7]));  // sources/rtl/test_camera.v(67)
  binary_mux_s1_w1 mux1_b0 (
    .i0(1'b0),
    .i1(vga_rddat[5]),
    .sel(vga_rden),
    .o(vga_g[2]));  // sources/rtl/test_camera.v(68)
  binary_mux_s1_w1 mux1_b1 (
    .i0(1'b0),
    .i1(vga_rddat[6]),
    .sel(vga_rden),
    .o(vga_g[3]));  // sources/rtl/test_camera.v(68)
  binary_mux_s1_w1 mux1_b2 (
    .i0(1'b0),
    .i1(vga_rddat[7]),
    .sel(vga_rden),
    .o(vga_g[4]));  // sources/rtl/test_camera.v(68)
  binary_mux_s1_w1 mux1_b3 (
    .i0(1'b0),
    .i1(vga_rddat[8]),
    .sel(vga_rden),
    .o(vga_g[5]));  // sources/rtl/test_camera.v(68)
  binary_mux_s1_w1 mux1_b4 (
    .i0(1'b0),
    .i1(vga_rddat[9]),
    .sel(vga_rden),
    .o(vga_g[6]));  // sources/rtl/test_camera.v(68)
  binary_mux_s1_w1 mux1_b5 (
    .i0(1'b0),
    .i1(vga_rddat[10]),
    .sel(vga_rden),
    .o(vga_g[7]));  // sources/rtl/test_camera.v(68)
  binary_mux_s1_w1 mux2_b0 (
    .i0(1'b0),
    .i1(vga_rddat[0]),
    .sel(vga_rden),
    .o(vga_b[3]));  // sources/rtl/test_camera.v(69)
  binary_mux_s1_w1 mux2_b1 (
    .i0(1'b0),
    .i1(vga_rddat[1]),
    .sel(vga_rden),
    .o(vga_b[4]));  // sources/rtl/test_camera.v(69)
  binary_mux_s1_w1 mux2_b2 (
    .i0(1'b0),
    .i1(vga_rddat[2]),
    .sel(vga_rden),
    .o(vga_b[5]));  // sources/rtl/test_camera.v(69)
  binary_mux_s1_w1 mux2_b3 (
    .i0(1'b0),
    .i1(vga_rddat[3]),
    .sel(vga_rden),
    .o(vga_b[6]));  // sources/rtl/test_camera.v(69)
  binary_mux_s1_w1 mux2_b4 (
    .i0(1'b0),
    .i1(vga_rddat[4]),
    .sel(vga_rden),
    .o(vga_b[7]));  // sources/rtl/test_camera.v(69)
  not u13 (n0, cam_vsync);  // sources/rtl/test_camera.v(124)
  not u14 (n1, cam_rst);  // sources/rtl/test_camera.v(139)
  bufif1 u6 (cam_soid, sda, sda_oe);  // sources/rtl/test_camera.v(61)
  camera_init u_camera_init (
    .clk(clk_sccb),
    .reset_n(cam_rst),
    .sda_in(cam_soid),
    .scl(cam_soic),
    .sda(sda),
    .sda_oe(sda_oe));  // sources/rtl/test_camera.v(84)
  add_pu20_pu20_o20 \u_camera_reader/add0  (
    .i0(\u_camera_reader/pixel_counter ),
    .i1(20'b00000000000000000001),
    .o(\u_camera_reader/n8 ));  // sources/rtl/camera_reader.v(78)
  add_pu16_pu16_o16 \u_camera_reader/add1  (
    .i0(camera_addr[15:0]),
    .i1(16'b0000000000000001),
    .o(\u_camera_reader/n9 [15:0]));  // sources/rtl/camera_reader.v(85)
  eq_w1 \u_camera_reader/eq0  (
    .i0(cam_rst),
    .i1(1'b1),
    .o(\u_camera_reader/n0 ));  // sources/rtl/camera_reader.v(33)
  eq_w1 \u_camera_reader/eq1  (
    .i0(cam_href),
    .i1(1'b1),
    .o(\u_camera_reader/n2 ));  // sources/rtl/camera_reader.v(47)
  eq_w1 \u_camera_reader/eq2  (
    .i0(cam_rst),
    .i1(1'b0),
    .o(\u_camera_reader/n3 ));  // sources/rtl/camera_reader.v(60)
  eq_w1 \u_camera_reader/eq3  (
    .i0(n0),
    .i1(1'b1),
    .o(\u_camera_reader/n4 ));  // sources/rtl/camera_reader.v(67)
  eq_w1 \u_camera_reader/eq4  (
    .i0(\u_camera_reader/vsync_passed ),
    .i1(1'b1),
    .o(\u_camera_reader/n5 ));  // sources/rtl/camera_reader.v(74)
  eq_w1 \u_camera_reader/eq5  (
    .i0(\u_camera_reader/pixel_counter [0]),
    .i1(1'b0),
    .o(\u_camera_reader/n7 ));  // sources/rtl/camera_reader.v(76)
  eq_w1 \u_camera_reader/eq6  (
    .i0(\u_camera_reader/write_pixel ),
    .i1(1'b1),
    .o(\u_camera_reader/n13 ));  // sources/rtl/camera_reader.v(90)
  lt_u20_u20 \u_camera_reader/lt0  (
    .ci(1'b0),
    .i0(20'b00000000000000000010),
    .i1(\u_camera_reader/pixel_counter ),
    .o(\u_camera_reader/n27 ));  // sources/rtl/camera_reader.v(98)
  and \u_camera_reader/mux10_b0_sel_is_2  (\u_camera_reader/mux10_b0_sel_is_2_o , \u_camera_reader/n4_neg , \u_camera_reader/mux5_b0_sel_is_3_o );
  and \u_camera_reader/mux11_b0_sel_is_2  (\u_camera_reader/mux11_b0_sel_is_2_o , \u_camera_reader/n4_neg , \u_camera_reader/mux6_b0_sel_is_1_o );
  and \u_camera_reader/mux13_b0_sel_is_2  (\u_camera_reader/mux13_b0_sel_is_2_o , \u_camera_reader/n3_neg , \u_camera_reader/mux10_b0_sel_is_2_o );
  and \u_camera_reader/mux14_b0_sel_is_2  (\u_camera_reader/mux14_b0_sel_is_2_o , \u_camera_reader/n3_neg , \u_camera_reader/mux11_b0_sel_is_2_o );
  and \u_camera_reader/mux4_b0_sel_is_0  (\u_camera_reader/mux4_b0_sel_is_0_o , \u_camera_reader/n6_neg , \u_camera_reader/n13_neg );
  not \u_camera_reader/mux4_b0_sel_is_0_o_inv  (\u_camera_reader/mux4_b0_sel_is_0_o_neg , \u_camera_reader/mux4_b0_sel_is_0_o );
  and \u_camera_reader/mux5_b0_sel_is_3  (\u_camera_reader/mux5_b0_sel_is_3_o , \u_camera_reader/n6 , \u_camera_reader/n7 );
  and \u_camera_reader/mux6_b0_sel_is_1  (\u_camera_reader/mux6_b0_sel_is_1_o , \u_camera_reader/n6 , \u_camera_reader/n7_neg );
  AL_MUX \u_camera_reader/mux7_b0  (
    .i0(camera_addr[0]),
    .i1(\u_camera_reader/n9 [0]),
    .sel(\u_camera_reader/mux6_b0_sel_is_1_o ),
    .o(\u_camera_reader/n18 [0]));
  AL_MUX \u_camera_reader/mux7_b1  (
    .i0(camera_addr[1]),
    .i1(\u_camera_reader/n9 [1]),
    .sel(\u_camera_reader/mux6_b0_sel_is_1_o ),
    .o(\u_camera_reader/n18 [1]));
  AL_MUX \u_camera_reader/mux7_b10  (
    .i0(camera_addr[10]),
    .i1(\u_camera_reader/n9 [10]),
    .sel(\u_camera_reader/mux6_b0_sel_is_1_o ),
    .o(\u_camera_reader/n18 [10]));
  AL_MUX \u_camera_reader/mux7_b11  (
    .i0(camera_addr[11]),
    .i1(\u_camera_reader/n9 [11]),
    .sel(\u_camera_reader/mux6_b0_sel_is_1_o ),
    .o(\u_camera_reader/n18 [11]));
  AL_MUX \u_camera_reader/mux7_b12  (
    .i0(camera_addr[12]),
    .i1(\u_camera_reader/n9 [12]),
    .sel(\u_camera_reader/mux6_b0_sel_is_1_o ),
    .o(\u_camera_reader/n18 [12]));
  AL_MUX \u_camera_reader/mux7_b13  (
    .i0(camera_addr[13]),
    .i1(\u_camera_reader/n9 [13]),
    .sel(\u_camera_reader/mux6_b0_sel_is_1_o ),
    .o(\u_camera_reader/n18 [13]));
  AL_MUX \u_camera_reader/mux7_b14  (
    .i0(camera_addr[14]),
    .i1(\u_camera_reader/n9 [14]),
    .sel(\u_camera_reader/mux6_b0_sel_is_1_o ),
    .o(\u_camera_reader/n18 [14]));
  AL_MUX \u_camera_reader/mux7_b15  (
    .i0(camera_addr[15]),
    .i1(\u_camera_reader/n9 [15]),
    .sel(\u_camera_reader/mux6_b0_sel_is_1_o ),
    .o(\u_camera_reader/n18 [15]));
  AL_MUX \u_camera_reader/mux7_b2  (
    .i0(camera_addr[2]),
    .i1(\u_camera_reader/n9 [2]),
    .sel(\u_camera_reader/mux6_b0_sel_is_1_o ),
    .o(\u_camera_reader/n18 [2]));
  AL_MUX \u_camera_reader/mux7_b3  (
    .i0(camera_addr[3]),
    .i1(\u_camera_reader/n9 [3]),
    .sel(\u_camera_reader/mux6_b0_sel_is_1_o ),
    .o(\u_camera_reader/n18 [3]));
  AL_MUX \u_camera_reader/mux7_b4  (
    .i0(camera_addr[4]),
    .i1(\u_camera_reader/n9 [4]),
    .sel(\u_camera_reader/mux6_b0_sel_is_1_o ),
    .o(\u_camera_reader/n18 [4]));
  AL_MUX \u_camera_reader/mux7_b5  (
    .i0(camera_addr[5]),
    .i1(\u_camera_reader/n9 [5]),
    .sel(\u_camera_reader/mux6_b0_sel_is_1_o ),
    .o(\u_camera_reader/n18 [5]));
  AL_MUX \u_camera_reader/mux7_b6  (
    .i0(camera_addr[6]),
    .i1(\u_camera_reader/n9 [6]),
    .sel(\u_camera_reader/mux6_b0_sel_is_1_o ),
    .o(\u_camera_reader/n18 [6]));
  AL_MUX \u_camera_reader/mux7_b7  (
    .i0(camera_addr[7]),
    .i1(\u_camera_reader/n9 [7]),
    .sel(\u_camera_reader/mux6_b0_sel_is_1_o ),
    .o(\u_camera_reader/n18 [7]));
  AL_MUX \u_camera_reader/mux7_b8  (
    .i0(camera_addr[8]),
    .i1(\u_camera_reader/n9 [8]),
    .sel(\u_camera_reader/mux6_b0_sel_is_1_o ),
    .o(\u_camera_reader/n18 [8]));
  AL_MUX \u_camera_reader/mux7_b9  (
    .i0(camera_addr[9]),
    .i1(\u_camera_reader/n9 [9]),
    .sel(\u_camera_reader/mux6_b0_sel_is_1_o ),
    .o(\u_camera_reader/n18 [9]));
  AL_MUX \u_camera_reader/mux8_b0  (
    .i0(1'b0),
    .i1(\u_camera_reader/n8 [0]),
    .sel(\u_camera_reader/mux8_b0_sel_is_0_o ),
    .o(\u_camera_reader/n19 [0]));
  and \u_camera_reader/mux8_b0_sel_is_0  (\u_camera_reader/mux8_b0_sel_is_0_o , \u_camera_reader/n4_neg , \u_camera_reader/mux4_b0_sel_is_0_o_neg );
  AL_MUX \u_camera_reader/mux8_b1  (
    .i0(1'b0),
    .i1(\u_camera_reader/n8 [1]),
    .sel(\u_camera_reader/mux8_b0_sel_is_0_o ),
    .o(\u_camera_reader/n19 [1]));
  AL_MUX \u_camera_reader/mux8_b10  (
    .i0(1'b0),
    .i1(\u_camera_reader/n8 [10]),
    .sel(\u_camera_reader/mux8_b0_sel_is_0_o ),
    .o(\u_camera_reader/n19 [10]));
  AL_MUX \u_camera_reader/mux8_b11  (
    .i0(1'b0),
    .i1(\u_camera_reader/n8 [11]),
    .sel(\u_camera_reader/mux8_b0_sel_is_0_o ),
    .o(\u_camera_reader/n19 [11]));
  AL_MUX \u_camera_reader/mux8_b12  (
    .i0(1'b0),
    .i1(\u_camera_reader/n8 [12]),
    .sel(\u_camera_reader/mux8_b0_sel_is_0_o ),
    .o(\u_camera_reader/n19 [12]));
  AL_MUX \u_camera_reader/mux8_b13  (
    .i0(1'b0),
    .i1(\u_camera_reader/n8 [13]),
    .sel(\u_camera_reader/mux8_b0_sel_is_0_o ),
    .o(\u_camera_reader/n19 [13]));
  AL_MUX \u_camera_reader/mux8_b14  (
    .i0(1'b0),
    .i1(\u_camera_reader/n8 [14]),
    .sel(\u_camera_reader/mux8_b0_sel_is_0_o ),
    .o(\u_camera_reader/n19 [14]));
  AL_MUX \u_camera_reader/mux8_b15  (
    .i0(1'b0),
    .i1(\u_camera_reader/n8 [15]),
    .sel(\u_camera_reader/mux8_b0_sel_is_0_o ),
    .o(\u_camera_reader/n19 [15]));
  AL_MUX \u_camera_reader/mux8_b16  (
    .i0(1'b0),
    .i1(\u_camera_reader/n8 [16]),
    .sel(\u_camera_reader/mux8_b0_sel_is_0_o ),
    .o(\u_camera_reader/n19 [16]));
  AL_MUX \u_camera_reader/mux8_b17  (
    .i0(1'b0),
    .i1(\u_camera_reader/n8 [17]),
    .sel(\u_camera_reader/mux8_b0_sel_is_0_o ),
    .o(\u_camera_reader/n19 [17]));
  AL_MUX \u_camera_reader/mux8_b18  (
    .i0(1'b0),
    .i1(\u_camera_reader/n8 [18]),
    .sel(\u_camera_reader/mux8_b0_sel_is_0_o ),
    .o(\u_camera_reader/n19 [18]));
  AL_MUX \u_camera_reader/mux8_b19  (
    .i0(1'b0),
    .i1(\u_camera_reader/n8 [19]),
    .sel(\u_camera_reader/mux8_b0_sel_is_0_o ),
    .o(\u_camera_reader/n19 [19]));
  AL_MUX \u_camera_reader/mux8_b2  (
    .i0(1'b0),
    .i1(\u_camera_reader/n8 [2]),
    .sel(\u_camera_reader/mux8_b0_sel_is_0_o ),
    .o(\u_camera_reader/n19 [2]));
  AL_MUX \u_camera_reader/mux8_b3  (
    .i0(1'b0),
    .i1(\u_camera_reader/n8 [3]),
    .sel(\u_camera_reader/mux8_b0_sel_is_0_o ),
    .o(\u_camera_reader/n19 [3]));
  AL_MUX \u_camera_reader/mux8_b4  (
    .i0(1'b0),
    .i1(\u_camera_reader/n8 [4]),
    .sel(\u_camera_reader/mux8_b0_sel_is_0_o ),
    .o(\u_camera_reader/n19 [4]));
  AL_MUX \u_camera_reader/mux8_b5  (
    .i0(1'b0),
    .i1(\u_camera_reader/n8 [5]),
    .sel(\u_camera_reader/mux8_b0_sel_is_0_o ),
    .o(\u_camera_reader/n19 [5]));
  AL_MUX \u_camera_reader/mux8_b6  (
    .i0(1'b0),
    .i1(\u_camera_reader/n8 [6]),
    .sel(\u_camera_reader/mux8_b0_sel_is_0_o ),
    .o(\u_camera_reader/n19 [6]));
  AL_MUX \u_camera_reader/mux8_b7  (
    .i0(1'b0),
    .i1(\u_camera_reader/n8 [7]),
    .sel(\u_camera_reader/mux8_b0_sel_is_0_o ),
    .o(\u_camera_reader/n19 [7]));
  AL_MUX \u_camera_reader/mux8_b8  (
    .i0(1'b0),
    .i1(\u_camera_reader/n8 [8]),
    .sel(\u_camera_reader/mux8_b0_sel_is_0_o ),
    .o(\u_camera_reader/n19 [8]));
  AL_MUX \u_camera_reader/mux8_b9  (
    .i0(1'b0),
    .i1(\u_camera_reader/n8 [9]),
    .sel(\u_camera_reader/mux8_b0_sel_is_0_o ),
    .o(\u_camera_reader/n19 [9]));
  binary_mux_s1_w1 \u_camera_reader/mux9_b0  (
    .i0(\u_camera_reader/n18 [0]),
    .i1(1'b0),
    .sel(\u_camera_reader/n4 ),
    .o(\u_camera_reader/n21 [0]));  // sources/rtl/camera_reader.v(94)
  binary_mux_s1_w1 \u_camera_reader/mux9_b1  (
    .i0(\u_camera_reader/n18 [1]),
    .i1(1'b0),
    .sel(\u_camera_reader/n4 ),
    .o(\u_camera_reader/n21 [1]));  // sources/rtl/camera_reader.v(94)
  binary_mux_s1_w1 \u_camera_reader/mux9_b10  (
    .i0(\u_camera_reader/n18 [10]),
    .i1(1'b0),
    .sel(\u_camera_reader/n4 ),
    .o(\u_camera_reader/n21 [10]));  // sources/rtl/camera_reader.v(94)
  binary_mux_s1_w1 \u_camera_reader/mux9_b11  (
    .i0(\u_camera_reader/n18 [11]),
    .i1(1'b0),
    .sel(\u_camera_reader/n4 ),
    .o(\u_camera_reader/n21 [11]));  // sources/rtl/camera_reader.v(94)
  binary_mux_s1_w1 \u_camera_reader/mux9_b12  (
    .i0(\u_camera_reader/n18 [12]),
    .i1(1'b0),
    .sel(\u_camera_reader/n4 ),
    .o(\u_camera_reader/n21 [12]));  // sources/rtl/camera_reader.v(94)
  binary_mux_s1_w1 \u_camera_reader/mux9_b13  (
    .i0(\u_camera_reader/n18 [13]),
    .i1(1'b0),
    .sel(\u_camera_reader/n4 ),
    .o(\u_camera_reader/n21 [13]));  // sources/rtl/camera_reader.v(94)
  binary_mux_s1_w1 \u_camera_reader/mux9_b14  (
    .i0(\u_camera_reader/n18 [14]),
    .i1(1'b0),
    .sel(\u_camera_reader/n4 ),
    .o(\u_camera_reader/n21 [14]));  // sources/rtl/camera_reader.v(94)
  binary_mux_s1_w1 \u_camera_reader/mux9_b15  (
    .i0(\u_camera_reader/n18 [15]),
    .i1(1'b0),
    .sel(\u_camera_reader/n4 ),
    .o(\u_camera_reader/n21 [15]));  // sources/rtl/camera_reader.v(94)
  binary_mux_s1_w1 \u_camera_reader/mux9_b2  (
    .i0(\u_camera_reader/n18 [2]),
    .i1(1'b0),
    .sel(\u_camera_reader/n4 ),
    .o(\u_camera_reader/n21 [2]));  // sources/rtl/camera_reader.v(94)
  binary_mux_s1_w1 \u_camera_reader/mux9_b3  (
    .i0(\u_camera_reader/n18 [3]),
    .i1(1'b0),
    .sel(\u_camera_reader/n4 ),
    .o(\u_camera_reader/n21 [3]));  // sources/rtl/camera_reader.v(94)
  binary_mux_s1_w1 \u_camera_reader/mux9_b4  (
    .i0(\u_camera_reader/n18 [4]),
    .i1(1'b0),
    .sel(\u_camera_reader/n4 ),
    .o(\u_camera_reader/n21 [4]));  // sources/rtl/camera_reader.v(94)
  binary_mux_s1_w1 \u_camera_reader/mux9_b5  (
    .i0(\u_camera_reader/n18 [5]),
    .i1(1'b0),
    .sel(\u_camera_reader/n4 ),
    .o(\u_camera_reader/n21 [5]));  // sources/rtl/camera_reader.v(94)
  binary_mux_s1_w1 \u_camera_reader/mux9_b6  (
    .i0(\u_camera_reader/n18 [6]),
    .i1(1'b0),
    .sel(\u_camera_reader/n4 ),
    .o(\u_camera_reader/n21 [6]));  // sources/rtl/camera_reader.v(94)
  binary_mux_s1_w1 \u_camera_reader/mux9_b7  (
    .i0(\u_camera_reader/n18 [7]),
    .i1(1'b0),
    .sel(\u_camera_reader/n4 ),
    .o(\u_camera_reader/n21 [7]));  // sources/rtl/camera_reader.v(94)
  binary_mux_s1_w1 \u_camera_reader/mux9_b8  (
    .i0(\u_camera_reader/n18 [8]),
    .i1(1'b0),
    .sel(\u_camera_reader/n4 ),
    .o(\u_camera_reader/n21 [8]));  // sources/rtl/camera_reader.v(94)
  binary_mux_s1_w1 \u_camera_reader/mux9_b9  (
    .i0(\u_camera_reader/n18 [9]),
    .i1(1'b0),
    .sel(\u_camera_reader/n4 ),
    .o(\u_camera_reader/n21 [9]));  // sources/rtl/camera_reader.v(94)
  not \u_camera_reader/n13_inv  (\u_camera_reader/n13_neg , \u_camera_reader/n13 );
  not \u_camera_reader/n3_inv  (\u_camera_reader/n3_neg , \u_camera_reader/n3 );
  not \u_camera_reader/n4_inv  (\u_camera_reader/n4_neg , \u_camera_reader/n4 );
  not \u_camera_reader/n6_inv  (\u_camera_reader/n6_neg , \u_camera_reader/n6 );
  not \u_camera_reader/n7_inv  (\u_camera_reader/n7_neg , \u_camera_reader/n7 );
  reg_ar_as_w1 \u_camera_reader/reg0_b0  (
    .clk(camera_wrreq),
    .d(\u_camera_reader/current_pixel [0]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(camera_wrdat[0]));  // sources/rtl/camera_reader.v(56)
  reg_ar_as_w1 \u_camera_reader/reg0_b1  (
    .clk(camera_wrreq),
    .d(\u_camera_reader/current_pixel [1]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(camera_wrdat[1]));  // sources/rtl/camera_reader.v(56)
  reg_ar_as_w1 \u_camera_reader/reg0_b10  (
    .clk(camera_wrreq),
    .d(\u_camera_reader/current_pixel [10]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(camera_wrdat[10]));  // sources/rtl/camera_reader.v(56)
  reg_ar_as_w1 \u_camera_reader/reg0_b11  (
    .clk(camera_wrreq),
    .d(\u_camera_reader/current_pixel [11]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(camera_wrdat[11]));  // sources/rtl/camera_reader.v(56)
  reg_ar_as_w1 \u_camera_reader/reg0_b12  (
    .clk(camera_wrreq),
    .d(\u_camera_reader/current_pixel [12]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(camera_wrdat[12]));  // sources/rtl/camera_reader.v(56)
  reg_ar_as_w1 \u_camera_reader/reg0_b13  (
    .clk(camera_wrreq),
    .d(\u_camera_reader/current_pixel [13]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(camera_wrdat[13]));  // sources/rtl/camera_reader.v(56)
  reg_ar_as_w1 \u_camera_reader/reg0_b14  (
    .clk(camera_wrreq),
    .d(\u_camera_reader/current_pixel [14]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(camera_wrdat[14]));  // sources/rtl/camera_reader.v(56)
  reg_ar_as_w1 \u_camera_reader/reg0_b15  (
    .clk(camera_wrreq),
    .d(\u_camera_reader/current_pixel [15]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(camera_wrdat[15]));  // sources/rtl/camera_reader.v(56)
  reg_ar_as_w1 \u_camera_reader/reg0_b2  (
    .clk(camera_wrreq),
    .d(\u_camera_reader/current_pixel [2]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(camera_wrdat[2]));  // sources/rtl/camera_reader.v(56)
  reg_ar_as_w1 \u_camera_reader/reg0_b3  (
    .clk(camera_wrreq),
    .d(\u_camera_reader/current_pixel [3]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(camera_wrdat[3]));  // sources/rtl/camera_reader.v(56)
  reg_ar_as_w1 \u_camera_reader/reg0_b4  (
    .clk(camera_wrreq),
    .d(\u_camera_reader/current_pixel [4]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(camera_wrdat[4]));  // sources/rtl/camera_reader.v(56)
  reg_ar_as_w1 \u_camera_reader/reg0_b5  (
    .clk(camera_wrreq),
    .d(\u_camera_reader/current_pixel [5]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(camera_wrdat[5]));  // sources/rtl/camera_reader.v(56)
  reg_ar_as_w1 \u_camera_reader/reg0_b6  (
    .clk(camera_wrreq),
    .d(\u_camera_reader/current_pixel [6]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(camera_wrdat[6]));  // sources/rtl/camera_reader.v(56)
  reg_ar_as_w1 \u_camera_reader/reg0_b7  (
    .clk(camera_wrreq),
    .d(\u_camera_reader/current_pixel [7]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(camera_wrdat[7]));  // sources/rtl/camera_reader.v(56)
  reg_ar_as_w1 \u_camera_reader/reg0_b8  (
    .clk(camera_wrreq),
    .d(\u_camera_reader/current_pixel [8]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(camera_wrdat[8]));  // sources/rtl/camera_reader.v(56)
  reg_ar_as_w1 \u_camera_reader/reg0_b9  (
    .clk(camera_wrreq),
    .d(\u_camera_reader/current_pixel [9]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(camera_wrdat[9]));  // sources/rtl/camera_reader.v(56)
  reg_ar_as_w1 \u_camera_reader/reg1_b0  (
    .clk(cam_pclk),
    .d(\u_camera_reader/n19 [0]),
    .en(1'b1),
    .reset(\u_camera_reader/n3 ),
    .set(1'b0),
    .q(\u_camera_reader/pixel_counter [0]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg1_b1  (
    .clk(cam_pclk),
    .d(\u_camera_reader/n19 [1]),
    .en(1'b1),
    .reset(\u_camera_reader/n3 ),
    .set(1'b0),
    .q(\u_camera_reader/pixel_counter [1]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg1_b10  (
    .clk(cam_pclk),
    .d(\u_camera_reader/n19 [10]),
    .en(1'b1),
    .reset(\u_camera_reader/n3 ),
    .set(1'b0),
    .q(\u_camera_reader/pixel_counter [10]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg1_b11  (
    .clk(cam_pclk),
    .d(\u_camera_reader/n19 [11]),
    .en(1'b1),
    .reset(\u_camera_reader/n3 ),
    .set(1'b0),
    .q(\u_camera_reader/pixel_counter [11]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg1_b12  (
    .clk(cam_pclk),
    .d(\u_camera_reader/n19 [12]),
    .en(1'b1),
    .reset(\u_camera_reader/n3 ),
    .set(1'b0),
    .q(\u_camera_reader/pixel_counter [12]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg1_b13  (
    .clk(cam_pclk),
    .d(\u_camera_reader/n19 [13]),
    .en(1'b1),
    .reset(\u_camera_reader/n3 ),
    .set(1'b0),
    .q(\u_camera_reader/pixel_counter [13]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg1_b14  (
    .clk(cam_pclk),
    .d(\u_camera_reader/n19 [14]),
    .en(1'b1),
    .reset(\u_camera_reader/n3 ),
    .set(1'b0),
    .q(\u_camera_reader/pixel_counter [14]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg1_b15  (
    .clk(cam_pclk),
    .d(\u_camera_reader/n19 [15]),
    .en(1'b1),
    .reset(\u_camera_reader/n3 ),
    .set(1'b0),
    .q(\u_camera_reader/pixel_counter [15]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg1_b16  (
    .clk(cam_pclk),
    .d(\u_camera_reader/n19 [16]),
    .en(1'b1),
    .reset(\u_camera_reader/n3 ),
    .set(1'b0),
    .q(\u_camera_reader/pixel_counter [16]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg1_b17  (
    .clk(cam_pclk),
    .d(\u_camera_reader/n19 [17]),
    .en(1'b1),
    .reset(\u_camera_reader/n3 ),
    .set(1'b0),
    .q(\u_camera_reader/pixel_counter [17]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg1_b18  (
    .clk(cam_pclk),
    .d(\u_camera_reader/n19 [18]),
    .en(1'b1),
    .reset(\u_camera_reader/n3 ),
    .set(1'b0),
    .q(\u_camera_reader/pixel_counter [18]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg1_b19  (
    .clk(cam_pclk),
    .d(\u_camera_reader/n19 [19]),
    .en(1'b1),
    .reset(\u_camera_reader/n3 ),
    .set(1'b0),
    .q(\u_camera_reader/pixel_counter [19]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg1_b2  (
    .clk(cam_pclk),
    .d(\u_camera_reader/n19 [2]),
    .en(1'b1),
    .reset(\u_camera_reader/n3 ),
    .set(1'b0),
    .q(\u_camera_reader/pixel_counter [2]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg1_b3  (
    .clk(cam_pclk),
    .d(\u_camera_reader/n19 [3]),
    .en(1'b1),
    .reset(\u_camera_reader/n3 ),
    .set(1'b0),
    .q(\u_camera_reader/pixel_counter [3]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg1_b4  (
    .clk(cam_pclk),
    .d(\u_camera_reader/n19 [4]),
    .en(1'b1),
    .reset(\u_camera_reader/n3 ),
    .set(1'b0),
    .q(\u_camera_reader/pixel_counter [4]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg1_b5  (
    .clk(cam_pclk),
    .d(\u_camera_reader/n19 [5]),
    .en(1'b1),
    .reset(\u_camera_reader/n3 ),
    .set(1'b0),
    .q(\u_camera_reader/pixel_counter [5]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg1_b6  (
    .clk(cam_pclk),
    .d(\u_camera_reader/n19 [6]),
    .en(1'b1),
    .reset(\u_camera_reader/n3 ),
    .set(1'b0),
    .q(\u_camera_reader/pixel_counter [6]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg1_b7  (
    .clk(cam_pclk),
    .d(\u_camera_reader/n19 [7]),
    .en(1'b1),
    .reset(\u_camera_reader/n3 ),
    .set(1'b0),
    .q(\u_camera_reader/pixel_counter [7]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg1_b8  (
    .clk(cam_pclk),
    .d(\u_camera_reader/n19 [8]),
    .en(1'b1),
    .reset(\u_camera_reader/n3 ),
    .set(1'b0),
    .q(\u_camera_reader/pixel_counter [8]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg1_b9  (
    .clk(cam_pclk),
    .d(\u_camera_reader/n19 [9]),
    .en(1'b1),
    .reset(\u_camera_reader/n3 ),
    .set(1'b0),
    .q(\u_camera_reader/pixel_counter [9]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg2_b0  (
    .clk(cam_pclk),
    .d(\u_camera_reader/n21 [0]),
    .en(~\u_camera_reader/n3 ),
    .reset(1'b0),
    .set(1'b0),
    .q(camera_addr[0]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg2_b1  (
    .clk(cam_pclk),
    .d(\u_camera_reader/n21 [1]),
    .en(~\u_camera_reader/n3 ),
    .reset(1'b0),
    .set(1'b0),
    .q(camera_addr[1]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg2_b10  (
    .clk(cam_pclk),
    .d(\u_camera_reader/n21 [10]),
    .en(~\u_camera_reader/n3 ),
    .reset(1'b0),
    .set(1'b0),
    .q(camera_addr[10]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg2_b11  (
    .clk(cam_pclk),
    .d(\u_camera_reader/n21 [11]),
    .en(~\u_camera_reader/n3 ),
    .reset(1'b0),
    .set(1'b0),
    .q(camera_addr[11]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg2_b12  (
    .clk(cam_pclk),
    .d(\u_camera_reader/n21 [12]),
    .en(~\u_camera_reader/n3 ),
    .reset(1'b0),
    .set(1'b0),
    .q(camera_addr[12]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg2_b13  (
    .clk(cam_pclk),
    .d(\u_camera_reader/n21 [13]),
    .en(~\u_camera_reader/n3 ),
    .reset(1'b0),
    .set(1'b0),
    .q(camera_addr[13]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg2_b14  (
    .clk(cam_pclk),
    .d(\u_camera_reader/n21 [14]),
    .en(~\u_camera_reader/n3 ),
    .reset(1'b0),
    .set(1'b0),
    .q(camera_addr[14]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg2_b15  (
    .clk(cam_pclk),
    .d(\u_camera_reader/n21 [15]),
    .en(~\u_camera_reader/n3 ),
    .reset(1'b0),
    .set(1'b0),
    .q(camera_addr[15]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg2_b2  (
    .clk(cam_pclk),
    .d(\u_camera_reader/n21 [2]),
    .en(~\u_camera_reader/n3 ),
    .reset(1'b0),
    .set(1'b0),
    .q(camera_addr[2]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg2_b3  (
    .clk(cam_pclk),
    .d(\u_camera_reader/n21 [3]),
    .en(~\u_camera_reader/n3 ),
    .reset(1'b0),
    .set(1'b0),
    .q(camera_addr[3]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg2_b4  (
    .clk(cam_pclk),
    .d(\u_camera_reader/n21 [4]),
    .en(~\u_camera_reader/n3 ),
    .reset(1'b0),
    .set(1'b0),
    .q(camera_addr[4]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg2_b5  (
    .clk(cam_pclk),
    .d(\u_camera_reader/n21 [5]),
    .en(~\u_camera_reader/n3 ),
    .reset(1'b0),
    .set(1'b0),
    .q(camera_addr[5]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg2_b6  (
    .clk(cam_pclk),
    .d(\u_camera_reader/n21 [6]),
    .en(~\u_camera_reader/n3 ),
    .reset(1'b0),
    .set(1'b0),
    .q(camera_addr[6]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg2_b7  (
    .clk(cam_pclk),
    .d(\u_camera_reader/n21 [7]),
    .en(~\u_camera_reader/n3 ),
    .reset(1'b0),
    .set(1'b0),
    .q(camera_addr[7]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg2_b8  (
    .clk(cam_pclk),
    .d(\u_camera_reader/n21 [8]),
    .en(~\u_camera_reader/n3 ),
    .reset(1'b0),
    .set(1'b0),
    .q(camera_addr[8]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg2_b9  (
    .clk(cam_pclk),
    .d(\u_camera_reader/n21 [9]),
    .en(~\u_camera_reader/n3 ),
    .reset(1'b0),
    .set(1'b0),
    .q(camera_addr[9]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg3_b0  (
    .clk(cam_pclk),
    .d(cam_data[0]),
    .en(\u_camera_reader/mux13_b0_sel_is_2_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_camera_reader/subpixel [0]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg3_b1  (
    .clk(cam_pclk),
    .d(cam_data[1]),
    .en(\u_camera_reader/mux13_b0_sel_is_2_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_camera_reader/subpixel [1]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg3_b2  (
    .clk(cam_pclk),
    .d(cam_data[2]),
    .en(\u_camera_reader/mux13_b0_sel_is_2_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_camera_reader/subpixel [2]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg3_b3  (
    .clk(cam_pclk),
    .d(cam_data[3]),
    .en(\u_camera_reader/mux13_b0_sel_is_2_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_camera_reader/subpixel [3]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg3_b4  (
    .clk(cam_pclk),
    .d(cam_data[4]),
    .en(\u_camera_reader/mux13_b0_sel_is_2_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_camera_reader/subpixel [4]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg3_b5  (
    .clk(cam_pclk),
    .d(cam_data[5]),
    .en(\u_camera_reader/mux13_b0_sel_is_2_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_camera_reader/subpixel [5]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg3_b6  (
    .clk(cam_pclk),
    .d(cam_data[6]),
    .en(\u_camera_reader/mux13_b0_sel_is_2_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_camera_reader/subpixel [6]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg3_b7  (
    .clk(cam_pclk),
    .d(cam_data[7]),
    .en(\u_camera_reader/mux13_b0_sel_is_2_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_camera_reader/subpixel [7]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg4_b0  (
    .clk(cam_pclk),
    .d(cam_data[0]),
    .en(\u_camera_reader/mux14_b0_sel_is_2_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_camera_reader/current_pixel [0]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg4_b1  (
    .clk(cam_pclk),
    .d(cam_data[1]),
    .en(\u_camera_reader/mux14_b0_sel_is_2_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_camera_reader/current_pixel [1]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg4_b10  (
    .clk(cam_pclk),
    .d(\u_camera_reader/subpixel [2]),
    .en(\u_camera_reader/mux14_b0_sel_is_2_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_camera_reader/current_pixel [10]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg4_b11  (
    .clk(cam_pclk),
    .d(\u_camera_reader/subpixel [3]),
    .en(\u_camera_reader/mux14_b0_sel_is_2_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_camera_reader/current_pixel [11]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg4_b12  (
    .clk(cam_pclk),
    .d(\u_camera_reader/subpixel [4]),
    .en(\u_camera_reader/mux14_b0_sel_is_2_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_camera_reader/current_pixel [12]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg4_b13  (
    .clk(cam_pclk),
    .d(\u_camera_reader/subpixel [5]),
    .en(\u_camera_reader/mux14_b0_sel_is_2_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_camera_reader/current_pixel [13]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg4_b14  (
    .clk(cam_pclk),
    .d(\u_camera_reader/subpixel [6]),
    .en(\u_camera_reader/mux14_b0_sel_is_2_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_camera_reader/current_pixel [14]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg4_b15  (
    .clk(cam_pclk),
    .d(\u_camera_reader/subpixel [7]),
    .en(\u_camera_reader/mux14_b0_sel_is_2_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_camera_reader/current_pixel [15]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg4_b2  (
    .clk(cam_pclk),
    .d(cam_data[2]),
    .en(\u_camera_reader/mux14_b0_sel_is_2_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_camera_reader/current_pixel [2]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg4_b3  (
    .clk(cam_pclk),
    .d(cam_data[3]),
    .en(\u_camera_reader/mux14_b0_sel_is_2_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_camera_reader/current_pixel [3]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg4_b4  (
    .clk(cam_pclk),
    .d(cam_data[4]),
    .en(\u_camera_reader/mux14_b0_sel_is_2_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_camera_reader/current_pixel [4]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg4_b5  (
    .clk(cam_pclk),
    .d(cam_data[5]),
    .en(\u_camera_reader/mux14_b0_sel_is_2_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_camera_reader/current_pixel [5]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg4_b6  (
    .clk(cam_pclk),
    .d(cam_data[6]),
    .en(\u_camera_reader/mux14_b0_sel_is_2_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_camera_reader/current_pixel [6]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg4_b7  (
    .clk(cam_pclk),
    .d(cam_data[7]),
    .en(\u_camera_reader/mux14_b0_sel_is_2_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_camera_reader/current_pixel [7]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg4_b8  (
    .clk(cam_pclk),
    .d(\u_camera_reader/subpixel [0]),
    .en(\u_camera_reader/mux14_b0_sel_is_2_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_camera_reader/current_pixel [8]));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/reg4_b9  (
    .clk(cam_pclk),
    .d(\u_camera_reader/subpixel [1]),
    .en(\u_camera_reader/mux14_b0_sel_is_2_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_camera_reader/current_pixel [9]));  // sources/rtl/camera_reader.v(95)
  AL_MUX \u_camera_reader/u2  (
    .i0(1'b0),
    .i1(clk_cam),
    .sel(\u_camera_reader/n0 ),
    .o(cam_xclk));  // sources/rtl/camera_reader.v(33)
  not \u_camera_reader/u3  (\u_camera_reader/n1 , \u_camera_reader/wrclk1 );  // sources/rtl/camera_reader.v(42)
  and \u_camera_reader/u4  (\u_camera_reader/n6 , \u_camera_reader/n2 , \u_camera_reader/n5 );  // sources/rtl/camera_reader.v(74)
  and \u_camera_reader/u6  (\u_camera_reader/n28 , \u_camera_reader/n13 , \u_camera_reader/n27 );  // sources/rtl/camera_reader.v(98)
  AL_MUX \u_camera_reader/u7  (
    .i0(1'b0),
    .i1(\u_camera_reader/wrclk1 ),
    .sel(\u_camera_reader/n28 ),
    .o(camera_wrreq));  // sources/rtl/camera_reader.v(98)
  reg_ar_ss_w1 \u_camera_reader/vsync_passed_reg  (
    .clk(cam_pclk),
    .d(\u_camera_reader/vsync_passed ),
    .en(1'b1),
    .reset(\u_camera_reader/n3 ),
    .set(\u_camera_reader/n4 ),
    .q(\u_camera_reader/vsync_passed ));  // sources/rtl/camera_reader.v(95)
  reg_ar_as_w1 \u_camera_reader/wrclk1_reg  (
    .clk(cam_pclk),
    .d(\u_camera_reader/n1 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_camera_reader/wrclk1 ));  // sources/rtl/camera_reader.v(43)
  reg_ar_as_w1 \u_camera_reader/write_pixel_reg  (
    .clk(~\u_camera_reader/wrclk1 ),
    .d(\u_camera_reader/n2 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\u_camera_reader/write_pixel ));  // sources/rtl/camera_reader.v(51)
  EG_LOGIC_BRAM #(
    //.FORCE_KEEP("OFF"),
    //.INIT_FILE("NONE"),
    .ADDR_WIDTH_A(16),
    .ADDR_WIDTH_B(16),
    .BYTE_A(1),
    .BYTE_B(1),
    .BYTE_ENABLE(0),
    .DATA_DEPTH_A(32800),
    .DATA_DEPTH_B(32800),
    .DATA_WIDTH_A(16),
    .DATA_WIDTH_B(16),
    .DEBUGGABLE("NO"),
    .FILL_ALL("NONE"),
    .IMPLEMENT("9K"),
    .MODE("PDPW"),
    .PACKABLE("NO"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("OUTREG"),
    .RESETMODE("SYNC"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_img/inst  (
    .addra(camera_addr[15:0]),
    .addrb(vga_rdaddr),
    .bea(1'b0),
    .beb(1'b0),
    .cea(camera_wrreq),
    .ceb(vga_rden),
    .clka(cam_pclk),
    .clkb(clk_lcd),
    .dia(camera_wrdat),
    .dib(16'b0000000000000000),
    .ocea(1'b0),
    .oceb(1'b1),
    .rsta(n1),
    .rstb(n1),
    .wea(1'b1),
    .web(1'b0),
    .dob(vga_rddat));  // al_ip/ip_ram.v(46)
  EG_LOGIC_BUFG \u_pll/bufg_feedback  (
    .i(\u_pll/clk0_buf ),
    .o(clk_lcd));  // al_ip/ip_pll.v(36)
  EG_PHY_PLL #(
    .CLKC0_CPHASE(19),
    .CLKC0_DIV(20),
    .CLKC0_DIV2_ENABLE("DISABLE"),
    .CLKC0_ENABLE("ENABLE"),
    .CLKC0_FPHASE(0),
    .CLKC1_CPHASE(41),
    .CLKC1_DIV(42),
    .CLKC1_DIV2_ENABLE("DISABLE"),
    .CLKC1_ENABLE("ENABLE"),
    .CLKC1_FPHASE(0),
    .CLKC2_CPHASE(125),
    .CLKC2_DIV(126),
    .CLKC2_DIV2_ENABLE("DISABLE"),
    .CLKC2_ENABLE("ENABLE"),
    .CLKC2_FPHASE(0),
    .CLKC3_CPHASE(1),
    .CLKC3_DIV(1),
    .CLKC3_DIV2_ENABLE("DISABLE"),
    .CLKC3_ENABLE("DISABLE"),
    .CLKC3_FPHASE(0),
    .CLKC4_CPHASE(1),
    .CLKC4_DIV(1),
    .CLKC4_DIV2_ENABLE("DISABLE"),
    .CLKC4_ENABLE("DISABLE"),
    .CLKC4_FPHASE(0),
    .DERIVE_PLL_CLOCKS("DISABLE"),
    .DPHASE_SOURCE("DISABLE"),
    .DYNCFG("DISABLE"),
    .FBCLK_DIV(17),
    .FEEDBK_MODE("NORMAL"),
    .FEEDBK_PATH("CLKC0_EXT"),
    .FIN("24.000"),
    .FREQ_LOCK_ACCURACY(2),
    .GEN_BASIC_CLOCK("DISABLE"),
    .GMC_GAIN(6),
    .GMC_TEST(14),
    .ICP_CURRENT(3),
    .IF_ESCLKSTSW("DISABLE"),
    .INTFB_WAKE("DISABLE"),
    .KVCO(6),
    .LPF_CAPACITOR(3),
    .LPF_RESISTOR(2),
    .NORESET("DISABLE"),
    .ODIV_MUXC0("DIV"),
    .ODIV_MUXC1("DIV"),
    .ODIV_MUXC2("DIV"),
    .ODIV_MUXC3("DIV"),
    .ODIV_MUXC4("DIV"),
    .PLLC2RST_ENA("DISABLE"),
    .PLLC34RST_ENA("DISABLE"),
    .PLLMRST_ENA("DISABLE"),
    .PLLRST_ENA("DISABLE"),
    .PLL_LOCK_MODE(0),
    .PREDIV_MUXC0("VCO"),
    .PREDIV_MUXC1("VCO"),
    .PREDIV_MUXC2("VCO"),
    .PREDIV_MUXC3("VCO"),
    .PREDIV_MUXC4("VCO"),
    .REFCLK_DIV(16),
    .REFCLK_SEL("INTERNAL"),
    .STDBY_ENABLE("DISABLE"),
    .STDBY_VCO_ENA("DISABLE"),
    .SYNC_ENABLE("DISABLE"),
    .VCO_NORESET("DISABLE"))
    \u_pll/pll_inst  (
    .daddr(6'b000000),
    .dclk(1'b0),
    .dcs(1'b0),
    .di(8'b00000000),
    .dwe(1'b0),
    .fbclk(clk_lcd),
    .psclk(1'b0),
    .psclksel(3'b000),
    .psdown(1'b0),
    .psstep(1'b0),
    .refclk(clk_24m),
    .reset(1'b0),
    .stdby(1'b0),
    .clkc({open_n17,open_n18,clk_sccb,clk_cam,\u_pll/clk0_buf }));  // al_ip/ip_pll.v(67)
  \lcd_sync(IMG_Y=1)  u_vga_sync (
    .clk(clk_lcd),
    .rest_n(cam_rst),
    .addr(vga_rdaddr),
    .img_ack(vga_rden),
    .lcd_clk(vga_clk),
    .lcd_hsync(vga_hsync),
    .lcd_vsync(vga_vsync));  // sources/rtl/test_camera.v(102)

endmodule 

module binary_mux_s1_w1
  (
  i0,
  i1,
  sel,
  o
  );

  input i0;
  input i1;
  input sel;
  output o;


  AL_MUX al_mux_b0_0_0 (
    .i0(i0),
    .i1(i1),
    .sel(sel),
    .o(o));

endmodule 

module camera_init  // sources/rtl/camera_init.v(14)
  (
  clk,
  reset_n,
  sda_in,
  ready,
  scl,
  sda,
  sda_oe
  );

  input clk;  // sources/rtl/camera_init.v(15)
  input reset_n;  // sources/rtl/camera_init.v(16)
  input sda_in;  // sources/rtl/camera_init.v(20)
  output ready;  // sources/rtl/camera_init.v(17)
  output scl;  // sources/rtl/camera_init.v(21)
  output sda;  // sources/rtl/camera_init.v(19)
  output sda_oe;  // sources/rtl/camera_init.v(18)

  parameter REGS_TO_INIT = 178;
  // localparam CAMERA_IDLE = 18;
  // localparam CAMERA_INIT_1 = 11;
  // localparam CAMERA_INIT_2 = 12;
  // localparam CAMERA_INIT_3 = 13;
  // localparam CAMERA_INIT_4 = 14;
  // localparam CAMERA_INIT_5 = 15;
  // localparam CAMERA_INIT_6 = 16;
  // localparam CAMERA_INIT_7 = 17;
  // localparam CONTROL_REG = 3'b000;
  // localparam SLAVE_ADDRESS = 3'b001;
  // localparam SLAVE_DATA_1 = 3'b011;
  // localparam SLAVE_DATA_2 = 3'b100;
  // localparam SLAVE_REG_ADDRESS = 3'b010;
  wire [7:0] cnt;  // sources/rtl/camera_init.v(64)
  wire [7:0] counter;  // sources/rtl/camera_init.v(63)
  wire [7:0] data_in_bus;  // sources/rtl/camera_init.v(42)
  wire [8:0] divider2;  // sources/rtl/camera_init.v(67)
  wire [8:0] n0;
  wire [10:0] n178;
  wire [15:0] n181;
  wire [15:0] n182;
  wire [15:0] n183;
  wire [15:0] n184;
  wire [15:0] n185;
  wire [15:0] n186;
  wire [15:0] n187;
  wire [15:0] n188;
  wire [15:0] n189;
  wire [15:0] n190;
  wire [15:0] n191;
  wire [15:0] n192;
  wire [15:0] n193;
  wire [15:0] n194;
  wire [15:0] n195;
  wire [15:0] n196;
  wire [15:0] n197;
  wire [15:0] n198;
  wire [15:0] n199;
  wire [15:0] n200;
  wire [15:0] n201;
  wire [15:0] n202;
  wire [15:0] n203;
  wire [15:0] n204;
  wire [15:0] n205;
  wire [15:0] n206;
  wire [15:0] n207;
  wire [15:0] n208;
  wire [15:0] n209;
  wire [15:0] n210;
  wire [15:0] n211;
  wire [15:0] n212;
  wire [15:0] n213;
  wire [15:0] n214;
  wire [15:0] n215;
  wire [15:0] n216;
  wire [15:0] n217;
  wire [15:0] n218;
  wire [15:0] n219;
  wire [15:0] n221;
  wire [15:0] n222;
  wire [15:0] n223;
  wire [15:0] n224;
  wire [15:0] n225;
  wire [15:0] n226;
  wire [15:0] n227;
  wire [15:0] n228;
  wire [15:0] n229;
  wire [15:0] n230;
  wire [15:0] n231;
  wire [15:0] n232;
  wire [15:0] n233;
  wire [15:0] n240;
  wire [15:0] n241;
  wire [15:0] n242;
  wire [15:0] n244;
  wire [15:0] n245;
  wire [15:0] n246;
  wire [15:0] n247;
  wire [15:0] n248;
  wire [15:0] n249;
  wire [15:0] n250;
  wire [15:0] n251;
  wire [15:0] n252;
  wire [15:0] n253;
  wire [15:0] n254;
  wire [15:0] n255;
  wire [15:0] n256;
  wire [15:0] n257;
  wire [15:0] n258;
  wire [15:0] n259;
  wire [15:0] n260;
  wire [15:0] n261;
  wire [15:0] n262;
  wire [15:0] n263;
  wire [15:0] n264;
  wire [15:0] n265;
  wire [15:0] n266;
  wire [15:0] n267;
  wire [15:0] n268;
  wire [15:0] n270;
  wire [15:0] n271;
  wire [15:0] n272;
  wire [15:0] n273;
  wire [15:0] n274;
  wire [15:0] n275;
  wire [15:0] n276;
  wire [15:0] n277;
  wire [15:0] n278;
  wire [15:0] n279;
  wire [15:0] n280;
  wire [15:0] n281;
  wire [15:0] n282;
  wire [15:0] n283;
  wire [15:0] n284;
  wire [15:0] n285;
  wire [15:0] n286;
  wire [15:0] n287;
  wire [15:0] n288;
  wire [15:0] n289;
  wire [15:0] n290;
  wire [15:0] n291;
  wire [15:0] n292;
  wire [15:0] n293;
  wire [15:0] n294;
  wire [15:0] n295;
  wire [15:0] n296;
  wire [15:0] n297;
  wire [15:0] n298;
  wire [15:0] n299;
  wire [15:0] n300;
  wire [15:0] n301;
  wire [15:0] n302;
  wire [15:0] n303;
  wire [15:0] n304;
  wire [15:0] n305;
  wire [15:0] n306;
  wire [15:0] n307;
  wire [15:0] n308;
  wire [15:0] n309;
  wire [15:0] n310;
  wire [15:0] n311;
  wire [15:0] n312;
  wire [15:0] n313;
  wire [15:0] n314;
  wire [15:0] n315;
  wire [15:0] n316;
  wire [15:0] n317;
  wire [15:0] n318;
  wire [15:0] n319;
  wire [15:0] n320;
  wire [15:0] n321;
  wire [15:0] n322;
  wire [15:0] n323;
  wire [15:0] n324;
  wire [15:0] n325;
  wire [15:0] n326;
  wire [15:0] n327;
  wire [15:0] n328;
  wire [15:0] n329;
  wire [15:0] n330;
  wire [15:0] n331;
  wire [15:0] n332;
  wire [15:0] n333;
  wire [15:0] n334;
  wire [15:0] n335;
  wire [15:0] n336;
  wire [15:0] n337;
  wire [15:0] n338;
  wire [15:0] n339;
  wire [15:0] n340;
  wire [15:0] n341;
  wire [15:0] n342;
  wire [15:0] n343;
  wire [15:0] n344;
  wire [15:0] n345;
  wire [15:0] n346;
  wire [15:0] n347;
  wire [15:0] n348;
  wire [15:0] n349;
  wire [15:0] n350;
  wire [15:0] n351;
  wire [15:0] n352;
  wire [15:0] n353;
  wire [15:0] n354;
  wire [15:0] n355;
  wire [7:0] n357;
  wire [4:0] n359;
  wire [4:0] n361;
  wire [4:0] n362;
  wire [7:0] n363;
  wire [7:0] n369;
  wire [7:0] n371;
  wire [7:0] n372;
  wire [7:0] n374;
  wire [2:0] n384;
  wire [2:0] reg_address;  // sources/rtl/camera_init.v(43)
  wire [15:0] regs_data;  // sources/rtl/camera_init.v(76)
  wire  \sel0_b0/B0 ;
  wire  \sel0_b0/B3 ;
  wire  \sel0_b0/B4 ;
  wire  \sel0_b1/B0 ;
  wire  \sel0_b1/B3 ;
  wire  \sel0_b1/B4 ;
  wire  \sel0_b2/B0 ;
  wire  \sel0_b2/B3 ;
  wire  \sel0_b2/B4 ;
  wire  \sel0_b3/B0 ;
  wire  \sel0_b3/B3 ;
  wire  \sel0_b3/B4 ;
  wire  \sel0_b4/B0 ;
  wire  \sel0_b4/B3 ;
  wire  \sel0_b4/B4 ;
  wire  \sel0_b5/B0 ;
  wire  \sel0_b5/B3 ;
  wire  \sel0_b5/B4 ;
  wire  \sel0_b6/B0 ;
  wire  \sel0_b6/B3 ;
  wire  \sel0_b6/B4 ;
  wire  \sel0_b7/B0 ;
  wire  \sel0_b7/B3 ;
  wire  \sel0_b7/B4 ;
  wire  \sel2_b0/B6 ;
  wire  \sel2_b0/B7 ;
  wire  \sel2_b1/B6 ;
  wire  \sel2_b1/B7 ;
  wire  \sel2_b2/B6 ;
  wire  \sel2_b2/B7 ;
  wire  \sel2_b3/B6 ;
  wire  \sel2_b3/B7 ;
  wire  \sel2_b4/B6 ;
  wire  \sel2_b4/B7 ;
  wire  \sel2_b5/B6 ;
  wire  \sel2_b5/B7 ;
  wire  \sel2_b6/B6 ;
  wire  \sel2_b6/B7 ;
  wire  \sel2_b7/B6 ;
  wire  \sel2_b7/B7 ;
  wire [7:0] state_next;  // sources/rtl/camera_init.v(66)
  wire bus_write;  // sources/rtl/camera_init.v(44)
  wire mux100_b10_sel_is_0_o;
  wire mux100_b12_sel_is_2_o;
  wire mux100_b13_sel_is_2_o;
  wire mux100_b9_sel_is_0_o;
  wire mux100_b9_sel_is_0_o_neg;
  wire mux101_b0_sel_is_0_o;
  wire mux101_b12_sel_is_2_o;
  wire mux101_b13_sel_is_2_o;
  wire mux101_b1_sel_is_2_o;
  wire mux101_b9_sel_is_0_o;
  wire mux102_b0_sel_is_2_o;
  wire mux102_b10_sel_is_0_o;
  wire mux102_b12_sel_is_2_o;
  wire mux102_b13_sel_is_2_o;
  wire mux102_b13_sel_is_2_o_neg;
  wire mux102_b1_sel_is_2_o;
  wire mux102_b9_sel_is_2_o;
  wire mux103_b0_sel_is_2_o;
  wire mux103_b10_sel_is_2_o;
  wire mux103_b13_sel_is_0_o;
  wire mux103_b1_sel_is_2_o;
  wire mux103_b3_sel_is_0_o;
  wire mux103_b9_sel_is_2_o;
  wire mux104_b11_sel_is_2_o;
  wire mux104_b12_sel_is_0_o;
  wire mux104_b13_sel_is_2_o;
  wire mux104_b15_sel_is_2_o;
  wire mux104_b5_sel_is_2_o;
  wire mux104_b9_sel_is_2_o;
  wire mux104_b9_sel_is_2_o_neg;
  wire mux105_b11_sel_is_2_o;
  wire mux105_b13_sel_is_2_o;
  wire mux105_b13_sel_is_2_o_neg;
  wire mux105_b14_sel_is_0_o;
  wire mux105_b9_sel_is_0_o;
  wire mux106_b0_sel_is_0_o;
  wire mux106_b11_sel_is_2_o;
  wire mux106_b13_sel_is_0_o;
  wire mux106_b13_sel_is_0_o_neg;
  wire mux106_b14_sel_is_2_o;
  wire mux106_b9_sel_is_2_o;
  wire mux107_b0_sel_is_2_o;
  wire mux107_b13_sel_is_0_o;
  wire mux107_b14_sel_is_2_o;
  wire mux107_b4_sel_is_0_o;
  wire mux107_b9_sel_is_2_o;
  wire mux108_b13_sel_is_2_o;
  wire mux108_b14_sel_is_2_o;
  wire mux108_b15_sel_is_0_o;
  wire mux108_b8_sel_is_2_o;
  wire mux108_b9_sel_is_2_o;
  wire mux108_b9_sel_is_2_o_neg;
  wire mux109_b10_sel_is_0_o;
  wire mux109_b13_sel_is_2_o;
  wire mux109_b14_sel_is_2_o;
  wire mux109_b15_sel_is_2_o;
  wire mux109_b8_sel_is_2_o;
  wire mux109_b9_sel_is_0_o;
  wire mux109_b9_sel_is_0_o_neg;
  wire mux10_b10_sel_is_0_o;
  wire mux10_b11_sel_is_2_o;
  wire mux10_b12_sel_is_2_o;
  wire mux10_b13_sel_is_2_o;
  wire mux10_b14_sel_is_2_o;
  wire mux10_b9_sel_is_2_o;
  wire mux10_b9_sel_is_2_o_neg;
  wire mux110_b0_sel_is_0_o;
  wire mux110_b10_sel_is_2_o;
  wire mux110_b13_sel_is_2_o;
  wire mux110_b8_sel_is_2_o;
  wire mux110_b9_sel_is_0_o;
  wire mux111_b0_sel_is_2_o;
  wire mux111_b10_sel_is_2_o;
  wire mux111_b13_sel_is_2_o;
  wire mux111_b13_sel_is_2_o_neg;
  wire mux111_b15_sel_is_0_o;
  wire mux111_b8_sel_is_2_o;
  wire mux111_b9_sel_is_2_o;
  wire mux111_b9_sel_is_2_o_neg;
  wire mux112_b11_sel_is_2_o;
  wire mux112_b13_sel_is_0_o;
  wire mux112_b14_sel_is_0_o;
  wire mux112_b15_sel_is_2_o;
  wire mux112_b7_sel_is_2_o;
  wire mux112_b9_sel_is_0_o;
  wire mux112_b9_sel_is_0_o_neg;
  wire mux113_b10_sel_is_0_o;
  wire mux113_b13_sel_is_2_o;
  wire mux113_b14_sel_is_2_o;
  wire mux113_b15_sel_is_2_o;
  wire mux113_b2_sel_is_2_o;
  wire mux113_b9_sel_is_0_o;
  wire mux113_b9_sel_is_0_o_neg;
  wire mux114_b0_sel_is_0_o;
  wire mux114_b13_sel_is_2_o;
  wire mux114_b13_sel_is_2_o_neg;
  wire mux114_b14_sel_is_2_o;
  wire mux114_b15_sel_is_2_o;
  wire mux114_b2_sel_is_2_o;
  wire mux114_b9_sel_is_0_o;
  wire mux115_b0_sel_is_2_o;
  wire mux115_b10_sel_is_0_o;
  wire mux115_b13_sel_is_0_o;
  wire mux115_b15_sel_is_2_o;
  wire mux115_b2_sel_is_2_o;
  wire mux115_b4_sel_is_2_o;
  wire mux115_b9_sel_is_2_o;
  wire mux116_b11_sel_is_0_o;
  wire mux116_b13_sel_is_2_o;
  wire mux116_b13_sel_is_2_o_neg;
  wire mux116_b15_sel_is_2_o;
  wire mux116_b2_sel_is_2_o;
  wire mux116_b4_sel_is_2_o;
  wire mux116_b5_sel_is_2_o;
  wire mux116_b9_sel_is_2_o;
  wire mux117_b0_sel_is_0_o;
  wire mux117_b12_sel_is_2_o;
  wire mux117_b13_sel_is_0_o;
  wire mux117_b15_sel_is_2_o;
  wire mux117_b2_sel_is_2_o;
  wire mux117_b4_sel_is_2_o;
  wire mux117_b5_sel_is_2_o;
  wire mux117_b9_sel_is_2_o;
  wire mux117_b9_sel_is_2_o_neg;
  wire mux118_b10_sel_is_2_o;
  wire mux118_b11_sel_is_0_o;
  wire mux118_b12_sel_is_2_o;
  wire mux118_b13_sel_is_2_o;
  wire mux118_b15_sel_is_2_o;
  wire mux118_b2_sel_is_2_o;
  wire mux118_b4_sel_is_2_o;
  wire mux118_b5_sel_is_2_o;
  wire mux118_b9_sel_is_0_o;
  wire mux119_b10_sel_is_2_o;
  wire mux119_b11_sel_is_2_o;
  wire mux119_b12_sel_is_2_o;
  wire mux119_b13_sel_is_2_o;
  wire mux119_b15_sel_is_2_o;
  wire mux119_b2_sel_is_2_o;
  wire mux119_b3_sel_is_0_o;
  wire mux119_b4_sel_is_2_o;
  wire mux119_b5_sel_is_2_o;
  wire mux119_b9_sel_is_2_o;
  wire mux119_b9_sel_is_2_o_neg;
  wire mux11_b0_sel_is_0_o;
  wire mux11_b12_sel_is_2_o;
  wire mux11_b13_sel_is_2_o;
  wire mux11_b14_sel_is_2_o;
  wire mux11_b15_sel_is_2_o;
  wire mux11_b2_sel_is_2_o;
  wire mux11_b9_sel_is_0_o;
  wire mux120_b0_sel_is_0_o;
  wire mux120_b12_sel_is_2_o;
  wire mux120_b13_sel_is_2_o;
  wire mux120_b15_sel_is_2_o;
  wire mux120_b2_sel_is_2_o;
  wire mux120_b3_sel_is_2_o;
  wire mux120_b5_sel_is_2_o;
  wire mux120_b7_sel_is_2_o;
  wire mux120_b9_sel_is_0_o;
  wire mux121_b11_sel_is_0_o;
  wire mux121_b12_sel_is_2_o;
  wire mux121_b13_sel_is_2_o;
  wire mux121_b13_sel_is_2_o_neg;
  wire mux121_b15_sel_is_2_o;
  wire mux121_b2_sel_is_2_o;
  wire mux121_b3_sel_is_2_o;
  wire mux121_b5_sel_is_2_o;
  wire mux121_b7_sel_is_2_o;
  wire mux121_b9_sel_is_2_o;
  wire mux122_b10_sel_is_0_o;
  wire mux122_b11_sel_is_2_o;
  wire mux122_b12_sel_is_2_o;
  wire mux122_b13_sel_is_0_o;
  wire mux122_b15_sel_is_2_o;
  wire mux122_b2_sel_is_2_o;
  wire mux122_b3_sel_is_2_o;
  wire mux122_b5_sel_is_2_o;
  wire mux122_b9_sel_is_2_o;
  wire mux122_b9_sel_is_2_o_neg;
  wire mux123_b10_sel_is_2_o;
  wire mux123_b11_sel_is_2_o;
  wire mux123_b12_sel_is_2_o;
  wire mux123_b13_sel_is_2_o;
  wire mux123_b14_sel_is_0_o;
  wire mux123_b15_sel_is_2_o;
  wire mux123_b3_sel_is_2_o;
  wire mux123_b5_sel_is_2_o;
  wire mux123_b9_sel_is_0_o;
  wire mux124_b0_sel_is_0_o;
  wire mux124_b10_sel_is_2_o;
  wire mux124_b11_sel_is_2_o;
  wire mux124_b12_sel_is_2_o;
  wire mux124_b13_sel_is_2_o;
  wire mux124_b14_sel_is_2_o;
  wire mux124_b15_sel_is_2_o;
  wire mux124_b3_sel_is_2_o;
  wire mux124_b5_sel_is_2_o;
  wire mux124_b9_sel_is_2_o;
  wire mux124_b9_sel_is_2_o_neg;
  wire mux125_b0_sel_is_2_o;
  wire mux125_b13_sel_is_2_o;
  wire mux125_b14_sel_is_2_o;
  wire mux125_b15_sel_is_2_o;
  wire mux125_b2_sel_is_0_o;
  wire mux125_b3_sel_is_2_o;
  wire mux125_b5_sel_is_2_o;
  wire mux125_b9_sel_is_0_o;
  wire mux125_b9_sel_is_0_o_neg;
  wire mux126_b0_sel_is_2_o;
  wire mux126_b10_sel_is_0_o;
  wire mux126_b13_sel_is_2_o;
  wire mux126_b14_sel_is_2_o;
  wire mux126_b15_sel_is_2_o;
  wire mux126_b2_sel_is_2_o;
  wire mux126_b3_sel_is_2_o;
  wire mux126_b5_sel_is_2_o;
  wire mux126_b9_sel_is_0_o;
  wire mux127_b0_sel_is_2_o;
  wire mux127_b10_sel_is_2_o;
  wire mux127_b13_sel_is_2_o;
  wire mux127_b14_sel_is_2_o;
  wire mux127_b15_sel_is_2_o;
  wire mux127_b2_sel_is_2_o;
  wire mux127_b3_sel_is_2_o;
  wire mux127_b5_sel_is_2_o;
  wire mux127_b9_sel_is_2_o;
  wire mux128_b0_sel_is_2_o;
  wire mux128_b11_sel_is_2_o;
  wire mux128_b13_sel_is_2_o;
  wire mux128_b15_sel_is_2_o;
  wire mux128_b2_sel_is_2_o;
  wire mux128_b3_sel_is_2_o;
  wire mux128_b7_sel_is_0_o;
  wire mux128_b9_sel_is_2_o;
  wire mux129_b0_sel_is_2_o;
  wire mux129_b10_sel_is_0_o;
  wire mux129_b12_sel_is_2_o;
  wire mux129_b13_sel_is_2_o;
  wire mux129_b15_sel_is_2_o;
  wire mux129_b2_sel_is_2_o;
  wire mux129_b3_sel_is_2_o;
  wire mux129_b8_sel_is_2_o;
  wire mux129_b9_sel_is_2_o;
  wire mux12_b0_sel_is_2_o;
  wire mux12_b10_sel_is_0_o;
  wire mux12_b12_sel_is_2_o;
  wire mux12_b13_sel_is_2_o;
  wire mux12_b14_sel_is_2_o;
  wire mux12_b15_sel_is_2_o;
  wire mux12_b2_sel_is_2_o;
  wire mux12_b9_sel_is_2_o;
  wire mux12_b9_sel_is_2_o_neg;
  wire mux130_b13_sel_is_2_o;
  wire mux130_b15_sel_is_2_o;
  wire mux130_b1_sel_is_2_o;
  wire mux130_b3_sel_is_2_o;
  wire mux130_b4_sel_is_0_o;
  wire mux130_b6_sel_is_2_o;
  wire mux130_b8_sel_is_2_o;
  wire mux130_b9_sel_is_2_o;
  wire mux130_b9_sel_is_2_o_neg;
  wire mux131_b13_sel_is_2_o;
  wire mux131_b14_sel_is_0_o;
  wire mux131_b15_sel_is_2_o;
  wire mux131_b1_sel_is_2_o;
  wire mux131_b3_sel_is_2_o;
  wire mux131_b4_sel_is_2_o;
  wire mux131_b6_sel_is_2_o;
  wire mux131_b8_sel_is_2_o;
  wire mux131_b9_sel_is_0_o;
  wire mux131_b9_sel_is_0_o_neg;
  wire mux132_b0_sel_is_0_o;
  wire mux132_b13_sel_is_2_o;
  wire mux132_b13_sel_is_2_o_neg;
  wire mux132_b14_sel_is_2_o;
  wire mux132_b15_sel_is_2_o;
  wire mux132_b1_sel_is_2_o;
  wire mux132_b3_sel_is_2_o;
  wire mux132_b9_sel_is_0_o;
  wire mux133_b0_sel_is_2_o;
  wire mux133_b13_sel_is_0_o;
  wire mux133_b15_sel_is_2_o;
  wire mux133_b1_sel_is_2_o;
  wire mux133_b4_sel_is_0_o;
  wire mux133_b9_sel_is_2_o;
  wire mux133_b9_sel_is_2_o_neg;
  wire mux134_b0_sel_is_2_o;
  wire mux134_b10_sel_is_0_o;
  wire mux134_b13_sel_is_2_o;
  wire mux134_b13_sel_is_2_o_neg;
  wire mux134_b15_sel_is_2_o;
  wire mux134_b5_sel_is_2_o;
  wire mux134_b9_sel_is_0_o;
  wire mux135_b0_sel_is_2_o;
  wire mux135_b11_sel_is_0_o;
  wire mux135_b13_sel_is_0_o;
  wire mux135_b13_sel_is_0_o_neg;
  wire mux135_b15_sel_is_2_o;
  wire mux135_b6_sel_is_2_o;
  wire mux135_b7_sel_is_2_o;
  wire mux135_b9_sel_is_2_o;
  wire mux135_b9_sel_is_2_o_neg;
  wire mux136_b0_sel_is_2_o;
  wire mux136_b13_sel_is_0_o;
  wire mux136_b13_sel_is_0_o_neg;
  wire mux136_b14_sel_is_2_o;
  wire mux136_b15_sel_is_2_o;
  wire mux136_b1_sel_is_0_o;
  wire mux136_b6_sel_is_2_o;
  wire mux136_b7_sel_is_2_o;
  wire mux136_b9_sel_is_0_o;
  wire mux136_b9_sel_is_0_o_neg;
  wire mux137_b0_sel_is_2_o;
  wire mux137_b10_sel_is_0_o;
  wire mux137_b13_sel_is_0_o;
  wire mux137_b15_sel_is_2_o;
  wire mux137_b2_sel_is_2_o;
  wire mux137_b5_sel_is_2_o;
  wire mux137_b6_sel_is_2_o;
  wire mux137_b9_sel_is_0_o;
  wire mux137_b9_sel_is_0_o_neg;
  wire mux138_b0_sel_is_2_o;
  wire mux138_b10_sel_is_2_o;
  wire mux138_b11_sel_is_0_o;
  wire mux138_b13_sel_is_2_o;
  wire mux138_b15_sel_is_2_o;
  wire mux138_b2_sel_is_2_o;
  wire mux138_b6_sel_is_2_o;
  wire mux138_b9_sel_is_0_o;
  wire mux139_b0_sel_is_2_o;
  wire mux139_b10_sel_is_2_o;
  wire mux139_b11_sel_is_2_o;
  wire mux139_b13_sel_is_2_o;
  wire mux139_b15_sel_is_2_o;
  wire mux139_b1_sel_is_0_o;
  wire mux139_b2_sel_is_2_o;
  wire mux139_b9_sel_is_2_o;
  wire mux13_b0_sel_is_2_o;
  wire mux13_b11_sel_is_2_o;
  wire mux13_b12_sel_is_2_o;
  wire mux13_b13_sel_is_2_o;
  wire mux13_b14_sel_is_2_o;
  wire mux13_b15_sel_is_2_o;
  wire mux13_b2_sel_is_2_o;
  wire mux13_b9_sel_is_0_o;
  wire mux140_b11_sel_is_2_o;
  wire mux140_b13_sel_is_2_o;
  wire mux140_b13_sel_is_2_o_neg;
  wire mux140_b15_sel_is_2_o;
  wire mux140_b1_sel_is_2_o;
  wire mux140_b2_sel_is_2_o;
  wire mux140_b5_sel_is_0_o;
  wire mux140_b9_sel_is_2_o;
  wire mux140_b9_sel_is_2_o_neg;
  wire mux141_b0_sel_is_0_o;
  wire mux141_b12_sel_is_2_o;
  wire mux141_b13_sel_is_0_o;
  wire mux141_b15_sel_is_2_o;
  wire mux141_b1_sel_is_2_o;
  wire mux141_b2_sel_is_2_o;
  wire mux141_b5_sel_is_2_o;
  wire mux141_b9_sel_is_0_o;
  wire mux142_b0_sel_is_2_o;
  wire mux142_b12_sel_is_2_o;
  wire mux142_b13_sel_is_2_o;
  wire mux142_b14_sel_is_0_o;
  wire mux142_b15_sel_is_2_o;
  wire mux142_b2_sel_is_2_o;
  wire mux142_b5_sel_is_2_o;
  wire mux142_b9_sel_is_2_o;
  wire mux143_b10_sel_is_2_o;
  wire mux143_b13_sel_is_2_o;
  wire mux143_b14_sel_is_2_o;
  wire mux143_b15_sel_is_2_o;
  wire mux143_b2_sel_is_2_o;
  wire mux143_b5_sel_is_2_o;
  wire mux143_b7_sel_is_0_o;
  wire mux143_b9_sel_is_2_o;
  wire mux143_b9_sel_is_2_o_neg;
  wire mux144_b0_sel_is_0_o;
  wire mux144_b10_sel_is_2_o;
  wire mux144_b13_sel_is_2_o;
  wire mux144_b14_sel_is_2_o;
  wire mux144_b15_sel_is_2_o;
  wire mux144_b2_sel_is_2_o;
  wire mux144_b5_sel_is_2_o;
  wire mux144_b7_sel_is_2_o;
  wire mux144_b9_sel_is_0_o;
  wire mux145_b0_sel_is_2_o;
  wire mux145_b12_sel_is_0_o;
  wire mux145_b13_sel_is_2_o;
  wire mux145_b14_sel_is_2_o;
  wire mux145_b15_sel_is_2_o;
  wire mux145_b2_sel_is_2_o;
  wire mux145_b5_sel_is_2_o;
  wire mux145_b6_sel_is_2_o;
  wire mux145_b7_sel_is_2_o;
  wire mux145_b9_sel_is_2_o;
  wire mux145_b9_sel_is_2_o_neg;
  wire mux146_b10_sel_is_0_o;
  wire mux146_b11_sel_is_2_o;
  wire mux146_b12_sel_is_2_o;
  wire mux146_b13_sel_is_2_o;
  wire mux146_b15_sel_is_2_o;
  wire mux146_b2_sel_is_2_o;
  wire mux146_b3_sel_is_2_o;
  wire mux146_b5_sel_is_2_o;
  wire mux146_b7_sel_is_2_o;
  wire mux146_b9_sel_is_0_o;
  wire mux146_b9_sel_is_0_o_neg;
  wire mux147_b0_sel_is_0_o;
  wire mux147_b10_sel_is_2_o;
  wire mux147_b11_sel_is_2_o;
  wire mux147_b12_sel_is_2_o;
  wire mux147_b13_sel_is_2_o;
  wire mux147_b15_sel_is_2_o;
  wire mux147_b3_sel_is_2_o;
  wire mux147_b5_sel_is_2_o;
  wire mux147_b9_sel_is_0_o;
  wire mux147_b9_sel_is_0_o_neg;
  wire mux148_b10_sel_is_2_o;
  wire mux148_b12_sel_is_2_o;
  wire mux148_b13_sel_is_2_o;
  wire mux148_b14_sel_is_2_o;
  wire mux148_b15_sel_is_2_o;
  wire mux148_b3_sel_is_2_o;
  wire mux148_b5_sel_is_2_o;
  wire mux148_b7_sel_is_0_o;
  wire mux148_b9_sel_is_0_o;
  wire mux149_b0_sel_is_0_o;
  wire mux149_b10_sel_is_2_o;
  wire mux149_b12_sel_is_2_o;
  wire mux149_b13_sel_is_2_o;
  wire mux149_b13_sel_is_2_o_neg;
  wire mux149_b14_sel_is_2_o;
  wire mux149_b15_sel_is_2_o;
  wire mux149_b4_sel_is_2_o;
  wire mux149_b5_sel_is_2_o;
  wire mux149_b7_sel_is_2_o;
  wire mux149_b9_sel_is_2_o;
  wire mux14_b0_sel_is_2_o;
  wire mux14_b10_sel_is_0_o;
  wire mux14_b11_sel_is_2_o;
  wire mux14_b12_sel_is_2_o;
  wire mux14_b13_sel_is_2_o;
  wire mux14_b14_sel_is_2_o;
  wire mux14_b15_sel_is_2_o;
  wire mux14_b6_sel_is_2_o;
  wire mux14_b9_sel_is_2_o;
  wire mux14_b9_sel_is_2_o_neg;
  wire mux150_b0_sel_is_2_o;
  wire mux150_b10_sel_is_2_o;
  wire mux150_b13_sel_is_0_o;
  wire mux150_b14_sel_is_2_o;
  wire mux150_b15_sel_is_2_o;
  wire mux150_b3_sel_is_0_o;
  wire mux150_b5_sel_is_2_o;
  wire mux150_b9_sel_is_2_o;
  wire mux150_b9_sel_is_2_o_neg;
  wire mux151_b0_sel_is_2_o;
  wire mux151_b10_sel_is_2_o;
  wire mux151_b12_sel_is_0_o;
  wire mux151_b13_sel_is_2_o;
  wire mux151_b14_sel_is_2_o;
  wire mux151_b15_sel_is_2_o;
  wire mux151_b5_sel_is_2_o;
  wire mux151_b8_sel_is_2_o;
  wire mux151_b9_sel_is_0_o;
  wire mux151_b9_sel_is_0_o_neg;
  wire mux152_b0_sel_is_2_o;
  wire mux152_b13_sel_is_2_o;
  wire mux152_b14_sel_is_2_o;
  wire mux152_b15_sel_is_2_o;
  wire mux152_b1_sel_is_0_o;
  wire mux152_b5_sel_is_2_o;
  wire mux152_b9_sel_is_0_o;
  wire mux153_b11_sel_is_2_o;
  wire mux153_b13_sel_is_2_o;
  wire mux153_b14_sel_is_2_o;
  wire mux153_b15_sel_is_2_o;
  wire mux153_b3_sel_is_2_o;
  wire mux153_b5_sel_is_2_o;
  wire mux153_b8_sel_is_0_o;
  wire mux153_b9_sel_is_2_o;
  wire mux154_b11_sel_is_2_o;
  wire mux154_b13_sel_is_2_o;
  wire mux154_b14_sel_is_2_o;
  wire mux154_b15_sel_is_2_o;
  wire mux154_b1_sel_is_0_o;
  wire mux154_b5_sel_is_2_o;
  wire mux154_b9_sel_is_2_o;
  wire mux154_b9_sel_is_2_o_neg;
  wire mux155_b0_sel_is_0_o;
  wire mux155_b11_sel_is_2_o;
  wire mux155_b13_sel_is_2_o;
  wire mux155_b14_sel_is_2_o;
  wire mux155_b15_sel_is_2_o;
  wire mux155_b1_sel_is_2_o;
  wire mux155_b5_sel_is_2_o;
  wire mux155_b9_sel_is_0_o;
  wire mux156_b0_sel_is_2_o;
  wire mux156_b12_sel_is_0_o;
  wire mux156_b13_sel_is_2_o;
  wire mux156_b13_sel_is_2_o_neg;
  wire mux156_b14_sel_is_2_o;
  wire mux156_b15_sel_is_2_o;
  wire mux156_b1_sel_is_2_o;
  wire mux156_b2_sel_is_2_o;
  wire mux156_b5_sel_is_2_o;
  wire mux156_b9_sel_is_2_o;
  wire mux156_b9_sel_is_2_o_neg;
  wire mux157_b0_sel_is_2_o;
  wire mux157_b12_sel_is_2_o;
  wire mux157_b13_sel_is_0_o;
  wire mux157_b14_sel_is_2_o;
  wire mux157_b15_sel_is_2_o;
  wire mux157_b2_sel_is_2_o;
  wire mux157_b3_sel_is_0_o;
  wire mux157_b5_sel_is_2_o;
  wire mux157_b9_sel_is_0_o;
  wire mux158_b11_sel_is_0_o;
  wire mux158_b13_sel_is_2_o;
  wire mux158_b13_sel_is_2_o_neg;
  wire mux158_b15_sel_is_2_o;
  wire mux158_b2_sel_is_2_o;
  wire mux158_b3_sel_is_2_o;
  wire mux158_b4_sel_is_2_o;
  wire mux158_b5_sel_is_2_o;
  wire mux158_b9_sel_is_2_o;
  wire mux159_b13_sel_is_0_o;
  wire mux159_b15_sel_is_2_o;
  wire mux159_b1_sel_is_2_o;
  wire mux159_b2_sel_is_2_o;
  wire mux159_b3_sel_is_2_o;
  wire mux159_b5_sel_is_2_o;
  wire mux159_b9_sel_is_2_o;
  wire mux15_b0_sel_is_2_o;
  wire mux15_b10_sel_is_2_o;
  wire mux15_b11_sel_is_2_o;
  wire mux15_b12_sel_is_2_o;
  wire mux15_b13_sel_is_2_o;
  wire mux15_b14_sel_is_2_o;
  wire mux15_b15_sel_is_2_o;
  wire mux15_b7_sel_is_0_o;
  wire mux15_b9_sel_is_0_o;
  wire mux160_b11_sel_is_0_o;
  wire mux160_b13_sel_is_2_o;
  wire mux160_b15_sel_is_2_o;
  wire mux160_b2_sel_is_2_o;
  wire mux160_b9_sel_is_2_o;
  wire mux161_b0_sel_is_0_o;
  wire mux161_b11_sel_is_2_o;
  wire mux161_b13_sel_is_2_o;
  wire mux161_b15_sel_is_2_o;
  wire mux161_b2_sel_is_2_o;
  wire mux161_b9_sel_is_2_o;
  wire mux162_b10_sel_is_2_o;
  wire mux162_b12_sel_is_2_o;
  wire mux162_b13_sel_is_2_o;
  wire mux162_b15_sel_is_2_o;
  wire mux162_b2_sel_is_2_o;
  wire mux162_b7_sel_is_0_o;
  wire mux162_b9_sel_is_2_o;
  wire mux162_b9_sel_is_2_o_neg;
  wire mux163_b0_sel_is_0_o;
  wire mux163_b13_sel_is_2_o;
  wire mux163_b13_sel_is_2_o_neg;
  wire mux163_b14_sel_is_2_o;
  wire mux163_b15_sel_is_2_o;
  wire mux163_b7_sel_is_2_o;
  wire mux163_b9_sel_is_0_o;
  wire mux164_b0_sel_is_2_o;
  wire mux164_b10_sel_is_0_o;
  wire mux164_b13_sel_is_0_o;
  wire mux164_b14_sel_is_2_o;
  wire mux164_b15_sel_is_2_o;
  wire mux164_b7_sel_is_2_o;
  wire mux164_b9_sel_is_2_o;
  wire mux164_b9_sel_is_2_o_neg;
  wire mux165_b11_sel_is_0_o;
  wire mux165_b13_sel_is_2_o;
  wire mux165_b14_sel_is_2_o;
  wire mux165_b15_sel_is_2_o;
  wire mux165_b1_sel_is_2_o;
  wire mux165_b4_sel_is_2_o;
  wire mux165_b9_sel_is_0_o;
  wire mux165_b9_sel_is_0_o_neg;
  wire mux166_b11_sel_is_2_o;
  wire mux166_b13_sel_is_2_o;
  wire mux166_b14_sel_is_2_o;
  wire mux166_b15_sel_is_2_o;
  wire mux166_b1_sel_is_2_o;
  wire mux166_b4_sel_is_2_o;
  wire mux166_b5_sel_is_0_o;
  wire mux166_b9_sel_is_0_o;
  wire mux167_b0_sel_is_0_o;
  wire mux167_b13_sel_is_2_o;
  wire mux167_b14_sel_is_2_o;
  wire mux167_b15_sel_is_2_o;
  wire mux167_b4_sel_is_2_o;
  wire mux167_b9_sel_is_2_o;
  wire mux168_b0_sel_is_2_o;
  wire mux168_b10_sel_is_0_o;
  wire mux168_b13_sel_is_2_o;
  wire mux168_b13_sel_is_2_o_neg;
  wire mux168_b14_sel_is_2_o;
  wire mux168_b15_sel_is_2_o;
  wire mux168_b4_sel_is_2_o;
  wire mux168_b9_sel_is_2_o;
  wire mux169_b0_sel_is_2_o;
  wire mux169_b12_sel_is_0_o;
  wire mux169_b13_sel_is_0_o;
  wire mux169_b14_sel_is_2_o;
  wire mux169_b15_sel_is_2_o;
  wire mux169_b3_sel_is_2_o;
  wire mux169_b9_sel_is_2_o;
  wire mux169_b9_sel_is_2_o_neg;
  wire mux16_b0_sel_is_2_o;
  wire mux16_b10_sel_is_2_o;
  wire mux16_b11_sel_is_2_o;
  wire mux16_b12_sel_is_2_o;
  wire mux16_b13_sel_is_2_o;
  wire mux16_b14_sel_is_2_o;
  wire mux16_b15_sel_is_2_o;
  wire mux16_b1_sel_is_0_o;
  wire mux16_b9_sel_is_2_o;
  wire mux16_b9_sel_is_2_o_neg;
  wire mux170_b10_sel_is_0_o;
  wire mux170_b12_sel_is_2_o;
  wire mux170_b13_sel_is_2_o;
  wire mux170_b2_sel_is_2_o;
  wire mux170_b3_sel_is_2_o;
  wire mux170_b9_sel_is_0_o;
  wire mux171_b0_sel_is_0_o;
  wire mux171_b10_sel_is_2_o;
  wire mux171_b13_sel_is_2_o;
  wire mux171_b9_sel_is_2_o;
  wire mux171_b9_sel_is_2_o_neg;
  wire mux172_b0_sel_is_2_o;
  wire mux172_b10_sel_is_2_o;
  wire mux172_b12_sel_is_0_o;
  wire mux172_b13_sel_is_2_o;
  wire mux172_b9_sel_is_0_o;
  wire mux172_b9_sel_is_0_o_neg;
  wire mux173_b10_sel_is_2_o;
  wire mux173_b13_sel_is_2_o;
  wire mux173_b13_sel_is_2_o_neg;
  wire mux173_b9_sel_is_0_o;
  wire mux174_b0_sel_is_0_o;
  wire mux174_b13_sel_is_0_o;
  wire mux174_b13_sel_is_0_o_neg;
  wire mux174_b9_sel_is_2_o;
  wire mux175_b12_sel_is_2_o;
  wire mux175_b13_sel_is_0_o;
  wire mux175_b9_sel_is_2_o;
  wire mux177_b1_sel_is_3_o;
  wire mux17_b11_sel_is_2_o;
  wire mux17_b13_sel_is_2_o;
  wire mux17_b1_sel_is_2_o;
  wire mux17_b6_sel_is_0_o;
  wire mux17_b9_sel_is_0_o;
  wire mux17_b9_sel_is_0_o_neg;
  wire mux181_b0_sel_is_2_o;
  wire mux18_b10_sel_is_0_o;
  wire mux18_b13_sel_is_2_o;
  wire mux18_b1_sel_is_2_o;
  wire mux18_b6_sel_is_2_o;
  wire mux18_b9_sel_is_0_o;
  wire mux19_b12_sel_is_2_o;
  wire mux19_b13_sel_is_2_o;
  wire mux19_b2_sel_is_0_o;
  wire mux19_b7_sel_is_2_o;
  wire mux19_b9_sel_is_2_o;
  wire mux1_b7_sel_is_0_o;
  wire mux20_b10_sel_is_0_o;
  wire mux20_b12_sel_is_2_o;
  wire mux20_b13_sel_is_2_o;
  wire mux20_b4_sel_is_2_o;
  wire mux20_b7_sel_is_2_o;
  wire mux20_b9_sel_is_2_o;
  wire mux21_b0_sel_is_0_o;
  wire mux21_b11_sel_is_2_o;
  wire mux21_b12_sel_is_2_o;
  wire mux21_b13_sel_is_2_o;
  wire mux21_b13_sel_is_2_o_neg;
  wire mux21_b7_sel_is_2_o;
  wire mux21_b9_sel_is_2_o;
  wire mux21_b9_sel_is_2_o_neg;
  wire mux22_b11_sel_is_2_o;
  wire mux22_b13_sel_is_0_o;
  wire mux22_b15_sel_is_2_o;
  wire mux22_b2_sel_is_2_o;
  wire mux22_b3_sel_is_0_o;
  wire mux22_b7_sel_is_2_o;
  wire mux22_b9_sel_is_0_o;
  wire mux22_b9_sel_is_0_o_neg;
  wire mux23_b10_sel_is_0_o;
  wire mux23_b11_sel_is_2_o;
  wire mux23_b13_sel_is_2_o;
  wire mux23_b15_sel_is_2_o;
  wire mux23_b2_sel_is_2_o;
  wire mux23_b5_sel_is_2_o;
  wire mux23_b9_sel_is_0_o;
  wire mux24_b10_sel_is_2_o;
  wire mux24_b11_sel_is_2_o;
  wire mux24_b13_sel_is_2_o;
  wire mux24_b15_sel_is_2_o;
  wire mux24_b1_sel_is_0_o;
  wire mux24_b2_sel_is_2_o;
  wire mux24_b5_sel_is_2_o;
  wire mux24_b9_sel_is_2_o;
  wire mux25_b0_sel_is_0_o;
  wire mux25_b11_sel_is_2_o;
  wire mux25_b12_sel_is_2_o;
  wire mux25_b13_sel_is_2_o;
  wire mux25_b15_sel_is_2_o;
  wire mux25_b2_sel_is_2_o;
  wire mux25_b7_sel_is_2_o;
  wire mux25_b9_sel_is_2_o;
  wire mux26_b0_sel_is_2_o;
  wire mux26_b10_sel_is_0_o;
  wire mux26_b11_sel_is_2_o;
  wire mux26_b12_sel_is_2_o;
  wire mux26_b13_sel_is_2_o;
  wire mux26_b15_sel_is_2_o;
  wire mux26_b2_sel_is_2_o;
  wire mux26_b7_sel_is_2_o;
  wire mux26_b9_sel_is_2_o;
  wire mux26_b9_sel_is_2_o_neg;
  wire mux27_b0_sel_is_2_o;
  wire mux27_b11_sel_is_2_o;
  wire mux27_b12_sel_is_2_o;
  wire mux27_b13_sel_is_2_o;
  wire mux27_b15_sel_is_2_o;
  wire mux27_b1_sel_is_2_o;
  wire mux27_b2_sel_is_2_o;
  wire mux27_b6_sel_is_0_o;
  wire mux27_b7_sel_is_2_o;
  wire mux27_b9_sel_is_0_o;
  wire mux27_b9_sel_is_0_o_neg;
  wire mux28_b10_sel_is_0_o;
  wire mux28_b12_sel_is_2_o;
  wire mux28_b13_sel_is_2_o;
  wire mux28_b15_sel_is_2_o;
  wire mux28_b2_sel_is_2_o;
  wire mux28_b9_sel_is_0_o;
  wire mux28_b9_sel_is_0_o_neg;
  wire mux29_b0_sel_is_0_o;
  wire mux29_b12_sel_is_2_o;
  wire mux29_b13_sel_is_2_o;
  wire mux29_b15_sel_is_2_o;
  wire mux29_b2_sel_is_2_o;
  wire mux29_b5_sel_is_2_o;
  wire mux29_b9_sel_is_0_o;
  wire mux29_b9_sel_is_0_o_neg;
  wire mux2_b11_sel_is_0_o;
  wire mux2_b7_sel_is_2_o;
  wire mux30_b12_sel_is_2_o;
  wire mux30_b13_sel_is_2_o;
  wire mux30_b15_sel_is_2_o;
  wire mux30_b1_sel_is_2_o;
  wire mux30_b2_sel_is_2_o;
  wire mux30_b3_sel_is_0_o;
  wire mux30_b5_sel_is_2_o;
  wire mux30_b9_sel_is_0_o;
  wire mux30_b9_sel_is_0_o_neg;
  wire mux31_b12_sel_is_2_o;
  wire mux31_b13_sel_is_2_o;
  wire mux31_b13_sel_is_2_o_neg;
  wire mux31_b15_sel_is_2_o;
  wire mux31_b2_sel_is_2_o;
  wire mux31_b3_sel_is_2_o;
  wire mux31_b5_sel_is_2_o;
  wire mux31_b8_sel_is_0_o;
  wire mux31_b9_sel_is_0_o;
  wire mux32_b0_sel_is_0_o;
  wire mux32_b13_sel_is_0_o;
  wire mux32_b13_sel_is_0_o_neg;
  wire mux32_b15_sel_is_2_o;
  wire mux32_b3_sel_is_2_o;
  wire mux32_b9_sel_is_2_o;
  wire mux33_b0_sel_is_2_o;
  wire mux33_b13_sel_is_0_o;
  wire mux33_b13_sel_is_0_o_neg;
  wire mux33_b15_sel_is_2_o;
  wire mux33_b1_sel_is_0_o;
  wire mux33_b3_sel_is_2_o;
  wire mux33_b9_sel_is_2_o;
  wire mux34_b10_sel_is_2_o;
  wire mux34_b13_sel_is_0_o;
  wire mux34_b15_sel_is_2_o;
  wire mux34_b1_sel_is_2_o;
  wire mux34_b3_sel_is_2_o;
  wire mux34_b9_sel_is_2_o;
  wire mux34_b9_sel_is_2_o_neg;
  wire mux35_b0_sel_is_0_o;
  wire mux35_b10_sel_is_2_o;
  wire mux35_b13_sel_is_2_o;
  wire mux35_b13_sel_is_2_o_neg;
  wire mux35_b15_sel_is_2_o;
  wire mux35_b1_sel_is_2_o;
  wire mux35_b3_sel_is_2_o;
  wire mux35_b9_sel_is_0_o;
  wire mux36_b12_sel_is_2_o;
  wire mux36_b13_sel_is_0_o;
  wire mux36_b15_sel_is_2_o;
  wire mux36_b1_sel_is_2_o;
  wire mux36_b3_sel_is_2_o;
  wire mux36_b6_sel_is_0_o;
  wire mux36_b9_sel_is_2_o;
  wire mux37_b0_sel_is_0_o;
  wire mux37_b12_sel_is_2_o;
  wire mux37_b13_sel_is_2_o;
  wire mux37_b13_sel_is_2_o_neg;
  wire mux37_b15_sel_is_2_o;
  wire mux37_b1_sel_is_2_o;
  wire mux37_b3_sel_is_2_o;
  wire mux37_b6_sel_is_2_o;
  wire mux37_b9_sel_is_2_o;
  wire mux37_b9_sel_is_2_o_neg;
  wire mux38_b11_sel_is_0_o;
  wire mux38_b12_sel_is_2_o;
  wire mux38_b13_sel_is_0_o;
  wire mux38_b15_sel_is_2_o;
  wire mux38_b1_sel_is_2_o;
  wire mux38_b4_sel_is_2_o;
  wire mux38_b9_sel_is_0_o;
  wire mux39_b11_sel_is_2_o;
  wire mux39_b13_sel_is_2_o;
  wire mux39_b15_sel_is_2_o;
  wire mux39_b1_sel_is_2_o;
  wire mux39_b4_sel_is_2_o;
  wire mux39_b8_sel_is_0_o;
  wire mux39_b9_sel_is_2_o;
  wire mux3_b11_sel_is_2_o;
  wire mux3_b13_sel_is_2_o_neg;
  wire mux3_b7_sel_is_2_o;
  wire mux3_b8_sel_is_0_o;
  wire mux40_b0_sel_is_0_o;
  wire mux40_b11_sel_is_2_o;
  wire mux40_b13_sel_is_2_o;
  wire mux40_b15_sel_is_2_o;
  wire mux40_b1_sel_is_2_o;
  wire mux40_b4_sel_is_2_o;
  wire mux40_b8_sel_is_2_o;
  wire mux40_b9_sel_is_2_o;
  wire mux41_b0_sel_is_2_o;
  wire mux41_b11_sel_is_2_o;
  wire mux41_b13_sel_is_2_o;
  wire mux41_b15_sel_is_2_o;
  wire mux41_b1_sel_is_2_o;
  wire mux41_b4_sel_is_2_o;
  wire mux41_b8_sel_is_2_o;
  wire mux41_b9_sel_is_2_o;
  wire mux42_b0_sel_is_2_o;
  wire mux42_b11_sel_is_2_o;
  wire mux42_b13_sel_is_2_o;
  wire mux42_b15_sel_is_2_o;
  wire mux42_b1_sel_is_2_o;
  wire mux42_b7_sel_is_0_o;
  wire mux42_b8_sel_is_2_o;
  wire mux42_b9_sel_is_2_o;
  wire mux43_b0_sel_is_2_o;
  wire mux43_b11_sel_is_2_o;
  wire mux43_b13_sel_is_2_o;
  wire mux43_b15_sel_is_2_o;
  wire mux43_b8_sel_is_2_o;
  wire mux43_b9_sel_is_2_o;
  wire mux44_b0_sel_is_2_o;
  wire mux44_b11_sel_is_2_o;
  wire mux44_b13_sel_is_2_o;
  wire mux44_b15_sel_is_2_o;
  wire mux44_b1_sel_is_0_o;
  wire mux44_b8_sel_is_2_o;
  wire mux44_b9_sel_is_2_o;
  wire mux45_b0_sel_is_2_o;
  wire mux45_b11_sel_is_2_o;
  wire mux45_b13_sel_is_2_o;
  wire mux45_b15_sel_is_2_o;
  wire mux45_b4_sel_is_2_o;
  wire mux45_b5_sel_is_0_o;
  wire mux45_b8_sel_is_2_o;
  wire mux45_b9_sel_is_2_o;
  wire mux46_b0_sel_is_2_o;
  wire mux46_b11_sel_is_2_o;
  wire mux46_b13_sel_is_2_o;
  wire mux46_b15_sel_is_2_o;
  wire mux46_b1_sel_is_0_o;
  wire mux46_b5_sel_is_2_o;
  wire mux46_b7_sel_is_2_o;
  wire mux46_b8_sel_is_2_o;
  wire mux46_b9_sel_is_2_o;
  wire mux47_b0_sel_is_2_o;
  wire mux47_b11_sel_is_2_o;
  wire mux47_b13_sel_is_2_o;
  wire mux47_b15_sel_is_2_o;
  wire mux47_b1_sel_is_2_o;
  wire mux47_b3_sel_is_0_o;
  wire mux47_b5_sel_is_2_o;
  wire mux47_b7_sel_is_2_o;
  wire mux47_b8_sel_is_2_o;
  wire mux47_b9_sel_is_2_o;
  wire mux48_b0_sel_is_2_o;
  wire mux48_b11_sel_is_2_o;
  wire mux48_b13_sel_is_2_o;
  wire mux48_b15_sel_is_2_o;
  wire mux48_b1_sel_is_2_o;
  wire mux48_b2_sel_is_0_o;
  wire mux48_b7_sel_is_2_o;
  wire mux48_b8_sel_is_2_o;
  wire mux48_b9_sel_is_2_o;
  wire mux49_b0_sel_is_2_o;
  wire mux49_b11_sel_is_2_o;
  wire mux49_b13_sel_is_2_o;
  wire mux49_b15_sel_is_2_o;
  wire mux49_b4_sel_is_2_o;
  wire mux49_b5_sel_is_0_o;
  wire mux49_b7_sel_is_2_o;
  wire mux49_b8_sel_is_2_o;
  wire mux49_b9_sel_is_2_o;
  wire mux4_b13_sel_is_0_o;
  wire mux4_b13_sel_is_0_o_neg;
  wire mux4_b14_sel_is_2_o;
  wire mux4_b5_sel_is_0_o;
  wire mux4_b7_sel_is_2_o;
  wire mux50_b10_sel_is_2_o;
  wire mux50_b11_sel_is_2_o;
  wire mux50_b13_sel_is_2_o;
  wire mux50_b15_sel_is_2_o;
  wire mux50_b2_sel_is_0_o;
  wire mux50_b5_sel_is_2_o;
  wire mux50_b7_sel_is_2_o;
  wire mux50_b8_sel_is_2_o;
  wire mux50_b9_sel_is_2_o;
  wire mux51_b10_sel_is_2_o;
  wire mux51_b11_sel_is_2_o;
  wire mux51_b13_sel_is_2_o;
  wire mux51_b15_sel_is_2_o;
  wire mux51_b1_sel_is_0_o;
  wire mux51_b2_sel_is_2_o;
  wire mux51_b5_sel_is_2_o;
  wire mux51_b7_sel_is_2_o;
  wire mux51_b8_sel_is_2_o;
  wire mux51_b9_sel_is_2_o;
  wire mux52_b0_sel_is_0_o;
  wire mux52_b10_sel_is_2_o;
  wire mux52_b11_sel_is_2_o;
  wire mux52_b13_sel_is_2_o;
  wire mux52_b15_sel_is_2_o;
  wire mux52_b1_sel_is_2_o;
  wire mux52_b2_sel_is_2_o;
  wire mux52_b5_sel_is_2_o;
  wire mux52_b7_sel_is_2_o;
  wire mux52_b9_sel_is_2_o;
  wire mux53_b0_sel_is_2_o;
  wire mux53_b11_sel_is_2_o;
  wire mux53_b12_sel_is_2_o;
  wire mux53_b13_sel_is_2_o;
  wire mux53_b15_sel_is_2_o;
  wire mux53_b1_sel_is_2_o;
  wire mux53_b2_sel_is_2_o;
  wire mux53_b3_sel_is_0_o;
  wire mux53_b5_sel_is_2_o;
  wire mux53_b7_sel_is_2_o;
  wire mux53_b9_sel_is_2_o;
  wire mux54_b0_sel_is_2_o;
  wire mux54_b10_sel_is_0_o;
  wire mux54_b11_sel_is_2_o;
  wire mux54_b12_sel_is_2_o;
  wire mux54_b13_sel_is_2_o;
  wire mux54_b15_sel_is_2_o;
  wire mux54_b1_sel_is_2_o;
  wire mux54_b2_sel_is_2_o;
  wire mux54_b3_sel_is_2_o;
  wire mux54_b5_sel_is_2_o;
  wire mux54_b7_sel_is_2_o;
  wire mux54_b9_sel_is_2_o;
  wire mux55_b0_sel_is_2_o;
  wire mux55_b10_sel_is_2_o;
  wire mux55_b11_sel_is_2_o;
  wire mux55_b12_sel_is_2_o;
  wire mux55_b13_sel_is_2_o;
  wire mux55_b15_sel_is_2_o;
  wire mux55_b1_sel_is_2_o;
  wire mux55_b2_sel_is_2_o;
  wire mux55_b3_sel_is_2_o;
  wire mux55_b5_sel_is_2_o;
  wire mux55_b7_sel_is_2_o;
  wire mux55_b9_sel_is_2_o;
  wire mux56_b0_sel_is_2_o;
  wire mux56_b10_sel_is_2_o;
  wire mux56_b11_sel_is_2_o;
  wire mux56_b12_sel_is_2_o;
  wire mux56_b13_sel_is_2_o;
  wire mux56_b15_sel_is_2_o;
  wire mux56_b1_sel_is_2_o;
  wire mux56_b2_sel_is_2_o;
  wire mux56_b3_sel_is_2_o;
  wire mux56_b5_sel_is_2_o;
  wire mux56_b7_sel_is_2_o;
  wire mux56_b9_sel_is_2_o;
  wire mux57_b0_sel_is_2_o;
  wire mux57_b10_sel_is_2_o;
  wire mux57_b11_sel_is_2_o;
  wire mux57_b12_sel_is_2_o;
  wire mux57_b13_sel_is_2_o;
  wire mux57_b15_sel_is_2_o;
  wire mux57_b1_sel_is_2_o;
  wire mux57_b2_sel_is_2_o;
  wire mux57_b3_sel_is_2_o;
  wire mux57_b5_sel_is_2_o;
  wire mux57_b7_sel_is_2_o;
  wire mux57_b9_sel_is_2_o;
  wire mux58_b0_sel_is_2_o;
  wire mux58_b10_sel_is_2_o;
  wire mux58_b11_sel_is_2_o;
  wire mux58_b12_sel_is_2_o;
  wire mux58_b13_sel_is_2_o;
  wire mux58_b15_sel_is_2_o;
  wire mux58_b1_sel_is_2_o;
  wire mux58_b2_sel_is_2_o;
  wire mux58_b3_sel_is_2_o;
  wire mux58_b5_sel_is_2_o;
  wire mux58_b7_sel_is_2_o;
  wire mux58_b9_sel_is_2_o;
  wire mux59_b0_sel_is_2_o;
  wire mux59_b10_sel_is_2_o;
  wire mux59_b11_sel_is_2_o;
  wire mux59_b12_sel_is_2_o;
  wire mux59_b13_sel_is_2_o;
  wire mux59_b15_sel_is_2_o;
  wire mux59_b1_sel_is_2_o;
  wire mux59_b2_sel_is_2_o;
  wire mux59_b3_sel_is_2_o;
  wire mux59_b5_sel_is_2_o;
  wire mux59_b7_sel_is_2_o;
  wire mux59_b9_sel_is_2_o;
  wire mux5_b0_sel_is_0_o;
  wire mux5_b13_sel_is_0_o;
  wire mux5_b13_sel_is_0_o_neg;
  wire mux5_b5_sel_is_2_o;
  wire mux5_b7_sel_is_2_o;
  wire mux60_b0_sel_is_2_o;
  wire mux60_b10_sel_is_2_o;
  wire mux60_b11_sel_is_2_o;
  wire mux60_b12_sel_is_2_o;
  wire mux60_b13_sel_is_2_o;
  wire mux60_b15_sel_is_2_o;
  wire mux60_b1_sel_is_2_o;
  wire mux60_b3_sel_is_2_o;
  wire mux60_b5_sel_is_2_o;
  wire mux60_b7_sel_is_2_o;
  wire mux60_b9_sel_is_2_o;
  wire mux61_b0_sel_is_2_o;
  wire mux61_b10_sel_is_2_o;
  wire mux61_b11_sel_is_2_o;
  wire mux61_b12_sel_is_2_o;
  wire mux61_b13_sel_is_2_o;
  wire mux61_b15_sel_is_2_o;
  wire mux61_b1_sel_is_2_o;
  wire mux61_b3_sel_is_2_o;
  wire mux61_b5_sel_is_2_o;
  wire mux61_b7_sel_is_2_o;
  wire mux61_b9_sel_is_2_o;
  wire mux62_b10_sel_is_2_o;
  wire mux62_b11_sel_is_2_o;
  wire mux62_b12_sel_is_2_o;
  wire mux62_b13_sel_is_2_o;
  wire mux62_b15_sel_is_2_o;
  wire mux62_b1_sel_is_2_o;
  wire mux62_b3_sel_is_2_o;
  wire mux62_b4_sel_is_2_o;
  wire mux62_b5_sel_is_2_o;
  wire mux62_b7_sel_is_2_o;
  wire mux62_b9_sel_is_2_o;
  wire mux63_b0_sel_is_0_o;
  wire mux63_b10_sel_is_2_o;
  wire mux63_b11_sel_is_2_o;
  wire mux63_b12_sel_is_2_o;
  wire mux63_b13_sel_is_2_o;
  wire mux63_b15_sel_is_2_o;
  wire mux63_b1_sel_is_2_o;
  wire mux63_b3_sel_is_2_o;
  wire mux63_b4_sel_is_2_o;
  wire mux63_b5_sel_is_2_o;
  wire mux63_b7_sel_is_2_o;
  wire mux63_b9_sel_is_2_o;
  wire mux64_b0_sel_is_2_o;
  wire mux64_b10_sel_is_2_o;
  wire mux64_b11_sel_is_2_o;
  wire mux64_b12_sel_is_2_o;
  wire mux64_b13_sel_is_2_o;
  wire mux64_b15_sel_is_2_o;
  wire mux64_b3_sel_is_2_o;
  wire mux64_b4_sel_is_2_o;
  wire mux64_b9_sel_is_2_o;
  wire mux65_b10_sel_is_2_o;
  wire mux65_b11_sel_is_2_o;
  wire mux65_b12_sel_is_2_o;
  wire mux65_b13_sel_is_2_o;
  wire mux65_b15_sel_is_2_o;
  wire mux65_b1_sel_is_0_o;
  wire mux65_b3_sel_is_2_o;
  wire mux65_b4_sel_is_2_o;
  wire mux65_b9_sel_is_2_o;
  wire mux66_b0_sel_is_0_o;
  wire mux66_b10_sel_is_2_o;
  wire mux66_b11_sel_is_2_o;
  wire mux66_b12_sel_is_2_o;
  wire mux66_b13_sel_is_2_o;
  wire mux66_b15_sel_is_2_o;
  wire mux66_b3_sel_is_2_o;
  wire mux66_b4_sel_is_2_o;
  wire mux66_b9_sel_is_2_o;
  wire mux66_b9_sel_is_2_o_neg;
  wire mux67_b0_sel_is_2_o;
  wire mux67_b10_sel_is_2_o;
  wire mux67_b11_sel_is_2_o;
  wire mux67_b12_sel_is_2_o;
  wire mux67_b13_sel_is_2_o;
  wire mux67_b15_sel_is_2_o;
  wire mux67_b1_sel_is_0_o;
  wire mux67_b3_sel_is_2_o;
  wire mux67_b4_sel_is_2_o;
  wire mux67_b9_sel_is_0_o;
  wire mux68_b0_sel_is_2_o;
  wire mux68_b10_sel_is_2_o;
  wire mux68_b11_sel_is_2_o;
  wire mux68_b12_sel_is_2_o;
  wire mux68_b13_sel_is_2_o;
  wire mux68_b15_sel_is_2_o;
  wire mux68_b1_sel_is_2_o;
  wire mux68_b4_sel_is_2_o;
  wire mux68_b5_sel_is_0_o;
  wire mux68_b9_sel_is_2_o;
  wire mux69_b10_sel_is_2_o;
  wire mux69_b11_sel_is_2_o;
  wire mux69_b12_sel_is_2_o;
  wire mux69_b13_sel_is_2_o;
  wire mux69_b15_sel_is_2_o;
  wire mux69_b6_sel_is_0_o;
  wire mux69_b8_sel_is_2_o;
  wire mux69_b9_sel_is_2_o;
  wire mux6_b13_sel_is_0_o;
  wire mux6_b14_sel_is_0_o;
  wire mux6_b4_sel_is_2_o;
  wire mux70_b10_sel_is_2_o;
  wire mux70_b11_sel_is_2_o;
  wire mux70_b12_sel_is_2_o;
  wire mux70_b13_sel_is_2_o;
  wire mux70_b15_sel_is_2_o;
  wire mux70_b2_sel_is_0_o;
  wire mux70_b6_sel_is_2_o;
  wire mux70_b8_sel_is_2_o;
  wire mux70_b9_sel_is_2_o;
  wire mux71_b10_sel_is_2_o;
  wire mux71_b11_sel_is_2_o;
  wire mux71_b12_sel_is_2_o;
  wire mux71_b13_sel_is_2_o;
  wire mux71_b15_sel_is_2_o;
  wire mux71_b2_sel_is_2_o;
  wire mux71_b4_sel_is_0_o;
  wire mux71_b7_sel_is_2_o;
  wire mux71_b8_sel_is_2_o;
  wire mux71_b9_sel_is_2_o;
  wire mux72_b0_sel_is_0_o;
  wire mux72_b10_sel_is_2_o;
  wire mux72_b11_sel_is_2_o;
  wire mux72_b12_sel_is_2_o;
  wire mux72_b13_sel_is_2_o;
  wire mux72_b15_sel_is_2_o;
  wire mux72_b4_sel_is_2_o;
  wire mux72_b7_sel_is_2_o;
  wire mux72_b8_sel_is_2_o;
  wire mux72_b9_sel_is_2_o;
  wire mux73_b10_sel_is_2_o;
  wire mux73_b11_sel_is_2_o;
  wire mux73_b12_sel_is_2_o;
  wire mux73_b13_sel_is_2_o;
  wire mux73_b15_sel_is_2_o;
  wire mux73_b1_sel_is_2_o;
  wire mux73_b3_sel_is_0_o;
  wire mux73_b7_sel_is_2_o;
  wire mux73_b8_sel_is_2_o;
  wire mux73_b9_sel_is_2_o;
  wire mux74_b10_sel_is_2_o;
  wire mux74_b11_sel_is_2_o;
  wire mux74_b12_sel_is_2_o;
  wire mux74_b13_sel_is_2_o;
  wire mux74_b15_sel_is_2_o;
  wire mux74_b1_sel_is_2_o;
  wire mux74_b2_sel_is_0_o;
  wire mux74_b7_sel_is_2_o;
  wire mux74_b8_sel_is_2_o;
  wire mux74_b9_sel_is_2_o;
  wire mux75_b10_sel_is_2_o;
  wire mux75_b11_sel_is_2_o;
  wire mux75_b12_sel_is_2_o;
  wire mux75_b13_sel_is_2_o;
  wire mux75_b15_sel_is_2_o;
  wire mux75_b3_sel_is_0_o;
  wire mux75_b5_sel_is_2_o;
  wire mux75_b6_sel_is_2_o;
  wire mux75_b7_sel_is_2_o;
  wire mux75_b8_sel_is_2_o;
  wire mux75_b9_sel_is_2_o;
  wire mux76_b0_sel_is_0_o;
  wire mux76_b10_sel_is_2_o;
  wire mux76_b11_sel_is_2_o;
  wire mux76_b12_sel_is_2_o;
  wire mux76_b13_sel_is_2_o;
  wire mux76_b15_sel_is_2_o;
  wire mux76_b3_sel_is_2_o;
  wire mux76_b8_sel_is_2_o;
  wire mux76_b9_sel_is_2_o;
  wire mux77_b10_sel_is_2_o;
  wire mux77_b11_sel_is_2_o;
  wire mux77_b12_sel_is_2_o;
  wire mux77_b13_sel_is_2_o;
  wire mux77_b15_sel_is_2_o;
  wire mux77_b2_sel_is_0_o;
  wire mux77_b8_sel_is_2_o;
  wire mux77_b9_sel_is_2_o;
  wire mux78_b0_sel_is_0_o;
  wire mux78_b10_sel_is_2_o;
  wire mux78_b11_sel_is_2_o;
  wire mux78_b12_sel_is_2_o;
  wire mux78_b13_sel_is_2_o;
  wire mux78_b15_sel_is_2_o;
  wire mux78_b5_sel_is_2_o;
  wire mux78_b8_sel_is_2_o;
  wire mux78_b9_sel_is_2_o;
  wire mux79_b10_sel_is_2_o;
  wire mux79_b11_sel_is_2_o;
  wire mux79_b12_sel_is_2_o;
  wire mux79_b13_sel_is_2_o;
  wire mux79_b15_sel_is_2_o;
  wire mux79_b2_sel_is_0_o;
  wire mux79_b6_sel_is_2_o;
  wire mux79_b8_sel_is_2_o;
  wire mux79_b9_sel_is_2_o;
  wire mux7_b10_sel_is_0_o;
  wire mux7_b13_sel_is_2_o;
  wire mux7_b14_sel_is_2_o;
  wire mux7_b4_sel_is_2_o;
  wire mux7_b9_sel_is_2_o_neg;
  wire mux80_b10_sel_is_2_o;
  wire mux80_b11_sel_is_2_o;
  wire mux80_b12_sel_is_2_o;
  wire mux80_b13_sel_is_2_o;
  wire mux80_b15_sel_is_2_o;
  wire mux80_b2_sel_is_2_o;
  wire mux80_b4_sel_is_0_o;
  wire mux80_b7_sel_is_2_o;
  wire mux80_b8_sel_is_2_o;
  wire mux80_b9_sel_is_2_o;
  wire mux81_b10_sel_is_2_o;
  wire mux81_b11_sel_is_2_o;
  wire mux81_b12_sel_is_2_o;
  wire mux81_b13_sel_is_2_o;
  wire mux81_b15_sel_is_2_o;
  wire mux81_b2_sel_is_2_o;
  wire mux81_b4_sel_is_2_o;
  wire mux81_b6_sel_is_0_o;
  wire mux81_b7_sel_is_2_o;
  wire mux81_b8_sel_is_2_o;
  wire mux81_b9_sel_is_2_o;
  wire mux82_b0_sel_is_0_o;
  wire mux82_b10_sel_is_2_o;
  wire mux82_b11_sel_is_2_o;
  wire mux82_b12_sel_is_2_o;
  wire mux82_b13_sel_is_2_o;
  wire mux82_b15_sel_is_2_o;
  wire mux82_b6_sel_is_2_o;
  wire mux82_b7_sel_is_2_o;
  wire mux82_b8_sel_is_2_o;
  wire mux82_b9_sel_is_2_o;
  wire mux83_b0_sel_is_2_o;
  wire mux83_b10_sel_is_2_o;
  wire mux83_b11_sel_is_2_o;
  wire mux83_b12_sel_is_2_o;
  wire mux83_b13_sel_is_2_o;
  wire mux83_b13_sel_is_2_o_neg;
  wire mux83_b15_sel_is_2_o;
  wire mux83_b4_sel_is_0_o;
  wire mux83_b6_sel_is_2_o;
  wire mux83_b7_sel_is_2_o;
  wire mux83_b9_sel_is_2_o;
  wire mux84_b0_sel_is_2_o;
  wire mux84_b12_sel_is_2_o;
  wire mux84_b13_sel_is_0_o;
  wire mux84_b4_sel_is_2_o;
  wire mux84_b6_sel_is_2_o;
  wire mux84_b7_sel_is_2_o;
  wire mux84_b9_sel_is_2_o;
  wire mux85_b0_sel_is_2_o;
  wire mux85_b10_sel_is_0_o;
  wire mux85_b12_sel_is_2_o;
  wire mux85_b13_sel_is_2_o;
  wire mux85_b6_sel_is_2_o;
  wire mux85_b7_sel_is_2_o;
  wire mux85_b9_sel_is_2_o;
  wire mux86_b0_sel_is_2_o;
  wire mux86_b10_sel_is_2_o;
  wire mux86_b12_sel_is_2_o;
  wire mux86_b13_sel_is_2_o;
  wire mux86_b1_sel_is_0_o;
  wire mux86_b6_sel_is_2_o;
  wire mux86_b7_sel_is_2_o;
  wire mux86_b9_sel_is_2_o;
  wire mux87_b0_sel_is_2_o;
  wire mux87_b10_sel_is_2_o;
  wire mux87_b12_sel_is_2_o;
  wire mux87_b13_sel_is_2_o;
  wire mux87_b1_sel_is_2_o;
  wire mux87_b4_sel_is_0_o;
  wire mux87_b6_sel_is_2_o;
  wire mux87_b7_sel_is_2_o;
  wire mux87_b9_sel_is_2_o;
  wire mux88_b0_sel_is_2_o;
  wire mux88_b10_sel_is_2_o;
  wire mux88_b12_sel_is_2_o;
  wire mux88_b13_sel_is_2_o;
  wire mux88_b1_sel_is_2_o;
  wire mux88_b3_sel_is_0_o;
  wire mux88_b4_sel_is_2_o;
  wire mux88_b7_sel_is_2_o;
  wire mux88_b9_sel_is_2_o;
  wire mux89_b0_sel_is_2_o;
  wire mux89_b10_sel_is_2_o;
  wire mux89_b12_sel_is_2_o;
  wire mux89_b13_sel_is_2_o;
  wire mux89_b1_sel_is_2_o;
  wire mux89_b3_sel_is_2_o;
  wire mux89_b4_sel_is_2_o;
  wire mux89_b6_sel_is_0_o;
  wire mux89_b7_sel_is_2_o;
  wire mux89_b9_sel_is_2_o;
  wire mux8_b0_sel_is_0_o;
  wire mux8_b13_sel_is_2_o;
  wire mux8_b14_sel_is_2_o;
  wire mux8_b4_sel_is_2_o;
  wire mux8_b9_sel_is_0_o;
  wire mux8_b9_sel_is_0_o_neg;
  wire mux90_b10_sel_is_2_o;
  wire mux90_b12_sel_is_2_o;
  wire mux90_b13_sel_is_2_o;
  wire mux90_b2_sel_is_2_o;
  wire mux90_b4_sel_is_2_o;
  wire mux90_b5_sel_is_2_o;
  wire mux90_b7_sel_is_2_o;
  wire mux90_b9_sel_is_2_o;
  wire mux91_b10_sel_is_2_o;
  wire mux91_b12_sel_is_2_o;
  wire mux91_b13_sel_is_2_o;
  wire mux91_b2_sel_is_2_o;
  wire mux91_b3_sel_is_0_o;
  wire mux91_b4_sel_is_2_o;
  wire mux91_b5_sel_is_2_o;
  wire mux91_b7_sel_is_2_o;
  wire mux91_b9_sel_is_2_o;
  wire mux92_b0_sel_is_0_o;
  wire mux92_b10_sel_is_2_o;
  wire mux92_b12_sel_is_2_o;
  wire mux92_b13_sel_is_2_o;
  wire mux92_b13_sel_is_2_o_neg;
  wire mux92_b2_sel_is_2_o;
  wire mux92_b3_sel_is_2_o;
  wire mux92_b4_sel_is_2_o;
  wire mux92_b5_sel_is_2_o;
  wire mux92_b7_sel_is_2_o;
  wire mux92_b9_sel_is_2_o;
  wire mux93_b0_sel_is_2_o;
  wire mux93_b11_sel_is_2_o;
  wire mux93_b13_sel_is_0_o;
  wire mux93_b2_sel_is_2_o;
  wire mux93_b3_sel_is_2_o;
  wire mux93_b4_sel_is_2_o;
  wire mux93_b5_sel_is_2_o;
  wire mux93_b9_sel_is_2_o;
  wire mux94_b0_sel_is_2_o;
  wire mux94_b10_sel_is_0_o;
  wire mux94_b11_sel_is_2_o;
  wire mux94_b13_sel_is_2_o;
  wire mux94_b2_sel_is_2_o;
  wire mux94_b4_sel_is_2_o;
  wire mux94_b5_sel_is_2_o;
  wire mux94_b6_sel_is_2_o;
  wire mux94_b9_sel_is_2_o;
  wire mux94_b9_sel_is_2_o_neg;
  wire mux95_b0_sel_is_2_o;
  wire mux95_b10_sel_is_2_o;
  wire mux95_b13_sel_is_2_o;
  wire mux95_b14_sel_is_2_o;
  wire mux95_b2_sel_is_2_o;
  wire mux95_b4_sel_is_2_o;
  wire mux95_b5_sel_is_2_o;
  wire mux95_b6_sel_is_2_o;
  wire mux95_b9_sel_is_0_o;
  wire mux95_b9_sel_is_0_o_neg;
  wire mux96_b0_sel_is_2_o;
  wire mux96_b10_sel_is_2_o;
  wire mux96_b12_sel_is_0_o;
  wire mux96_b13_sel_is_2_o;
  wire mux96_b14_sel_is_2_o;
  wire mux96_b2_sel_is_2_o;
  wire mux96_b5_sel_is_2_o;
  wire mux96_b6_sel_is_2_o;
  wire mux96_b9_sel_is_0_o;
  wire mux96_b9_sel_is_0_o_neg;
  wire mux97_b12_sel_is_2_o;
  wire mux97_b13_sel_is_2_o;
  wire mux97_b14_sel_is_2_o;
  wire mux97_b15_sel_is_2_o;
  wire mux97_b2_sel_is_2_o;
  wire mux97_b5_sel_is_2_o;
  wire mux97_b6_sel_is_2_o;
  wire mux97_b7_sel_is_0_o;
  wire mux97_b9_sel_is_0_o;
  wire mux97_b9_sel_is_0_o_neg;
  wire mux98_b0_sel_is_0_o;
  wire mux98_b13_sel_is_2_o;
  wire mux98_b15_sel_is_2_o;
  wire mux98_b6_sel_is_2_o;
  wire mux98_b7_sel_is_2_o;
  wire mux98_b9_sel_is_0_o;
  wire mux98_b9_sel_is_0_o_neg;
  wire mux99_b0_sel_is_2_o;
  wire mux99_b12_sel_is_0_o;
  wire mux99_b13_sel_is_2_o;
  wire mux99_b15_sel_is_2_o;
  wire mux99_b9_sel_is_0_o;
  wire mux99_b9_sel_is_0_o_neg;
  wire mux9_b11_sel_is_0_o;
  wire mux9_b12_sel_is_2_o;
  wire mux9_b13_sel_is_2_o;
  wire mux9_b14_sel_is_2_o;
  wire mux9_b4_sel_is_2_o;
  wire mux9_b9_sel_is_0_o;
  wire n1;
  wire n10;
  wire n100;
  wire n100_neg;
  wire n101;
  wire n101_neg;
  wire n102;
  wire n102_neg;
  wire n103;
  wire n103_neg;
  wire n104;
  wire n104_neg;
  wire n105;
  wire n105_neg;
  wire n106;
  wire n106_neg;
  wire n107;
  wire n107_neg;
  wire n108;
  wire n108_neg;
  wire n109;
  wire n109_neg;
  wire n10_neg;
  wire n11;
  wire n110;
  wire n110_neg;
  wire n111;
  wire n111_neg;
  wire n112;
  wire n112_neg;
  wire n113;
  wire n113_neg;
  wire n114;
  wire n114_neg;
  wire n115;
  wire n115_neg;
  wire n116;
  wire n116_neg;
  wire n117;
  wire n117_neg;
  wire n118;
  wire n118_neg;
  wire n119;
  wire n119_neg;
  wire n11_neg;
  wire n12;
  wire n120;
  wire n120_neg;
  wire n121;
  wire n121_neg;
  wire n122;
  wire n122_neg;
  wire n123;
  wire n123_neg;
  wire n124;
  wire n124_neg;
  wire n125;
  wire n125_neg;
  wire n126;
  wire n126_neg;
  wire n127;
  wire n127_neg;
  wire n128;
  wire n128_neg;
  wire n129;
  wire n129_neg;
  wire n12_neg;
  wire n13;
  wire n130;
  wire n130_neg;
  wire n131;
  wire n131_neg;
  wire n132;
  wire n132_neg;
  wire n133;
  wire n133_neg;
  wire n134;
  wire n134_neg;
  wire n135;
  wire n135_neg;
  wire n136;
  wire n136_neg;
  wire n137;
  wire n137_neg;
  wire n138;
  wire n138_neg;
  wire n139;
  wire n139_neg;
  wire n13_neg;
  wire n14;
  wire n140;
  wire n140_neg;
  wire n141;
  wire n141_neg;
  wire n142;
  wire n142_neg;
  wire n143;
  wire n143_neg;
  wire n144;
  wire n144_neg;
  wire n145;
  wire n145_neg;
  wire n146;
  wire n146_neg;
  wire n147;
  wire n147_neg;
  wire n148;
  wire n148_neg;
  wire n149;
  wire n149_neg;
  wire n14_neg;
  wire n15;
  wire n150;
  wire n150_neg;
  wire n151;
  wire n151_neg;
  wire n152;
  wire n152_neg;
  wire n153;
  wire n153_neg;
  wire n154;
  wire n154_neg;
  wire n155;
  wire n155_neg;
  wire n156;
  wire n156_neg;
  wire n157;
  wire n157_neg;
  wire n158;
  wire n158_neg;
  wire n159;
  wire n159_neg;
  wire n15_neg;
  wire n16;
  wire n160;
  wire n160_neg;
  wire n161;
  wire n161_neg;
  wire n162;
  wire n162_neg;
  wire n163;
  wire n163_neg;
  wire n164;
  wire n164_neg;
  wire n165;
  wire n165_neg;
  wire n166;
  wire n166_neg;
  wire n167;
  wire n167_neg;
  wire n168;
  wire n168_neg;
  wire n169;
  wire n169_neg;
  wire n16_neg;
  wire n17;
  wire n170;
  wire n170_neg;
  wire n171;
  wire n171_neg;
  wire n172;
  wire n172_neg;
  wire n173;
  wire n173_neg;
  wire n174;
  wire n174_neg;
  wire n175;
  wire n175_neg;
  wire n176;
  wire n176_neg;
  wire n177;
  wire n179;
  wire n17_neg;
  wire n18;
  wire n180;
  wire n18_neg;
  wire n19;
  wire n19_neg;
  wire n1_neg;
  wire n2;
  wire n20;
  wire n20_neg;
  wire n21;
  wire n21_neg;
  wire n22;
  wire n22_neg;
  wire n23;
  wire n23_neg;
  wire n24;
  wire n24_neg;
  wire n25;
  wire n25_neg;
  wire n26;
  wire n26_neg;
  wire n27;
  wire n27_neg;
  wire n28;
  wire n28_neg;
  wire n29;
  wire n29_neg;
  wire n2_neg;
  wire n3;
  wire n30;
  wire n30_neg;
  wire n31;
  wire n31_neg;
  wire n32;
  wire n32_neg;
  wire n33;
  wire n33_neg;
  wire n34;
  wire n34_neg;
  wire n35;
  wire n356;
  wire n358;
  wire n35_neg;
  wire n36;
  wire n364;
  wire n365;
  wire n366;
  wire n36_neg;
  wire n37;
  wire n375;
  wire n376;
  wire n377;
  wire n378;
  wire n379;
  wire n37_neg;
  wire n38;
  wire n380;
  wire n381;
  wire n382;
  wire n383;
  wire n38_neg;
  wire n39;
  wire n39_neg;
  wire n3_neg;
  wire n4;
  wire n40;
  wire n40_neg;
  wire n41;
  wire n41_neg;
  wire n42;
  wire n42_neg;
  wire n43;
  wire n43_neg;
  wire n44;
  wire n44_neg;
  wire n45;
  wire n45_neg;
  wire n46;
  wire n46_neg;
  wire n47;
  wire n47_neg;
  wire n48;
  wire n48_neg;
  wire n49;
  wire n49_neg;
  wire n4_neg;
  wire n5;
  wire n50;
  wire n50_neg;
  wire n51;
  wire n51_neg;
  wire n52;
  wire n52_neg;
  wire n53;
  wire n53_neg;
  wire n54;
  wire n54_neg;
  wire n55;
  wire n55_neg;
  wire n56;
  wire n56_neg;
  wire n57;
  wire n57_neg;
  wire n58;
  wire n58_neg;
  wire n59;
  wire n59_neg;
  wire n5_neg;
  wire n6;
  wire n60;
  wire n60_neg;
  wire n61;
  wire n61_neg;
  wire n62;
  wire n62_neg;
  wire n63;
  wire n63_neg;
  wire n64;
  wire n64_neg;
  wire n65;
  wire n65_neg;
  wire n66;
  wire n66_neg;
  wire n67;
  wire n67_neg;
  wire n68;
  wire n68_neg;
  wire n69;
  wire n69_neg;
  wire n6_neg;
  wire n7;
  wire n70;
  wire n70_neg;
  wire n71;
  wire n71_neg;
  wire n72;
  wire n72_neg;
  wire n73;
  wire n73_neg;
  wire n74;
  wire n74_neg;
  wire n75;
  wire n75_neg;
  wire n76;
  wire n76_neg;
  wire n77;
  wire n77_neg;
  wire n78;
  wire n78_neg;
  wire n79;
  wire n79_neg;
  wire n7_neg;
  wire n8;
  wire n80;
  wire n80_neg;
  wire n81;
  wire n81_neg;
  wire n82;
  wire n82_neg;
  wire n83;
  wire n83_neg;
  wire n84;
  wire n84_neg;
  wire n85;
  wire n85_neg;
  wire n86;
  wire n86_neg;
  wire n87;
  wire n87_neg;
  wire n88;
  wire n88_neg;
  wire n89;
  wire n89_neg;
  wire n8_neg;
  wire n9;
  wire n90;
  wire n90_neg;
  wire n91;
  wire n91_neg;
  wire n92;
  wire n92_neg;
  wire n93;
  wire n93_neg;
  wire n94;
  wire n94_neg;
  wire n95;
  wire n95_neg;
  wire n96;
  wire n96_neg;
  wire n97;
  wire n97_neg;
  wire n98;
  wire n98_neg;
  wire n99;
  wire n99_neg;
  wire n9_neg;
  wire ready_out;  // sources/rtl/camera_init.v(45)
  wire \sel0_b0/or_B4_B5_o ;
  wire \sel0_b0/or_or_B0_B1_o_or_B2__o ;
  wire \sel0_b0/or_or_B4_B5_o_or_B6__o ;
  wire \sel0_b1/or_B0_B1_o ;
  wire \sel0_b1/or_or_B0_B1_o_or_B2__o ;
  wire \sel0_b1/or_or_B4_B5_o_or_B6__o ;
  wire \sel0_b2/or_B2_B3_o ;
  wire \sel0_b2/or_B6_or_B7_B8_o_o ;
  wire \sel0_b2/or_B7_B8_o ;
  wire \sel0_b2/or_or_B0_B1_o_or_B2__o ;
  wire \sel0_b2/or_or_B4_B5_o_or_B6__o ;
  wire \sel0_b3/or_B2_B3_o ;
  wire \sel0_b3/or_or_B0_B1_o_or_B2__o ;
  wire \sel0_b3/or_or_B4_B5_o_or_B6__o ;
  wire \sel0_b4/or_B0_B1_o ;
  wire \sel0_b4/or_B4_B5_o ;
  wire \sel0_b4/or_or_B0_B1_o_or_B2__o ;
  wire \sel0_b5/or_or_B0_B1_o_or_B2__o ;
  wire \sel0_b6/or_or_B0_B1_o_or_B2__o ;
  wire \sel0_b7/or_or_B0_B1_o_or_B2__o ;
  wire sel1_b0_sel_o;  // sources/rtl/camera_init.v(388)
  wire sel1_b1_sel_o;  // sources/rtl/camera_init.v(388)
  wire \sel2_b0/or_B6_or_B7_B8_o_o ;
  wire \sel2_b0/or_or_B4_B5_o_or_B6__o ;
  wire \sel2_b1/or_B6_or_B7_B8_o_o ;
  wire \sel2_b2/or_B6_or_B7_B8_o_o ;
  wire \sel2_b3/or_B6_or_B7_B8_o_o ;
  wire \sel2_b4/or_B6_or_B7_B8_o_o ;
  wire \sel2_b5/or_B6_or_B7_B8_o_o ;
  wire \sel2_b5/or_B7_B8_o ;
  wire \sel2_b6/or_B6_or_B7_B8_o_o ;
  wire \sel2_b6/or_B7_B8_o ;
  wire \sel2_b7/or_B6_or_B7_B8_o_o ;
  wire sel3_b0_sel_is_3_o;
  wire success_out;  // sources/rtl/camera_init.v(46)

  add_pu9_pu9_o9 add0 (
    .i0(divider2),
    .i1(9'b000000001),
    .o(n0));  // sources/rtl/camera_init.v(71)
  add_pu8_pu8_o8 add1 (
    .i0(cnt),
    .i1(8'b00000001),
    .o(n371));  // sources/rtl/camera_init.v(364)
  add_pu8_pu8_o8 add2 (
    .i0(counter),
    .i1(8'b00000001),
    .o(n372));  // sources/rtl/camera_init.v(368)
  reg_ar_as_w1 bus_write_reg (
    .clk(divider2[8]),
    .d(n366),
    .en(1'b1),
    .reset(~reset_n),
    .set(1'b0),
    .q(bus_write));  // sources/rtl/camera_init.v(389)
  eq_w8 eq0 (
    .i0(counter),
    .i1(8'b00000000),
    .o(n1));  // sources/rtl/camera_init.v(77)
  eq_w8 eq1 (
    .i0(counter),
    .i1(8'b00000001),
    .o(n2));  // sources/rtl/camera_init.v(78)
  eq_w8 eq10 (
    .i0(counter),
    .i1(8'b00001010),
    .o(n11));  // sources/rtl/camera_init.v(88)
  eq_w8 eq100 (
    .i0(counter),
    .i1(8'b01100100),
    .o(n101));  // sources/rtl/camera_init.v(178)
  eq_w8 eq101 (
    .i0(counter),
    .i1(8'b01100101),
    .o(n102));  // sources/rtl/camera_init.v(179)
  eq_w8 eq102 (
    .i0(counter),
    .i1(8'b01100110),
    .o(n103));  // sources/rtl/camera_init.v(180)
  eq_w8 eq103 (
    .i0(counter),
    .i1(8'b01100111),
    .o(n104));  // sources/rtl/camera_init.v(181)
  eq_w8 eq104 (
    .i0(counter),
    .i1(8'b01101000),
    .o(n105));  // sources/rtl/camera_init.v(182)
  eq_w8 eq105 (
    .i0(counter),
    .i1(8'b01101001),
    .o(n106));  // sources/rtl/camera_init.v(183)
  eq_w8 eq106 (
    .i0(counter),
    .i1(8'b01101010),
    .o(n107));  // sources/rtl/camera_init.v(184)
  eq_w8 eq107 (
    .i0(counter),
    .i1(8'b01101011),
    .o(n108));  // sources/rtl/camera_init.v(185)
  eq_w8 eq108 (
    .i0(counter),
    .i1(8'b01101100),
    .o(n109));  // sources/rtl/camera_init.v(186)
  eq_w8 eq109 (
    .i0(counter),
    .i1(8'b01101101),
    .o(n110));  // sources/rtl/camera_init.v(187)
  eq_w8 eq11 (
    .i0(counter),
    .i1(8'b00001011),
    .o(n12));  // sources/rtl/camera_init.v(89)
  eq_w8 eq110 (
    .i0(counter),
    .i1(8'b01101110),
    .o(n111));  // sources/rtl/camera_init.v(188)
  eq_w8 eq111 (
    .i0(counter),
    .i1(8'b01101111),
    .o(n112));  // sources/rtl/camera_init.v(189)
  eq_w8 eq112 (
    .i0(counter),
    .i1(8'b01110000),
    .o(n113));  // sources/rtl/camera_init.v(190)
  eq_w8 eq113 (
    .i0(counter),
    .i1(8'b01110001),
    .o(n114));  // sources/rtl/camera_init.v(191)
  eq_w8 eq114 (
    .i0(counter),
    .i1(8'b01110010),
    .o(n115));  // sources/rtl/camera_init.v(192)
  eq_w8 eq115 (
    .i0(counter),
    .i1(8'b01110011),
    .o(n116));  // sources/rtl/camera_init.v(193)
  eq_w8 eq116 (
    .i0(counter),
    .i1(8'b01110100),
    .o(n117));  // sources/rtl/camera_init.v(194)
  eq_w8 eq117 (
    .i0(counter),
    .i1(8'b01110101),
    .o(n118));  // sources/rtl/camera_init.v(195)
  eq_w8 eq118 (
    .i0(counter),
    .i1(8'b01110110),
    .o(n119));  // sources/rtl/camera_init.v(196)
  eq_w8 eq119 (
    .i0(counter),
    .i1(8'b01110111),
    .o(n120));  // sources/rtl/camera_init.v(197)
  eq_w8 eq12 (
    .i0(counter),
    .i1(8'b00001100),
    .o(n13));  // sources/rtl/camera_init.v(90)
  eq_w8 eq120 (
    .i0(counter),
    .i1(8'b01111000),
    .o(n121));  // sources/rtl/camera_init.v(198)
  eq_w8 eq121 (
    .i0(counter),
    .i1(8'b01111001),
    .o(n122));  // sources/rtl/camera_init.v(199)
  eq_w8 eq122 (
    .i0(counter),
    .i1(8'b01111010),
    .o(n123));  // sources/rtl/camera_init.v(200)
  eq_w8 eq123 (
    .i0(counter),
    .i1(8'b01111011),
    .o(n124));  // sources/rtl/camera_init.v(201)
  eq_w8 eq124 (
    .i0(counter),
    .i1(8'b01111100),
    .o(n125));  // sources/rtl/camera_init.v(202)
  eq_w8 eq125 (
    .i0(counter),
    .i1(8'b01111101),
    .o(n126));  // sources/rtl/camera_init.v(203)
  eq_w8 eq126 (
    .i0(counter),
    .i1(8'b01111110),
    .o(n127));  // sources/rtl/camera_init.v(204)
  eq_w8 eq127 (
    .i0(counter),
    .i1(8'b01111111),
    .o(n128));  // sources/rtl/camera_init.v(205)
  eq_w8 eq128 (
    .i0(counter),
    .i1(8'b10000000),
    .o(n129));  // sources/rtl/camera_init.v(206)
  eq_w8 eq129 (
    .i0(counter),
    .i1(8'b10000001),
    .o(n130));  // sources/rtl/camera_init.v(207)
  eq_w8 eq13 (
    .i0(counter),
    .i1(8'b00001101),
    .o(n14));  // sources/rtl/camera_init.v(91)
  eq_w8 eq130 (
    .i0(counter),
    .i1(8'b10000010),
    .o(n131));  // sources/rtl/camera_init.v(208)
  eq_w8 eq131 (
    .i0(counter),
    .i1(8'b10000011),
    .o(n132));  // sources/rtl/camera_init.v(209)
  eq_w8 eq132 (
    .i0(counter),
    .i1(8'b10000100),
    .o(n133));  // sources/rtl/camera_init.v(210)
  eq_w8 eq133 (
    .i0(counter),
    .i1(8'b10000101),
    .o(n134));  // sources/rtl/camera_init.v(211)
  eq_w8 eq134 (
    .i0(counter),
    .i1(8'b10000110),
    .o(n135));  // sources/rtl/camera_init.v(212)
  eq_w8 eq135 (
    .i0(counter),
    .i1(8'b10000111),
    .o(n136));  // sources/rtl/camera_init.v(213)
  eq_w8 eq136 (
    .i0(counter),
    .i1(8'b10001000),
    .o(n137));  // sources/rtl/camera_init.v(214)
  eq_w8 eq137 (
    .i0(counter),
    .i1(8'b10001001),
    .o(n138));  // sources/rtl/camera_init.v(215)
  eq_w8 eq138 (
    .i0(counter),
    .i1(8'b10001010),
    .o(n139));  // sources/rtl/camera_init.v(216)
  eq_w8 eq139 (
    .i0(counter),
    .i1(8'b10001011),
    .o(n140));  // sources/rtl/camera_init.v(217)
  eq_w8 eq14 (
    .i0(counter),
    .i1(8'b00001110),
    .o(n15));  // sources/rtl/camera_init.v(92)
  eq_w8 eq140 (
    .i0(counter),
    .i1(8'b10001100),
    .o(n141));  // sources/rtl/camera_init.v(218)
  eq_w8 eq141 (
    .i0(counter),
    .i1(8'b10001101),
    .o(n142));  // sources/rtl/camera_init.v(219)
  eq_w8 eq142 (
    .i0(counter),
    .i1(8'b10001110),
    .o(n143));  // sources/rtl/camera_init.v(220)
  eq_w8 eq143 (
    .i0(counter),
    .i1(8'b10001111),
    .o(n144));  // sources/rtl/camera_init.v(221)
  eq_w8 eq144 (
    .i0(counter),
    .i1(8'b10010000),
    .o(n145));  // sources/rtl/camera_init.v(222)
  eq_w8 eq145 (
    .i0(counter),
    .i1(8'b10010001),
    .o(n146));  // sources/rtl/camera_init.v(223)
  eq_w8 eq146 (
    .i0(counter),
    .i1(8'b10010010),
    .o(n147));  // sources/rtl/camera_init.v(224)
  eq_w8 eq147 (
    .i0(counter),
    .i1(8'b10010011),
    .o(n148));  // sources/rtl/camera_init.v(225)
  eq_w8 eq148 (
    .i0(counter),
    .i1(8'b10010100),
    .o(n149));  // sources/rtl/camera_init.v(226)
  eq_w8 eq149 (
    .i0(counter),
    .i1(8'b10010101),
    .o(n150));  // sources/rtl/camera_init.v(227)
  eq_w8 eq15 (
    .i0(counter),
    .i1(8'b00001111),
    .o(n16));  // sources/rtl/camera_init.v(93)
  eq_w8 eq150 (
    .i0(counter),
    .i1(8'b10010110),
    .o(n151));  // sources/rtl/camera_init.v(228)
  eq_w8 eq151 (
    .i0(counter),
    .i1(8'b10010111),
    .o(n152));  // sources/rtl/camera_init.v(229)
  eq_w8 eq152 (
    .i0(counter),
    .i1(8'b10011000),
    .o(n153));  // sources/rtl/camera_init.v(230)
  eq_w8 eq153 (
    .i0(counter),
    .i1(8'b10011001),
    .o(n154));  // sources/rtl/camera_init.v(231)
  eq_w8 eq154 (
    .i0(counter),
    .i1(8'b10011010),
    .o(n155));  // sources/rtl/camera_init.v(232)
  eq_w8 eq155 (
    .i0(counter),
    .i1(8'b10011011),
    .o(n156));  // sources/rtl/camera_init.v(233)
  eq_w8 eq156 (
    .i0(counter),
    .i1(8'b10011100),
    .o(n157));  // sources/rtl/camera_init.v(234)
  eq_w8 eq157 (
    .i0(counter),
    .i1(8'b10011101),
    .o(n158));  // sources/rtl/camera_init.v(235)
  eq_w8 eq158 (
    .i0(counter),
    .i1(8'b10011110),
    .o(n159));  // sources/rtl/camera_init.v(236)
  eq_w8 eq159 (
    .i0(counter),
    .i1(8'b10011111),
    .o(n160));  // sources/rtl/camera_init.v(237)
  eq_w8 eq16 (
    .i0(counter),
    .i1(8'b00010000),
    .o(n17));  // sources/rtl/camera_init.v(94)
  eq_w8 eq160 (
    .i0(counter),
    .i1(8'b10100000),
    .o(n161));  // sources/rtl/camera_init.v(238)
  eq_w8 eq161 (
    .i0(counter),
    .i1(8'b10100001),
    .o(n162));  // sources/rtl/camera_init.v(239)
  eq_w8 eq162 (
    .i0(counter),
    .i1(8'b10100010),
    .o(n163));  // sources/rtl/camera_init.v(240)
  eq_w8 eq163 (
    .i0(counter),
    .i1(8'b10100011),
    .o(n164));  // sources/rtl/camera_init.v(241)
  eq_w8 eq164 (
    .i0(counter),
    .i1(8'b10100100),
    .o(n165));  // sources/rtl/camera_init.v(242)
  eq_w8 eq165 (
    .i0(counter),
    .i1(8'b10100101),
    .o(n166));  // sources/rtl/camera_init.v(243)
  eq_w8 eq166 (
    .i0(counter),
    .i1(8'b10100110),
    .o(n167));  // sources/rtl/camera_init.v(244)
  eq_w8 eq167 (
    .i0(counter),
    .i1(8'b10100111),
    .o(n168));  // sources/rtl/camera_init.v(245)
  eq_w8 eq168 (
    .i0(counter),
    .i1(8'b10101000),
    .o(n169));  // sources/rtl/camera_init.v(246)
  eq_w8 eq169 (
    .i0(counter),
    .i1(8'b10101001),
    .o(n170));  // sources/rtl/camera_init.v(247)
  eq_w8 eq17 (
    .i0(counter),
    .i1(8'b00010001),
    .o(n18));  // sources/rtl/camera_init.v(95)
  eq_w8 eq170 (
    .i0(counter),
    .i1(8'b10101010),
    .o(n171));  // sources/rtl/camera_init.v(248)
  eq_w8 eq171 (
    .i0(counter),
    .i1(8'b10101011),
    .o(n172));  // sources/rtl/camera_init.v(249)
  eq_w8 eq172 (
    .i0(counter),
    .i1(8'b10101101),
    .o(n173));  // sources/rtl/camera_init.v(251)
  eq_w8 eq173 (
    .i0(counter),
    .i1(8'b10101110),
    .o(n174));  // sources/rtl/camera_init.v(252)
  eq_w8 eq174 (
    .i0(counter),
    .i1(8'b10101111),
    .o(n175));  // sources/rtl/camera_init.v(253)
  eq_w8 eq175 (
    .i0(counter),
    .i1(8'b10110000),
    .o(n176));  // sources/rtl/camera_init.v(254)
  eq_w8 eq176 (
    .i0(counter),
    .i1(8'b10110001),
    .o(n177));  // sources/rtl/camera_init.v(255)
  eq_w8 eq177 (
    .i0(state_next),
    .i1(8'b00010010),
    .o(n382));  // sources/rtl/camera_init.v(261)
  eq_w8 eq178 (
    .i0(cnt),
    .i1(8'b00000100),
    .o(n358));  // sources/rtl/camera_init.v(294)
  eq_w8 eq179 (
    .i0(state_next),
    .i1(8'b00001011),
    .o(n375));  // sources/rtl/camera_init.v(277)
  eq_w8 eq18 (
    .i0(counter),
    .i1(8'b00010010),
    .o(n19));  // sources/rtl/camera_init.v(96)
  eq_w8 eq180 (
    .i0(state_next),
    .i1(8'b00001100),
    .o(n376));  // sources/rtl/camera_init.v(278)
  eq_w8 eq181 (
    .i0(state_next),
    .i1(8'b00001101),
    .o(n377));  // sources/rtl/camera_init.v(279)
  eq_w8 eq182 (
    .i0(state_next),
    .i1(8'b00001110),
    .o(n378));  // sources/rtl/camera_init.v(280)
  eq_w8 eq183 (
    .i0(state_next),
    .i1(8'b00010001),
    .o(n381));  // sources/rtl/camera_init.v(281)
  eq_w8 eq184 (
    .i0(state_next),
    .i1(8'b00001111),
    .o(n379));  // sources/rtl/camera_init.v(286)
  eq_w8 eq185 (
    .i0(state_next),
    .i1(8'b00010000),
    .o(n380));  // sources/rtl/camera_init.v(308)
  eq_w8 eq19 (
    .i0(counter),
    .i1(8'b00010011),
    .o(n20));  // sources/rtl/camera_init.v(97)
  eq_w8 eq2 (
    .i0(counter),
    .i1(8'b00000010),
    .o(n3));  // sources/rtl/camera_init.v(80)
  eq_w8 eq20 (
    .i0(counter),
    .i1(8'b00010100),
    .o(n21));  // sources/rtl/camera_init.v(98)
  eq_w8 eq21 (
    .i0(counter),
    .i1(8'b00010101),
    .o(n22));  // sources/rtl/camera_init.v(99)
  eq_w8 eq22 (
    .i0(counter),
    .i1(8'b00010110),
    .o(n23));  // sources/rtl/camera_init.v(100)
  eq_w8 eq23 (
    .i0(counter),
    .i1(8'b00010111),
    .o(n24));  // sources/rtl/camera_init.v(101)
  eq_w8 eq24 (
    .i0(counter),
    .i1(8'b00011000),
    .o(n25));  // sources/rtl/camera_init.v(102)
  eq_w8 eq25 (
    .i0(counter),
    .i1(8'b00011001),
    .o(n26));  // sources/rtl/camera_init.v(103)
  eq_w8 eq26 (
    .i0(counter),
    .i1(8'b00011010),
    .o(n27));  // sources/rtl/camera_init.v(104)
  eq_w8 eq27 (
    .i0(counter),
    .i1(8'b00011011),
    .o(n28));  // sources/rtl/camera_init.v(105)
  eq_w8 eq28 (
    .i0(counter),
    .i1(8'b00011100),
    .o(n29));  // sources/rtl/camera_init.v(106)
  eq_w8 eq29 (
    .i0(counter),
    .i1(8'b00011101),
    .o(n30));  // sources/rtl/camera_init.v(107)
  eq_w8 eq3 (
    .i0(counter),
    .i1(8'b00000011),
    .o(n4));  // sources/rtl/camera_init.v(81)
  eq_w8 eq30 (
    .i0(counter),
    .i1(8'b00011110),
    .o(n31));  // sources/rtl/camera_init.v(108)
  eq_w8 eq31 (
    .i0(counter),
    .i1(8'b00011111),
    .o(n32));  // sources/rtl/camera_init.v(109)
  eq_w8 eq32 (
    .i0(counter),
    .i1(8'b00100000),
    .o(n33));  // sources/rtl/camera_init.v(110)
  eq_w8 eq33 (
    .i0(counter),
    .i1(8'b00100001),
    .o(n34));  // sources/rtl/camera_init.v(111)
  eq_w8 eq34 (
    .i0(counter),
    .i1(8'b00100010),
    .o(n35));  // sources/rtl/camera_init.v(112)
  eq_w8 eq35 (
    .i0(counter),
    .i1(8'b00100011),
    .o(n36));  // sources/rtl/camera_init.v(113)
  eq_w8 eq36 (
    .i0(counter),
    .i1(8'b00100100),
    .o(n37));  // sources/rtl/camera_init.v(114)
  eq_w8 eq37 (
    .i0(counter),
    .i1(8'b00100101),
    .o(n38));  // sources/rtl/camera_init.v(115)
  eq_w8 eq38 (
    .i0(counter),
    .i1(8'b00100110),
    .o(n39));  // sources/rtl/camera_init.v(116)
  eq_w8 eq39 (
    .i0(counter),
    .i1(8'b00100111),
    .o(n40));  // sources/rtl/camera_init.v(117)
  eq_w8 eq4 (
    .i0(counter),
    .i1(8'b00000100),
    .o(n5));  // sources/rtl/camera_init.v(82)
  eq_w8 eq40 (
    .i0(counter),
    .i1(8'b00101000),
    .o(n41));  // sources/rtl/camera_init.v(118)
  eq_w8 eq41 (
    .i0(counter),
    .i1(8'b00101001),
    .o(n42));  // sources/rtl/camera_init.v(119)
  eq_w8 eq42 (
    .i0(counter),
    .i1(8'b00101010),
    .o(n43));  // sources/rtl/camera_init.v(120)
  eq_w8 eq43 (
    .i0(counter),
    .i1(8'b00101011),
    .o(n44));  // sources/rtl/camera_init.v(121)
  eq_w8 eq44 (
    .i0(counter),
    .i1(8'b00101100),
    .o(n45));  // sources/rtl/camera_init.v(122)
  eq_w8 eq45 (
    .i0(counter),
    .i1(8'b00101101),
    .o(n46));  // sources/rtl/camera_init.v(123)
  eq_w8 eq46 (
    .i0(counter),
    .i1(8'b00101110),
    .o(n47));  // sources/rtl/camera_init.v(124)
  eq_w8 eq47 (
    .i0(counter),
    .i1(8'b00101111),
    .o(n48));  // sources/rtl/camera_init.v(125)
  eq_w8 eq48 (
    .i0(counter),
    .i1(8'b00110000),
    .o(n49));  // sources/rtl/camera_init.v(126)
  eq_w8 eq49 (
    .i0(counter),
    .i1(8'b00110001),
    .o(n50));  // sources/rtl/camera_init.v(127)
  eq_w8 eq5 (
    .i0(counter),
    .i1(8'b00000101),
    .o(n6));  // sources/rtl/camera_init.v(83)
  eq_w8 eq50 (
    .i0(counter),
    .i1(8'b00110010),
    .o(n51));  // sources/rtl/camera_init.v(128)
  eq_w8 eq51 (
    .i0(counter),
    .i1(8'b00110011),
    .o(n52));  // sources/rtl/camera_init.v(129)
  eq_w8 eq52 (
    .i0(counter),
    .i1(8'b00110100),
    .o(n53));  // sources/rtl/camera_init.v(130)
  eq_w8 eq53 (
    .i0(counter),
    .i1(8'b00110101),
    .o(n54));  // sources/rtl/camera_init.v(131)
  eq_w8 eq54 (
    .i0(counter),
    .i1(8'b00110110),
    .o(n55));  // sources/rtl/camera_init.v(132)
  eq_w8 eq55 (
    .i0(counter),
    .i1(8'b00110111),
    .o(n56));  // sources/rtl/camera_init.v(133)
  eq_w8 eq56 (
    .i0(counter),
    .i1(8'b00111000),
    .o(n57));  // sources/rtl/camera_init.v(134)
  eq_w8 eq57 (
    .i0(counter),
    .i1(8'b00111001),
    .o(n58));  // sources/rtl/camera_init.v(135)
  eq_w8 eq58 (
    .i0(counter),
    .i1(8'b00111010),
    .o(n59));  // sources/rtl/camera_init.v(136)
  eq_w8 eq59 (
    .i0(counter),
    .i1(8'b00111011),
    .o(n60));  // sources/rtl/camera_init.v(137)
  eq_w8 eq6 (
    .i0(counter),
    .i1(8'b00000110),
    .o(n7));  // sources/rtl/camera_init.v(84)
  eq_w8 eq60 (
    .i0(counter),
    .i1(8'b00111100),
    .o(n61));  // sources/rtl/camera_init.v(138)
  eq_w8 eq61 (
    .i0(counter),
    .i1(8'b00111101),
    .o(n62));  // sources/rtl/camera_init.v(139)
  eq_w8 eq62 (
    .i0(counter),
    .i1(8'b00111110),
    .o(n63));  // sources/rtl/camera_init.v(140)
  eq_w8 eq63 (
    .i0(counter),
    .i1(8'b00111111),
    .o(n64));  // sources/rtl/camera_init.v(141)
  eq_w8 eq64 (
    .i0(counter),
    .i1(8'b01000000),
    .o(n65));  // sources/rtl/camera_init.v(142)
  eq_w8 eq65 (
    .i0(counter),
    .i1(8'b01000001),
    .o(n66));  // sources/rtl/camera_init.v(143)
  eq_w8 eq66 (
    .i0(counter),
    .i1(8'b01000010),
    .o(n67));  // sources/rtl/camera_init.v(144)
  eq_w8 eq67 (
    .i0(counter),
    .i1(8'b01000011),
    .o(n68));  // sources/rtl/camera_init.v(145)
  eq_w8 eq68 (
    .i0(counter),
    .i1(8'b01000100),
    .o(n69));  // sources/rtl/camera_init.v(146)
  eq_w8 eq69 (
    .i0(counter),
    .i1(8'b01000101),
    .o(n70));  // sources/rtl/camera_init.v(147)
  eq_w8 eq7 (
    .i0(counter),
    .i1(8'b00000111),
    .o(n8));  // sources/rtl/camera_init.v(85)
  eq_w8 eq70 (
    .i0(counter),
    .i1(8'b01000110),
    .o(n71));  // sources/rtl/camera_init.v(148)
  eq_w8 eq71 (
    .i0(counter),
    .i1(8'b01000111),
    .o(n72));  // sources/rtl/camera_init.v(149)
  eq_w8 eq72 (
    .i0(counter),
    .i1(8'b01001000),
    .o(n73));  // sources/rtl/camera_init.v(150)
  eq_w8 eq73 (
    .i0(counter),
    .i1(8'b01001001),
    .o(n74));  // sources/rtl/camera_init.v(151)
  eq_w8 eq74 (
    .i0(counter),
    .i1(8'b01001010),
    .o(n75));  // sources/rtl/camera_init.v(152)
  eq_w8 eq75 (
    .i0(counter),
    .i1(8'b01001011),
    .o(n76));  // sources/rtl/camera_init.v(153)
  eq_w8 eq76 (
    .i0(counter),
    .i1(8'b01001100),
    .o(n77));  // sources/rtl/camera_init.v(154)
  eq_w8 eq77 (
    .i0(counter),
    .i1(8'b01001101),
    .o(n78));  // sources/rtl/camera_init.v(155)
  eq_w8 eq78 (
    .i0(counter),
    .i1(8'b01001110),
    .o(n79));  // sources/rtl/camera_init.v(156)
  eq_w8 eq79 (
    .i0(counter),
    .i1(8'b01001111),
    .o(n80));  // sources/rtl/camera_init.v(157)
  eq_w8 eq8 (
    .i0(counter),
    .i1(8'b00001000),
    .o(n9));  // sources/rtl/camera_init.v(86)
  eq_w8 eq80 (
    .i0(counter),
    .i1(8'b01010000),
    .o(n81));  // sources/rtl/camera_init.v(158)
  eq_w8 eq81 (
    .i0(counter),
    .i1(8'b01010001),
    .o(n82));  // sources/rtl/camera_init.v(159)
  eq_w8 eq82 (
    .i0(counter),
    .i1(8'b01010010),
    .o(n83));  // sources/rtl/camera_init.v(160)
  eq_w8 eq83 (
    .i0(counter),
    .i1(8'b01010011),
    .o(n84));  // sources/rtl/camera_init.v(161)
  eq_w8 eq84 (
    .i0(counter),
    .i1(8'b01010100),
    .o(n85));  // sources/rtl/camera_init.v(162)
  eq_w8 eq85 (
    .i0(counter),
    .i1(8'b01010101),
    .o(n86));  // sources/rtl/camera_init.v(163)
  eq_w8 eq86 (
    .i0(counter),
    .i1(8'b01010110),
    .o(n87));  // sources/rtl/camera_init.v(164)
  eq_w8 eq87 (
    .i0(counter),
    .i1(8'b01010111),
    .o(n88));  // sources/rtl/camera_init.v(165)
  eq_w8 eq88 (
    .i0(counter),
    .i1(8'b01011000),
    .o(n89));  // sources/rtl/camera_init.v(166)
  eq_w8 eq89 (
    .i0(counter),
    .i1(8'b01011001),
    .o(n90));  // sources/rtl/camera_init.v(167)
  eq_w8 eq9 (
    .i0(counter),
    .i1(8'b00001001),
    .o(n10));  // sources/rtl/camera_init.v(87)
  eq_w8 eq90 (
    .i0(counter),
    .i1(8'b01011010),
    .o(n91));  // sources/rtl/camera_init.v(168)
  eq_w8 eq91 (
    .i0(counter),
    .i1(8'b01011011),
    .o(n92));  // sources/rtl/camera_init.v(169)
  eq_w8 eq92 (
    .i0(counter),
    .i1(8'b01011100),
    .o(n93));  // sources/rtl/camera_init.v(170)
  eq_w8 eq93 (
    .i0(counter),
    .i1(8'b01011101),
    .o(n94));  // sources/rtl/camera_init.v(171)
  eq_w8 eq94 (
    .i0(counter),
    .i1(8'b01011110),
    .o(n95));  // sources/rtl/camera_init.v(172)
  eq_w8 eq95 (
    .i0(counter),
    .i1(8'b01011111),
    .o(n96));  // sources/rtl/camera_init.v(173)
  eq_w8 eq96 (
    .i0(counter),
    .i1(8'b01100000),
    .o(n97));  // sources/rtl/camera_init.v(174)
  eq_w8 eq97 (
    .i0(counter),
    .i1(8'b01100001),
    .o(n98));  // sources/rtl/camera_init.v(175)
  eq_w8 eq98 (
    .i0(counter),
    .i1(8'b01100010),
    .o(n99));  // sources/rtl/camera_init.v(176)
  eq_w8 eq99 (
    .i0(counter),
    .i1(8'b01100011),
    .o(n100));  // sources/rtl/camera_init.v(177)
  binary_mux_s1_w1 mux0_b0 (
    .i0(n178[2]),
    .i1(1'b1),
    .sel(n176),
    .o(n181[0]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux0_b10 (
    .i0(n177),
    .i1(1'b1),
    .sel(n176),
    .o(n181[10]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux0_b11 (
    .i0(1'b0),
    .i1(1'b1),
    .sel(n176),
    .o(n181[11]));  // sources/rtl/camera_init.v(256)
  AL_MUX mux100_b10 (
    .i0(1'b1),
    .i1(n279[10]),
    .sel(mux100_b10_sel_is_0_o),
    .o(n281[10]));
  and mux100_b10_sel_is_0 (mux100_b10_sel_is_0_o, n76_neg, n77_neg);
  binary_mux_s1_w1 mux100_b11 (
    .i0(n280[11]),
    .i1(1'b1),
    .sel(n76),
    .o(n281[11]));  // sources/rtl/camera_init.v(256)
  and mux100_b12_sel_is_2 (mux100_b12_sel_is_2_o, n76_neg, mux99_b12_sel_is_0_o);
  and mux100_b13_sel_is_2 (mux100_b13_sel_is_2_o, n76_neg, mux99_b13_sel_is_2_o);
  AL_MUX mux100_b3 (
    .i0(1'b0),
    .i1(n279[3]),
    .sel(mux100_b10_sel_is_0_o),
    .o(n281[3]));
  binary_mux_s1_w1 mux100_b4 (
    .i0(n280[4]),
    .i1(1'b0),
    .sel(n76),
    .o(n281[4]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux100_b8 (
    .i0(n280[8]),
    .i1(1'b0),
    .sel(n76),
    .o(n281[8]));  // sources/rtl/camera_init.v(256)
  and mux100_b9_sel_is_0 (mux100_b9_sel_is_0_o, n76_neg, mux99_b9_sel_is_0_o_neg);
  not mux100_b9_sel_is_0_o_inv (mux100_b9_sel_is_0_o_neg, mux100_b9_sel_is_0_o);
  and mux101_b0_sel_is_0 (mux101_b0_sel_is_0_o, n75_neg, n76_neg);
  and mux101_b12_sel_is_2 (mux101_b12_sel_is_2_o, n75_neg, mux100_b12_sel_is_2_o);
  and mux101_b13_sel_is_2 (mux101_b13_sel_is_2_o, n75_neg, mux100_b13_sel_is_2_o);
  and mux101_b1_sel_is_2 (mux101_b1_sel_is_2_o, n75_neg, mux100_b10_sel_is_0_o);
  binary_mux_s1_w1 mux101_b3 (
    .i0(n281[3]),
    .i1(1'b1),
    .sel(n75),
    .o(n282[3]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux101_b4 (
    .i0(n281[4]),
    .i1(1'b1),
    .sel(n75),
    .o(n282[4]));  // sources/rtl/camera_init.v(256)
  AL_MUX mux101_b5 (
    .i0(1'b0),
    .i1(n279[5]),
    .sel(mux101_b1_sel_is_2_o),
    .o(n282[5]));
  binary_mux_s1_w1 mux101_b8 (
    .i0(n281[8]),
    .i1(1'b1),
    .sel(n75),
    .o(n282[8]));  // sources/rtl/camera_init.v(256)
  and mux101_b9_sel_is_0 (mux101_b9_sel_is_0_o, n75_neg, mux100_b9_sel_is_0_o_neg);
  and mux102_b0_sel_is_2 (mux102_b0_sel_is_2_o, n74_neg, mux101_b0_sel_is_0_o);
  and mux102_b10_sel_is_0 (mux102_b10_sel_is_0_o, n74_neg, n75_neg);
  AL_MUX mux102_b12 (
    .i0(1'b0),
    .i1(n278[12]),
    .sel(mux102_b12_sel_is_2_o),
    .o(n283[12]));
  and mux102_b12_sel_is_2 (mux102_b12_sel_is_2_o, n74_neg, mux101_b12_sel_is_2_o);
  and mux102_b13_sel_is_2 (mux102_b13_sel_is_2_o, n74_neg, mux101_b13_sel_is_2_o);
  not mux102_b13_sel_is_2_o_inv (mux102_b13_sel_is_2_o_neg, mux102_b13_sel_is_2_o);
  AL_MUX mux102_b14 (
    .i0(1'b1),
    .i1(n280[14]),
    .sel(mux102_b0_sel_is_2_o),
    .o(n283[14]));
  and mux102_b1_sel_is_2 (mux102_b1_sel_is_2_o, n74_neg, mux101_b1_sel_is_2_o);
  AL_MUX mux102_b7 (
    .i0(1'b0),
    .i1(n280[7]),
    .sel(mux102_b0_sel_is_2_o),
    .o(n283[7]));
  binary_mux_s1_w1 mux102_b8 (
    .i0(n282[8]),
    .i1(1'b0),
    .sel(n74),
    .o(n283[8]));  // sources/rtl/camera_init.v(256)
  and mux102_b9_sel_is_2 (mux102_b9_sel_is_2_o, n74_neg, mux101_b9_sel_is_0_o);
  AL_MUX mux103_b0 (
    .i0(1'b0),
    .i1(n280[0]),
    .sel(mux103_b0_sel_is_2_o),
    .o(n284[0]));
  and mux103_b0_sel_is_2 (mux103_b0_sel_is_2_o, n73_neg, mux102_b0_sel_is_2_o);
  AL_MUX mux103_b1 (
    .i0(1'b0),
    .i1(n279[1]),
    .sel(mux103_b1_sel_is_2_o),
    .o(n284[1]));
  AL_MUX mux103_b10 (
    .i0(1'b0),
    .i1(n281[10]),
    .sel(mux103_b10_sel_is_2_o),
    .o(n284[10]));
  and mux103_b10_sel_is_2 (mux103_b10_sel_is_2_o, n73_neg, mux102_b10_sel_is_0_o);
  and mux103_b13_sel_is_0 (mux103_b13_sel_is_0_o, n73_neg, mux102_b13_sel_is_2_o_neg);
  binary_mux_s1_w1 mux103_b14 (
    .i0(n283[14]),
    .i1(1'b0),
    .sel(n73),
    .o(n284[14]));  // sources/rtl/camera_init.v(256)
  and mux103_b1_sel_is_2 (mux103_b1_sel_is_2_o, n73_neg, mux102_b1_sel_is_2_o);
  AL_MUX mux103_b2 (
    .i0(1'b0),
    .i1(n280[2]),
    .sel(mux103_b0_sel_is_2_o),
    .o(n284[2]));
  AL_MUX mux103_b3 (
    .i0(1'b0),
    .i1(n282[3]),
    .sel(mux103_b3_sel_is_0_o),
    .o(n284[3]));
  and mux103_b3_sel_is_0 (mux103_b3_sel_is_0_o, n73_neg, n74_neg);
  AL_MUX mux103_b4 (
    .i0(1'b0),
    .i1(n282[4]),
    .sel(mux103_b3_sel_is_0_o),
    .o(n284[4]));
  AL_MUX mux103_b6 (
    .i0(1'b0),
    .i1(n280[6]),
    .sel(mux103_b0_sel_is_2_o),
    .o(n284[6]));
  binary_mux_s1_w1 mux103_b8 (
    .i0(n283[8]),
    .i1(1'b1),
    .sel(n73),
    .o(n284[8]));  // sources/rtl/camera_init.v(256)
  and mux103_b9_sel_is_2 (mux103_b9_sel_is_2_o, n73_neg, mux102_b9_sel_is_2_o);
  binary_mux_s1_w1 mux104_b0 (
    .i0(n284[0]),
    .i1(1'b1),
    .sel(n72),
    .o(n285[0]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux104_b1 (
    .i0(n284[1]),
    .i1(1'b1),
    .sel(n72),
    .o(n285[1]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux104_b10 (
    .i0(n284[10]),
    .i1(1'b1),
    .sel(n72),
    .o(n285[10]));  // sources/rtl/camera_init.v(256)
  and mux104_b11_sel_is_2 (mux104_b11_sel_is_2_o, n72_neg, mux103_b10_sel_is_2_o);
  AL_MUX mux104_b12 (
    .i0(1'b1),
    .i1(n283[12]),
    .sel(mux104_b12_sel_is_0_o),
    .o(n285[12]));
  and mux104_b12_sel_is_0 (mux104_b12_sel_is_0_o, n72_neg, n73_neg);
  and mux104_b13_sel_is_2 (mux104_b13_sel_is_2_o, n72_neg, mux103_b13_sel_is_0_o);
  AL_MUX mux104_b15 (
    .i0(1'b0),
    .i1(n280[15]),
    .sel(mux104_b15_sel_is_2_o),
    .o(n285[15]));
  and mux104_b15_sel_is_2 (mux104_b15_sel_is_2_o, n72_neg, mux103_b0_sel_is_2_o);
  binary_mux_s1_w1 mux104_b3 (
    .i0(n284[3]),
    .i1(1'b1),
    .sel(n72),
    .o(n285[3]));  // sources/rtl/camera_init.v(256)
  AL_MUX mux104_b5 (
    .i0(1'b1),
    .i1(n282[5]),
    .sel(mux104_b5_sel_is_2_o),
    .o(n285[5]));
  and mux104_b5_sel_is_2 (mux104_b5_sel_is_2_o, n72_neg, mux103_b3_sel_is_0_o);
  binary_mux_s1_w1 mux104_b6 (
    .i0(n284[6]),
    .i1(1'b1),
    .sel(n72),
    .o(n285[6]));  // sources/rtl/camera_init.v(256)
  AL_MUX mux104_b7 (
    .i0(1'b1),
    .i1(n283[7]),
    .sel(mux104_b12_sel_is_0_o),
    .o(n285[7]));
  and mux104_b9_sel_is_2 (mux104_b9_sel_is_2_o, n72_neg, mux103_b9_sel_is_2_o);
  not mux104_b9_sel_is_2_o_inv (mux104_b9_sel_is_2_o_neg, mux104_b9_sel_is_2_o);
  and mux105_b11_sel_is_2 (mux105_b11_sel_is_2_o, n71_neg, mux104_b11_sel_is_2_o);
  and mux105_b13_sel_is_2 (mux105_b13_sel_is_2_o, n71_neg, mux104_b13_sel_is_2_o);
  not mux105_b13_sel_is_2_o_inv (mux105_b13_sel_is_2_o_neg, mux105_b13_sel_is_2_o);
  and mux105_b14_sel_is_0 (mux105_b14_sel_is_0_o, n71_neg, n72_neg);
  binary_mux_s1_w1 mux105_b15 (
    .i0(n285[15]),
    .i1(1'b1),
    .sel(n71),
    .o(n286[15]));  // sources/rtl/camera_init.v(256)
  AL_MUX mux105_b4 (
    .i0(1'b1),
    .i1(n284[4]),
    .sel(mux105_b14_sel_is_0_o),
    .o(n286[4]));
  binary_mux_s1_w1 mux105_b5 (
    .i0(n285[5]),
    .i1(1'b0),
    .sel(n71),
    .o(n286[5]));  // sources/rtl/camera_init.v(256)
  AL_MUX mux105_b8 (
    .i0(1'b0),
    .i1(n284[8]),
    .sel(mux105_b14_sel_is_0_o),
    .o(n286[8]));
  and mux105_b9_sel_is_0 (mux105_b9_sel_is_0_o, n71_neg, mux104_b9_sel_is_2_o_neg);
  and mux106_b0_sel_is_0 (mux106_b0_sel_is_0_o, n70_neg, n71_neg);
  AL_MUX mux106_b11 (
    .i0(1'b0),
    .i1(n281[11]),
    .sel(mux106_b11_sel_is_2_o),
    .o(n287[11]));
  and mux106_b11_sel_is_2 (mux106_b11_sel_is_2_o, n70_neg, mux105_b11_sel_is_2_o);
  AL_MUX mux106_b12 (
    .i0(1'b0),
    .i1(n285[12]),
    .sel(mux106_b0_sel_is_0_o),
    .o(n287[12]));
  and mux106_b13_sel_is_0 (mux106_b13_sel_is_0_o, n70_neg, mux105_b13_sel_is_2_o_neg);
  not mux106_b13_sel_is_0_o_inv (mux106_b13_sel_is_0_o_neg, mux106_b13_sel_is_0_o);
  and mux106_b14_sel_is_2 (mux106_b14_sel_is_2_o, n70_neg, mux105_b14_sel_is_0_o);
  binary_mux_s1_w1 mux106_b15 (
    .i0(n286[15]),
    .i1(1'b0),
    .sel(n70),
    .o(n287[15]));  // sources/rtl/camera_init.v(256)
  AL_MUX mux106_b2 (
    .i0(1'b1),
    .i1(n284[2]),
    .sel(mux106_b14_sel_is_2_o),
    .o(n287[2]));
  binary_mux_s1_w1 mux106_b5 (
    .i0(n286[5]),
    .i1(1'b1),
    .sel(n70),
    .o(n287[5]));  // sources/rtl/camera_init.v(256)
  AL_MUX mux106_b6 (
    .i0(1'b0),
    .i1(n285[6]),
    .sel(mux106_b0_sel_is_0_o),
    .o(n287[6]));
  AL_MUX mux106_b7 (
    .i0(1'b0),
    .i1(n285[7]),
    .sel(mux106_b0_sel_is_0_o),
    .o(n287[7]));
  and mux106_b9_sel_is_2 (mux106_b9_sel_is_2_o, n70_neg, mux105_b9_sel_is_0_o);
  AL_MUX mux107_b0 (
    .i0(1'b0),
    .i1(n285[0]),
    .sel(mux107_b0_sel_is_2_o),
    .o(n288[0]));
  and mux107_b0_sel_is_2 (mux107_b0_sel_is_2_o, n69_neg, mux106_b0_sel_is_0_o);
  AL_MUX mux107_b1 (
    .i0(1'b0),
    .i1(n285[1]),
    .sel(mux107_b0_sel_is_2_o),
    .o(n288[1]));
  AL_MUX mux107_b10 (
    .i0(1'b0),
    .i1(n285[10]),
    .sel(mux107_b0_sel_is_2_o),
    .o(n288[10]));
  binary_mux_s1_w1 mux107_b11 (
    .i0(n287[11]),
    .i1(1'b1),
    .sel(n69),
    .o(n288[11]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux107_b12 (
    .i0(n287[12]),
    .i1(1'b1),
    .sel(n69),
    .o(n288[12]));  // sources/rtl/camera_init.v(256)
  and mux107_b13_sel_is_0 (mux107_b13_sel_is_0_o, n69_neg, mux106_b13_sel_is_0_o_neg);
  and mux107_b14_sel_is_2 (mux107_b14_sel_is_2_o, n69_neg, mux106_b14_sel_is_2_o);
  binary_mux_s1_w1 mux107_b2 (
    .i0(n287[2]),
    .i1(1'b0),
    .sel(n69),
    .o(n288[2]));  // sources/rtl/camera_init.v(256)
  AL_MUX mux107_b3 (
    .i0(1'b0),
    .i1(n285[3]),
    .sel(mux107_b0_sel_is_2_o),
    .o(n288[3]));
  AL_MUX mux107_b4 (
    .i0(1'b0),
    .i1(n286[4]),
    .sel(mux107_b4_sel_is_0_o),
    .o(n288[4]));
  and mux107_b4_sel_is_0 (mux107_b4_sel_is_0_o, n69_neg, n70_neg);
  binary_mux_s1_w1 mux107_b5 (
    .i0(n287[5]),
    .i1(1'b0),
    .sel(n69),
    .o(n288[5]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux107_b7 (
    .i0(n287[7]),
    .i1(1'b1),
    .sel(n69),
    .o(n288[7]));  // sources/rtl/camera_init.v(256)
  and mux107_b9_sel_is_2 (mux107_b9_sel_is_2_o, n69_neg, mux106_b9_sel_is_2_o);
  binary_mux_s1_w1 mux108_b0 (
    .i0(n288[0]),
    .i1(1'b1),
    .sel(n68),
    .o(n289[0]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux108_b1 (
    .i0(n288[1]),
    .i1(1'b1),
    .sel(n68),
    .o(n289[1]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux108_b11 (
    .i0(n288[11]),
    .i1(1'b0),
    .sel(n68),
    .o(n289[11]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux108_b12 (
    .i0(n288[12]),
    .i1(1'b0),
    .sel(n68),
    .o(n289[12]));  // sources/rtl/camera_init.v(256)
  and mux108_b13_sel_is_2 (mux108_b13_sel_is_2_o, n68_neg, mux107_b13_sel_is_0_o);
  and mux108_b14_sel_is_2 (mux108_b14_sel_is_2_o, n68_neg, mux107_b14_sel_is_2_o);
  and mux108_b15_sel_is_0 (mux108_b15_sel_is_0_o, n68_neg, n69_neg);
  binary_mux_s1_w1 mux108_b2 (
    .i0(n288[2]),
    .i1(1'b1),
    .sel(n68),
    .o(n289[2]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux108_b3 (
    .i0(n288[3]),
    .i1(1'b1),
    .sel(n68),
    .o(n289[3]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux108_b4 (
    .i0(n288[4]),
    .i1(1'b1),
    .sel(n68),
    .o(n289[4]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux108_b5 (
    .i0(n288[5]),
    .i1(1'b1),
    .sel(n68),
    .o(n289[5]));  // sources/rtl/camera_init.v(256)
  AL_MUX mux108_b6 (
    .i0(1'b1),
    .i1(n287[6]),
    .sel(mux108_b15_sel_is_0_o),
    .o(n289[6]));
  and mux108_b8_sel_is_2 (mux108_b8_sel_is_2_o, n68_neg, mux107_b4_sel_is_0_o);
  and mux108_b9_sel_is_2 (mux108_b9_sel_is_2_o, n68_neg, mux107_b9_sel_is_2_o);
  not mux108_b9_sel_is_2_o_inv (mux108_b9_sel_is_2_o_neg, mux108_b9_sel_is_2_o);
  and mux109_b10_sel_is_0 (mux109_b10_sel_is_0_o, n67_neg, n68_neg);
  and mux109_b13_sel_is_2 (mux109_b13_sel_is_2_o, n67_neg, mux108_b13_sel_is_2_o);
  AL_MUX mux109_b14 (
    .i0(1'b1),
    .i1(n284[14]),
    .sel(mux109_b14_sel_is_2_o),
    .o(n290[14]));
  and mux109_b14_sel_is_2 (mux109_b14_sel_is_2_o, n67_neg, mux108_b14_sel_is_2_o);
  AL_MUX mux109_b15 (
    .i0(1'b1),
    .i1(n287[15]),
    .sel(mux109_b15_sel_is_2_o),
    .o(n290[15]));
  and mux109_b15_sel_is_2 (mux109_b15_sel_is_2_o, n67_neg, mux108_b15_sel_is_0_o);
  binary_mux_s1_w1 mux109_b3 (
    .i0(n289[3]),
    .i1(1'b0),
    .sel(n67),
    .o(n290[3]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux109_b4 (
    .i0(n289[4]),
    .i1(1'b0),
    .sel(n67),
    .o(n290[4]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux109_b5 (
    .i0(n289[5]),
    .i1(1'b0),
    .sel(n67),
    .o(n290[5]));  // sources/rtl/camera_init.v(256)
  and mux109_b8_sel_is_2 (mux109_b8_sel_is_2_o, n67_neg, mux108_b8_sel_is_2_o);
  and mux109_b9_sel_is_0 (mux109_b9_sel_is_0_o, n67_neg, mux108_b9_sel_is_2_o_neg);
  not mux109_b9_sel_is_0_o_inv (mux109_b9_sel_is_0_o_neg, mux109_b9_sel_is_0_o);
  binary_mux_s1_w1 mux10_b1 (
    .i0(n190[1]),
    .i1(1'b1),
    .sel(n166),
    .o(n191[1]));  // sources/rtl/camera_init.v(256)
  AL_MUX mux10_b10 (
    .i0(1'b0),
    .i1(n189[10]),
    .sel(mux10_b10_sel_is_0_o),
    .o(n191[10]));
  and mux10_b10_sel_is_0 (mux10_b10_sel_is_0_o, n166_neg, n167_neg);
  AL_MUX mux10_b11 (
    .i0(1'b1),
    .i1(n188[11]),
    .sel(mux10_b11_sel_is_2_o),
    .o(n191[11]));
  and mux10_b11_sel_is_2 (mux10_b11_sel_is_2_o, n166_neg, mux9_b11_sel_is_0_o);
  and mux10_b12_sel_is_2 (mux10_b12_sel_is_2_o, n166_neg, mux9_b12_sel_is_2_o);
  and mux10_b13_sel_is_2 (mux10_b13_sel_is_2_o, n166_neg, mux9_b13_sel_is_2_o);
  and mux10_b14_sel_is_2 (mux10_b14_sel_is_2_o, n166_neg, mux9_b14_sel_is_2_o);
  binary_mux_s1_w1 mux10_b4 (
    .i0(n190[4]),
    .i1(1'b1),
    .sel(n166),
    .o(n191[4]));  // sources/rtl/camera_init.v(256)
  AL_MUX mux10_b5 (
    .i0(1'b1),
    .i1(n189[5]),
    .sel(mux10_b10_sel_is_0_o),
    .o(n191[5]));
  binary_mux_s1_w1 mux10_b8 (
    .i0(n190[8]),
    .i1(1'b0),
    .sel(n166),
    .o(n191[8]));  // sources/rtl/camera_init.v(256)
  and mux10_b9_sel_is_2 (mux10_b9_sel_is_2_o, n166_neg, mux9_b9_sel_is_0_o);
  not mux10_b9_sel_is_2_o_inv (mux10_b9_sel_is_2_o_neg, mux10_b9_sel_is_2_o);
  and mux110_b0_sel_is_0 (mux110_b0_sel_is_0_o, n66_neg, n67_neg);
  and mux110_b10_sel_is_2 (mux110_b10_sel_is_2_o, n66_neg, mux109_b10_sel_is_0_o);
  AL_MUX mux110_b12 (
    .i0(1'b1),
    .i1(n289[12]),
    .sel(mux110_b0_sel_is_0_o),
    .o(n291[12]));
  and mux110_b13_sel_is_2 (mux110_b13_sel_is_2_o, n66_neg, mux109_b13_sel_is_2_o);
  binary_mux_s1_w1 mux110_b14 (
    .i0(n290[14]),
    .i1(1'b0),
    .sel(n66),
    .o(n291[14]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux110_b3 (
    .i0(n290[3]),
    .i1(1'b1),
    .sel(n66),
    .o(n291[3]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux110_b4 (
    .i0(n290[4]),
    .i1(1'b1),
    .sel(n66),
    .o(n291[4]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux110_b5 (
    .i0(n290[5]),
    .i1(1'b1),
    .sel(n66),
    .o(n291[5]));  // sources/rtl/camera_init.v(256)
  and mux110_b8_sel_is_2 (mux110_b8_sel_is_2_o, n66_neg, mux109_b8_sel_is_2_o);
  and mux110_b9_sel_is_0 (mux110_b9_sel_is_0_o, n66_neg, mux109_b9_sel_is_0_o_neg);
  AL_MUX mux111_b0 (
    .i0(1'b0),
    .i1(n289[0]),
    .sel(mux111_b0_sel_is_2_o),
    .o(n292[0]));
  and mux111_b0_sel_is_2 (mux111_b0_sel_is_2_o, n65_neg, mux110_b0_sel_is_0_o);
  AL_MUX mux111_b1 (
    .i0(1'b0),
    .i1(n289[1]),
    .sel(mux111_b0_sel_is_2_o),
    .o(n292[1]));
  AL_MUX mux111_b10 (
    .i0(1'b1),
    .i1(n288[10]),
    .sel(mux111_b10_sel_is_2_o),
    .o(n292[10]));
  and mux111_b10_sel_is_2 (mux111_b10_sel_is_2_o, n65_neg, mux110_b10_sel_is_2_o);
  binary_mux_s1_w1 mux111_b12 (
    .i0(n291[12]),
    .i1(1'b0),
    .sel(n65),
    .o(n292[12]));  // sources/rtl/camera_init.v(256)
  and mux111_b13_sel_is_2 (mux111_b13_sel_is_2_o, n65_neg, mux110_b13_sel_is_2_o);
  not mux111_b13_sel_is_2_o_inv (mux111_b13_sel_is_2_o_neg, mux111_b13_sel_is_2_o);
  and mux111_b15_sel_is_0 (mux111_b15_sel_is_0_o, n65_neg, n66_neg);
  binary_mux_s1_w1 mux111_b5 (
    .i0(n291[5]),
    .i1(1'b0),
    .sel(n65),
    .o(n292[5]));  // sources/rtl/camera_init.v(256)
  AL_MUX mux111_b8 (
    .i0(1'b1),
    .i1(n286[8]),
    .sel(mux111_b8_sel_is_2_o),
    .o(n292[8]));
  and mux111_b8_sel_is_2 (mux111_b8_sel_is_2_o, n65_neg, mux110_b8_sel_is_2_o);
  and mux111_b9_sel_is_2 (mux111_b9_sel_is_2_o, n65_neg, mux110_b9_sel_is_0_o);
  not mux111_b9_sel_is_2_o_inv (mux111_b9_sel_is_2_o_neg, mux111_b9_sel_is_2_o);
  binary_mux_s1_w1 mux112_b0 (
    .i0(n292[0]),
    .i1(1'b1),
    .sel(n64),
    .o(n293[0]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux112_b1 (
    .i0(n292[1]),
    .i1(1'b1),
    .sel(n64),
    .o(n293[1]));  // sources/rtl/camera_init.v(256)
  AL_MUX mux112_b11 (
    .i0(1'b1),
    .i1(n289[11]),
    .sel(mux112_b11_sel_is_2_o),
    .o(n293[11]));
  and mux112_b11_sel_is_2 (mux112_b11_sel_is_2_o, n64_neg, mux111_b0_sel_is_2_o);
  and mux112_b13_sel_is_0 (mux112_b13_sel_is_0_o, n64_neg, mux111_b13_sel_is_2_o_neg);
  and mux112_b14_sel_is_0 (mux112_b14_sel_is_0_o, n64_neg, n65_neg);
  and mux112_b15_sel_is_2 (mux112_b15_sel_is_2_o, n64_neg, mux111_b15_sel_is_0_o);
  AL_MUX mux112_b3 (
    .i0(1'b0),
    .i1(n291[3]),
    .sel(mux112_b14_sel_is_0_o),
    .o(n293[3]));
  AL_MUX mux112_b7 (
    .i0(1'b0),
    .i1(n288[7]),
    .sel(mux112_b7_sel_is_2_o),
    .o(n293[7]));
  and mux112_b7_sel_is_2 (mux112_b7_sel_is_2_o, n64_neg, mux111_b10_sel_is_2_o);
  and mux112_b9_sel_is_0 (mux112_b9_sel_is_0_o, n64_neg, mux111_b9_sel_is_2_o_neg);
  not mux112_b9_sel_is_0_o_inv (mux112_b9_sel_is_0_o_neg, mux112_b9_sel_is_0_o);
  binary_mux_s1_w1 mux113_b1 (
    .i0(n293[1]),
    .i1(1'b0),
    .sel(n63),
    .o(n294[1]));  // sources/rtl/camera_init.v(256)
  AL_MUX mux113_b10 (
    .i0(1'b0),
    .i1(n292[10]),
    .sel(mux113_b10_sel_is_0_o),
    .o(n294[10]));
  and mux113_b10_sel_is_0 (mux113_b10_sel_is_0_o, n63_neg, n64_neg);
  binary_mux_s1_w1 mux113_b11 (
    .i0(n293[11]),
    .i1(1'b0),
    .sel(n63),
    .o(n294[11]));  // sources/rtl/camera_init.v(256)
  AL_MUX mux113_b12 (
    .i0(1'b1),
    .i1(n292[12]),
    .sel(mux113_b10_sel_is_0_o),
    .o(n294[12]));
  and mux113_b13_sel_is_2 (mux113_b13_sel_is_2_o, n63_neg, mux112_b13_sel_is_0_o);
  and mux113_b14_sel_is_2 (mux113_b14_sel_is_2_o, n63_neg, mux112_b14_sel_is_0_o);
  and mux113_b15_sel_is_2 (mux113_b15_sel_is_2_o, n63_neg, mux112_b15_sel_is_2_o);
  and mux113_b2_sel_is_2 (mux113_b2_sel_is_2_o, n63_neg, mux112_b11_sel_is_2_o);
  AL_MUX mux113_b5 (
    .i0(1'b1),
    .i1(n292[5]),
    .sel(mux113_b10_sel_is_0_o),
    .o(n294[5]));
  AL_MUX mux113_b6 (
    .i0(1'b0),
    .i1(n289[6]),
    .sel(mux113_b2_sel_is_2_o),
    .o(n294[6]));
  AL_MUX mux113_b8 (
    .i0(1'b0),
    .i1(n292[8]),
    .sel(mux113_b10_sel_is_0_o),
    .o(n294[8]));
  and mux113_b9_sel_is_0 (mux113_b9_sel_is_0_o, n63_neg, mux112_b9_sel_is_0_o_neg);
  not mux113_b9_sel_is_0_o_inv (mux113_b9_sel_is_0_o_neg, mux113_b9_sel_is_0_o);
  and mux114_b0_sel_is_0 (mux114_b0_sel_is_0_o, n62_neg, n63_neg);
  binary_mux_s1_w1 mux114_b1 (
    .i0(n294[1]),
    .i1(1'b1),
    .sel(n62),
    .o(n295[1]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux114_b11 (
    .i0(n294[11]),
    .i1(1'b1),
    .sel(n62),
    .o(n295[11]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux114_b12 (
    .i0(n294[12]),
    .i1(1'b0),
    .sel(n62),
    .o(n295[12]));  // sources/rtl/camera_init.v(256)
  and mux114_b13_sel_is_2 (mux114_b13_sel_is_2_o, n62_neg, mux113_b13_sel_is_2_o);
  not mux114_b13_sel_is_2_o_inv (mux114_b13_sel_is_2_o_neg, mux114_b13_sel_is_2_o);
  AL_MUX mux114_b14 (
    .i0(1'b1),
    .i1(n291[14]),
    .sel(mux114_b14_sel_is_2_o),
    .o(n295[14]));
  and mux114_b14_sel_is_2 (mux114_b14_sel_is_2_o, n62_neg, mux113_b14_sel_is_2_o);
  and mux114_b15_sel_is_2 (mux114_b15_sel_is_2_o, n62_neg, mux113_b15_sel_is_2_o);
  and mux114_b2_sel_is_2 (mux114_b2_sel_is_2_o, n62_neg, mux113_b2_sel_is_2_o);
  AL_MUX mux114_b3 (
    .i0(1'b1),
    .i1(n293[3]),
    .sel(mux114_b0_sel_is_0_o),
    .o(n295[3]));
  and mux114_b9_sel_is_0 (mux114_b9_sel_is_0_o, n62_neg, mux113_b9_sel_is_0_o_neg);
  AL_MUX mux115_b0 (
    .i0(1'b0),
    .i1(n293[0]),
    .sel(mux115_b0_sel_is_2_o),
    .o(n296[0]));
  and mux115_b0_sel_is_2 (mux115_b0_sel_is_2_o, n61_neg, mux114_b0_sel_is_0_o);
  AL_MUX mux115_b10 (
    .i0(1'b1),
    .i1(n294[10]),
    .sel(mux115_b10_sel_is_0_o),
    .o(n296[10]));
  and mux115_b10_sel_is_0 (mux115_b10_sel_is_0_o, n61_neg, n62_neg);
  and mux115_b13_sel_is_0 (mux115_b13_sel_is_0_o, n61_neg, mux114_b13_sel_is_2_o_neg);
  and mux115_b15_sel_is_2 (mux115_b15_sel_is_2_o, n61_neg, mux114_b15_sel_is_2_o);
  and mux115_b2_sel_is_2 (mux115_b2_sel_is_2_o, n61_neg, mux114_b2_sel_is_2_o);
  binary_mux_s1_w1 mux115_b3 (
    .i0(n295[3]),
    .i1(1'b0),
    .sel(n61),
    .o(n296[3]));  // sources/rtl/camera_init.v(256)
  and mux115_b4_sel_is_2 (mux115_b4_sel_is_2_o, n61_neg, mux114_b14_sel_is_2_o);
  AL_MUX mux115_b6 (
    .i0(1'b1),
    .i1(n294[6]),
    .sel(mux115_b10_sel_is_0_o),
    .o(n296[6]));
  AL_MUX mux115_b7 (
    .i0(1'b1),
    .i1(n293[7]),
    .sel(mux115_b0_sel_is_2_o),
    .o(n296[7]));
  AL_MUX mux115_b8 (
    .i0(1'b1),
    .i1(n294[8]),
    .sel(mux115_b10_sel_is_0_o),
    .o(n296[8]));
  and mux115_b9_sel_is_2 (mux115_b9_sel_is_2_o, n61_neg, mux114_b9_sel_is_0_o);
  AL_MUX mux116_b1 (
    .i0(1'b0),
    .i1(n295[1]),
    .sel(mux116_b11_sel_is_0_o),
    .o(n297[1]));
  AL_MUX mux116_b11 (
    .i0(1'b0),
    .i1(n295[11]),
    .sel(mux116_b11_sel_is_0_o),
    .o(n297[11]));
  and mux116_b11_sel_is_0 (mux116_b11_sel_is_0_o, n60_neg, n61_neg);
  and mux116_b13_sel_is_2 (mux116_b13_sel_is_2_o, n60_neg, mux115_b13_sel_is_0_o);
  not mux116_b13_sel_is_2_o_inv (mux116_b13_sel_is_2_o_neg, mux116_b13_sel_is_2_o);
  and mux116_b15_sel_is_2 (mux116_b15_sel_is_2_o, n60_neg, mux115_b15_sel_is_2_o);
  and mux116_b2_sel_is_2 (mux116_b2_sel_is_2_o, n60_neg, mux115_b2_sel_is_2_o);
  and mux116_b4_sel_is_2 (mux116_b4_sel_is_2_o, n60_neg, mux115_b4_sel_is_2_o);
  and mux116_b5_sel_is_2 (mux116_b5_sel_is_2_o, n60_neg, mux115_b10_sel_is_0_o);
  binary_mux_s1_w1 mux116_b6 (
    .i0(n296[6]),
    .i1(1'b0),
    .sel(n60),
    .o(n297[6]));  // sources/rtl/camera_init.v(256)
  and mux116_b9_sel_is_2 (mux116_b9_sel_is_2_o, n60_neg, mux115_b9_sel_is_2_o);
  AL_MUX mux117_b0 (
    .i0(1'b1),
    .i1(n296[0]),
    .sel(mux117_b0_sel_is_0_o),
    .o(n298[0]));
  and mux117_b0_sel_is_0 (mux117_b0_sel_is_0_o, n59_neg, n60_neg);
  binary_mux_s1_w1 mux117_b1 (
    .i0(n297[1]),
    .i1(1'b1),
    .sel(n59),
    .o(n298[1]));  // sources/rtl/camera_init.v(256)
  and mux117_b12_sel_is_2 (mux117_b12_sel_is_2_o, n59_neg, mux116_b11_sel_is_0_o);
  and mux117_b13_sel_is_0 (mux117_b13_sel_is_0_o, n59_neg, mux116_b13_sel_is_2_o_neg);
  and mux117_b15_sel_is_2 (mux117_b15_sel_is_2_o, n59_neg, mux116_b15_sel_is_2_o);
  and mux117_b2_sel_is_2 (mux117_b2_sel_is_2_o, n59_neg, mux116_b2_sel_is_2_o);
  AL_MUX mux117_b3 (
    .i0(1'b1),
    .i1(n296[3]),
    .sel(mux117_b0_sel_is_0_o),
    .o(n298[3]));
  and mux117_b4_sel_is_2 (mux117_b4_sel_is_2_o, n59_neg, mux116_b4_sel_is_2_o);
  and mux117_b5_sel_is_2 (mux117_b5_sel_is_2_o, n59_neg, mux116_b5_sel_is_2_o);
  binary_mux_s1_w1 mux117_b6 (
    .i0(n297[6]),
    .i1(1'b1),
    .sel(n59),
    .o(n298[6]));  // sources/rtl/camera_init.v(256)
  AL_MUX mux117_b8 (
    .i0(1'b0),
    .i1(n296[8]),
    .sel(mux117_b0_sel_is_0_o),
    .o(n298[8]));
  and mux117_b9_sel_is_2 (mux117_b9_sel_is_2_o, n59_neg, mux116_b9_sel_is_2_o);
  not mux117_b9_sel_is_2_o_inv (mux117_b9_sel_is_2_o_neg, mux117_b9_sel_is_2_o);
  binary_mux_s1_w1 mux118_b0 (
    .i0(n298[0]),
    .i1(1'b0),
    .sel(n58),
    .o(n299[0]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux118_b1 (
    .i0(n298[1]),
    .i1(1'b0),
    .sel(n58),
    .o(n299[1]));  // sources/rtl/camera_init.v(256)
  and mux118_b10_sel_is_2 (mux118_b10_sel_is_2_o, n58_neg, mux117_b0_sel_is_0_o);
  and mux118_b11_sel_is_0 (mux118_b11_sel_is_0_o, n58_neg, n59_neg);
  and mux118_b12_sel_is_2 (mux118_b12_sel_is_2_o, n58_neg, mux117_b12_sel_is_2_o);
  and mux118_b13_sel_is_2 (mux118_b13_sel_is_2_o, n58_neg, mux117_b13_sel_is_0_o);
  and mux118_b15_sel_is_2 (mux118_b15_sel_is_2_o, n58_neg, mux117_b15_sel_is_2_o);
  and mux118_b2_sel_is_2 (mux118_b2_sel_is_2_o, n58_neg, mux117_b2_sel_is_2_o);
  and mux118_b4_sel_is_2 (mux118_b4_sel_is_2_o, n58_neg, mux117_b4_sel_is_2_o);
  and mux118_b5_sel_is_2 (mux118_b5_sel_is_2_o, n58_neg, mux117_b5_sel_is_2_o);
  binary_mux_s1_w1 mux118_b6 (
    .i0(n298[6]),
    .i1(1'b0),
    .sel(n58),
    .o(n299[6]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux118_b8 (
    .i0(n298[8]),
    .i1(1'b1),
    .sel(n58),
    .o(n299[8]));  // sources/rtl/camera_init.v(256)
  and mux118_b9_sel_is_0 (mux118_b9_sel_is_0_o, n58_neg, mux117_b9_sel_is_2_o_neg);
  binary_mux_s1_w1 mux119_b1 (
    .i0(n299[1]),
    .i1(1'b1),
    .sel(n57),
    .o(n300[1]));  // sources/rtl/camera_init.v(256)
  AL_MUX mux119_b10 (
    .i0(1'b0),
    .i1(n296[10]),
    .sel(mux119_b10_sel_is_2_o),
    .o(n300[10]));
  and mux119_b10_sel_is_2 (mux119_b10_sel_is_2_o, n57_neg, mux118_b10_sel_is_2_o);
  AL_MUX mux119_b11 (
    .i0(1'b1),
    .i1(n297[11]),
    .sel(mux119_b11_sel_is_2_o),
    .o(n300[11]));
  and mux119_b11_sel_is_2 (mux119_b11_sel_is_2_o, n57_neg, mux118_b11_sel_is_0_o);
  and mux119_b12_sel_is_2 (mux119_b12_sel_is_2_o, n57_neg, mux118_b12_sel_is_2_o);
  and mux119_b13_sel_is_2 (mux119_b13_sel_is_2_o, n57_neg, mux118_b13_sel_is_2_o);
  and mux119_b15_sel_is_2 (mux119_b15_sel_is_2_o, n57_neg, mux118_b15_sel_is_2_o);
  and mux119_b2_sel_is_2 (mux119_b2_sel_is_2_o, n57_neg, mux118_b2_sel_is_2_o);
  and mux119_b3_sel_is_0 (mux119_b3_sel_is_0_o, n57_neg, n58_neg);
  AL_MUX mux119_b4 (
    .i0(1'b0),
    .i1(n291[4]),
    .sel(mux119_b4_sel_is_2_o),
    .o(n300[4]));
  and mux119_b4_sel_is_2 (mux119_b4_sel_is_2_o, n57_neg, mux118_b4_sel_is_2_o);
  and mux119_b5_sel_is_2 (mux119_b5_sel_is_2_o, n57_neg, mux118_b5_sel_is_2_o);
  binary_mux_s1_w1 mux119_b6 (
    .i0(n299[6]),
    .i1(1'b1),
    .sel(n57),
    .o(n300[6]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux119_b8 (
    .i0(n299[8]),
    .i1(1'b0),
    .sel(n57),
    .o(n300[8]));  // sources/rtl/camera_init.v(256)
  and mux119_b9_sel_is_2 (mux119_b9_sel_is_2_o, n57_neg, mux118_b9_sel_is_0_o);
  not mux119_b9_sel_is_2_o_inv (mux119_b9_sel_is_2_o_neg, mux119_b9_sel_is_2_o);
  and mux11_b0_sel_is_0 (mux11_b0_sel_is_0_o, n165_neg, n166_neg);
  and mux11_b12_sel_is_2 (mux11_b12_sel_is_2_o, n165_neg, mux10_b12_sel_is_2_o);
  and mux11_b13_sel_is_2 (mux11_b13_sel_is_2_o, n165_neg, mux10_b13_sel_is_2_o);
  and mux11_b14_sel_is_2 (mux11_b14_sel_is_2_o, n165_neg, mux10_b14_sel_is_2_o);
  and mux11_b15_sel_is_2 (mux11_b15_sel_is_2_o, n165_neg, mux10_b11_sel_is_2_o);
  and mux11_b2_sel_is_2 (mux11_b2_sel_is_2_o, n165_neg, mux10_b10_sel_is_0_o);
  binary_mux_s1_w1 mux11_b8 (
    .i0(n191[8]),
    .i1(1'b1),
    .sel(n165),
    .o(n192[8]));  // sources/rtl/camera_init.v(256)
  and mux11_b9_sel_is_0 (mux11_b9_sel_is_0_o, n165_neg, mux10_b9_sel_is_2_o_neg);
  AL_MUX mux120_b0 (
    .i0(1'b1),
    .i1(n299[0]),
    .sel(mux120_b0_sel_is_0_o),
    .o(n301[0]));
  and mux120_b0_sel_is_0 (mux120_b0_sel_is_0_o, n56_neg, n57_neg);
  binary_mux_s1_w1 mux120_b10 (
    .i0(n300[10]),
    .i1(1'b1),
    .sel(n56),
    .o(n301[10]));  // sources/rtl/camera_init.v(256)
  and mux120_b12_sel_is_2 (mux120_b12_sel_is_2_o, n56_neg, mux119_b12_sel_is_2_o);
  and mux120_b13_sel_is_2 (mux120_b13_sel_is_2_o, n56_neg, mux119_b13_sel_is_2_o);
  and mux120_b15_sel_is_2 (mux120_b15_sel_is_2_o, n56_neg, mux119_b15_sel_is_2_o);
  and mux120_b2_sel_is_2 (mux120_b2_sel_is_2_o, n56_neg, mux119_b2_sel_is_2_o);
  and mux120_b3_sel_is_2 (mux120_b3_sel_is_2_o, n56_neg, mux119_b3_sel_is_0_o);
  binary_mux_s1_w1 mux120_b4 (
    .i0(n300[4]),
    .i1(1'b1),
    .sel(n56),
    .o(n301[4]));  // sources/rtl/camera_init.v(256)
  and mux120_b5_sel_is_2 (mux120_b5_sel_is_2_o, n56_neg, mux119_b5_sel_is_2_o);
  binary_mux_s1_w1 mux120_b6 (
    .i0(n300[6]),
    .i1(1'b0),
    .sel(n56),
    .o(n301[6]));  // sources/rtl/camera_init.v(256)
  and mux120_b7_sel_is_2 (mux120_b7_sel_is_2_o, n56_neg, mux119_b10_sel_is_2_o);
  binary_mux_s1_w1 mux120_b8 (
    .i0(n300[8]),
    .i1(1'b1),
    .sel(n56),
    .o(n301[8]));  // sources/rtl/camera_init.v(256)
  and mux120_b9_sel_is_0 (mux120_b9_sel_is_0_o, n56_neg, mux119_b9_sel_is_2_o_neg);
  binary_mux_s1_w1 mux121_b0 (
    .i0(n301[0]),
    .i1(1'b0),
    .sel(n55),
    .o(n302[0]));  // sources/rtl/camera_init.v(256)
  and mux121_b11_sel_is_0 (mux121_b11_sel_is_0_o, n55_neg, n56_neg);
  and mux121_b12_sel_is_2 (mux121_b12_sel_is_2_o, n55_neg, mux120_b12_sel_is_2_o);
  and mux121_b13_sel_is_2 (mux121_b13_sel_is_2_o, n55_neg, mux120_b13_sel_is_2_o);
  not mux121_b13_sel_is_2_o_inv (mux121_b13_sel_is_2_o_neg, mux121_b13_sel_is_2_o);
  AL_MUX mux121_b14 (
    .i0(1'b0),
    .i1(n295[14]),
    .sel(mux121_b12_sel_is_2_o),
    .o(n302[14]));
  and mux121_b15_sel_is_2 (mux121_b15_sel_is_2_o, n55_neg, mux120_b15_sel_is_2_o);
  and mux121_b2_sel_is_2 (mux121_b2_sel_is_2_o, n55_neg, mux120_b2_sel_is_2_o);
  and mux121_b3_sel_is_2 (mux121_b3_sel_is_2_o, n55_neg, mux120_b3_sel_is_2_o);
  and mux121_b5_sel_is_2 (mux121_b5_sel_is_2_o, n55_neg, mux120_b5_sel_is_2_o);
  AL_MUX mux121_b7 (
    .i0(1'b0),
    .i1(n296[7]),
    .sel(mux121_b7_sel_is_2_o),
    .o(n302[7]));
  and mux121_b7_sel_is_2 (mux121_b7_sel_is_2_o, n55_neg, mux120_b7_sel_is_2_o);
  binary_mux_s1_w1 mux121_b8 (
    .i0(n301[8]),
    .i1(1'b0),
    .sel(n55),
    .o(n302[8]));  // sources/rtl/camera_init.v(256)
  and mux121_b9_sel_is_2 (mux121_b9_sel_is_2_o, n55_neg, mux120_b9_sel_is_0_o);
  binary_mux_s1_w1 mux122_b0 (
    .i0(n302[0]),
    .i1(1'b1),
    .sel(n54),
    .o(n303[0]));  // sources/rtl/camera_init.v(256)
  and mux122_b10_sel_is_0 (mux122_b10_sel_is_0_o, n54_neg, n55_neg);
  and mux122_b11_sel_is_2 (mux122_b11_sel_is_2_o, n54_neg, mux121_b11_sel_is_0_o);
  and mux122_b12_sel_is_2 (mux122_b12_sel_is_2_o, n54_neg, mux121_b12_sel_is_2_o);
  and mux122_b13_sel_is_0 (mux122_b13_sel_is_0_o, n54_neg, mux121_b13_sel_is_2_o_neg);
  and mux122_b15_sel_is_2 (mux122_b15_sel_is_2_o, n54_neg, mux121_b15_sel_is_2_o);
  AL_MUX mux122_b2 (
    .i0(1'b0),
    .i1(n289[2]),
    .sel(mux122_b2_sel_is_2_o),
    .o(n303[2]));
  and mux122_b2_sel_is_2 (mux122_b2_sel_is_2_o, n54_neg, mux121_b2_sel_is_2_o);
  and mux122_b3_sel_is_2 (mux122_b3_sel_is_2_o, n54_neg, mux121_b3_sel_is_2_o);
  AL_MUX mux122_b4 (
    .i0(1'b0),
    .i1(n301[4]),
    .sel(mux122_b10_sel_is_0_o),
    .o(n303[4]));
  and mux122_b5_sel_is_2 (mux122_b5_sel_is_2_o, n54_neg, mux121_b5_sel_is_2_o);
  AL_MUX mux122_b6 (
    .i0(1'b1),
    .i1(n301[6]),
    .sel(mux122_b10_sel_is_0_o),
    .o(n303[6]));
  and mux122_b9_sel_is_2 (mux122_b9_sel_is_2_o, n54_neg, mux121_b9_sel_is_2_o);
  not mux122_b9_sel_is_2_o_inv (mux122_b9_sel_is_2_o_neg, mux122_b9_sel_is_2_o);
  AL_MUX mux123_b1 (
    .i0(1'b0),
    .i1(n300[1]),
    .sel(mux123_b11_sel_is_2_o),
    .o(n304[1]));
  and mux123_b10_sel_is_2 (mux123_b10_sel_is_2_o, n53_neg, mux122_b10_sel_is_0_o);
  and mux123_b11_sel_is_2 (mux123_b11_sel_is_2_o, n53_neg, mux122_b11_sel_is_2_o);
  and mux123_b12_sel_is_2 (mux123_b12_sel_is_2_o, n53_neg, mux122_b12_sel_is_2_o);
  and mux123_b13_sel_is_2 (mux123_b13_sel_is_2_o, n53_neg, mux122_b13_sel_is_0_o);
  and mux123_b14_sel_is_0 (mux123_b14_sel_is_0_o, n53_neg, n54_neg);
  and mux123_b15_sel_is_2 (mux123_b15_sel_is_2_o, n53_neg, mux122_b15_sel_is_2_o);
  binary_mux_s1_w1 mux123_b2 (
    .i0(n303[2]),
    .i1(1'b1),
    .sel(n53),
    .o(n304[2]));  // sources/rtl/camera_init.v(256)
  and mux123_b3_sel_is_2 (mux123_b3_sel_is_2_o, n53_neg, mux122_b3_sel_is_2_o);
  binary_mux_s1_w1 mux123_b4 (
    .i0(n303[4]),
    .i1(1'b1),
    .sel(n53),
    .o(n304[4]));  // sources/rtl/camera_init.v(256)
  and mux123_b5_sel_is_2 (mux123_b5_sel_is_2_o, n53_neg, mux122_b5_sel_is_2_o);
  AL_MUX mux123_b7 (
    .i0(1'b1),
    .i1(n302[7]),
    .sel(mux123_b14_sel_is_0_o),
    .o(n304[7]));
  AL_MUX mux123_b8 (
    .i0(1'b1),
    .i1(n302[8]),
    .sel(mux123_b14_sel_is_0_o),
    .o(n304[8]));
  and mux123_b9_sel_is_0 (mux123_b9_sel_is_0_o, n53_neg, mux122_b9_sel_is_2_o_neg);
  and mux124_b0_sel_is_0 (mux124_b0_sel_is_0_o, n52_neg, n53_neg);
  binary_mux_s1_w1 mux124_b1 (
    .i0(n304[1]),
    .i1(1'b1),
    .sel(n52),
    .o(n305[1]));  // sources/rtl/camera_init.v(256)
  AL_MUX mux124_b10 (
    .i0(1'b0),
    .i1(n301[10]),
    .sel(mux124_b10_sel_is_2_o),
    .o(n305[10]));
  and mux124_b10_sel_is_2 (mux124_b10_sel_is_2_o, n52_neg, mux123_b10_sel_is_2_o);
  AL_MUX mux124_b11 (
    .i0(1'b0),
    .i1(n300[11]),
    .sel(mux124_b11_sel_is_2_o),
    .o(n305[11]));
  and mux124_b11_sel_is_2 (mux124_b11_sel_is_2_o, n52_neg, mux123_b11_sel_is_2_o);
  AL_MUX mux124_b12 (
    .i0(1'b1),
    .i1(n295[12]),
    .sel(mux124_b12_sel_is_2_o),
    .o(n305[12]));
  and mux124_b12_sel_is_2 (mux124_b12_sel_is_2_o, n52_neg, mux123_b12_sel_is_2_o);
  and mux124_b13_sel_is_2 (mux124_b13_sel_is_2_o, n52_neg, mux123_b13_sel_is_2_o);
  and mux124_b14_sel_is_2 (mux124_b14_sel_is_2_o, n52_neg, mux123_b14_sel_is_0_o);
  and mux124_b15_sel_is_2 (mux124_b15_sel_is_2_o, n52_neg, mux123_b15_sel_is_2_o);
  and mux124_b3_sel_is_2 (mux124_b3_sel_is_2_o, n52_neg, mux123_b3_sel_is_2_o);
  and mux124_b5_sel_is_2 (mux124_b5_sel_is_2_o, n52_neg, mux123_b5_sel_is_2_o);
  and mux124_b9_sel_is_2 (mux124_b9_sel_is_2_o, n52_neg, mux123_b9_sel_is_0_o);
  not mux124_b9_sel_is_2_o_inv (mux124_b9_sel_is_2_o_neg, mux124_b9_sel_is_2_o);
  and mux125_b0_sel_is_2 (mux125_b0_sel_is_2_o, n51_neg, mux124_b0_sel_is_0_o);
  and mux125_b13_sel_is_2 (mux125_b13_sel_is_2_o, n51_neg, mux124_b13_sel_is_2_o);
  and mux125_b14_sel_is_2 (mux125_b14_sel_is_2_o, n51_neg, mux124_b14_sel_is_2_o);
  and mux125_b15_sel_is_2 (mux125_b15_sel_is_2_o, n51_neg, mux124_b15_sel_is_2_o);
  and mux125_b2_sel_is_0 (mux125_b2_sel_is_0_o, n51_neg, n52_neg);
  and mux125_b3_sel_is_2 (mux125_b3_sel_is_2_o, n51_neg, mux124_b3_sel_is_2_o);
  and mux125_b5_sel_is_2 (mux125_b5_sel_is_2_o, n51_neg, mux124_b5_sel_is_2_o);
  AL_MUX mux125_b7 (
    .i0(1'b0),
    .i1(n304[7]),
    .sel(mux125_b2_sel_is_0_o),
    .o(n306[7]));
  AL_MUX mux125_b8 (
    .i0(1'b0),
    .i1(n304[8]),
    .sel(mux125_b2_sel_is_0_o),
    .o(n306[8]));
  and mux125_b9_sel_is_0 (mux125_b9_sel_is_0_o, n51_neg, mux124_b9_sel_is_2_o_neg);
  not mux125_b9_sel_is_0_o_inv (mux125_b9_sel_is_0_o_neg, mux125_b9_sel_is_0_o);
  and mux126_b0_sel_is_2 (mux126_b0_sel_is_2_o, n50_neg, mux125_b0_sel_is_2_o);
  and mux126_b10_sel_is_0 (mux126_b10_sel_is_0_o, n50_neg, n51_neg);
  and mux126_b13_sel_is_2 (mux126_b13_sel_is_2_o, n50_neg, mux125_b13_sel_is_2_o);
  and mux126_b14_sel_is_2 (mux126_b14_sel_is_2_o, n50_neg, mux125_b14_sel_is_2_o);
  and mux126_b15_sel_is_2 (mux126_b15_sel_is_2_o, n50_neg, mux125_b15_sel_is_2_o);
  and mux126_b2_sel_is_2 (mux126_b2_sel_is_2_o, n50_neg, mux125_b2_sel_is_0_o);
  and mux126_b3_sel_is_2 (mux126_b3_sel_is_2_o, n50_neg, mux125_b3_sel_is_2_o);
  and mux126_b5_sel_is_2 (mux126_b5_sel_is_2_o, n50_neg, mux125_b5_sel_is_2_o);
  binary_mux_s1_w1 mux126_b7 (
    .i0(n306[7]),
    .i1(1'b1),
    .sel(n50),
    .o(n307[7]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux126_b8 (
    .i0(n306[8]),
    .i1(1'b1),
    .sel(n50),
    .o(n307[8]));  // sources/rtl/camera_init.v(256)
  and mux126_b9_sel_is_0 (mux126_b9_sel_is_0_o, n50_neg, mux125_b9_sel_is_0_o_neg);
  and mux127_b0_sel_is_2 (mux127_b0_sel_is_2_o, n49_neg, mux126_b0_sel_is_2_o);
  AL_MUX mux127_b10 (
    .i0(1'b1),
    .i1(n305[10]),
    .sel(mux127_b10_sel_is_2_o),
    .o(n308[10]));
  and mux127_b10_sel_is_2 (mux127_b10_sel_is_2_o, n49_neg, mux126_b10_sel_is_0_o);
  and mux127_b13_sel_is_2 (mux127_b13_sel_is_2_o, n49_neg, mux126_b13_sel_is_2_o);
  AL_MUX mux127_b14 (
    .i0(1'b1),
    .i1(n302[14]),
    .sel(mux127_b14_sel_is_2_o),
    .o(n308[14]));
  and mux127_b14_sel_is_2 (mux127_b14_sel_is_2_o, n49_neg, mux126_b14_sel_is_2_o);
  and mux127_b15_sel_is_2 (mux127_b15_sel_is_2_o, n49_neg, mux126_b15_sel_is_2_o);
  and mux127_b2_sel_is_2 (mux127_b2_sel_is_2_o, n49_neg, mux126_b2_sel_is_2_o);
  and mux127_b3_sel_is_2 (mux127_b3_sel_is_2_o, n49_neg, mux126_b3_sel_is_2_o);
  AL_MUX mux127_b4 (
    .i0(1'b0),
    .i1(n304[4]),
    .sel(mux127_b2_sel_is_2_o),
    .o(n308[4]));
  AL_MUX mux127_b5 (
    .i0(1'b0),
    .i1(n294[5]),
    .sel(mux127_b5_sel_is_2_o),
    .o(n308[5]));
  and mux127_b5_sel_is_2 (mux127_b5_sel_is_2_o, n49_neg, mux126_b5_sel_is_2_o);
  and mux127_b9_sel_is_2 (mux127_b9_sel_is_2_o, n49_neg, mux126_b9_sel_is_0_o);
  and mux128_b0_sel_is_2 (mux128_b0_sel_is_2_o, n48_neg, mux127_b0_sel_is_2_o);
  AL_MUX mux128_b11 (
    .i0(1'b1),
    .i1(n305[11]),
    .sel(mux128_b11_sel_is_2_o),
    .o(n309[11]));
  and mux128_b11_sel_is_2 (mux128_b11_sel_is_2_o, n48_neg, mux127_b10_sel_is_2_o);
  and mux128_b13_sel_is_2 (mux128_b13_sel_is_2_o, n48_neg, mux127_b13_sel_is_2_o);
  and mux128_b15_sel_is_2 (mux128_b15_sel_is_2_o, n48_neg, mux127_b15_sel_is_2_o);
  and mux128_b2_sel_is_2 (mux128_b2_sel_is_2_o, n48_neg, mux127_b2_sel_is_2_o);
  and mux128_b3_sel_is_2 (mux128_b3_sel_is_2_o, n48_neg, mux127_b3_sel_is_2_o);
  binary_mux_s1_w1 mux128_b4 (
    .i0(n308[4]),
    .i1(1'b1),
    .sel(n48),
    .o(n309[4]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux128_b5 (
    .i0(n308[5]),
    .i1(1'b1),
    .sel(n48),
    .o(n309[5]));  // sources/rtl/camera_init.v(256)
  AL_MUX mux128_b7 (
    .i0(1'b0),
    .i1(n307[7]),
    .sel(mux128_b7_sel_is_0_o),
    .o(n309[7]));
  and mux128_b7_sel_is_0 (mux128_b7_sel_is_0_o, n48_neg, n49_neg);
  and mux128_b9_sel_is_2 (mux128_b9_sel_is_2_o, n48_neg, mux127_b9_sel_is_2_o);
  AL_MUX mux129_b0 (
    .i0(1'b0),
    .i1(n303[0]),
    .sel(mux129_b0_sel_is_2_o),
    .o(n310[0]));
  and mux129_b0_sel_is_2 (mux129_b0_sel_is_2_o, n47_neg, mux128_b0_sel_is_2_o);
  AL_MUX mux129_b10 (
    .i0(1'b0),
    .i1(n308[10]),
    .sel(mux129_b10_sel_is_0_o),
    .o(n310[10]));
  and mux129_b10_sel_is_0 (mux129_b10_sel_is_0_o, n47_neg, n48_neg);
  binary_mux_s1_w1 mux129_b11 (
    .i0(n309[11]),
    .i1(1'b0),
    .sel(n47),
    .o(n310[11]));  // sources/rtl/camera_init.v(256)
  AL_MUX mux129_b12 (
    .i0(1'b0),
    .i1(n305[12]),
    .sel(mux129_b12_sel_is_2_o),
    .o(n310[12]));
  and mux129_b12_sel_is_2 (mux129_b12_sel_is_2_o, n47_neg, mux128_b11_sel_is_2_o);
  and mux129_b13_sel_is_2 (mux129_b13_sel_is_2_o, n47_neg, mux128_b13_sel_is_2_o);
  AL_MUX mux129_b14 (
    .i0(1'b0),
    .i1(n308[14]),
    .sel(mux129_b10_sel_is_0_o),
    .o(n310[14]));
  and mux129_b15_sel_is_2 (mux129_b15_sel_is_2_o, n47_neg, mux128_b15_sel_is_2_o);
  AL_MUX mux129_b2 (
    .i0(1'b0),
    .i1(n304[2]),
    .sel(mux129_b2_sel_is_2_o),
    .o(n310[2]));
  and mux129_b2_sel_is_2 (mux129_b2_sel_is_2_o, n47_neg, mux128_b2_sel_is_2_o);
  and mux129_b3_sel_is_2 (mux129_b3_sel_is_2_o, n47_neg, mux128_b3_sel_is_2_o);
  binary_mux_s1_w1 mux129_b7 (
    .i0(n309[7]),
    .i1(1'b1),
    .sel(n47),
    .o(n310[7]));  // sources/rtl/camera_init.v(256)
  and mux129_b8_sel_is_2 (mux129_b8_sel_is_2_o, n47_neg, mux128_b7_sel_is_0_o);
  and mux129_b9_sel_is_2 (mux129_b9_sel_is_2_o, n47_neg, mux128_b9_sel_is_2_o);
  and mux12_b0_sel_is_2 (mux12_b0_sel_is_2_o, n164_neg, mux11_b0_sel_is_0_o);
  AL_MUX mux12_b10 (
    .i0(1'b1),
    .i1(n191[10]),
    .sel(mux12_b10_sel_is_0_o),
    .o(n193[10]));
  and mux12_b10_sel_is_0 (mux12_b10_sel_is_0_o, n164_neg, n165_neg);
  and mux12_b12_sel_is_2 (mux12_b12_sel_is_2_o, n164_neg, mux11_b12_sel_is_2_o);
  and mux12_b13_sel_is_2 (mux12_b13_sel_is_2_o, n164_neg, mux11_b13_sel_is_2_o);
  and mux12_b14_sel_is_2 (mux12_b14_sel_is_2_o, n164_neg, mux11_b14_sel_is_2_o);
  and mux12_b15_sel_is_2 (mux12_b15_sel_is_2_o, n164_neg, mux11_b15_sel_is_2_o);
  and mux12_b2_sel_is_2 (mux12_b2_sel_is_2_o, n164_neg, mux11_b2_sel_is_2_o);
  binary_mux_s1_w1 mux12_b8 (
    .i0(n192[8]),
    .i1(1'b0),
    .sel(n164),
    .o(n193[8]));  // sources/rtl/camera_init.v(256)
  and mux12_b9_sel_is_2 (mux12_b9_sel_is_2_o, n164_neg, mux11_b9_sel_is_0_o);
  not mux12_b9_sel_is_2_o_inv (mux12_b9_sel_is_2_o_neg, mux12_b9_sel_is_2_o);
  binary_mux_s1_w1 mux130_b0 (
    .i0(n310[0]),
    .i1(1'b1),
    .sel(n46),
    .o(n311[0]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux130_b10 (
    .i0(n310[10]),
    .i1(1'b1),
    .sel(n46),
    .o(n311[10]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux130_b11 (
    .i0(n310[11]),
    .i1(1'b1),
    .sel(n46),
    .o(n311[11]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux130_b12 (
    .i0(n310[12]),
    .i1(1'b1),
    .sel(n46),
    .o(n311[12]));  // sources/rtl/camera_init.v(256)
  and mux130_b13_sel_is_2 (mux130_b13_sel_is_2_o, n46_neg, mux129_b13_sel_is_2_o);
  and mux130_b15_sel_is_2 (mux130_b15_sel_is_2_o, n46_neg, mux129_b15_sel_is_2_o);
  and mux130_b1_sel_is_2 (mux130_b1_sel_is_2_o, n46_neg, mux129_b12_sel_is_2_o);
  binary_mux_s1_w1 mux130_b2 (
    .i0(n310[2]),
    .i1(1'b1),
    .sel(n46),
    .o(n311[2]));  // sources/rtl/camera_init.v(256)
  and mux130_b3_sel_is_2 (mux130_b3_sel_is_2_o, n46_neg, mux129_b3_sel_is_2_o);
  and mux130_b4_sel_is_0 (mux130_b4_sel_is_0_o, n46_neg, n47_neg);
  and mux130_b6_sel_is_2 (mux130_b6_sel_is_2_o, n46_neg, mux129_b0_sel_is_2_o);
  binary_mux_s1_w1 mux130_b7 (
    .i0(n310[7]),
    .i1(1'b0),
    .sel(n46),
    .o(n311[7]));  // sources/rtl/camera_init.v(256)
  and mux130_b8_sel_is_2 (mux130_b8_sel_is_2_o, n46_neg, mux129_b8_sel_is_2_o);
  and mux130_b9_sel_is_2 (mux130_b9_sel_is_2_o, n46_neg, mux129_b9_sel_is_2_o);
  not mux130_b9_sel_is_2_o_inv (mux130_b9_sel_is_2_o_neg, mux130_b9_sel_is_2_o);
  and mux131_b13_sel_is_2 (mux131_b13_sel_is_2_o, n45_neg, mux130_b13_sel_is_2_o);
  and mux131_b14_sel_is_0 (mux131_b14_sel_is_0_o, n45_neg, n46_neg);
  and mux131_b15_sel_is_2 (mux131_b15_sel_is_2_o, n45_neg, mux130_b15_sel_is_2_o);
  and mux131_b1_sel_is_2 (mux131_b1_sel_is_2_o, n45_neg, mux130_b1_sel_is_2_o);
  and mux131_b3_sel_is_2 (mux131_b3_sel_is_2_o, n45_neg, mux130_b3_sel_is_2_o);
  AL_MUX mux131_b4 (
    .i0(1'b0),
    .i1(n309[4]),
    .sel(mux131_b4_sel_is_2_o),
    .o(n312[4]));
  and mux131_b4_sel_is_2 (mux131_b4_sel_is_2_o, n45_neg, mux130_b4_sel_is_0_o);
  AL_MUX mux131_b5 (
    .i0(1'b0),
    .i1(n309[5]),
    .sel(mux131_b4_sel_is_2_o),
    .o(n312[5]));
  AL_MUX mux131_b6 (
    .i0(1'b0),
    .i1(n303[6]),
    .sel(mux131_b6_sel_is_2_o),
    .o(n312[6]));
  and mux131_b6_sel_is_2 (mux131_b6_sel_is_2_o, n45_neg, mux130_b6_sel_is_2_o);
  binary_mux_s1_w1 mux131_b7 (
    .i0(n311[7]),
    .i1(1'b1),
    .sel(n45),
    .o(n312[7]));  // sources/rtl/camera_init.v(256)
  AL_MUX mux131_b8 (
    .i0(1'b0),
    .i1(n307[8]),
    .sel(mux131_b8_sel_is_2_o),
    .o(n312[8]));
  and mux131_b8_sel_is_2 (mux131_b8_sel_is_2_o, n45_neg, mux130_b8_sel_is_2_o);
  and mux131_b9_sel_is_0 (mux131_b9_sel_is_0_o, n45_neg, mux130_b9_sel_is_2_o_neg);
  not mux131_b9_sel_is_0_o_inv (mux131_b9_sel_is_0_o_neg, mux131_b9_sel_is_0_o);
  and mux132_b0_sel_is_0 (mux132_b0_sel_is_0_o, n44_neg, n45_neg);
  AL_MUX mux132_b10 (
    .i0(1'b0),
    .i1(n311[10]),
    .sel(mux132_b0_sel_is_0_o),
    .o(n313[10]));
  AL_MUX mux132_b11 (
    .i0(1'b0),
    .i1(n311[11]),
    .sel(mux132_b0_sel_is_0_o),
    .o(n313[11]));
  and mux132_b13_sel_is_2 (mux132_b13_sel_is_2_o, n44_neg, mux131_b13_sel_is_2_o);
  not mux132_b13_sel_is_2_o_inv (mux132_b13_sel_is_2_o_neg, mux132_b13_sel_is_2_o);
  AL_MUX mux132_b14 (
    .i0(1'b1),
    .i1(n310[14]),
    .sel(mux132_b14_sel_is_2_o),
    .o(n313[14]));
  and mux132_b14_sel_is_2 (mux132_b14_sel_is_2_o, n44_neg, mux131_b14_sel_is_0_o);
  and mux132_b15_sel_is_2 (mux132_b15_sel_is_2_o, n44_neg, mux131_b15_sel_is_2_o);
  and mux132_b1_sel_is_2 (mux132_b1_sel_is_2_o, n44_neg, mux131_b1_sel_is_2_o);
  AL_MUX mux132_b2 (
    .i0(1'b0),
    .i1(n311[2]),
    .sel(mux132_b0_sel_is_0_o),
    .o(n313[2]));
  AL_MUX mux132_b3 (
    .i0(1'b0),
    .i1(n298[3]),
    .sel(mux132_b3_sel_is_2_o),
    .o(n313[3]));
  and mux132_b3_sel_is_2 (mux132_b3_sel_is_2_o, n44_neg, mux131_b3_sel_is_2_o);
  binary_mux_s1_w1 mux132_b6 (
    .i0(n312[6]),
    .i1(1'b1),
    .sel(n44),
    .o(n313[6]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux132_b8 (
    .i0(n312[8]),
    .i1(1'b1),
    .sel(n44),
    .o(n313[8]));  // sources/rtl/camera_init.v(256)
  and mux132_b9_sel_is_0 (mux132_b9_sel_is_0_o, n44_neg, mux131_b9_sel_is_0_o_neg);
  and mux133_b0_sel_is_2 (mux133_b0_sel_is_2_o, n43_neg, mux132_b0_sel_is_0_o);
  AL_MUX mux133_b1 (
    .i0(1'b0),
    .i1(n305[1]),
    .sel(mux133_b1_sel_is_2_o),
    .o(n314[1]));
  binary_mux_s1_w1 mux133_b11 (
    .i0(n313[11]),
    .i1(1'b1),
    .sel(n43),
    .o(n314[11]));  // sources/rtl/camera_init.v(256)
  and mux133_b13_sel_is_0 (mux133_b13_sel_is_0_o, n43_neg, mux132_b13_sel_is_2_o_neg);
  binary_mux_s1_w1 mux133_b14 (
    .i0(n313[14]),
    .i1(1'b0),
    .sel(n43),
    .o(n314[14]));  // sources/rtl/camera_init.v(256)
  and mux133_b15_sel_is_2 (mux133_b15_sel_is_2_o, n43_neg, mux132_b15_sel_is_2_o);
  and mux133_b1_sel_is_2 (mux133_b1_sel_is_2_o, n43_neg, mux132_b1_sel_is_2_o);
  binary_mux_s1_w1 mux133_b2 (
    .i0(n313[2]),
    .i1(1'b1),
    .sel(n43),
    .o(n314[2]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux133_b3 (
    .i0(n313[3]),
    .i1(1'b1),
    .sel(n43),
    .o(n314[3]));  // sources/rtl/camera_init.v(256)
  AL_MUX mux133_b4 (
    .i0(1'b1),
    .i1(n312[4]),
    .sel(mux133_b4_sel_is_0_o),
    .o(n314[4]));
  and mux133_b4_sel_is_0 (mux133_b4_sel_is_0_o, n43_neg, n44_neg);
  and mux133_b9_sel_is_2 (mux133_b9_sel_is_2_o, n43_neg, mux132_b9_sel_is_0_o);
  not mux133_b9_sel_is_2_o_inv (mux133_b9_sel_is_2_o_neg, mux133_b9_sel_is_2_o);
  and mux134_b0_sel_is_2 (mux134_b0_sel_is_2_o, n42_neg, mux133_b0_sel_is_2_o);
  binary_mux_s1_w1 mux134_b1 (
    .i0(n314[1]),
    .i1(1'b1),
    .sel(n42),
    .o(n315[1]));  // sources/rtl/camera_init.v(256)
  AL_MUX mux134_b10 (
    .i0(1'b1),
    .i1(n313[10]),
    .sel(mux134_b10_sel_is_0_o),
    .o(n315[10]));
  and mux134_b10_sel_is_0 (mux134_b10_sel_is_0_o, n42_neg, n43_neg);
  and mux134_b13_sel_is_2 (mux134_b13_sel_is_2_o, n42_neg, mux133_b13_sel_is_0_o);
  not mux134_b13_sel_is_2_o_inv (mux134_b13_sel_is_2_o_neg, mux134_b13_sel_is_2_o);
  and mux134_b15_sel_is_2 (mux134_b15_sel_is_2_o, n42_neg, mux133_b15_sel_is_2_o);
  AL_MUX mux134_b5 (
    .i0(1'b1),
    .i1(n312[5]),
    .sel(mux134_b5_sel_is_2_o),
    .o(n315[5]));
  and mux134_b5_sel_is_2 (mux134_b5_sel_is_2_o, n42_neg, mux133_b4_sel_is_0_o);
  AL_MUX mux134_b8 (
    .i0(1'b0),
    .i1(n313[8]),
    .sel(mux134_b10_sel_is_0_o),
    .o(n315[8]));
  and mux134_b9_sel_is_0 (mux134_b9_sel_is_0_o, n42_neg, mux133_b9_sel_is_2_o_neg);
  and mux135_b0_sel_is_2 (mux135_b0_sel_is_2_o, n41_neg, mux134_b0_sel_is_2_o);
  binary_mux_s1_w1 mux135_b10 (
    .i0(n315[10]),
    .i1(1'b0),
    .sel(n41),
    .o(n316[10]));  // sources/rtl/camera_init.v(256)
  AL_MUX mux135_b11 (
    .i0(1'b0),
    .i1(n314[11]),
    .sel(mux135_b11_sel_is_0_o),
    .o(n316[11]));
  and mux135_b11_sel_is_0 (mux135_b11_sel_is_0_o, n41_neg, n42_neg);
  AL_MUX mux135_b12 (
    .i0(1'b0),
    .i1(n311[12]),
    .sel(mux135_b0_sel_is_2_o),
    .o(n316[12]));
  and mux135_b13_sel_is_0 (mux135_b13_sel_is_0_o, n41_neg, mux134_b13_sel_is_2_o_neg);
  not mux135_b13_sel_is_0_o_inv (mux135_b13_sel_is_0_o_neg, mux135_b13_sel_is_0_o);
  and mux135_b15_sel_is_2 (mux135_b15_sel_is_2_o, n41_neg, mux134_b15_sel_is_2_o);
  and mux135_b6_sel_is_2 (mux135_b6_sel_is_2_o, n41_neg, mux134_b10_sel_is_0_o);
  and mux135_b7_sel_is_2 (mux135_b7_sel_is_2_o, n41_neg, mux134_b5_sel_is_2_o);
  binary_mux_s1_w1 mux135_b8 (
    .i0(n315[8]),
    .i1(1'b1),
    .sel(n41),
    .o(n316[8]));  // sources/rtl/camera_init.v(256)
  and mux135_b9_sel_is_2 (mux135_b9_sel_is_2_o, n41_neg, mux134_b9_sel_is_0_o);
  not mux135_b9_sel_is_2_o_inv (mux135_b9_sel_is_2_o_neg, mux135_b9_sel_is_2_o);
  and mux136_b0_sel_is_2 (mux136_b0_sel_is_2_o, n40_neg, mux135_b0_sel_is_2_o);
  AL_MUX mux136_b1 (
    .i0(1'b0),
    .i1(n315[1]),
    .sel(mux136_b1_sel_is_0_o),
    .o(n317[1]));
  binary_mux_s1_w1 mux136_b11 (
    .i0(n316[11]),
    .i1(1'b1),
    .sel(n40),
    .o(n317[11]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux136_b12 (
    .i0(n316[12]),
    .i1(1'b1),
    .sel(n40),
    .o(n317[12]));  // sources/rtl/camera_init.v(256)
  and mux136_b13_sel_is_0 (mux136_b13_sel_is_0_o, n40_neg, mux135_b13_sel_is_0_o_neg);
  not mux136_b13_sel_is_0_o_inv (mux136_b13_sel_is_0_o_neg, mux136_b13_sel_is_0_o);
  AL_MUX mux136_b14 (
    .i0(1'b1),
    .i1(n314[14]),
    .sel(mux136_b14_sel_is_2_o),
    .o(n317[14]));
  and mux136_b14_sel_is_2 (mux136_b14_sel_is_2_o, n40_neg, mux135_b11_sel_is_0_o);
  and mux136_b15_sel_is_2 (mux136_b15_sel_is_2_o, n40_neg, mux135_b15_sel_is_2_o);
  and mux136_b1_sel_is_0 (mux136_b1_sel_is_0_o, n40_neg, n41_neg);
  and mux136_b6_sel_is_2 (mux136_b6_sel_is_2_o, n40_neg, mux135_b6_sel_is_2_o);
  AL_MUX mux136_b7 (
    .i0(1'b0),
    .i1(n312[7]),
    .sel(mux136_b7_sel_is_2_o),
    .o(n317[7]));
  and mux136_b7_sel_is_2 (mux136_b7_sel_is_2_o, n40_neg, mux135_b7_sel_is_2_o);
  and mux136_b9_sel_is_0 (mux136_b9_sel_is_0_o, n40_neg, mux135_b9_sel_is_2_o_neg);
  not mux136_b9_sel_is_0_o_inv (mux136_b9_sel_is_0_o_neg, mux136_b9_sel_is_0_o);
  and mux137_b0_sel_is_2 (mux137_b0_sel_is_2_o, n39_neg, mux136_b0_sel_is_2_o);
  binary_mux_s1_w1 mux137_b1 (
    .i0(n317[1]),
    .i1(1'b1),
    .sel(n39),
    .o(n318[1]));  // sources/rtl/camera_init.v(256)
  and mux137_b10_sel_is_0 (mux137_b10_sel_is_0_o, n39_neg, n40_neg);
  and mux137_b13_sel_is_0 (mux137_b13_sel_is_0_o, n39_neg, mux136_b13_sel_is_0_o_neg);
  and mux137_b15_sel_is_2 (mux137_b15_sel_is_2_o, n39_neg, mux136_b15_sel_is_2_o);
  and mux137_b2_sel_is_2 (mux137_b2_sel_is_2_o, n39_neg, mux136_b14_sel_is_2_o);
  AL_MUX mux137_b3 (
    .i0(1'b0),
    .i1(n314[3]),
    .sel(mux137_b2_sel_is_2_o),
    .o(n318[3]));
  AL_MUX mux137_b4 (
    .i0(1'b0),
    .i1(n314[4]),
    .sel(mux137_b2_sel_is_2_o),
    .o(n318[4]));
  AL_MUX mux137_b5 (
    .i0(1'b0),
    .i1(n315[5]),
    .sel(mux137_b5_sel_is_2_o),
    .o(n318[5]));
  and mux137_b5_sel_is_2 (mux137_b5_sel_is_2_o, n39_neg, mux136_b1_sel_is_0_o);
  and mux137_b6_sel_is_2 (mux137_b6_sel_is_2_o, n39_neg, mux136_b6_sel_is_2_o);
  binary_mux_s1_w1 mux137_b7 (
    .i0(n317[7]),
    .i1(1'b1),
    .sel(n39),
    .o(n318[7]));  // sources/rtl/camera_init.v(256)
  AL_MUX mux137_b8 (
    .i0(1'b0),
    .i1(n316[8]),
    .sel(mux137_b10_sel_is_0_o),
    .o(n318[8]));
  and mux137_b9_sel_is_0 (mux137_b9_sel_is_0_o, n39_neg, mux136_b9_sel_is_0_o_neg);
  not mux137_b9_sel_is_0_o_inv (mux137_b9_sel_is_0_o_neg, mux137_b9_sel_is_0_o);
  and mux138_b0_sel_is_2 (mux138_b0_sel_is_2_o, n38_neg, mux137_b0_sel_is_2_o);
  and mux138_b10_sel_is_2 (mux138_b10_sel_is_2_o, n38_neg, mux137_b10_sel_is_0_o);
  and mux138_b11_sel_is_0 (mux138_b11_sel_is_0_o, n38_neg, n39_neg);
  and mux138_b13_sel_is_2 (mux138_b13_sel_is_2_o, n38_neg, mux137_b13_sel_is_0_o);
  and mux138_b15_sel_is_2 (mux138_b15_sel_is_2_o, n38_neg, mux137_b15_sel_is_2_o);
  and mux138_b2_sel_is_2 (mux138_b2_sel_is_2_o, n38_neg, mux137_b2_sel_is_2_o);
  binary_mux_s1_w1 mux138_b3 (
    .i0(n318[3]),
    .i1(1'b1),
    .sel(n38),
    .o(n319[3]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux138_b4 (
    .i0(n318[4]),
    .i1(1'b1),
    .sel(n38),
    .o(n319[4]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux138_b5 (
    .i0(n318[5]),
    .i1(1'b1),
    .sel(n38),
    .o(n319[5]));  // sources/rtl/camera_init.v(256)
  AL_MUX mux138_b6 (
    .i0(1'b0),
    .i1(n313[6]),
    .sel(mux138_b6_sel_is_2_o),
    .o(n319[6]));
  and mux138_b6_sel_is_2 (mux138_b6_sel_is_2_o, n38_neg, mux137_b6_sel_is_2_o);
  binary_mux_s1_w1 mux138_b8 (
    .i0(n318[8]),
    .i1(1'b1),
    .sel(n38),
    .o(n319[8]));  // sources/rtl/camera_init.v(256)
  and mux138_b9_sel_is_0 (mux138_b9_sel_is_0_o, n38_neg, mux137_b9_sel_is_0_o_neg);
  AL_MUX mux139_b0 (
    .i0(1'b0),
    .i1(n311[0]),
    .sel(mux139_b0_sel_is_2_o),
    .o(n320[0]));
  and mux139_b0_sel_is_2 (mux139_b0_sel_is_2_o, n37_neg, mux138_b0_sel_is_2_o);
  AL_MUX mux139_b10 (
    .i0(1'b1),
    .i1(n316[10]),
    .sel(mux139_b10_sel_is_2_o),
    .o(n320[10]));
  and mux139_b10_sel_is_2 (mux139_b10_sel_is_2_o, n37_neg, mux138_b10_sel_is_2_o);
  and mux139_b11_sel_is_2 (mux139_b11_sel_is_2_o, n37_neg, mux138_b11_sel_is_0_o);
  and mux139_b13_sel_is_2 (mux139_b13_sel_is_2_o, n37_neg, mux138_b13_sel_is_2_o);
  and mux139_b15_sel_is_2 (mux139_b15_sel_is_2_o, n37_neg, mux138_b15_sel_is_2_o);
  and mux139_b1_sel_is_0 (mux139_b1_sel_is_0_o, n37_neg, n38_neg);
  and mux139_b2_sel_is_2 (mux139_b2_sel_is_2_o, n37_neg, mux138_b2_sel_is_2_o);
  binary_mux_s1_w1 mux139_b3 (
    .i0(n319[3]),
    .i1(1'b0),
    .sel(n37),
    .o(n320[3]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux139_b4 (
    .i0(n319[4]),
    .i1(1'b0),
    .sel(n37),
    .o(n320[4]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux139_b6 (
    .i0(n319[6]),
    .i1(1'b1),
    .sel(n37),
    .o(n320[6]));  // sources/rtl/camera_init.v(256)
  AL_MUX mux139_b7 (
    .i0(1'b0),
    .i1(n318[7]),
    .sel(mux139_b1_sel_is_0_o),
    .o(n320[7]));
  binary_mux_s1_w1 mux139_b8 (
    .i0(n319[8]),
    .i1(1'b0),
    .sel(n37),
    .o(n320[8]));  // sources/rtl/camera_init.v(256)
  and mux139_b9_sel_is_2 (mux139_b9_sel_is_2_o, n37_neg, mux138_b9_sel_is_0_o);
  and mux13_b0_sel_is_2 (mux13_b0_sel_is_2_o, n163_neg, mux12_b0_sel_is_2_o);
  AL_MUX mux13_b1 (
    .i0(1'b0),
    .i1(n191[1]),
    .sel(mux13_b11_sel_is_2_o),
    .o(n194[1]));
  and mux13_b11_sel_is_2 (mux13_b11_sel_is_2_o, n163_neg, mux12_b10_sel_is_0_o);
  and mux13_b12_sel_is_2 (mux13_b12_sel_is_2_o, n163_neg, mux12_b12_sel_is_2_o);
  and mux13_b13_sel_is_2 (mux13_b13_sel_is_2_o, n163_neg, mux12_b13_sel_is_2_o);
  and mux13_b14_sel_is_2 (mux13_b14_sel_is_2_o, n163_neg, mux12_b14_sel_is_2_o);
  and mux13_b15_sel_is_2 (mux13_b15_sel_is_2_o, n163_neg, mux12_b15_sel_is_2_o);
  AL_MUX mux13_b2 (
    .i0(1'b0),
    .i1(n189[0]),
    .sel(mux13_b2_sel_is_2_o),
    .o(n194[2]));
  and mux13_b2_sel_is_2 (mux13_b2_sel_is_2_o, n163_neg, mux12_b2_sel_is_2_o);
  AL_MUX mux13_b4 (
    .i0(1'b0),
    .i1(n191[4]),
    .sel(mux13_b11_sel_is_2_o),
    .o(n194[4]));
  AL_MUX mux13_b7 (
    .i0(1'b0),
    .i1(n188[7]),
    .sel(mux13_b15_sel_is_2_o),
    .o(n194[7]));
  binary_mux_s1_w1 mux13_b8 (
    .i0(n193[8]),
    .i1(1'b1),
    .sel(n163),
    .o(n194[8]));  // sources/rtl/camera_init.v(256)
  and mux13_b9_sel_is_0 (mux13_b9_sel_is_0_o, n163_neg, mux12_b9_sel_is_2_o_neg);
  AL_MUX mux140_b11 (
    .i0(1'b0),
    .i1(n317[11]),
    .sel(mux140_b11_sel_is_2_o),
    .o(n321[11]));
  and mux140_b11_sel_is_2 (mux140_b11_sel_is_2_o, n36_neg, mux139_b11_sel_is_2_o);
  and mux140_b13_sel_is_2 (mux140_b13_sel_is_2_o, n36_neg, mux139_b13_sel_is_2_o);
  not mux140_b13_sel_is_2_o_inv (mux140_b13_sel_is_2_o_neg, mux140_b13_sel_is_2_o);
  AL_MUX mux140_b14 (
    .i0(1'b0),
    .i1(n317[14]),
    .sel(mux140_b11_sel_is_2_o),
    .o(n321[14]));
  and mux140_b15_sel_is_2 (mux140_b15_sel_is_2_o, n36_neg, mux139_b15_sel_is_2_o);
  and mux140_b1_sel_is_2 (mux140_b1_sel_is_2_o, n36_neg, mux139_b1_sel_is_0_o);
  and mux140_b2_sel_is_2 (mux140_b2_sel_is_2_o, n36_neg, mux139_b2_sel_is_2_o);
  binary_mux_s1_w1 mux140_b3 (
    .i0(n320[3]),
    .i1(1'b1),
    .sel(n36),
    .o(n321[3]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux140_b4 (
    .i0(n320[4]),
    .i1(1'b1),
    .sel(n36),
    .o(n321[4]));  // sources/rtl/camera_init.v(256)
  and mux140_b5_sel_is_0 (mux140_b5_sel_is_0_o, n36_neg, n37_neg);
  binary_mux_s1_w1 mux140_b8 (
    .i0(n320[8]),
    .i1(1'b1),
    .sel(n36),
    .o(n321[8]));  // sources/rtl/camera_init.v(256)
  and mux140_b9_sel_is_2 (mux140_b9_sel_is_2_o, n36_neg, mux139_b9_sel_is_2_o);
  not mux140_b9_sel_is_2_o_inv (mux140_b9_sel_is_2_o_neg, mux140_b9_sel_is_2_o);
  and mux141_b0_sel_is_0 (mux141_b0_sel_is_0_o, n35_neg, n36_neg);
  AL_MUX mux141_b1 (
    .i0(1'b0),
    .i1(n318[1]),
    .sel(mux141_b1_sel_is_2_o),
    .o(n322[1]));
  binary_mux_s1_w1 mux141_b11 (
    .i0(n321[11]),
    .i1(1'b1),
    .sel(n35),
    .o(n322[11]));  // sources/rtl/camera_init.v(256)
  and mux141_b12_sel_is_2 (mux141_b12_sel_is_2_o, n35_neg, mux140_b11_sel_is_2_o);
  and mux141_b13_sel_is_0 (mux141_b13_sel_is_0_o, n35_neg, mux140_b13_sel_is_2_o_neg);
  and mux141_b15_sel_is_2 (mux141_b15_sel_is_2_o, n35_neg, mux140_b15_sel_is_2_o);
  and mux141_b1_sel_is_2 (mux141_b1_sel_is_2_o, n35_neg, mux140_b1_sel_is_2_o);
  and mux141_b2_sel_is_2 (mux141_b2_sel_is_2_o, n35_neg, mux140_b2_sel_is_2_o);
  and mux141_b5_sel_is_2 (mux141_b5_sel_is_2_o, n35_neg, mux140_b5_sel_is_0_o);
  AL_MUX mux141_b7 (
    .i0(1'b1),
    .i1(n320[7]),
    .sel(mux141_b0_sel_is_0_o),
    .o(n322[7]));
  and mux141_b9_sel_is_0 (mux141_b9_sel_is_0_o, n35_neg, mux140_b9_sel_is_2_o_neg);
  AL_MUX mux142_b0 (
    .i0(1'b1),
    .i1(n320[0]),
    .sel(mux142_b0_sel_is_2_o),
    .o(n323[0]));
  and mux142_b0_sel_is_2 (mux142_b0_sel_is_2_o, n34_neg, mux141_b0_sel_is_0_o);
  binary_mux_s1_w1 mux142_b1 (
    .i0(n322[1]),
    .i1(1'b1),
    .sel(n34),
    .o(n323[1]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux142_b11 (
    .i0(n322[11]),
    .i1(1'b0),
    .sel(n34),
    .o(n323[11]));  // sources/rtl/camera_init.v(256)
  AL_MUX mux142_b12 (
    .i0(1'b0),
    .i1(n317[12]),
    .sel(mux142_b12_sel_is_2_o),
    .o(n323[12]));
  and mux142_b12_sel_is_2 (mux142_b12_sel_is_2_o, n34_neg, mux141_b12_sel_is_2_o);
  and mux142_b13_sel_is_2 (mux142_b13_sel_is_2_o, n34_neg, mux141_b13_sel_is_0_o);
  and mux142_b14_sel_is_0 (mux142_b14_sel_is_0_o, n34_neg, n35_neg);
  and mux142_b15_sel_is_2 (mux142_b15_sel_is_2_o, n34_neg, mux141_b15_sel_is_2_o);
  and mux142_b2_sel_is_2 (mux142_b2_sel_is_2_o, n34_neg, mux141_b2_sel_is_2_o);
  and mux142_b5_sel_is_2 (mux142_b5_sel_is_2_o, n34_neg, mux141_b5_sel_is_2_o);
  AL_MUX mux142_b8 (
    .i0(1'b0),
    .i1(n321[8]),
    .sel(mux142_b14_sel_is_0_o),
    .o(n323[8]));
  and mux142_b9_sel_is_2 (mux142_b9_sel_is_2_o, n34_neg, mux141_b9_sel_is_0_o);
  and mux143_b10_sel_is_2 (mux143_b10_sel_is_2_o, n33_neg, mux142_b0_sel_is_2_o);
  binary_mux_s1_w1 mux143_b12 (
    .i0(n323[12]),
    .i1(1'b1),
    .sel(n33),
    .o(n324[12]));  // sources/rtl/camera_init.v(256)
  and mux143_b13_sel_is_2 (mux143_b13_sel_is_2_o, n33_neg, mux142_b13_sel_is_2_o);
  and mux143_b14_sel_is_2 (mux143_b14_sel_is_2_o, n33_neg, mux142_b14_sel_is_0_o);
  and mux143_b15_sel_is_2 (mux143_b15_sel_is_2_o, n33_neg, mux142_b15_sel_is_2_o);
  and mux143_b2_sel_is_2 (mux143_b2_sel_is_2_o, n33_neg, mux142_b2_sel_is_2_o);
  and mux143_b5_sel_is_2 (mux143_b5_sel_is_2_o, n33_neg, mux142_b5_sel_is_2_o);
  and mux143_b7_sel_is_0 (mux143_b7_sel_is_0_o, n33_neg, n34_neg);
  binary_mux_s1_w1 mux143_b8 (
    .i0(n323[8]),
    .i1(1'b1),
    .sel(n33),
    .o(n324[8]));  // sources/rtl/camera_init.v(256)
  and mux143_b9_sel_is_2 (mux143_b9_sel_is_2_o, n33_neg, mux142_b9_sel_is_2_o);
  not mux143_b9_sel_is_2_o_inv (mux143_b9_sel_is_2_o_neg, mux143_b9_sel_is_2_o);
  and mux144_b0_sel_is_0 (mux144_b0_sel_is_0_o, n32_neg, n33_neg);
  AL_MUX mux144_b10 (
    .i0(1'b0),
    .i1(n320[10]),
    .sel(mux144_b10_sel_is_2_o),
    .o(n325[10]));
  and mux144_b10_sel_is_2 (mux144_b10_sel_is_2_o, n32_neg, mux143_b10_sel_is_2_o);
  and mux144_b13_sel_is_2 (mux144_b13_sel_is_2_o, n32_neg, mux143_b13_sel_is_2_o);
  and mux144_b14_sel_is_2 (mux144_b14_sel_is_2_o, n32_neg, mux143_b14_sel_is_2_o);
  and mux144_b15_sel_is_2 (mux144_b15_sel_is_2_o, n32_neg, mux143_b15_sel_is_2_o);
  and mux144_b2_sel_is_2 (mux144_b2_sel_is_2_o, n32_neg, mux143_b2_sel_is_2_o);
  and mux144_b5_sel_is_2 (mux144_b5_sel_is_2_o, n32_neg, mux143_b5_sel_is_2_o);
  and mux144_b7_sel_is_2 (mux144_b7_sel_is_2_o, n32_neg, mux143_b7_sel_is_0_o);
  and mux144_b9_sel_is_0 (mux144_b9_sel_is_0_o, n32_neg, mux143_b9_sel_is_2_o_neg);
  AL_MUX mux145_b0 (
    .i0(1'b0),
    .i1(n323[0]),
    .sel(mux145_b0_sel_is_2_o),
    .o(n326[0]));
  and mux145_b0_sel_is_2 (mux145_b0_sel_is_2_o, n31_neg, mux144_b0_sel_is_0_o);
  and mux145_b12_sel_is_0 (mux145_b12_sel_is_0_o, n31_neg, n32_neg);
  and mux145_b13_sel_is_2 (mux145_b13_sel_is_2_o, n31_neg, mux144_b13_sel_is_2_o);
  AL_MUX mux145_b14 (
    .i0(1'b1),
    .i1(n321[14]),
    .sel(mux145_b14_sel_is_2_o),
    .o(n326[14]));
  and mux145_b14_sel_is_2 (mux145_b14_sel_is_2_o, n31_neg, mux144_b14_sel_is_2_o);
  and mux145_b15_sel_is_2 (mux145_b15_sel_is_2_o, n31_neg, mux144_b15_sel_is_2_o);
  and mux145_b2_sel_is_2 (mux145_b2_sel_is_2_o, n31_neg, mux144_b2_sel_is_2_o);
  and mux145_b5_sel_is_2 (mux145_b5_sel_is_2_o, n31_neg, mux144_b5_sel_is_2_o);
  AL_MUX mux145_b6 (
    .i0(1'b0),
    .i1(n320[6]),
    .sel(mux145_b6_sel_is_2_o),
    .o(n326[6]));
  and mux145_b6_sel_is_2 (mux145_b6_sel_is_2_o, n31_neg, mux144_b10_sel_is_2_o);
  and mux145_b7_sel_is_2 (mux145_b7_sel_is_2_o, n31_neg, mux144_b7_sel_is_2_o);
  and mux145_b9_sel_is_2 (mux145_b9_sel_is_2_o, n31_neg, mux144_b9_sel_is_0_o);
  not mux145_b9_sel_is_2_o_inv (mux145_b9_sel_is_2_o_neg, mux145_b9_sel_is_2_o);
  AL_MUX mux146_b1 (
    .i0(1'b0),
    .i1(n323[1]),
    .sel(mux146_b11_sel_is_2_o),
    .o(n327[1]));
  and mux146_b10_sel_is_0 (mux146_b10_sel_is_0_o, n30_neg, n31_neg);
  and mux146_b11_sel_is_2 (mux146_b11_sel_is_2_o, n30_neg, mux145_b0_sel_is_2_o);
  and mux146_b12_sel_is_2 (mux146_b12_sel_is_2_o, n30_neg, mux145_b12_sel_is_0_o);
  and mux146_b13_sel_is_2 (mux146_b13_sel_is_2_o, n30_neg, mux145_b13_sel_is_2_o);
  and mux146_b15_sel_is_2 (mux146_b15_sel_is_2_o, n30_neg, mux145_b15_sel_is_2_o);
  AL_MUX mux146_b2 (
    .i0(1'b0),
    .i1(n314[2]),
    .sel(mux146_b2_sel_is_2_o),
    .o(n327[2]));
  and mux146_b2_sel_is_2 (mux146_b2_sel_is_2_o, n30_neg, mux145_b2_sel_is_2_o);
  and mux146_b3_sel_is_2 (mux146_b3_sel_is_2_o, n30_neg, mux145_b14_sel_is_2_o);
  and mux146_b5_sel_is_2 (mux146_b5_sel_is_2_o, n30_neg, mux145_b5_sel_is_2_o);
  binary_mux_s1_w1 mux146_b6 (
    .i0(n326[6]),
    .i1(1'b1),
    .sel(n30),
    .o(n327[6]));  // sources/rtl/camera_init.v(256)
  AL_MUX mux146_b7 (
    .i0(1'b0),
    .i1(n322[7]),
    .sel(mux146_b7_sel_is_2_o),
    .o(n327[7]));
  and mux146_b7_sel_is_2 (mux146_b7_sel_is_2_o, n30_neg, mux145_b7_sel_is_2_o);
  AL_MUX mux146_b8 (
    .i0(1'b0),
    .i1(n324[8]),
    .sel(mux146_b12_sel_is_2_o),
    .o(n327[8]));
  and mux146_b9_sel_is_0 (mux146_b9_sel_is_0_o, n30_neg, mux145_b9_sel_is_2_o_neg);
  not mux146_b9_sel_is_0_o_inv (mux146_b9_sel_is_0_o_neg, mux146_b9_sel_is_0_o);
  AL_MUX mux147_b0 (
    .i0(1'b1),
    .i1(n326[0]),
    .sel(mux147_b0_sel_is_0_o),
    .o(n328[0]));
  and mux147_b0_sel_is_0 (mux147_b0_sel_is_0_o, n29_neg, n30_neg);
  binary_mux_s1_w1 mux147_b1 (
    .i0(n327[1]),
    .i1(1'b1),
    .sel(n29),
    .o(n328[1]));  // sources/rtl/camera_init.v(256)
  and mux147_b10_sel_is_2 (mux147_b10_sel_is_2_o, n29_neg, mux146_b10_sel_is_0_o);
  AL_MUX mux147_b11 (
    .i0(1'b1),
    .i1(n323[11]),
    .sel(mux147_b11_sel_is_2_o),
    .o(n328[11]));
  and mux147_b11_sel_is_2 (mux147_b11_sel_is_2_o, n29_neg, mux146_b11_sel_is_2_o);
  and mux147_b12_sel_is_2 (mux147_b12_sel_is_2_o, n29_neg, mux146_b12_sel_is_2_o);
  and mux147_b13_sel_is_2 (mux147_b13_sel_is_2_o, n29_neg, mux146_b13_sel_is_2_o);
  and mux147_b15_sel_is_2 (mux147_b15_sel_is_2_o, n29_neg, mux146_b15_sel_is_2_o);
  binary_mux_s1_w1 mux147_b2 (
    .i0(n327[2]),
    .i1(1'b1),
    .sel(n29),
    .o(n328[2]));  // sources/rtl/camera_init.v(256)
  and mux147_b3_sel_is_2 (mux147_b3_sel_is_2_o, n29_neg, mux146_b3_sel_is_2_o);
  and mux147_b5_sel_is_2 (mux147_b5_sel_is_2_o, n29_neg, mux146_b5_sel_is_2_o);
  binary_mux_s1_w1 mux147_b6 (
    .i0(n327[6]),
    .i1(1'b0),
    .sel(n29),
    .o(n328[6]));  // sources/rtl/camera_init.v(256)
  and mux147_b9_sel_is_0 (mux147_b9_sel_is_0_o, n29_neg, mux146_b9_sel_is_0_o_neg);
  not mux147_b9_sel_is_0_o_inv (mux147_b9_sel_is_0_o_neg, mux147_b9_sel_is_0_o);
  and mux148_b10_sel_is_2 (mux148_b10_sel_is_2_o, n28_neg, mux147_b10_sel_is_2_o);
  and mux148_b12_sel_is_2 (mux148_b12_sel_is_2_o, n28_neg, mux147_b12_sel_is_2_o);
  and mux148_b13_sel_is_2 (mux148_b13_sel_is_2_o, n28_neg, mux147_b13_sel_is_2_o);
  and mux148_b14_sel_is_2 (mux148_b14_sel_is_2_o, n28_neg, mux147_b0_sel_is_0_o);
  and mux148_b15_sel_is_2 (mux148_b15_sel_is_2_o, n28_neg, mux147_b15_sel_is_2_o);
  AL_MUX mux148_b3 (
    .i0(1'b0),
    .i1(n321[3]),
    .sel(mux148_b3_sel_is_2_o),
    .o(n329[3]));
  and mux148_b3_sel_is_2 (mux148_b3_sel_is_2_o, n28_neg, mux147_b3_sel_is_2_o);
  and mux148_b5_sel_is_2 (mux148_b5_sel_is_2_o, n28_neg, mux147_b5_sel_is_2_o);
  binary_mux_s1_w1 mux148_b6 (
    .i0(n328[6]),
    .i1(1'b1),
    .sel(n28),
    .o(n329[6]));  // sources/rtl/camera_init.v(256)
  and mux148_b7_sel_is_0 (mux148_b7_sel_is_0_o, n28_neg, n29_neg);
  AL_MUX mux148_b8 (
    .i0(1'b1),
    .i1(n327[8]),
    .sel(mux148_b7_sel_is_0_o),
    .o(n329[8]));
  and mux148_b9_sel_is_0 (mux148_b9_sel_is_0_o, n28_neg, mux147_b9_sel_is_0_o_neg);
  and mux149_b0_sel_is_0 (mux149_b0_sel_is_0_o, n27_neg, n28_neg);
  AL_MUX mux149_b1 (
    .i0(1'b0),
    .i1(n328[1]),
    .sel(mux149_b0_sel_is_0_o),
    .o(n330[1]));
  and mux149_b10_sel_is_2 (mux149_b10_sel_is_2_o, n27_neg, mux148_b10_sel_is_2_o);
  AL_MUX mux149_b12 (
    .i0(1'b0),
    .i1(n324[12]),
    .sel(mux149_b12_sel_is_2_o),
    .o(n330[12]));
  and mux149_b12_sel_is_2 (mux149_b12_sel_is_2_o, n27_neg, mux148_b12_sel_is_2_o);
  and mux149_b13_sel_is_2 (mux149_b13_sel_is_2_o, n27_neg, mux148_b13_sel_is_2_o);
  not mux149_b13_sel_is_2_o_inv (mux149_b13_sel_is_2_o_neg, mux149_b13_sel_is_2_o);
  and mux149_b14_sel_is_2 (mux149_b14_sel_is_2_o, n27_neg, mux148_b14_sel_is_2_o);
  and mux149_b15_sel_is_2 (mux149_b15_sel_is_2_o, n27_neg, mux148_b15_sel_is_2_o);
  AL_MUX mux149_b4 (
    .i0(1'b0),
    .i1(n321[4]),
    .sel(mux149_b4_sel_is_2_o),
    .o(n330[4]));
  and mux149_b4_sel_is_2 (mux149_b4_sel_is_2_o, n27_neg, mux148_b3_sel_is_2_o);
  and mux149_b5_sel_is_2 (mux149_b5_sel_is_2_o, n27_neg, mux148_b5_sel_is_2_o);
  AL_MUX mux149_b7 (
    .i0(1'b1),
    .i1(n327[7]),
    .sel(mux149_b7_sel_is_2_o),
    .o(n330[7]));
  and mux149_b7_sel_is_2 (mux149_b7_sel_is_2_o, n27_neg, mux148_b7_sel_is_0_o);
  and mux149_b9_sel_is_2 (mux149_b9_sel_is_2_o, n27_neg, mux148_b9_sel_is_0_o);
  and mux14_b0_sel_is_2 (mux14_b0_sel_is_2_o, n162_neg, mux13_b0_sel_is_2_o);
  binary_mux_s1_w1 mux14_b1 (
    .i0(n194[1]),
    .i1(1'b1),
    .sel(n162),
    .o(n195[1]));  // sources/rtl/camera_init.v(256)
  and mux14_b10_sel_is_0 (mux14_b10_sel_is_0_o, n162_neg, n163_neg);
  and mux14_b11_sel_is_2 (mux14_b11_sel_is_2_o, n162_neg, mux13_b11_sel_is_2_o);
  and mux14_b12_sel_is_2 (mux14_b12_sel_is_2_o, n162_neg, mux13_b12_sel_is_2_o);
  and mux14_b13_sel_is_2 (mux14_b13_sel_is_2_o, n162_neg, mux13_b13_sel_is_2_o);
  and mux14_b14_sel_is_2 (mux14_b14_sel_is_2_o, n162_neg, mux13_b14_sel_is_2_o);
  and mux14_b15_sel_is_2 (mux14_b15_sel_is_2_o, n162_neg, mux13_b15_sel_is_2_o);
  binary_mux_s1_w1 mux14_b2 (
    .i0(n194[2]),
    .i1(1'b1),
    .sel(n162),
    .o(n195[2]));  // sources/rtl/camera_init.v(256)
  AL_MUX mux14_b3 (
    .i0(1'b0),
    .i1(n190[3]),
    .sel(mux14_b0_sel_is_2_o),
    .o(n195[3]));
  binary_mux_s1_w1 mux14_b4 (
    .i0(n194[4]),
    .i1(1'b1),
    .sel(n162),
    .o(n195[4]));  // sources/rtl/camera_init.v(256)
  AL_MUX mux14_b6 (
    .i0(1'b0),
    .i1(n189[5]),
    .sel(mux14_b6_sel_is_2_o),
    .o(n195[6]));
  and mux14_b6_sel_is_2 (mux14_b6_sel_is_2_o, n162_neg, mux13_b2_sel_is_2_o);
  binary_mux_s1_w1 mux14_b8 (
    .i0(n194[8]),
    .i1(1'b0),
    .sel(n162),
    .o(n195[8]));  // sources/rtl/camera_init.v(256)
  and mux14_b9_sel_is_2 (mux14_b9_sel_is_2_o, n162_neg, mux13_b9_sel_is_0_o);
  not mux14_b9_sel_is_2_o_inv (mux14_b9_sel_is_2_o_neg, mux14_b9_sel_is_2_o);
  and mux150_b0_sel_is_2 (mux150_b0_sel_is_2_o, n26_neg, mux149_b0_sel_is_0_o);
  binary_mux_s1_w1 mux150_b1 (
    .i0(n330[1]),
    .i1(1'b1),
    .sel(n26),
    .o(n331[1]));  // sources/rtl/camera_init.v(256)
  and mux150_b10_sel_is_2 (mux150_b10_sel_is_2_o, n26_neg, mux149_b10_sel_is_2_o);
  and mux150_b13_sel_is_0 (mux150_b13_sel_is_0_o, n26_neg, mux149_b13_sel_is_2_o_neg);
  and mux150_b14_sel_is_2 (mux150_b14_sel_is_2_o, n26_neg, mux149_b14_sel_is_2_o);
  and mux150_b15_sel_is_2 (mux150_b15_sel_is_2_o, n26_neg, mux149_b15_sel_is_2_o);
  AL_MUX mux150_b3 (
    .i0(1'b1),
    .i1(n329[3]),
    .sel(mux150_b3_sel_is_0_o),
    .o(n331[3]));
  and mux150_b3_sel_is_0 (mux150_b3_sel_is_0_o, n26_neg, n27_neg);
  binary_mux_s1_w1 mux150_b4 (
    .i0(n330[4]),
    .i1(1'b1),
    .sel(n26),
    .o(n331[4]));  // sources/rtl/camera_init.v(256)
  and mux150_b5_sel_is_2 (mux150_b5_sel_is_2_o, n26_neg, mux149_b5_sel_is_2_o);
  AL_MUX mux150_b6 (
    .i0(1'b0),
    .i1(n329[6]),
    .sel(mux150_b3_sel_is_0_o),
    .o(n331[6]));
  binary_mux_s1_w1 mux150_b7 (
    .i0(n330[7]),
    .i1(1'b0),
    .sel(n26),
    .o(n331[7]));  // sources/rtl/camera_init.v(256)
  and mux150_b9_sel_is_2 (mux150_b9_sel_is_2_o, n26_neg, mux149_b9_sel_is_2_o);
  not mux150_b9_sel_is_2_o_inv (mux150_b9_sel_is_2_o_neg, mux150_b9_sel_is_2_o);
  and mux151_b0_sel_is_2 (mux151_b0_sel_is_2_o, n25_neg, mux150_b0_sel_is_2_o);
  AL_MUX mux151_b10 (
    .i0(1'b1),
    .i1(n325[10]),
    .sel(mux151_b10_sel_is_2_o),
    .o(n332[10]));
  and mux151_b10_sel_is_2 (mux151_b10_sel_is_2_o, n25_neg, mux150_b10_sel_is_2_o);
  AL_MUX mux151_b12 (
    .i0(1'b1),
    .i1(n330[12]),
    .sel(mux151_b12_sel_is_0_o),
    .o(n332[12]));
  and mux151_b12_sel_is_0 (mux151_b12_sel_is_0_o, n25_neg, n26_neg);
  and mux151_b13_sel_is_2 (mux151_b13_sel_is_2_o, n25_neg, mux150_b13_sel_is_0_o);
  and mux151_b14_sel_is_2 (mux151_b14_sel_is_2_o, n25_neg, mux150_b14_sel_is_2_o);
  and mux151_b15_sel_is_2 (mux151_b15_sel_is_2_o, n25_neg, mux150_b15_sel_is_2_o);
  and mux151_b5_sel_is_2 (mux151_b5_sel_is_2_o, n25_neg, mux150_b5_sel_is_2_o);
  binary_mux_s1_w1 mux151_b6 (
    .i0(n331[6]),
    .i1(1'b1),
    .sel(n25),
    .o(n332[6]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux151_b7 (
    .i0(n331[7]),
    .i1(1'b1),
    .sel(n25),
    .o(n332[7]));  // sources/rtl/camera_init.v(256)
  AL_MUX mux151_b8 (
    .i0(1'b0),
    .i1(n329[8]),
    .sel(mux151_b8_sel_is_2_o),
    .o(n332[8]));
  and mux151_b8_sel_is_2 (mux151_b8_sel_is_2_o, n25_neg, mux150_b3_sel_is_0_o);
  and mux151_b9_sel_is_0 (mux151_b9_sel_is_0_o, n25_neg, mux150_b9_sel_is_2_o_neg);
  not mux151_b9_sel_is_0_o_inv (mux151_b9_sel_is_0_o_neg, mux151_b9_sel_is_0_o);
  AL_MUX mux152_b0 (
    .i0(1'b0),
    .i1(n328[0]),
    .sel(mux152_b0_sel_is_2_o),
    .o(n333[0]));
  and mux152_b0_sel_is_2 (mux152_b0_sel_is_2_o, n24_neg, mux151_b0_sel_is_2_o);
  AL_MUX mux152_b1 (
    .i0(1'b0),
    .i1(n331[1]),
    .sel(mux152_b1_sel_is_0_o),
    .o(n333[1]));
  binary_mux_s1_w1 mux152_b10 (
    .i0(n332[10]),
    .i1(1'b0),
    .sel(n24),
    .o(n333[10]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux152_b12 (
    .i0(n332[12]),
    .i1(1'b0),
    .sel(n24),
    .o(n333[12]));  // sources/rtl/camera_init.v(256)
  and mux152_b13_sel_is_2 (mux152_b13_sel_is_2_o, n24_neg, mux151_b13_sel_is_2_o);
  and mux152_b14_sel_is_2 (mux152_b14_sel_is_2_o, n24_neg, mux151_b14_sel_is_2_o);
  and mux152_b15_sel_is_2 (mux152_b15_sel_is_2_o, n24_neg, mux151_b15_sel_is_2_o);
  and mux152_b1_sel_is_0 (mux152_b1_sel_is_0_o, n24_neg, n25_neg);
  and mux152_b5_sel_is_2 (mux152_b5_sel_is_2_o, n24_neg, mux151_b5_sel_is_2_o);
  binary_mux_s1_w1 mux152_b6 (
    .i0(n332[6]),
    .i1(1'b0),
    .sel(n24),
    .o(n333[6]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux152_b7 (
    .i0(n332[7]),
    .i1(1'b0),
    .sel(n24),
    .o(n333[7]));  // sources/rtl/camera_init.v(256)
  and mux152_b9_sel_is_0 (mux152_b9_sel_is_0_o, n24_neg, mux151_b9_sel_is_0_o_neg);
  binary_mux_s1_w1 mux153_b0 (
    .i0(n333[0]),
    .i1(1'b1),
    .sel(n23),
    .o(n334[0]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux153_b10 (
    .i0(n333[10]),
    .i1(1'b1),
    .sel(n23),
    .o(n334[10]));  // sources/rtl/camera_init.v(256)
  and mux153_b11_sel_is_2 (mux153_b11_sel_is_2_o, n23_neg, mux152_b0_sel_is_2_o);
  binary_mux_s1_w1 mux153_b12 (
    .i0(n333[12]),
    .i1(1'b1),
    .sel(n23),
    .o(n334[12]));  // sources/rtl/camera_init.v(256)
  and mux153_b13_sel_is_2 (mux153_b13_sel_is_2_o, n23_neg, mux152_b13_sel_is_2_o);
  and mux153_b14_sel_is_2 (mux153_b14_sel_is_2_o, n23_neg, mux152_b14_sel_is_2_o);
  and mux153_b15_sel_is_2 (mux153_b15_sel_is_2_o, n23_neg, mux152_b15_sel_is_2_o);
  AL_MUX mux153_b3 (
    .i0(1'b0),
    .i1(n331[3]),
    .sel(mux153_b3_sel_is_2_o),
    .o(n334[3]));
  and mux153_b3_sel_is_2 (mux153_b3_sel_is_2_o, n23_neg, mux152_b1_sel_is_0_o);
  AL_MUX mux153_b4 (
    .i0(1'b0),
    .i1(n331[4]),
    .sel(mux153_b3_sel_is_2_o),
    .o(n334[4]));
  and mux153_b5_sel_is_2 (mux153_b5_sel_is_2_o, n23_neg, mux152_b5_sel_is_2_o);
  binary_mux_s1_w1 mux153_b6 (
    .i0(n333[6]),
    .i1(1'b1),
    .sel(n23),
    .o(n334[6]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux153_b7 (
    .i0(n333[7]),
    .i1(1'b1),
    .sel(n23),
    .o(n334[7]));  // sources/rtl/camera_init.v(256)
  AL_MUX mux153_b8 (
    .i0(1'b1),
    .i1(n332[8]),
    .sel(mux153_b8_sel_is_0_o),
    .o(n334[8]));
  and mux153_b8_sel_is_0 (mux153_b8_sel_is_0_o, n23_neg, n24_neg);
  and mux153_b9_sel_is_2 (mux153_b9_sel_is_2_o, n23_neg, mux152_b9_sel_is_0_o);
  binary_mux_s1_w1 mux154_b10 (
    .i0(n334[10]),
    .i1(1'b0),
    .sel(n22),
    .o(n335[10]));  // sources/rtl/camera_init.v(256)
  and mux154_b11_sel_is_2 (mux154_b11_sel_is_2_o, n22_neg, mux153_b11_sel_is_2_o);
  binary_mux_s1_w1 mux154_b12 (
    .i0(n334[12]),
    .i1(1'b0),
    .sel(n22),
    .o(n335[12]));  // sources/rtl/camera_init.v(256)
  and mux154_b13_sel_is_2 (mux154_b13_sel_is_2_o, n22_neg, mux153_b13_sel_is_2_o);
  and mux154_b14_sel_is_2 (mux154_b14_sel_is_2_o, n22_neg, mux153_b14_sel_is_2_o);
  and mux154_b15_sel_is_2 (mux154_b15_sel_is_2_o, n22_neg, mux153_b15_sel_is_2_o);
  and mux154_b1_sel_is_0 (mux154_b1_sel_is_0_o, n22_neg, n23_neg);
  and mux154_b5_sel_is_2 (mux154_b5_sel_is_2_o, n22_neg, mux153_b5_sel_is_2_o);
  binary_mux_s1_w1 mux154_b6 (
    .i0(n334[6]),
    .i1(1'b0),
    .sel(n22),
    .o(n335[6]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux154_b7 (
    .i0(n334[7]),
    .i1(1'b0),
    .sel(n22),
    .o(n335[7]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux154_b8 (
    .i0(n334[8]),
    .i1(1'b0),
    .sel(n22),
    .o(n335[8]));  // sources/rtl/camera_init.v(256)
  and mux154_b9_sel_is_2 (mux154_b9_sel_is_2_o, n22_neg, mux153_b9_sel_is_2_o);
  not mux154_b9_sel_is_2_o_inv (mux154_b9_sel_is_2_o_neg, mux154_b9_sel_is_2_o);
  and mux155_b0_sel_is_0 (mux155_b0_sel_is_0_o, n21_neg, n22_neg);
  binary_mux_s1_w1 mux155_b10 (
    .i0(n335[10]),
    .i1(1'b1),
    .sel(n21),
    .o(n336[10]));  // sources/rtl/camera_init.v(256)
  AL_MUX mux155_b11 (
    .i0(1'b0),
    .i1(n328[11]),
    .sel(mux155_b11_sel_is_2_o),
    .o(n336[11]));
  and mux155_b11_sel_is_2 (mux155_b11_sel_is_2_o, n21_neg, mux154_b11_sel_is_2_o);
  and mux155_b13_sel_is_2 (mux155_b13_sel_is_2_o, n21_neg, mux154_b13_sel_is_2_o);
  and mux155_b14_sel_is_2 (mux155_b14_sel_is_2_o, n21_neg, mux154_b14_sel_is_2_o);
  and mux155_b15_sel_is_2 (mux155_b15_sel_is_2_o, n21_neg, mux154_b15_sel_is_2_o);
  and mux155_b1_sel_is_2 (mux155_b1_sel_is_2_o, n21_neg, mux154_b1_sel_is_0_o);
  AL_MUX mux155_b3 (
    .i0(1'b1),
    .i1(n334[3]),
    .sel(mux155_b0_sel_is_0_o),
    .o(n336[3]));
  and mux155_b5_sel_is_2 (mux155_b5_sel_is_2_o, n21_neg, mux154_b5_sel_is_2_o);
  binary_mux_s1_w1 mux155_b6 (
    .i0(n335[6]),
    .i1(1'b1),
    .sel(n21),
    .o(n336[6]));  // sources/rtl/camera_init.v(256)
  and mux155_b9_sel_is_0 (mux155_b9_sel_is_0_o, n21_neg, mux154_b9_sel_is_2_o_neg);
  and mux156_b0_sel_is_2 (mux156_b0_sel_is_2_o, n20_neg, mux155_b0_sel_is_0_o);
  AL_MUX mux156_b1 (
    .i0(1'b1),
    .i1(n333[1]),
    .sel(mux156_b1_sel_is_2_o),
    .o(n337[1]));
  binary_mux_s1_w1 mux156_b10 (
    .i0(n336[10]),
    .i1(1'b0),
    .sel(n20),
    .o(n337[10]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux156_b11 (
    .i0(n336[11]),
    .i1(1'b1),
    .sel(n20),
    .o(n337[11]));  // sources/rtl/camera_init.v(256)
  and mux156_b12_sel_is_0 (mux156_b12_sel_is_0_o, n20_neg, n21_neg);
  and mux156_b13_sel_is_2 (mux156_b13_sel_is_2_o, n20_neg, mux155_b13_sel_is_2_o);
  not mux156_b13_sel_is_2_o_inv (mux156_b13_sel_is_2_o_neg, mux156_b13_sel_is_2_o);
  and mux156_b14_sel_is_2 (mux156_b14_sel_is_2_o, n20_neg, mux155_b14_sel_is_2_o);
  and mux156_b15_sel_is_2 (mux156_b15_sel_is_2_o, n20_neg, mux155_b15_sel_is_2_o);
  and mux156_b1_sel_is_2 (mux156_b1_sel_is_2_o, n20_neg, mux155_b1_sel_is_2_o);
  and mux156_b2_sel_is_2 (mux156_b2_sel_is_2_o, n20_neg, mux155_b11_sel_is_2_o);
  and mux156_b5_sel_is_2 (mux156_b5_sel_is_2_o, n20_neg, mux155_b5_sel_is_2_o);
  AL_MUX mux156_b7 (
    .i0(1'b1),
    .i1(n335[7]),
    .sel(mux156_b12_sel_is_0_o),
    .o(n337[7]));
  AL_MUX mux156_b8 (
    .i0(1'b1),
    .i1(n335[8]),
    .sel(mux156_b12_sel_is_0_o),
    .o(n337[8]));
  and mux156_b9_sel_is_2 (mux156_b9_sel_is_2_o, n20_neg, mux155_b9_sel_is_0_o);
  not mux156_b9_sel_is_2_o_inv (mux156_b9_sel_is_2_o_neg, mux156_b9_sel_is_2_o);
  AL_MUX mux157_b0 (
    .i0(1'b0),
    .i1(n334[0]),
    .sel(mux157_b0_sel_is_2_o),
    .o(n338[0]));
  and mux157_b0_sel_is_2 (mux157_b0_sel_is_2_o, n19_neg, mux156_b0_sel_is_2_o);
  binary_mux_s1_w1 mux157_b10 (
    .i0(n337[10]),
    .i1(1'b1),
    .sel(n19),
    .o(n338[10]));  // sources/rtl/camera_init.v(256)
  AL_MUX mux157_b12 (
    .i0(1'b1),
    .i1(n335[12]),
    .sel(mux157_b12_sel_is_2_o),
    .o(n338[12]));
  and mux157_b12_sel_is_2 (mux157_b12_sel_is_2_o, n19_neg, mux156_b12_sel_is_0_o);
  and mux157_b13_sel_is_0 (mux157_b13_sel_is_0_o, n19_neg, mux156_b13_sel_is_2_o_neg);
  AL_MUX mux157_b14 (
    .i0(1'b0),
    .i1(n326[14]),
    .sel(mux157_b14_sel_is_2_o),
    .o(n338[14]));
  and mux157_b14_sel_is_2 (mux157_b14_sel_is_2_o, n19_neg, mux156_b14_sel_is_2_o);
  and mux157_b15_sel_is_2 (mux157_b15_sel_is_2_o, n19_neg, mux156_b15_sel_is_2_o);
  and mux157_b2_sel_is_2 (mux157_b2_sel_is_2_o, n19_neg, mux156_b2_sel_is_2_o);
  and mux157_b3_sel_is_0 (mux157_b3_sel_is_0_o, n19_neg, n20_neg);
  and mux157_b5_sel_is_2 (mux157_b5_sel_is_2_o, n19_neg, mux156_b5_sel_is_2_o);
  binary_mux_s1_w1 mux157_b8 (
    .i0(n337[8]),
    .i1(1'b0),
    .sel(n19),
    .o(n338[8]));  // sources/rtl/camera_init.v(256)
  and mux157_b9_sel_is_0 (mux157_b9_sel_is_0_o, n19_neg, mux156_b9_sel_is_2_o_neg);
  binary_mux_s1_w1 mux158_b0 (
    .i0(n338[0]),
    .i1(1'b1),
    .sel(n18),
    .o(n339[0]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux158_b10 (
    .i0(n338[10]),
    .i1(1'b0),
    .sel(n18),
    .o(n339[10]));  // sources/rtl/camera_init.v(256)
  AL_MUX mux158_b11 (
    .i0(1'b0),
    .i1(n337[11]),
    .sel(mux158_b11_sel_is_0_o),
    .o(n339[11]));
  and mux158_b11_sel_is_0 (mux158_b11_sel_is_0_o, n18_neg, n19_neg);
  binary_mux_s1_w1 mux158_b12 (
    .i0(n338[12]),
    .i1(1'b0),
    .sel(n18),
    .o(n339[12]));  // sources/rtl/camera_init.v(256)
  and mux158_b13_sel_is_2 (mux158_b13_sel_is_2_o, n18_neg, mux157_b13_sel_is_0_o);
  not mux158_b13_sel_is_2_o_inv (mux158_b13_sel_is_2_o_neg, mux158_b13_sel_is_2_o);
  binary_mux_s1_w1 mux158_b14 (
    .i0(n338[14]),
    .i1(1'b1),
    .sel(n18),
    .o(n339[14]));  // sources/rtl/camera_init.v(256)
  and mux158_b15_sel_is_2 (mux158_b15_sel_is_2_o, n18_neg, mux157_b15_sel_is_2_o);
  and mux158_b2_sel_is_2 (mux158_b2_sel_is_2_o, n18_neg, mux157_b2_sel_is_2_o);
  and mux158_b3_sel_is_2 (mux158_b3_sel_is_2_o, n18_neg, mux157_b3_sel_is_0_o);
  AL_MUX mux158_b4 (
    .i0(1'b1),
    .i1(n334[4]),
    .sel(mux158_b4_sel_is_2_o),
    .o(n339[4]));
  and mux158_b4_sel_is_2 (mux158_b4_sel_is_2_o, n18_neg, mux157_b0_sel_is_2_o);
  and mux158_b5_sel_is_2 (mux158_b5_sel_is_2_o, n18_neg, mux157_b5_sel_is_2_o);
  binary_mux_s1_w1 mux158_b8 (
    .i0(n338[8]),
    .i1(1'b1),
    .sel(n18),
    .o(n339[8]));  // sources/rtl/camera_init.v(256)
  and mux158_b9_sel_is_2 (mux158_b9_sel_is_2_o, n18_neg, mux157_b9_sel_is_0_o);
  binary_mux_s1_w1 mux159_b0 (
    .i0(n339[0]),
    .i1(1'b0),
    .sel(n17),
    .o(n340[0]));  // sources/rtl/camera_init.v(256)
  AL_MUX mux159_b1 (
    .i0(1'b0),
    .i1(n337[1]),
    .sel(mux159_b1_sel_is_2_o),
    .o(n340[1]));
  binary_mux_s1_w1 mux159_b10 (
    .i0(n339[10]),
    .i1(1'b1),
    .sel(n17),
    .o(n340[10]));  // sources/rtl/camera_init.v(256)
  and mux159_b13_sel_is_0 (mux159_b13_sel_is_0_o, n17_neg, mux158_b13_sel_is_2_o_neg);
  and mux159_b15_sel_is_2 (mux159_b15_sel_is_2_o, n17_neg, mux158_b15_sel_is_2_o);
  and mux159_b1_sel_is_2 (mux159_b1_sel_is_2_o, n17_neg, mux158_b11_sel_is_0_o);
  and mux159_b2_sel_is_2 (mux159_b2_sel_is_2_o, n17_neg, mux158_b2_sel_is_2_o);
  AL_MUX mux159_b3 (
    .i0(1'b0),
    .i1(n336[3]),
    .sel(mux159_b3_sel_is_2_o),
    .o(n340[3]));
  and mux159_b3_sel_is_2 (mux159_b3_sel_is_2_o, n17_neg, mux158_b3_sel_is_2_o);
  binary_mux_s1_w1 mux159_b4 (
    .i0(n339[4]),
    .i1(1'b0),
    .sel(n17),
    .o(n340[4]));  // sources/rtl/camera_init.v(256)
  AL_MUX mux159_b5 (
    .i0(1'b0),
    .i1(n319[5]),
    .sel(mux159_b5_sel_is_2_o),
    .o(n340[5]));
  and mux159_b5_sel_is_2 (mux159_b5_sel_is_2_o, n17_neg, mux158_b5_sel_is_2_o);
  AL_MUX mux159_b6 (
    .i0(1'b0),
    .i1(n336[6]),
    .sel(mux159_b3_sel_is_2_o),
    .o(n340[6]));
  AL_MUX mux159_b7 (
    .i0(1'b0),
    .i1(n337[7]),
    .sel(mux159_b1_sel_is_2_o),
    .o(n340[7]));
  binary_mux_s1_w1 mux159_b8 (
    .i0(n339[8]),
    .i1(1'b0),
    .sel(n17),
    .o(n340[8]));  // sources/rtl/camera_init.v(256)
  and mux159_b9_sel_is_2 (mux159_b9_sel_is_2_o, n17_neg, mux158_b9_sel_is_2_o);
  and mux15_b0_sel_is_2 (mux15_b0_sel_is_2_o, n161_neg, mux14_b0_sel_is_2_o);
  and mux15_b10_sel_is_2 (mux15_b10_sel_is_2_o, n161_neg, mux14_b10_sel_is_0_o);
  and mux15_b11_sel_is_2 (mux15_b11_sel_is_2_o, n161_neg, mux14_b11_sel_is_2_o);
  and mux15_b12_sel_is_2 (mux15_b12_sel_is_2_o, n161_neg, mux14_b12_sel_is_2_o);
  and mux15_b13_sel_is_2 (mux15_b13_sel_is_2_o, n161_neg, mux14_b13_sel_is_2_o);
  and mux15_b14_sel_is_2 (mux15_b14_sel_is_2_o, n161_neg, mux14_b14_sel_is_2_o);
  and mux15_b15_sel_is_2 (mux15_b15_sel_is_2_o, n161_neg, mux14_b15_sel_is_2_o);
  binary_mux_s1_w1 mux15_b3 (
    .i0(n195[3]),
    .i1(1'b1),
    .sel(n161),
    .o(n196[3]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux15_b6 (
    .i0(n195[6]),
    .i1(1'b1),
    .sel(n161),
    .o(n196[6]));  // sources/rtl/camera_init.v(256)
  AL_MUX mux15_b7 (
    .i0(1'b1),
    .i1(n194[7]),
    .sel(mux15_b7_sel_is_0_o),
    .o(n196[7]));
  and mux15_b7_sel_is_0 (mux15_b7_sel_is_0_o, n161_neg, n162_neg);
  binary_mux_s1_w1 mux15_b8 (
    .i0(n195[8]),
    .i1(1'b1),
    .sel(n161),
    .o(n196[8]));  // sources/rtl/camera_init.v(256)
  and mux15_b9_sel_is_0 (mux15_b9_sel_is_0_o, n161_neg, mux14_b9_sel_is_2_o_neg);
  and mux160_b11_sel_is_0 (mux160_b11_sel_is_0_o, n16_neg, n17_neg);
  and mux160_b13_sel_is_2 (mux160_b13_sel_is_2_o, n16_neg, mux159_b13_sel_is_0_o);
  and mux160_b15_sel_is_2 (mux160_b15_sel_is_2_o, n16_neg, mux159_b15_sel_is_2_o);
  and mux160_b2_sel_is_2 (mux160_b2_sel_is_2_o, n16_neg, mux159_b2_sel_is_2_o);
  binary_mux_s1_w1 mux160_b3 (
    .i0(n340[3]),
    .i1(1'b1),
    .sel(n16),
    .o(n341[3]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux160_b6 (
    .i0(n340[6]),
    .i1(1'b1),
    .sel(n16),
    .o(n341[6]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux160_b7 (
    .i0(n340[7]),
    .i1(1'b1),
    .sel(n16),
    .o(n341[7]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux160_b8 (
    .i0(n340[8]),
    .i1(1'b1),
    .sel(n16),
    .o(n341[8]));  // sources/rtl/camera_init.v(256)
  and mux160_b9_sel_is_2 (mux160_b9_sel_is_2_o, n16_neg, mux159_b9_sel_is_2_o);
  AL_MUX mux161_b0 (
    .i0(1'b1),
    .i1(n340[0]),
    .sel(mux161_b0_sel_is_0_o),
    .o(n342[0]));
  and mux161_b0_sel_is_0 (mux161_b0_sel_is_0_o, n15_neg, n16_neg);
  AL_MUX mux161_b1 (
    .i0(1'b1),
    .i1(n340[1]),
    .sel(mux161_b0_sel_is_0_o),
    .o(n342[1]));
  AL_MUX mux161_b11 (
    .i0(1'b1),
    .i1(n339[11]),
    .sel(mux161_b11_sel_is_2_o),
    .o(n342[11]));
  and mux161_b11_sel_is_2 (mux161_b11_sel_is_2_o, n15_neg, mux160_b11_sel_is_0_o);
  and mux161_b13_sel_is_2 (mux161_b13_sel_is_2_o, n15_neg, mux160_b13_sel_is_2_o);
  and mux161_b15_sel_is_2 (mux161_b15_sel_is_2_o, n15_neg, mux160_b15_sel_is_2_o);
  and mux161_b2_sel_is_2 (mux161_b2_sel_is_2_o, n15_neg, mux160_b2_sel_is_2_o);
  binary_mux_s1_w1 mux161_b3 (
    .i0(n341[3]),
    .i1(1'b0),
    .sel(n15),
    .o(n342[3]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux161_b6 (
    .i0(n341[6]),
    .i1(1'b0),
    .sel(n15),
    .o(n342[6]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux161_b8 (
    .i0(n341[8]),
    .i1(1'b0),
    .sel(n15),
    .o(n342[8]));  // sources/rtl/camera_init.v(256)
  and mux161_b9_sel_is_2 (mux161_b9_sel_is_2_o, n15_neg, mux160_b9_sel_is_2_o);
  AL_MUX mux162_b10 (
    .i0(1'b0),
    .i1(n340[10]),
    .sel(mux162_b10_sel_is_2_o),
    .o(n343[10]));
  and mux162_b10_sel_is_2 (mux162_b10_sel_is_2_o, n14_neg, mux161_b0_sel_is_0_o);
  binary_mux_s1_w1 mux162_b11 (
    .i0(n342[11]),
    .i1(1'b0),
    .sel(n14),
    .o(n343[11]));  // sources/rtl/camera_init.v(256)
  AL_MUX mux162_b12 (
    .i0(1'b1),
    .i1(n339[12]),
    .sel(mux162_b12_sel_is_2_o),
    .o(n343[12]));
  and mux162_b12_sel_is_2 (mux162_b12_sel_is_2_o, n14_neg, mux161_b11_sel_is_2_o);
  and mux162_b13_sel_is_2 (mux162_b13_sel_is_2_o, n14_neg, mux161_b13_sel_is_2_o);
  and mux162_b15_sel_is_2 (mux162_b15_sel_is_2_o, n14_neg, mux161_b15_sel_is_2_o);
  AL_MUX mux162_b2 (
    .i0(1'b0),
    .i1(n328[2]),
    .sel(mux162_b2_sel_is_2_o),
    .o(n343[2]));
  and mux162_b2_sel_is_2 (mux162_b2_sel_is_2_o, n14_neg, mux161_b2_sel_is_2_o);
  AL_MUX mux162_b4 (
    .i0(1'b1),
    .i1(n340[4]),
    .sel(mux162_b10_sel_is_2_o),
    .o(n343[4]));
  AL_MUX mux162_b5 (
    .i0(1'b1),
    .i1(n340[5]),
    .sel(mux162_b10_sel_is_2_o),
    .o(n343[5]));
  binary_mux_s1_w1 mux162_b6 (
    .i0(n342[6]),
    .i1(1'b1),
    .sel(n14),
    .o(n343[6]));  // sources/rtl/camera_init.v(256)
  and mux162_b7_sel_is_0 (mux162_b7_sel_is_0_o, n14_neg, n15_neg);
  binary_mux_s1_w1 mux162_b8 (
    .i0(n342[8]),
    .i1(1'b1),
    .sel(n14),
    .o(n343[8]));  // sources/rtl/camera_init.v(256)
  and mux162_b9_sel_is_2 (mux162_b9_sel_is_2_o, n14_neg, mux161_b9_sel_is_2_o);
  not mux162_b9_sel_is_2_o_inv (mux162_b9_sel_is_2_o_neg, mux162_b9_sel_is_2_o);
  and mux163_b0_sel_is_0 (mux163_b0_sel_is_0_o, n13_neg, n14_neg);
  binary_mux_s1_w1 mux163_b11 (
    .i0(n343[11]),
    .i1(1'b1),
    .sel(n13),
    .o(n344[11]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux163_b12 (
    .i0(n343[12]),
    .i1(1'b0),
    .sel(n13),
    .o(n344[12]));  // sources/rtl/camera_init.v(256)
  and mux163_b13_sel_is_2 (mux163_b13_sel_is_2_o, n13_neg, mux162_b13_sel_is_2_o);
  not mux163_b13_sel_is_2_o_inv (mux163_b13_sel_is_2_o_neg, mux163_b13_sel_is_2_o);
  and mux163_b14_sel_is_2 (mux163_b14_sel_is_2_o, n13_neg, mux162_b12_sel_is_2_o);
  and mux163_b15_sel_is_2 (mux163_b15_sel_is_2_o, n13_neg, mux162_b15_sel_is_2_o);
  binary_mux_s1_w1 mux163_b2 (
    .i0(n343[2]),
    .i1(1'b1),
    .sel(n13),
    .o(n344[2]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux163_b6 (
    .i0(n343[6]),
    .i1(1'b0),
    .sel(n13),
    .o(n344[6]));  // sources/rtl/camera_init.v(256)
  and mux163_b7_sel_is_2 (mux163_b7_sel_is_2_o, n13_neg, mux162_b7_sel_is_0_o);
  and mux163_b9_sel_is_0 (mux163_b9_sel_is_0_o, n13_neg, mux162_b9_sel_is_2_o_neg);
  AL_MUX mux164_b0 (
    .i0(1'b0),
    .i1(n342[0]),
    .sel(mux164_b0_sel_is_2_o),
    .o(n345[0]));
  and mux164_b0_sel_is_2 (mux164_b0_sel_is_2_o, n12_neg, mux163_b0_sel_is_0_o);
  AL_MUX mux164_b10 (
    .i0(1'b1),
    .i1(n343[10]),
    .sel(mux164_b10_sel_is_0_o),
    .o(n345[10]));
  and mux164_b10_sel_is_0 (mux164_b10_sel_is_0_o, n12_neg, n13_neg);
  and mux164_b13_sel_is_0 (mux164_b13_sel_is_0_o, n12_neg, mux163_b13_sel_is_2_o_neg);
  and mux164_b14_sel_is_2 (mux164_b14_sel_is_2_o, n12_neg, mux163_b14_sel_is_2_o);
  and mux164_b15_sel_is_2 (mux164_b15_sel_is_2_o, n12_neg, mux163_b15_sel_is_2_o);
  binary_mux_s1_w1 mux164_b2 (
    .i0(n344[2]),
    .i1(1'b0),
    .sel(n12),
    .o(n345[2]));  // sources/rtl/camera_init.v(256)
  AL_MUX mux164_b3 (
    .i0(1'b1),
    .i1(n342[3]),
    .sel(mux164_b0_sel_is_2_o),
    .o(n345[3]));
  AL_MUX mux164_b5 (
    .i0(1'b0),
    .i1(n343[5]),
    .sel(mux164_b10_sel_is_0_o),
    .o(n345[5]));
  AL_MUX mux164_b7 (
    .i0(1'b0),
    .i1(n341[7]),
    .sel(mux164_b7_sel_is_2_o),
    .o(n345[7]));
  and mux164_b7_sel_is_2 (mux164_b7_sel_is_2_o, n12_neg, mux163_b7_sel_is_2_o);
  AL_MUX mux164_b8 (
    .i0(1'b0),
    .i1(n343[8]),
    .sel(mux164_b10_sel_is_0_o),
    .o(n345[8]));
  and mux164_b9_sel_is_2 (mux164_b9_sel_is_2_o, n12_neg, mux163_b9_sel_is_0_o);
  not mux164_b9_sel_is_2_o_inv (mux164_b9_sel_is_2_o_neg, mux164_b9_sel_is_2_o);
  binary_mux_s1_w1 mux165_b0 (
    .i0(n345[0]),
    .i1(1'b1),
    .sel(n11),
    .o(n346[0]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux165_b10 (
    .i0(n345[10]),
    .i1(1'b0),
    .sel(n11),
    .o(n346[10]));  // sources/rtl/camera_init.v(256)
  and mux165_b11_sel_is_0 (mux165_b11_sel_is_0_o, n11_neg, n12_neg);
  AL_MUX mux165_b12 (
    .i0(1'b1),
    .i1(n344[12]),
    .sel(mux165_b11_sel_is_0_o),
    .o(n346[12]));
  and mux165_b13_sel_is_2 (mux165_b13_sel_is_2_o, n11_neg, mux164_b13_sel_is_0_o);
  and mux165_b14_sel_is_2 (mux165_b14_sel_is_2_o, n11_neg, mux164_b14_sel_is_2_o);
  and mux165_b15_sel_is_2 (mux165_b15_sel_is_2_o, n11_neg, mux164_b15_sel_is_2_o);
  and mux165_b1_sel_is_2 (mux165_b1_sel_is_2_o, n11_neg, mux164_b0_sel_is_2_o);
  binary_mux_s1_w1 mux165_b2 (
    .i0(n345[2]),
    .i1(1'b1),
    .sel(n11),
    .o(n346[2]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux165_b3 (
    .i0(n345[3]),
    .i1(1'b0),
    .sel(n11),
    .o(n346[3]));  // sources/rtl/camera_init.v(256)
  and mux165_b4_sel_is_2 (mux165_b4_sel_is_2_o, n11_neg, mux164_b10_sel_is_0_o);
  AL_MUX mux165_b6 (
    .i0(1'b1),
    .i1(n344[6]),
    .sel(mux165_b11_sel_is_0_o),
    .o(n346[6]));
  binary_mux_s1_w1 mux165_b7 (
    .i0(n345[7]),
    .i1(1'b1),
    .sel(n11),
    .o(n346[7]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux165_b8 (
    .i0(n345[8]),
    .i1(1'b1),
    .sel(n11),
    .o(n346[8]));  // sources/rtl/camera_init.v(256)
  and mux165_b9_sel_is_0 (mux165_b9_sel_is_0_o, n11_neg, mux164_b9_sel_is_2_o_neg);
  not mux165_b9_sel_is_0_o_inv (mux165_b9_sel_is_0_o_neg, mux165_b9_sel_is_0_o);
  AL_MUX mux166_b1 (
    .i0(1'b0),
    .i1(n342[1]),
    .sel(mux166_b1_sel_is_2_o),
    .o(n347[1]));
  binary_mux_s1_w1 mux166_b10 (
    .i0(n346[10]),
    .i1(1'b1),
    .sel(n10),
    .o(n347[10]));  // sources/rtl/camera_init.v(256)
  AL_MUX mux166_b11 (
    .i0(1'b0),
    .i1(n344[11]),
    .sel(mux166_b11_sel_is_2_o),
    .o(n347[11]));
  and mux166_b11_sel_is_2 (mux166_b11_sel_is_2_o, n10_neg, mux165_b11_sel_is_0_o);
  and mux166_b13_sel_is_2 (mux166_b13_sel_is_2_o, n10_neg, mux165_b13_sel_is_2_o);
  and mux166_b14_sel_is_2 (mux166_b14_sel_is_2_o, n10_neg, mux165_b14_sel_is_2_o);
  and mux166_b15_sel_is_2 (mux166_b15_sel_is_2_o, n10_neg, mux165_b15_sel_is_2_o);
  and mux166_b1_sel_is_2 (mux166_b1_sel_is_2_o, n10_neg, mux165_b1_sel_is_2_o);
  binary_mux_s1_w1 mux166_b3 (
    .i0(n346[3]),
    .i1(1'b1),
    .sel(n10),
    .o(n347[3]));  // sources/rtl/camera_init.v(256)
  and mux166_b4_sel_is_2 (mux166_b4_sel_is_2_o, n10_neg, mux165_b4_sel_is_2_o);
  AL_MUX mux166_b5 (
    .i0(1'b1),
    .i1(n345[5]),
    .sel(mux166_b5_sel_is_0_o),
    .o(n347[5]));
  and mux166_b5_sel_is_0 (mux166_b5_sel_is_0_o, n10_neg, n11_neg);
  binary_mux_s1_w1 mux166_b8 (
    .i0(n346[8]),
    .i1(1'b0),
    .sel(n10),
    .o(n347[8]));  // sources/rtl/camera_init.v(256)
  and mux166_b9_sel_is_0 (mux166_b9_sel_is_0_o, n10_neg, mux165_b9_sel_is_0_o_neg);
  and mux167_b0_sel_is_0 (mux167_b0_sel_is_0_o, n9_neg, n10_neg);
  binary_mux_s1_w1 mux167_b1 (
    .i0(n347[1]),
    .i1(1'b1),
    .sel(n9),
    .o(n348[1]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux167_b11 (
    .i0(n347[11]),
    .i1(1'b1),
    .sel(n9),
    .o(n348[11]));  // sources/rtl/camera_init.v(256)
  AL_MUX mux167_b12 (
    .i0(1'b0),
    .i1(n346[12]),
    .sel(mux167_b0_sel_is_0_o),
    .o(n348[12]));
  and mux167_b13_sel_is_2 (mux167_b13_sel_is_2_o, n9_neg, mux166_b13_sel_is_2_o);
  and mux167_b14_sel_is_2 (mux167_b14_sel_is_2_o, n9_neg, mux166_b14_sel_is_2_o);
  and mux167_b15_sel_is_2 (mux167_b15_sel_is_2_o, n9_neg, mux166_b15_sel_is_2_o);
  and mux167_b4_sel_is_2 (mux167_b4_sel_is_2_o, n9_neg, mux166_b4_sel_is_2_o);
  and mux167_b9_sel_is_2 (mux167_b9_sel_is_2_o, n9_neg, mux166_b9_sel_is_0_o);
  and mux168_b0_sel_is_2 (mux168_b0_sel_is_2_o, n8_neg, mux167_b0_sel_is_0_o);
  binary_mux_s1_w1 mux168_b1 (
    .i0(n348[1]),
    .i1(1'b0),
    .sel(n8),
    .o(n349[1]));  // sources/rtl/camera_init.v(256)
  AL_MUX mux168_b10 (
    .i0(1'b0),
    .i1(n347[10]),
    .sel(mux168_b10_sel_is_0_o),
    .o(n349[10]));
  and mux168_b10_sel_is_0 (mux168_b10_sel_is_0_o, n8_neg, n9_neg);
  binary_mux_s1_w1 mux168_b11 (
    .i0(n348[11]),
    .i1(1'b0),
    .sel(n8),
    .o(n349[11]));  // sources/rtl/camera_init.v(256)
  and mux168_b13_sel_is_2 (mux168_b13_sel_is_2_o, n8_neg, mux167_b13_sel_is_2_o);
  not mux168_b13_sel_is_2_o_inv (mux168_b13_sel_is_2_o_neg, mux168_b13_sel_is_2_o);
  and mux168_b14_sel_is_2 (mux168_b14_sel_is_2_o, n8_neg, mux167_b14_sel_is_2_o);
  and mux168_b15_sel_is_2 (mux168_b15_sel_is_2_o, n8_neg, mux167_b15_sel_is_2_o);
  AL_MUX mux168_b4 (
    .i0(1'b0),
    .i1(n343[4]),
    .sel(mux168_b4_sel_is_2_o),
    .o(n349[4]));
  and mux168_b4_sel_is_2 (mux168_b4_sel_is_2_o, n8_neg, mux167_b4_sel_is_2_o);
  AL_MUX mux168_b5 (
    .i0(1'b0),
    .i1(n347[5]),
    .sel(mux168_b10_sel_is_0_o),
    .o(n349[5]));
  AL_MUX mux168_b8 (
    .i0(1'b1),
    .i1(n347[8]),
    .sel(mux168_b10_sel_is_0_o),
    .o(n349[8]));
  and mux168_b9_sel_is_2 (mux168_b9_sel_is_2_o, n8_neg, mux167_b9_sel_is_2_o);
  AL_MUX mux169_b0 (
    .i0(1'b0),
    .i1(n346[0]),
    .sel(mux169_b0_sel_is_2_o),
    .o(n350[0]));
  and mux169_b0_sel_is_2 (mux169_b0_sel_is_2_o, n7_neg, mux168_b0_sel_is_2_o);
  binary_mux_s1_w1 mux169_b1 (
    .i0(n349[1]),
    .i1(1'b1),
    .sel(n7),
    .o(n350[1]));  // sources/rtl/camera_init.v(256)
  and mux169_b12_sel_is_0 (mux169_b12_sel_is_0_o, n7_neg, n8_neg);
  and mux169_b13_sel_is_0 (mux169_b13_sel_is_0_o, n7_neg, mux168_b13_sel_is_2_o_neg);
  AL_MUX mux169_b14 (
    .i0(1'b0),
    .i1(n339[14]),
    .sel(mux169_b14_sel_is_2_o),
    .o(n350[14]));
  and mux169_b14_sel_is_2 (mux169_b14_sel_is_2_o, n7_neg, mux168_b14_sel_is_2_o);
  AL_MUX mux169_b15 (
    .i0(1'b0),
    .i1(n290[15]),
    .sel(mux169_b15_sel_is_2_o),
    .o(n350[15]));
  and mux169_b15_sel_is_2 (mux169_b15_sel_is_2_o, n7_neg, mux168_b15_sel_is_2_o);
  and mux169_b3_sel_is_2 (mux169_b3_sel_is_2_o, n7_neg, mux168_b10_sel_is_0_o);
  binary_mux_s1_w1 mux169_b4 (
    .i0(n349[4]),
    .i1(1'b1),
    .sel(n7),
    .o(n350[4]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux169_b5 (
    .i0(n349[5]),
    .i1(1'b1),
    .sel(n7),
    .o(n350[5]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux169_b8 (
    .i0(n349[8]),
    .i1(1'b0),
    .sel(n7),
    .o(n350[8]));  // sources/rtl/camera_init.v(256)
  and mux169_b9_sel_is_2 (mux169_b9_sel_is_2_o, n7_neg, mux168_b9_sel_is_2_o);
  not mux169_b9_sel_is_2_o_inv (mux169_b9_sel_is_2_o_neg, mux169_b9_sel_is_2_o);
  AL_MUX mux16_b0 (
    .i0(1'b0),
    .i1(n190[0]),
    .sel(mux16_b0_sel_is_2_o),
    .o(n197[0]));
  and mux16_b0_sel_is_2 (mux16_b0_sel_is_2_o, n160_neg, mux15_b0_sel_is_2_o);
  AL_MUX mux16_b10 (
    .i0(1'b0),
    .i1(n193[10]),
    .sel(mux16_b10_sel_is_2_o),
    .o(n197[10]));
  and mux16_b10_sel_is_2 (mux16_b10_sel_is_2_o, n160_neg, mux15_b10_sel_is_2_o);
  and mux16_b11_sel_is_2 (mux16_b11_sel_is_2_o, n160_neg, mux15_b11_sel_is_2_o);
  AL_MUX mux16_b12 (
    .i0(1'b1),
    .i1(n187[11]),
    .sel(mux16_b12_sel_is_2_o),
    .o(n197[12]));
  and mux16_b12_sel_is_2 (mux16_b12_sel_is_2_o, n160_neg, mux15_b12_sel_is_2_o);
  and mux16_b13_sel_is_2 (mux16_b13_sel_is_2_o, n160_neg, mux15_b13_sel_is_2_o);
  AL_MUX mux16_b14 (
    .i0(1'b1),
    .i1(n185[14]),
    .sel(mux16_b14_sel_is_2_o),
    .o(n197[14]));
  and mux16_b14_sel_is_2 (mux16_b14_sel_is_2_o, n160_neg, mux15_b14_sel_is_2_o);
  AL_MUX mux16_b15 (
    .i0(1'b0),
    .i1(n188[15]),
    .sel(mux16_b15_sel_is_2_o),
    .o(n197[15]));
  and mux16_b15_sel_is_2 (mux16_b15_sel_is_2_o, n160_neg, mux15_b15_sel_is_2_o);
  and mux16_b1_sel_is_0 (mux16_b1_sel_is_0_o, n160_neg, n161_neg);
  AL_MUX mux16_b2 (
    .i0(1'b0),
    .i1(n195[2]),
    .sel(mux16_b1_sel_is_0_o),
    .o(n197[2]));
  binary_mux_s1_w1 mux16_b3 (
    .i0(n196[3]),
    .i1(1'b0),
    .sel(n160),
    .o(n197[3]));  // sources/rtl/camera_init.v(256)
  AL_MUX mux16_b4 (
    .i0(1'b0),
    .i1(n195[4]),
    .sel(mux16_b1_sel_is_0_o),
    .o(n197[4]));
  AL_MUX mux16_b5 (
    .i0(1'b0),
    .i1(n191[5]),
    .sel(mux16_b11_sel_is_2_o),
    .o(n197[5]));
  and mux16_b9_sel_is_2 (mux16_b9_sel_is_2_o, n160_neg, mux15_b9_sel_is_0_o);
  not mux16_b9_sel_is_2_o_inv (mux16_b9_sel_is_2_o_neg, mux16_b9_sel_is_2_o);
  binary_mux_s1_w1 mux170_b1 (
    .i0(n350[1]),
    .i1(1'b0),
    .sel(n6),
    .o(n351[1]));  // sources/rtl/camera_init.v(256)
  and mux170_b10_sel_is_0 (mux170_b10_sel_is_0_o, n6_neg, n7_neg);
  AL_MUX mux170_b12 (
    .i0(1'b1),
    .i1(n348[12]),
    .sel(mux170_b12_sel_is_2_o),
    .o(n351[12]));
  and mux170_b12_sel_is_2 (mux170_b12_sel_is_2_o, n6_neg, mux169_b12_sel_is_0_o);
  and mux170_b13_sel_is_2 (mux170_b13_sel_is_2_o, n6_neg, mux169_b13_sel_is_0_o);
  binary_mux_s1_w1 mux170_b14 (
    .i0(n350[14]),
    .i1(1'b1),
    .sel(n6),
    .o(n351[14]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux170_b15 (
    .i0(n350[15]),
    .i1(1'b1),
    .sel(n6),
    .o(n351[15]));  // sources/rtl/camera_init.v(256)
  AL_MUX mux170_b2 (
    .i0(1'b0),
    .i1(n346[2]),
    .sel(mux170_b2_sel_is_2_o),
    .o(n351[2]));
  and mux170_b2_sel_is_2 (mux170_b2_sel_is_2_o, n6_neg, mux169_b0_sel_is_2_o);
  AL_MUX mux170_b3 (
    .i0(1'b0),
    .i1(n347[3]),
    .sel(mux170_b3_sel_is_2_o),
    .o(n351[3]));
  and mux170_b3_sel_is_2 (mux170_b3_sel_is_2_o, n6_neg, mux169_b3_sel_is_2_o);
  binary_mux_s1_w1 mux170_b4 (
    .i0(n350[4]),
    .i1(1'b0),
    .sel(n6),
    .o(n351[4]));  // sources/rtl/camera_init.v(256)
  AL_MUX mux170_b6 (
    .i0(1'b0),
    .i1(n346[6]),
    .sel(mux170_b2_sel_is_2_o),
    .o(n351[6]));
  AL_MUX mux170_b7 (
    .i0(1'b0),
    .i1(n346[7]),
    .sel(mux170_b2_sel_is_2_o),
    .o(n351[7]));
  binary_mux_s1_w1 mux170_b8 (
    .i0(n350[8]),
    .i1(1'b1),
    .sel(n6),
    .o(n351[8]));  // sources/rtl/camera_init.v(256)
  and mux170_b9_sel_is_0 (mux170_b9_sel_is_0_o, n6_neg, mux169_b9_sel_is_2_o_neg);
  and mux171_b0_sel_is_0 (mux171_b0_sel_is_0_o, n5_neg, n6_neg);
  and mux171_b10_sel_is_2 (mux171_b10_sel_is_2_o, n5_neg, mux170_b10_sel_is_0_o);
  and mux171_b13_sel_is_2 (mux171_b13_sel_is_2_o, n5_neg, mux170_b13_sel_is_2_o);
  AL_MUX mux171_b5 (
    .i0(1'b0),
    .i1(n350[5]),
    .sel(mux171_b0_sel_is_0_o),
    .o(n352[5]));
  and mux171_b9_sel_is_2 (mux171_b9_sel_is_2_o, n5_neg, mux170_b9_sel_is_0_o);
  not mux171_b9_sel_is_2_o_inv (mux171_b9_sel_is_2_o_neg, mux171_b9_sel_is_2_o);
  AL_MUX mux172_b0 (
    .i0(1'b1),
    .i1(n350[0]),
    .sel(mux172_b0_sel_is_2_o),
    .o(n353[0]));
  and mux172_b0_sel_is_2 (mux172_b0_sel_is_2_o, n4_neg, mux171_b0_sel_is_0_o);
  AL_MUX mux172_b1 (
    .i0(1'b1),
    .i1(n351[1]),
    .sel(mux172_b12_sel_is_0_o),
    .o(n353[1]));
  and mux172_b10_sel_is_2 (mux172_b10_sel_is_2_o, n4_neg, mux171_b10_sel_is_2_o);
  AL_MUX mux172_b12 (
    .i0(1'b0),
    .i1(n351[12]),
    .sel(mux172_b12_sel_is_0_o),
    .o(n353[12]));
  and mux172_b12_sel_is_0 (mux172_b12_sel_is_0_o, n4_neg, n5_neg);
  and mux172_b13_sel_is_2 (mux172_b13_sel_is_2_o, n4_neg, mux171_b13_sel_is_2_o);
  AL_MUX mux172_b14 (
    .i0(1'b0),
    .i1(n351[14]),
    .sel(mux172_b12_sel_is_0_o),
    .o(n353[14]));
  AL_MUX mux172_b15 (
    .i0(1'b0),
    .i1(n351[15]),
    .sel(mux172_b12_sel_is_0_o),
    .o(n353[15]));
  AL_MUX mux172_b2 (
    .i0(1'b1),
    .i1(n351[2]),
    .sel(mux172_b12_sel_is_0_o),
    .o(n353[2]));
  AL_MUX mux172_b3 (
    .i0(1'b1),
    .i1(n351[3]),
    .sel(mux172_b12_sel_is_0_o),
    .o(n353[3]));
  AL_MUX mux172_b4 (
    .i0(1'b1),
    .i1(n351[4]),
    .sel(mux172_b12_sel_is_0_o),
    .o(n353[4]));
  binary_mux_s1_w1 mux172_b5 (
    .i0(n352[5]),
    .i1(1'b1),
    .sel(n4),
    .o(n353[5]));  // sources/rtl/camera_init.v(256)
  AL_MUX mux172_b6 (
    .i0(1'b1),
    .i1(n351[6]),
    .sel(mux172_b12_sel_is_0_o),
    .o(n353[6]));
  AL_MUX mux172_b7 (
    .i0(1'b1),
    .i1(n351[7]),
    .sel(mux172_b12_sel_is_0_o),
    .o(n353[7]));
  AL_MUX mux172_b8 (
    .i0(1'b0),
    .i1(n351[8]),
    .sel(mux172_b12_sel_is_0_o),
    .o(n353[8]));
  and mux172_b9_sel_is_0 (mux172_b9_sel_is_0_o, n4_neg, mux171_b9_sel_is_2_o_neg);
  not mux172_b9_sel_is_0_o_inv (mux172_b9_sel_is_0_o_neg, mux172_b9_sel_is_0_o);
  AL_MUX mux173_b10 (
    .i0(1'b1),
    .i1(n349[10]),
    .sel(mux173_b10_sel_is_2_o),
    .o(n354[10]));
  and mux173_b10_sel_is_2 (mux173_b10_sel_is_2_o, n3_neg, mux172_b10_sel_is_2_o);
  AL_MUX mux173_b11 (
    .i0(1'b1),
    .i1(n349[11]),
    .sel(mux173_b10_sel_is_2_o),
    .o(n354[11]));
  and mux173_b13_sel_is_2 (mux173_b13_sel_is_2_o, n3_neg, mux172_b13_sel_is_2_o);
  not mux173_b13_sel_is_2_o_inv (mux173_b13_sel_is_2_o_neg, mux173_b13_sel_is_2_o);
  binary_mux_s1_w1 mux173_b14 (
    .i0(n353[14]),
    .i1(1'b1),
    .sel(n3),
    .o(n354[14]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux173_b15 (
    .i0(n353[15]),
    .i1(1'b1),
    .sel(n3),
    .o(n354[15]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux173_b7 (
    .i0(n353[7]),
    .i1(1'b0),
    .sel(n3),
    .o(n354[7]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux173_b8 (
    .i0(n353[8]),
    .i1(1'b1),
    .sel(n3),
    .o(n354[8]));  // sources/rtl/camera_init.v(256)
  and mux173_b9_sel_is_0 (mux173_b9_sel_is_0_o, n3_neg, mux172_b9_sel_is_0_o_neg);
  AL_MUX mux174_b0 (
    .i0(1'b0),
    .i1(n353[0]),
    .sel(mux174_b0_sel_is_0_o),
    .o(n355[0]));
  and mux174_b0_sel_is_0 (mux174_b0_sel_is_0_o, n2_neg, n3_neg);
  binary_mux_s1_w1 mux174_b10 (
    .i0(n354[10]),
    .i1(1'b0),
    .sel(n2),
    .o(n355[10]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux174_b11 (
    .i0(n354[11]),
    .i1(1'b0),
    .sel(n2),
    .o(n355[11]));  // sources/rtl/camera_init.v(256)
  and mux174_b13_sel_is_0 (mux174_b13_sel_is_0_o, n2_neg, mux173_b13_sel_is_2_o_neg);
  not mux174_b13_sel_is_0_o_inv (mux174_b13_sel_is_0_o_neg, mux174_b13_sel_is_0_o);
  binary_mux_s1_w1 mux174_b14 (
    .i0(n354[14]),
    .i1(1'b0),
    .sel(n2),
    .o(n355[14]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux174_b15 (
    .i0(n354[15]),
    .i1(1'b0),
    .sel(n2),
    .o(n355[15]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux174_b7 (
    .i0(n354[7]),
    .i1(1'b1),
    .sel(n2),
    .o(n355[7]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux174_b8 (
    .i0(n354[8]),
    .i1(1'b0),
    .sel(n2),
    .o(n355[8]));  // sources/rtl/camera_init.v(256)
  and mux174_b9_sel_is_2 (mux174_b9_sel_is_2_o, n2_neg, mux173_b9_sel_is_0_o);
  binary_mux_s1_w1 mux175_b0 (
    .i0(n355[0]),
    .i1(1'b1),
    .sel(n1),
    .o(regs_data[0]));  // sources/rtl/camera_init.v(256)
  AL_MUX mux175_b1 (
    .i0(1'b0),
    .i1(n353[1]),
    .sel(mux175_b12_sel_is_2_o),
    .o(regs_data[1]));
  binary_mux_s1_w1 mux175_b10 (
    .i0(n355[10]),
    .i1(1'b1),
    .sel(n1),
    .o(regs_data[10]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux175_b11 (
    .i0(n355[11]),
    .i1(1'b1),
    .sel(n1),
    .o(regs_data[11]));  // sources/rtl/camera_init.v(256)
  AL_MUX mux175_b12 (
    .i0(1'b1),
    .i1(n353[12]),
    .sel(mux175_b12_sel_is_2_o),
    .o(regs_data[12]));
  and mux175_b12_sel_is_2 (mux175_b12_sel_is_2_o, n1_neg, mux174_b0_sel_is_0_o);
  AL_MUX mux175_b13 (
    .i0(1'b1),
    .i1(1'b0),
    .sel(mux175_b13_sel_is_0_o),
    .o(regs_data[13]));
  and mux175_b13_sel_is_0 (mux175_b13_sel_is_0_o, n1_neg, mux174_b13_sel_is_0_o_neg);
  binary_mux_s1_w1 mux175_b14 (
    .i0(n355[14]),
    .i1(1'b1),
    .sel(n1),
    .o(regs_data[14]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux175_b15 (
    .i0(n355[15]),
    .i1(1'b1),
    .sel(n1),
    .o(regs_data[15]));  // sources/rtl/camera_init.v(256)
  AL_MUX mux175_b2 (
    .i0(1'b0),
    .i1(n353[2]),
    .sel(mux175_b12_sel_is_2_o),
    .o(regs_data[2]));
  AL_MUX mux175_b3 (
    .i0(1'b0),
    .i1(n353[3]),
    .sel(mux175_b12_sel_is_2_o),
    .o(regs_data[3]));
  AL_MUX mux175_b4 (
    .i0(1'b0),
    .i1(n353[4]),
    .sel(mux175_b12_sel_is_2_o),
    .o(regs_data[4]));
  AL_MUX mux175_b5 (
    .i0(1'b0),
    .i1(n353[5]),
    .sel(mux175_b12_sel_is_2_o),
    .o(regs_data[5]));
  AL_MUX mux175_b6 (
    .i0(1'b0),
    .i1(n353[6]),
    .sel(mux175_b12_sel_is_2_o),
    .o(regs_data[6]));
  binary_mux_s1_w1 mux175_b7 (
    .i0(n355[7]),
    .i1(1'b0),
    .sel(n1),
    .o(regs_data[7]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux175_b8 (
    .i0(n355[8]),
    .i1(1'b1),
    .sel(n1),
    .o(regs_data[8]));  // sources/rtl/camera_init.v(256)
  AL_MUX mux175_b9 (
    .i0(1'b1),
    .i1(1'b0),
    .sel(mux175_b9_sel_is_2_o),
    .o(regs_data[9]));
  and mux175_b9_sel_is_2 (mux175_b9_sel_is_2_o, n1_neg, mux174_b9_sel_is_2_o);
  binary_mux_s1_w1 mux176_b0 (
    .i0(1'b0),
    .i1(n359[3]),
    .sel(n177),
    .o(n361[0]));  // sources/rtl/camera_init.v(302)
  binary_mux_s1_w1 mux176_b4 (
    .i0(1'b1),
    .i1(n358),
    .sel(n177),
    .o(n361[4]));  // sources/rtl/camera_init.v(302)
  binary_mux_s1_w1 mux177_b0 (
    .i0(1'b0),
    .i1(n361[0]),
    .sel(success_out),
    .o(n362[0]));  // sources/rtl/camera_init.v(305)
  AL_MUX mux177_b1 (
    .i0(1'b0),
    .i1(1'b1),
    .sel(mux177_b1_sel_is_3_o),
    .o(n362[1]));
  and mux177_b1_sel_is_3 (mux177_b1_sel_is_3_o, success_out, n177);
  binary_mux_s1_w1 mux177_b2 (
    .i0(1'b1),
    .i1(1'b0),
    .sel(success_out),
    .o(n362[2]));  // sources/rtl/camera_init.v(305)
  binary_mux_s1_w1 mux177_b3 (
    .i0(1'b1),
    .i1(n361[0]),
    .sel(success_out),
    .o(n362[3]));  // sources/rtl/camera_init.v(305)
  binary_mux_s1_w1 mux177_b4 (
    .i0(1'b0),
    .i1(n361[4]),
    .sel(success_out),
    .o(n362[4]));  // sources/rtl/camera_init.v(305)
  binary_mux_s1_w1 mux178_b0 (
    .i0(state_next[0]),
    .i1(n362[0]),
    .sel(ready_out),
    .o(n363[0]));  // sources/rtl/camera_init.v(284)
  binary_mux_s1_w1 mux178_b1 (
    .i0(state_next[1]),
    .i1(n362[1]),
    .sel(ready_out),
    .o(n363[1]));  // sources/rtl/camera_init.v(284)
  binary_mux_s1_w1 mux178_b10 (
    .i0(1'b1),
    .i1(state_next[2]),
    .sel(ready_out),
    .o(n357[2]));  // sources/rtl/camera_init.v(284)
  binary_mux_s1_w1 mux178_b11 (
    .i0(1'b1),
    .i1(state_next[3]),
    .sel(ready_out),
    .o(n357[3]));  // sources/rtl/camera_init.v(284)
  binary_mux_s1_w1 mux178_b12 (
    .i0(1'b0),
    .i1(state_next[4]),
    .sel(ready_out),
    .o(n357[4]));  // sources/rtl/camera_init.v(284)
  binary_mux_s1_w1 mux178_b13 (
    .i0(1'b0),
    .i1(state_next[5]),
    .sel(ready_out),
    .o(n357[5]));  // sources/rtl/camera_init.v(284)
  binary_mux_s1_w1 mux178_b14 (
    .i0(1'b0),
    .i1(state_next[6]),
    .sel(ready_out),
    .o(n357[6]));  // sources/rtl/camera_init.v(284)
  binary_mux_s1_w1 mux178_b15 (
    .i0(1'b0),
    .i1(state_next[7]),
    .sel(ready_out),
    .o(n357[7]));  // sources/rtl/camera_init.v(284)
  binary_mux_s1_w1 mux178_b2 (
    .i0(state_next[2]),
    .i1(n362[2]),
    .sel(ready_out),
    .o(n363[2]));  // sources/rtl/camera_init.v(284)
  binary_mux_s1_w1 mux178_b3 (
    .i0(state_next[3]),
    .i1(n362[3]),
    .sel(ready_out),
    .o(n363[3]));  // sources/rtl/camera_init.v(284)
  binary_mux_s1_w1 mux178_b4 (
    .i0(state_next[4]),
    .i1(n362[4]),
    .sel(ready_out),
    .o(n363[4]));  // sources/rtl/camera_init.v(284)
  binary_mux_s1_w1 mux178_b5 (
    .i0(state_next[5]),
    .i1(1'b0),
    .sel(ready_out),
    .o(n363[5]));  // sources/rtl/camera_init.v(284)
  binary_mux_s1_w1 mux178_b6 (
    .i0(state_next[6]),
    .i1(1'b0),
    .sel(ready_out),
    .o(n363[6]));  // sources/rtl/camera_init.v(284)
  binary_mux_s1_w1 mux178_b7 (
    .i0(state_next[7]),
    .i1(1'b0),
    .sel(ready_out),
    .o(n363[7]));  // sources/rtl/camera_init.v(284)
  binary_mux_s1_w1 mux178_b8 (
    .i0(1'b1),
    .i1(state_next[0]),
    .sel(ready_out),
    .o(n357[0]));  // sources/rtl/camera_init.v(284)
  binary_mux_s1_w1 mux178_b9 (
    .i0(1'b1),
    .i1(state_next[1]),
    .sel(ready_out),
    .o(n357[1]));  // sources/rtl/camera_init.v(284)
  binary_mux_s1_w1 mux17_b0 (
    .i0(n197[0]),
    .i1(1'b1),
    .sel(n159),
    .o(n198[0]));  // sources/rtl/camera_init.v(256)
  AL_MUX mux17_b11 (
    .i0(1'b0),
    .i1(n191[11]),
    .sel(mux17_b11_sel_is_2_o),
    .o(n198[11]));
  and mux17_b11_sel_is_2 (mux17_b11_sel_is_2_o, n159_neg, mux16_b11_sel_is_2_o);
  and mux17_b13_sel_is_2 (mux17_b13_sel_is_2_o, n159_neg, mux16_b13_sel_is_2_o);
  and mux17_b1_sel_is_2 (mux17_b1_sel_is_2_o, n159_neg, mux16_b1_sel_is_0_o);
  binary_mux_s1_w1 mux17_b2 (
    .i0(n197[2]),
    .i1(1'b1),
    .sel(n159),
    .o(n198[2]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux17_b3 (
    .i0(n197[3]),
    .i1(1'b1),
    .sel(n159),
    .o(n198[3]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux17_b4 (
    .i0(n197[4]),
    .i1(1'b1),
    .sel(n159),
    .o(n198[4]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux17_b5 (
    .i0(n197[5]),
    .i1(1'b1),
    .sel(n159),
    .o(n198[5]));  // sources/rtl/camera_init.v(256)
  and mux17_b6_sel_is_0 (mux17_b6_sel_is_0_o, n159_neg, n160_neg);
  and mux17_b9_sel_is_0 (mux17_b9_sel_is_0_o, n159_neg, mux16_b9_sel_is_2_o_neg);
  not mux17_b9_sel_is_0_o_inv (mux17_b9_sel_is_0_o_neg, mux17_b9_sel_is_0_o);
  binary_mux_s1_w1 mux180_b0 (
    .i0(n372[0]),
    .i1(1'b1),
    .sel(n177),
    .o(n374[0]));  // sources/rtl/camera_init.v(368)
  binary_mux_s1_w1 mux180_b1 (
    .i0(n372[1]),
    .i1(1'b1),
    .sel(n177),
    .o(n374[1]));  // sources/rtl/camera_init.v(368)
  binary_mux_s1_w1 mux180_b2 (
    .i0(n372[2]),
    .i1(1'b0),
    .sel(n177),
    .o(n374[2]));  // sources/rtl/camera_init.v(368)
  binary_mux_s1_w1 mux180_b3 (
    .i0(n372[3]),
    .i1(1'b0),
    .sel(n177),
    .o(n374[3]));  // sources/rtl/camera_init.v(368)
  binary_mux_s1_w1 mux180_b4 (
    .i0(n372[4]),
    .i1(1'b0),
    .sel(n177),
    .o(n374[4]));  // sources/rtl/camera_init.v(368)
  binary_mux_s1_w1 mux180_b5 (
    .i0(n372[5]),
    .i1(1'b0),
    .sel(n177),
    .o(n374[5]));  // sources/rtl/camera_init.v(368)
  binary_mux_s1_w1 mux180_b6 (
    .i0(n372[6]),
    .i1(1'b0),
    .sel(n177),
    .o(n374[6]));  // sources/rtl/camera_init.v(368)
  binary_mux_s1_w1 mux180_b7 (
    .i0(n372[7]),
    .i1(1'b0),
    .sel(n177),
    .o(n374[7]));  // sources/rtl/camera_init.v(368)
  and mux181_b0_sel_is_2 (mux181_b0_sel_is_2_o, reset_n, sel3_b0_sel_is_3_o);
  binary_mux_s1_w1 mux18_b0 (
    .i0(n198[0]),
    .i1(1'b0),
    .sel(n158),
    .o(n199[0]));  // sources/rtl/camera_init.v(256)
  AL_MUX mux18_b1 (
    .i0(1'b0),
    .i1(n195[1]),
    .sel(mux18_b1_sel_is_2_o),
    .o(n199[1]));
  AL_MUX mux18_b10 (
    .i0(1'b1),
    .i1(n197[10]),
    .sel(mux18_b10_sel_is_0_o),
    .o(n199[10]));
  and mux18_b10_sel_is_0 (mux18_b10_sel_is_0_o, n158_neg, n159_neg);
  binary_mux_s1_w1 mux18_b11 (
    .i0(n198[11]),
    .i1(1'b1),
    .sel(n158),
    .o(n199[11]));  // sources/rtl/camera_init.v(256)
  and mux18_b13_sel_is_2 (mux18_b13_sel_is_2_o, n158_neg, mux17_b13_sel_is_2_o);
  AL_MUX mux18_b14 (
    .i0(1'b0),
    .i1(n197[14]),
    .sel(mux18_b10_sel_is_0_o),
    .o(n199[14]));
  and mux18_b1_sel_is_2 (mux18_b1_sel_is_2_o, n158_neg, mux17_b1_sel_is_2_o);
  binary_mux_s1_w1 mux18_b3 (
    .i0(n198[3]),
    .i1(1'b0),
    .sel(n158),
    .o(n199[3]));  // sources/rtl/camera_init.v(256)
  AL_MUX mux18_b6 (
    .i0(1'b0),
    .i1(n196[6]),
    .sel(mux18_b6_sel_is_2_o),
    .o(n199[6]));
  and mux18_b6_sel_is_2 (mux18_b6_sel_is_2_o, n158_neg, mux17_b6_sel_is_0_o);
  AL_MUX mux18_b8 (
    .i0(1'b0),
    .i1(n196[8]),
    .sel(mux18_b6_sel_is_2_o),
    .o(n199[8]));
  and mux18_b9_sel_is_0 (mux18_b9_sel_is_0_o, n158_neg, mux17_b9_sel_is_0_o_neg);
  binary_mux_s1_w1 mux19_b0 (
    .i0(n199[0]),
    .i1(1'b1),
    .sel(n157),
    .o(n200[0]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux19_b1 (
    .i0(n199[1]),
    .i1(1'b1),
    .sel(n157),
    .o(n200[1]));  // sources/rtl/camera_init.v(256)
  and mux19_b12_sel_is_2 (mux19_b12_sel_is_2_o, n157_neg, mux18_b10_sel_is_0_o);
  and mux19_b13_sel_is_2 (mux19_b13_sel_is_2_o, n157_neg, mux18_b13_sel_is_2_o);
  AL_MUX mux19_b2 (
    .i0(1'b0),
    .i1(n198[2]),
    .sel(mux19_b2_sel_is_0_o),
    .o(n200[2]));
  and mux19_b2_sel_is_0 (mux19_b2_sel_is_0_o, n157_neg, n158_neg);
  binary_mux_s1_w1 mux19_b3 (
    .i0(n199[3]),
    .i1(1'b1),
    .sel(n157),
    .o(n200[3]));  // sources/rtl/camera_init.v(256)
  AL_MUX mux19_b5 (
    .i0(1'b0),
    .i1(n198[5]),
    .sel(mux19_b2_sel_is_0_o),
    .o(n200[5]));
  and mux19_b7_sel_is_2 (mux19_b7_sel_is_2_o, n157_neg, mux18_b6_sel_is_2_o);
  binary_mux_s1_w1 mux19_b8 (
    .i0(n199[8]),
    .i1(1'b1),
    .sel(n157),
    .o(n200[8]));  // sources/rtl/camera_init.v(256)
  and mux19_b9_sel_is_2 (mux19_b9_sel_is_2_o, n157_neg, mux18_b9_sel_is_0_o);
  binary_mux_s1_w1 mux1_b0 (
    .i0(n181[0]),
    .i1(1'b0),
    .sel(n175),
    .o(n182[0]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux1_b10 (
    .i0(n181[10]),
    .i1(1'b0),
    .sel(n175),
    .o(n182[10]));  // sources/rtl/camera_init.v(256)
  and mux1_b7_sel_is_0 (mux1_b7_sel_is_0_o, n175_neg, n176_neg);
  AL_MUX mux20_b10 (
    .i0(1'b0),
    .i1(n199[10]),
    .sel(mux20_b10_sel_is_0_o),
    .o(n201[10]));
  and mux20_b10_sel_is_0 (mux20_b10_sel_is_0_o, n156_neg, n157_neg);
  and mux20_b12_sel_is_2 (mux20_b12_sel_is_2_o, n156_neg, mux19_b12_sel_is_2_o);
  and mux20_b13_sel_is_2 (mux20_b13_sel_is_2_o, n156_neg, mux19_b13_sel_is_2_o);
  binary_mux_s1_w1 mux20_b3 (
    .i0(n200[3]),
    .i1(1'b0),
    .sel(n156),
    .o(n201[3]));  // sources/rtl/camera_init.v(256)
  AL_MUX mux20_b4 (
    .i0(1'b0),
    .i1(n198[4]),
    .sel(mux20_b4_sel_is_2_o),
    .o(n201[4]));
  and mux20_b4_sel_is_2 (mux20_b4_sel_is_2_o, n156_neg, mux19_b2_sel_is_0_o);
  binary_mux_s1_w1 mux20_b5 (
    .i0(n200[5]),
    .i1(1'b1),
    .sel(n156),
    .o(n201[5]));  // sources/rtl/camera_init.v(256)
  and mux20_b7_sel_is_2 (mux20_b7_sel_is_2_o, n156_neg, mux19_b7_sel_is_2_o);
  and mux20_b9_sel_is_2 (mux20_b9_sel_is_2_o, n156_neg, mux19_b9_sel_is_2_o);
  AL_MUX mux21_b0 (
    .i0(1'b0),
    .i1(n200[0]),
    .sel(mux21_b0_sel_is_0_o),
    .o(n202[0]));
  and mux21_b0_sel_is_0 (mux21_b0_sel_is_0_o, n155_neg, n156_neg);
  AL_MUX mux21_b1 (
    .i0(1'b0),
    .i1(n200[1]),
    .sel(mux21_b0_sel_is_0_o),
    .o(n202[1]));
  binary_mux_s1_w1 mux21_b10 (
    .i0(n201[10]),
    .i1(1'b1),
    .sel(n155),
    .o(n202[10]));  // sources/rtl/camera_init.v(256)
  and mux21_b11_sel_is_2 (mux21_b11_sel_is_2_o, n155_neg, mux20_b10_sel_is_0_o);
  AL_MUX mux21_b12 (
    .i0(1'b0),
    .i1(n197[12]),
    .sel(mux21_b12_sel_is_2_o),
    .o(n202[12]));
  and mux21_b12_sel_is_2 (mux21_b12_sel_is_2_o, n155_neg, mux20_b12_sel_is_2_o);
  and mux21_b13_sel_is_2 (mux21_b13_sel_is_2_o, n155_neg, mux20_b13_sel_is_2_o);
  not mux21_b13_sel_is_2_o_inv (mux21_b13_sel_is_2_o_neg, mux21_b13_sel_is_2_o);
  AL_MUX mux21_b14 (
    .i0(1'b1),
    .i1(n199[14]),
    .sel(mux21_b11_sel_is_2_o),
    .o(n202[14]));
  binary_mux_s1_w1 mux21_b4 (
    .i0(n201[4]),
    .i1(1'b1),
    .sel(n155),
    .o(n202[4]));  // sources/rtl/camera_init.v(256)
  AL_MUX mux21_b6 (
    .i0(1'b1),
    .i1(n199[6]),
    .sel(mux21_b11_sel_is_2_o),
    .o(n202[6]));
  and mux21_b7_sel_is_2 (mux21_b7_sel_is_2_o, n155_neg, mux20_b7_sel_is_2_o);
  and mux21_b9_sel_is_2 (mux21_b9_sel_is_2_o, n155_neg, mux20_b9_sel_is_2_o);
  not mux21_b9_sel_is_2_o_inv (mux21_b9_sel_is_2_o_neg, mux21_b9_sel_is_2_o);
  binary_mux_s1_w1 mux22_b0 (
    .i0(n202[0]),
    .i1(1'b1),
    .sel(n154),
    .o(n203[0]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux22_b1 (
    .i0(n202[1]),
    .i1(1'b1),
    .sel(n154),
    .o(n203[1]));  // sources/rtl/camera_init.v(256)
  and mux22_b11_sel_is_2 (mux22_b11_sel_is_2_o, n154_neg, mux21_b11_sel_is_2_o);
  and mux22_b13_sel_is_0 (mux22_b13_sel_is_0_o, n154_neg, mux21_b13_sel_is_2_o_neg);
  and mux22_b15_sel_is_2 (mux22_b15_sel_is_2_o, n154_neg, mux21_b12_sel_is_2_o);
  and mux22_b2_sel_is_2 (mux22_b2_sel_is_2_o, n154_neg, mux21_b0_sel_is_0_o);
  AL_MUX mux22_b3 (
    .i0(1'b1),
    .i1(n201[3]),
    .sel(mux22_b3_sel_is_0_o),
    .o(n203[3]));
  and mux22_b3_sel_is_0 (mux22_b3_sel_is_0_o, n154_neg, n155_neg);
  binary_mux_s1_w1 mux22_b4 (
    .i0(n202[4]),
    .i1(1'b0),
    .sel(n154),
    .o(n203[4]));  // sources/rtl/camera_init.v(256)
  AL_MUX mux22_b7 (
    .i0(1'b0),
    .i1(n196[7]),
    .sel(mux22_b7_sel_is_2_o),
    .o(n203[7]));
  and mux22_b7_sel_is_2 (mux22_b7_sel_is_2_o, n154_neg, mux21_b7_sel_is_2_o);
  AL_MUX mux22_b8 (
    .i0(1'b0),
    .i1(n200[8]),
    .sel(mux22_b2_sel_is_2_o),
    .o(n203[8]));
  and mux22_b9_sel_is_0 (mux22_b9_sel_is_0_o, n154_neg, mux21_b9_sel_is_2_o_neg);
  not mux22_b9_sel_is_0_o_inv (mux22_b9_sel_is_0_o_neg, mux22_b9_sel_is_0_o);
  binary_mux_s1_w1 mux23_b0 (
    .i0(n203[0]),
    .i1(1'b0),
    .sel(n153),
    .o(n204[0]));  // sources/rtl/camera_init.v(256)
  and mux23_b10_sel_is_0 (mux23_b10_sel_is_0_o, n153_neg, n154_neg);
  and mux23_b11_sel_is_2 (mux23_b11_sel_is_2_o, n153_neg, mux22_b11_sel_is_2_o);
  and mux23_b13_sel_is_2 (mux23_b13_sel_is_2_o, n153_neg, mux22_b13_sel_is_0_o);
  and mux23_b15_sel_is_2 (mux23_b15_sel_is_2_o, n153_neg, mux22_b15_sel_is_2_o);
  and mux23_b2_sel_is_2 (mux23_b2_sel_is_2_o, n153_neg, mux22_b2_sel_is_2_o);
  binary_mux_s1_w1 mux23_b4 (
    .i0(n203[4]),
    .i1(1'b1),
    .sel(n153),
    .o(n204[4]));  // sources/rtl/camera_init.v(256)
  and mux23_b5_sel_is_2 (mux23_b5_sel_is_2_o, n153_neg, mux22_b3_sel_is_0_o);
  AL_MUX mux23_b6 (
    .i0(1'b0),
    .i1(n202[6]),
    .sel(mux23_b10_sel_is_0_o),
    .o(n204[6]));
  binary_mux_s1_w1 mux23_b8 (
    .i0(n203[8]),
    .i1(1'b1),
    .sel(n153),
    .o(n204[8]));  // sources/rtl/camera_init.v(256)
  and mux23_b9_sel_is_0 (mux23_b9_sel_is_0_o, n153_neg, mux22_b9_sel_is_0_o_neg);
  AL_MUX mux24_b1 (
    .i0(1'b0),
    .i1(n203[1]),
    .sel(mux24_b1_sel_is_0_o),
    .o(n205[1]));
  AL_MUX mux24_b10 (
    .i0(1'b0),
    .i1(n202[10]),
    .sel(mux24_b10_sel_is_2_o),
    .o(n205[10]));
  and mux24_b10_sel_is_2 (mux24_b10_sel_is_2_o, n152_neg, mux23_b10_sel_is_0_o);
  and mux24_b11_sel_is_2 (mux24_b11_sel_is_2_o, n152_neg, mux23_b11_sel_is_2_o);
  and mux24_b13_sel_is_2 (mux24_b13_sel_is_2_o, n152_neg, mux23_b13_sel_is_2_o);
  and mux24_b15_sel_is_2 (mux24_b15_sel_is_2_o, n152_neg, mux23_b15_sel_is_2_o);
  and mux24_b1_sel_is_0 (mux24_b1_sel_is_0_o, n152_neg, n153_neg);
  and mux24_b2_sel_is_2 (mux24_b2_sel_is_2_o, n152_neg, mux23_b2_sel_is_2_o);
  AL_MUX mux24_b3 (
    .i0(1'b0),
    .i1(n203[3]),
    .sel(mux24_b1_sel_is_0_o),
    .o(n205[3]));
  binary_mux_s1_w1 mux24_b4 (
    .i0(n204[4]),
    .i1(1'b0),
    .sel(n152),
    .o(n205[4]));  // sources/rtl/camera_init.v(256)
  AL_MUX mux24_b5 (
    .i0(1'b0),
    .i1(n201[5]),
    .sel(mux24_b5_sel_is_2_o),
    .o(n205[5]));
  and mux24_b5_sel_is_2 (mux24_b5_sel_is_2_o, n152_neg, mux23_b5_sel_is_2_o);
  binary_mux_s1_w1 mux24_b8 (
    .i0(n204[8]),
    .i1(1'b0),
    .sel(n152),
    .o(n205[8]));  // sources/rtl/camera_init.v(256)
  and mux24_b9_sel_is_2 (mux24_b9_sel_is_2_o, n152_neg, mux23_b9_sel_is_0_o);
  and mux25_b0_sel_is_0 (mux25_b0_sel_is_0_o, n151_neg, n152_neg);
  and mux25_b11_sel_is_2 (mux25_b11_sel_is_2_o, n151_neg, mux24_b11_sel_is_2_o);
  and mux25_b12_sel_is_2 (mux25_b12_sel_is_2_o, n151_neg, mux24_b10_sel_is_2_o);
  and mux25_b13_sel_is_2 (mux25_b13_sel_is_2_o, n151_neg, mux24_b13_sel_is_2_o);
  and mux25_b15_sel_is_2 (mux25_b15_sel_is_2_o, n151_neg, mux24_b15_sel_is_2_o);
  and mux25_b2_sel_is_2 (mux25_b2_sel_is_2_o, n151_neg, mux24_b2_sel_is_2_o);
  binary_mux_s1_w1 mux25_b3 (
    .i0(n205[3]),
    .i1(1'b1),
    .sel(n151),
    .o(n206[3]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux25_b5 (
    .i0(n205[5]),
    .i1(1'b1),
    .sel(n151),
    .o(n206[5]));  // sources/rtl/camera_init.v(256)
  AL_MUX mux25_b6 (
    .i0(1'b1),
    .i1(n204[6]),
    .sel(mux25_b0_sel_is_0_o),
    .o(n206[6]));
  and mux25_b7_sel_is_2 (mux25_b7_sel_is_2_o, n151_neg, mux24_b1_sel_is_0_o);
  binary_mux_s1_w1 mux25_b8 (
    .i0(n205[8]),
    .i1(1'b1),
    .sel(n151),
    .o(n206[8]));  // sources/rtl/camera_init.v(256)
  and mux25_b9_sel_is_2 (mux25_b9_sel_is_2_o, n151_neg, mux24_b9_sel_is_2_o);
  and mux26_b0_sel_is_2 (mux26_b0_sel_is_2_o, n150_neg, mux25_b0_sel_is_0_o);
  AL_MUX mux26_b10 (
    .i0(1'b1),
    .i1(n205[10]),
    .sel(mux26_b10_sel_is_0_o),
    .o(n207[10]));
  and mux26_b10_sel_is_0 (mux26_b10_sel_is_0_o, n150_neg, n151_neg);
  and mux26_b11_sel_is_2 (mux26_b11_sel_is_2_o, n150_neg, mux25_b11_sel_is_2_o);
  and mux26_b12_sel_is_2 (mux26_b12_sel_is_2_o, n150_neg, mux25_b12_sel_is_2_o);
  and mux26_b13_sel_is_2 (mux26_b13_sel_is_2_o, n150_neg, mux25_b13_sel_is_2_o);
  and mux26_b15_sel_is_2 (mux26_b15_sel_is_2_o, n150_neg, mux25_b15_sel_is_2_o);
  and mux26_b2_sel_is_2 (mux26_b2_sel_is_2_o, n150_neg, mux25_b2_sel_is_2_o);
  binary_mux_s1_w1 mux26_b3 (
    .i0(n206[3]),
    .i1(1'b0),
    .sel(n150),
    .o(n207[3]));  // sources/rtl/camera_init.v(256)
  AL_MUX mux26_b4 (
    .i0(1'b1),
    .i1(n205[4]),
    .sel(mux26_b10_sel_is_0_o),
    .o(n207[4]));
  binary_mux_s1_w1 mux26_b5 (
    .i0(n206[5]),
    .i1(1'b0),
    .sel(n150),
    .o(n207[5]));  // sources/rtl/camera_init.v(256)
  and mux26_b7_sel_is_2 (mux26_b7_sel_is_2_o, n150_neg, mux25_b7_sel_is_2_o);
  binary_mux_s1_w1 mux26_b8 (
    .i0(n206[8]),
    .i1(1'b0),
    .sel(n150),
    .o(n207[8]));  // sources/rtl/camera_init.v(256)
  and mux26_b9_sel_is_2 (mux26_b9_sel_is_2_o, n150_neg, mux25_b9_sel_is_2_o);
  not mux26_b9_sel_is_2_o_inv (mux26_b9_sel_is_2_o_neg, mux26_b9_sel_is_2_o);
  AL_MUX mux27_b0 (
    .i0(1'b1),
    .i1(n204[0]),
    .sel(mux27_b0_sel_is_2_o),
    .o(n208[0]));
  and mux27_b0_sel_is_2 (mux27_b0_sel_is_2_o, n149_neg, mux26_b0_sel_is_2_o);
  AL_MUX mux27_b1 (
    .i0(1'b1),
    .i1(n205[1]),
    .sel(mux27_b1_sel_is_2_o),
    .o(n208[1]));
  AL_MUX mux27_b11 (
    .i0(1'b0),
    .i1(n199[11]),
    .sel(mux27_b11_sel_is_2_o),
    .o(n208[11]));
  and mux27_b11_sel_is_2 (mux27_b11_sel_is_2_o, n149_neg, mux26_b11_sel_is_2_o);
  and mux27_b12_sel_is_2 (mux27_b12_sel_is_2_o, n149_neg, mux26_b12_sel_is_2_o);
  and mux27_b13_sel_is_2 (mux27_b13_sel_is_2_o, n149_neg, mux26_b13_sel_is_2_o);
  and mux27_b15_sel_is_2 (mux27_b15_sel_is_2_o, n149_neg, mux26_b15_sel_is_2_o);
  and mux27_b1_sel_is_2 (mux27_b1_sel_is_2_o, n149_neg, mux26_b10_sel_is_0_o);
  and mux27_b2_sel_is_2 (mux27_b2_sel_is_2_o, n149_neg, mux26_b2_sel_is_2_o);
  binary_mux_s1_w1 mux27_b4 (
    .i0(n207[4]),
    .i1(1'b0),
    .sel(n149),
    .o(n208[4]));  // sources/rtl/camera_init.v(256)
  AL_MUX mux27_b6 (
    .i0(1'b0),
    .i1(n206[6]),
    .sel(mux27_b6_sel_is_0_o),
    .o(n208[6]));
  and mux27_b6_sel_is_0 (mux27_b6_sel_is_0_o, n149_neg, n150_neg);
  AL_MUX mux27_b7 (
    .i0(1'b1),
    .i1(n203[7]),
    .sel(mux27_b7_sel_is_2_o),
    .o(n208[7]));
  and mux27_b7_sel_is_2 (mux27_b7_sel_is_2_o, n149_neg, mux26_b7_sel_is_2_o);
  and mux27_b9_sel_is_0 (mux27_b9_sel_is_0_o, n149_neg, mux26_b9_sel_is_2_o_neg);
  not mux27_b9_sel_is_0_o_inv (mux27_b9_sel_is_0_o_neg, mux27_b9_sel_is_0_o);
  AL_MUX mux28_b10 (
    .i0(1'b0),
    .i1(n207[10]),
    .sel(mux28_b10_sel_is_0_o),
    .o(n209[10]));
  and mux28_b10_sel_is_0 (mux28_b10_sel_is_0_o, n148_neg, n149_neg);
  binary_mux_s1_w1 mux28_b11 (
    .i0(n208[11]),
    .i1(1'b1),
    .sel(n148),
    .o(n209[11]));  // sources/rtl/camera_init.v(256)
  and mux28_b12_sel_is_2 (mux28_b12_sel_is_2_o, n148_neg, mux27_b12_sel_is_2_o);
  and mux28_b13_sel_is_2 (mux28_b13_sel_is_2_o, n148_neg, mux27_b13_sel_is_2_o);
  and mux28_b15_sel_is_2 (mux28_b15_sel_is_2_o, n148_neg, mux27_b15_sel_is_2_o);
  and mux28_b2_sel_is_2 (mux28_b2_sel_is_2_o, n148_neg, mux27_b2_sel_is_2_o);
  AL_MUX mux28_b3 (
    .i0(1'b1),
    .i1(n207[3]),
    .sel(mux28_b10_sel_is_0_o),
    .o(n209[3]));
  binary_mux_s1_w1 mux28_b4 (
    .i0(n208[4]),
    .i1(1'b1),
    .sel(n148),
    .o(n209[4]));  // sources/rtl/camera_init.v(256)
  and mux28_b9_sel_is_0 (mux28_b9_sel_is_0_o, n148_neg, mux27_b9_sel_is_0_o_neg);
  not mux28_b9_sel_is_0_o_inv (mux28_b9_sel_is_0_o_neg, mux28_b9_sel_is_0_o);
  AL_MUX mux29_b0 (
    .i0(1'b0),
    .i1(n208[0]),
    .sel(mux29_b0_sel_is_0_o),
    .o(n210[0]));
  and mux29_b0_sel_is_0 (mux29_b0_sel_is_0_o, n147_neg, n148_neg);
  binary_mux_s1_w1 mux29_b10 (
    .i0(n209[10]),
    .i1(1'b1),
    .sel(n147),
    .o(n210[10]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux29_b11 (
    .i0(n209[11]),
    .i1(1'b0),
    .sel(n147),
    .o(n210[11]));  // sources/rtl/camera_init.v(256)
  and mux29_b12_sel_is_2 (mux29_b12_sel_is_2_o, n147_neg, mux28_b12_sel_is_2_o);
  and mux29_b13_sel_is_2 (mux29_b13_sel_is_2_o, n147_neg, mux28_b13_sel_is_2_o);
  and mux29_b15_sel_is_2 (mux29_b15_sel_is_2_o, n147_neg, mux28_b15_sel_is_2_o);
  and mux29_b2_sel_is_2 (mux29_b2_sel_is_2_o, n147_neg, mux28_b2_sel_is_2_o);
  and mux29_b5_sel_is_2 (mux29_b5_sel_is_2_o, n147_neg, mux28_b10_sel_is_0_o);
  AL_MUX mux29_b6 (
    .i0(1'b1),
    .i1(n208[6]),
    .sel(mux29_b0_sel_is_0_o),
    .o(n210[6]));
  AL_MUX mux29_b7 (
    .i0(1'b0),
    .i1(n208[7]),
    .sel(mux29_b0_sel_is_0_o),
    .o(n210[7]));
  AL_MUX mux29_b8 (
    .i0(1'b1),
    .i1(n207[8]),
    .sel(mux29_b5_sel_is_2_o),
    .o(n210[8]));
  and mux29_b9_sel_is_0 (mux29_b9_sel_is_0_o, n147_neg, mux28_b9_sel_is_0_o_neg);
  not mux29_b9_sel_is_0_o_inv (mux29_b9_sel_is_0_o_neg, mux29_b9_sel_is_0_o);
  binary_mux_s1_w1 mux2_b0 (
    .i0(n182[0]),
    .i1(1'b1),
    .sel(n174),
    .o(n183[0]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux2_b10 (
    .i0(n182[10]),
    .i1(1'b0),
    .sel(n174),
    .o(n183[10]));  // sources/rtl/camera_init.v(256)
  and mux2_b11_sel_is_0 (mux2_b11_sel_is_0_o, n174_neg, n175_neg);
  binary_mux_s1_w1 mux2_b3 (
    .i0(n182[0]),
    .i1(1'b0),
    .sel(n174),
    .o(n183[3]));  // sources/rtl/camera_init.v(256)
  and mux2_b7_sel_is_2 (mux2_b7_sel_is_2_o, n174_neg, mux1_b7_sel_is_0_o);
  binary_mux_s1_w1 mux30_b0 (
    .i0(n210[0]),
    .i1(1'b1),
    .sel(n146),
    .o(n211[0]));  // sources/rtl/camera_init.v(256)
  AL_MUX mux30_b1 (
    .i0(1'b0),
    .i1(n208[1]),
    .sel(mux30_b1_sel_is_2_o),
    .o(n211[1]));
  binary_mux_s1_w1 mux30_b10 (
    .i0(n210[10]),
    .i1(1'b0),
    .sel(n146),
    .o(n211[10]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux30_b11 (
    .i0(n210[11]),
    .i1(1'b1),
    .sel(n146),
    .o(n211[11]));  // sources/rtl/camera_init.v(256)
  and mux30_b12_sel_is_2 (mux30_b12_sel_is_2_o, n146_neg, mux29_b12_sel_is_2_o);
  and mux30_b13_sel_is_2 (mux30_b13_sel_is_2_o, n146_neg, mux29_b13_sel_is_2_o);
  and mux30_b15_sel_is_2 (mux30_b15_sel_is_2_o, n146_neg, mux29_b15_sel_is_2_o);
  and mux30_b1_sel_is_2 (mux30_b1_sel_is_2_o, n146_neg, mux29_b0_sel_is_0_o);
  and mux30_b2_sel_is_2 (mux30_b2_sel_is_2_o, n146_neg, mux29_b2_sel_is_2_o);
  and mux30_b3_sel_is_0 (mux30_b3_sel_is_0_o, n146_neg, n147_neg);
  and mux30_b5_sel_is_2 (mux30_b5_sel_is_2_o, n146_neg, mux29_b5_sel_is_2_o);
  binary_mux_s1_w1 mux30_b6 (
    .i0(n210[6]),
    .i1(1'b0),
    .sel(n146),
    .o(n211[6]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux30_b7 (
    .i0(n210[7]),
    .i1(1'b1),
    .sel(n146),
    .o(n211[7]));  // sources/rtl/camera_init.v(256)
  and mux30_b9_sel_is_0 (mux30_b9_sel_is_0_o, n146_neg, mux29_b9_sel_is_0_o_neg);
  not mux30_b9_sel_is_0_o_inv (mux30_b9_sel_is_0_o_neg, mux30_b9_sel_is_0_o);
  binary_mux_s1_w1 mux31_b1 (
    .i0(n211[1]),
    .i1(1'b1),
    .sel(n145),
    .o(n212[1]));  // sources/rtl/camera_init.v(256)
  AL_MUX mux31_b12 (
    .i0(1'b1),
    .i1(n202[12]),
    .sel(mux31_b12_sel_is_2_o),
    .o(n212[12]));
  and mux31_b12_sel_is_2 (mux31_b12_sel_is_2_o, n145_neg, mux30_b12_sel_is_2_o);
  and mux31_b13_sel_is_2 (mux31_b13_sel_is_2_o, n145_neg, mux30_b13_sel_is_2_o);
  not mux31_b13_sel_is_2_o_inv (mux31_b13_sel_is_2_o_neg, mux31_b13_sel_is_2_o);
  AL_MUX mux31_b14 (
    .i0(1'b0),
    .i1(n202[14]),
    .sel(mux31_b12_sel_is_2_o),
    .o(n212[14]));
  and mux31_b15_sel_is_2 (mux31_b15_sel_is_2_o, n145_neg, mux30_b15_sel_is_2_o);
  AL_MUX mux31_b2 (
    .i0(1'b1),
    .i1(n200[2]),
    .sel(mux31_b2_sel_is_2_o),
    .o(n212[2]));
  and mux31_b2_sel_is_2 (mux31_b2_sel_is_2_o, n145_neg, mux30_b2_sel_is_2_o);
  and mux31_b3_sel_is_2 (mux31_b3_sel_is_2_o, n145_neg, mux30_b3_sel_is_0_o);
  AL_MUX mux31_b4 (
    .i0(1'b0),
    .i1(n209[4]),
    .sel(mux31_b3_sel_is_2_o),
    .o(n212[4]));
  AL_MUX mux31_b5 (
    .i0(1'b1),
    .i1(n207[5]),
    .sel(mux31_b5_sel_is_2_o),
    .o(n212[5]));
  and mux31_b5_sel_is_2 (mux31_b5_sel_is_2_o, n145_neg, mux30_b5_sel_is_2_o);
  binary_mux_s1_w1 mux31_b6 (
    .i0(n211[6]),
    .i1(1'b1),
    .sel(n145),
    .o(n212[6]));  // sources/rtl/camera_init.v(256)
  AL_MUX mux31_b8 (
    .i0(1'b0),
    .i1(n210[8]),
    .sel(mux31_b8_sel_is_0_o),
    .o(n212[8]));
  and mux31_b8_sel_is_0 (mux31_b8_sel_is_0_o, n145_neg, n146_neg);
  and mux31_b9_sel_is_0 (mux31_b9_sel_is_0_o, n145_neg, mux30_b9_sel_is_0_o_neg);
  and mux32_b0_sel_is_0 (mux32_b0_sel_is_0_o, n144_neg, n145_neg);
  AL_MUX mux32_b11 (
    .i0(1'b0),
    .i1(n211[11]),
    .sel(mux32_b0_sel_is_0_o),
    .o(n213[11]));
  binary_mux_s1_w1 mux32_b12 (
    .i0(n212[12]),
    .i1(1'b0),
    .sel(n144),
    .o(n213[12]));  // sources/rtl/camera_init.v(256)
  and mux32_b13_sel_is_0 (mux32_b13_sel_is_0_o, n144_neg, mux31_b13_sel_is_2_o_neg);
  not mux32_b13_sel_is_0_o_inv (mux32_b13_sel_is_0_o_neg, mux32_b13_sel_is_0_o);
  binary_mux_s1_w1 mux32_b14 (
    .i0(n212[14]),
    .i1(1'b1),
    .sel(n144),
    .o(n213[14]));  // sources/rtl/camera_init.v(256)
  and mux32_b15_sel_is_2 (mux32_b15_sel_is_2_o, n144_neg, mux31_b15_sel_is_2_o);
  and mux32_b3_sel_is_2 (mux32_b3_sel_is_2_o, n144_neg, mux31_b3_sel_is_2_o);
  binary_mux_s1_w1 mux32_b4 (
    .i0(n212[4]),
    .i1(1'b1),
    .sel(n144),
    .o(n213[4]));  // sources/rtl/camera_init.v(256)
  AL_MUX mux32_b7 (
    .i0(1'b0),
    .i1(n211[7]),
    .sel(mux32_b0_sel_is_0_o),
    .o(n213[7]));
  and mux32_b9_sel_is_2 (mux32_b9_sel_is_2_o, n144_neg, mux31_b9_sel_is_0_o);
  AL_MUX mux33_b0 (
    .i0(1'b0),
    .i1(n211[0]),
    .sel(mux33_b0_sel_is_2_o),
    .o(n214[0]));
  and mux33_b0_sel_is_2 (mux33_b0_sel_is_2_o, n143_neg, mux32_b0_sel_is_0_o);
  binary_mux_s1_w1 mux33_b11 (
    .i0(n213[11]),
    .i1(1'b1),
    .sel(n143),
    .o(n214[11]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux33_b12 (
    .i0(n213[12]),
    .i1(1'b1),
    .sel(n143),
    .o(n214[12]));  // sources/rtl/camera_init.v(256)
  and mux33_b13_sel_is_0 (mux33_b13_sel_is_0_o, n143_neg, mux32_b13_sel_is_0_o_neg);
  not mux33_b13_sel_is_0_o_inv (mux33_b13_sel_is_0_o_neg, mux33_b13_sel_is_0_o);
  binary_mux_s1_w1 mux33_b14 (
    .i0(n213[14]),
    .i1(1'b0),
    .sel(n143),
    .o(n214[14]));  // sources/rtl/camera_init.v(256)
  and mux33_b15_sel_is_2 (mux33_b15_sel_is_2_o, n143_neg, mux32_b15_sel_is_2_o);
  and mux33_b1_sel_is_0 (mux33_b1_sel_is_0_o, n143_neg, n144_neg);
  and mux33_b3_sel_is_2 (mux33_b3_sel_is_2_o, n143_neg, mux32_b3_sel_is_2_o);
  binary_mux_s1_w1 mux33_b4 (
    .i0(n213[4]),
    .i1(1'b0),
    .sel(n143),
    .o(n214[4]));  // sources/rtl/camera_init.v(256)
  AL_MUX mux33_b6 (
    .i0(1'b0),
    .i1(n212[6]),
    .sel(mux33_b1_sel_is_0_o),
    .o(n214[6]));
  binary_mux_s1_w1 mux33_b7 (
    .i0(n213[7]),
    .i1(1'b1),
    .sel(n143),
    .o(n214[7]));  // sources/rtl/camera_init.v(256)
  AL_MUX mux33_b8 (
    .i0(1'b1),
    .i1(n212[8]),
    .sel(mux33_b1_sel_is_0_o),
    .o(n214[8]));
  and mux33_b9_sel_is_2 (mux33_b9_sel_is_2_o, n143_neg, mux32_b9_sel_is_2_o);
  and mux34_b10_sel_is_2 (mux34_b10_sel_is_2_o, n142_neg, mux33_b0_sel_is_2_o);
  and mux34_b13_sel_is_0 (mux34_b13_sel_is_0_o, n142_neg, mux33_b13_sel_is_0_o_neg);
  and mux34_b15_sel_is_2 (mux34_b15_sel_is_2_o, n142_neg, mux33_b15_sel_is_2_o);
  and mux34_b1_sel_is_2 (mux34_b1_sel_is_2_o, n142_neg, mux33_b1_sel_is_0_o);
  and mux34_b3_sel_is_2 (mux34_b3_sel_is_2_o, n142_neg, mux33_b3_sel_is_2_o);
  binary_mux_s1_w1 mux34_b6 (
    .i0(n214[6]),
    .i1(1'b1),
    .sel(n142),
    .o(n215[6]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux34_b8 (
    .i0(n214[8]),
    .i1(1'b0),
    .sel(n142),
    .o(n215[8]));  // sources/rtl/camera_init.v(256)
  and mux34_b9_sel_is_2 (mux34_b9_sel_is_2_o, n142_neg, mux33_b9_sel_is_2_o);
  not mux34_b9_sel_is_2_o_inv (mux34_b9_sel_is_2_o_neg, mux34_b9_sel_is_2_o);
  AL_MUX mux35_b0 (
    .i0(1'b1),
    .i1(n214[0]),
    .sel(mux35_b0_sel_is_0_o),
    .o(n216[0]));
  and mux35_b0_sel_is_0 (mux35_b0_sel_is_0_o, n141_neg, n142_neg);
  AL_MUX mux35_b10 (
    .i0(1'b1),
    .i1(n211[10]),
    .sel(mux35_b10_sel_is_2_o),
    .o(n216[10]));
  and mux35_b10_sel_is_2 (mux35_b10_sel_is_2_o, n141_neg, mux34_b10_sel_is_2_o);
  AL_MUX mux35_b11 (
    .i0(1'b0),
    .i1(n214[11]),
    .sel(mux35_b0_sel_is_0_o),
    .o(n216[11]));
  and mux35_b13_sel_is_2 (mux35_b13_sel_is_2_o, n141_neg, mux34_b13_sel_is_0_o);
  not mux35_b13_sel_is_2_o_inv (mux35_b13_sel_is_2_o_neg, mux35_b13_sel_is_2_o);
  AL_MUX mux35_b14 (
    .i0(1'b1),
    .i1(n214[14]),
    .sel(mux35_b0_sel_is_0_o),
    .o(n216[14]));
  and mux35_b15_sel_is_2 (mux35_b15_sel_is_2_o, n141_neg, mux34_b15_sel_is_2_o);
  and mux35_b1_sel_is_2 (mux35_b1_sel_is_2_o, n141_neg, mux34_b1_sel_is_2_o);
  and mux35_b3_sel_is_2 (mux35_b3_sel_is_2_o, n141_neg, mux34_b3_sel_is_2_o);
  AL_MUX mux35_b4 (
    .i0(1'b1),
    .i1(n214[4]),
    .sel(mux35_b0_sel_is_0_o),
    .o(n216[4]));
  binary_mux_s1_w1 mux35_b8 (
    .i0(n215[8]),
    .i1(1'b1),
    .sel(n141),
    .o(n216[8]));  // sources/rtl/camera_init.v(256)
  and mux35_b9_sel_is_0 (mux35_b9_sel_is_0_o, n141_neg, mux34_b9_sel_is_2_o_neg);
  binary_mux_s1_w1 mux36_b10 (
    .i0(n216[10]),
    .i1(1'b0),
    .sel(n140),
    .o(n217[10]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux36_b11 (
    .i0(n216[11]),
    .i1(1'b1),
    .sel(n140),
    .o(n217[11]));  // sources/rtl/camera_init.v(256)
  and mux36_b12_sel_is_2 (mux36_b12_sel_is_2_o, n140_neg, mux35_b0_sel_is_0_o);
  and mux36_b13_sel_is_0 (mux36_b13_sel_is_0_o, n140_neg, mux35_b13_sel_is_2_o_neg);
  and mux36_b15_sel_is_2 (mux36_b15_sel_is_2_o, n140_neg, mux35_b15_sel_is_2_o);
  and mux36_b1_sel_is_2 (mux36_b1_sel_is_2_o, n140_neg, mux35_b1_sel_is_2_o);
  and mux36_b3_sel_is_2 (mux36_b3_sel_is_2_o, n140_neg, mux35_b3_sel_is_2_o);
  and mux36_b6_sel_is_0 (mux36_b6_sel_is_0_o, n140_neg, n141_neg);
  and mux36_b9_sel_is_2 (mux36_b9_sel_is_2_o, n140_neg, mux35_b9_sel_is_0_o);
  AL_MUX mux37_b0 (
    .i0(1'b0),
    .i1(n216[0]),
    .sel(mux37_b0_sel_is_0_o),
    .o(n218[0]));
  and mux37_b0_sel_is_0 (mux37_b0_sel_is_0_o, n139_neg, n140_neg);
  binary_mux_s1_w1 mux37_b10 (
    .i0(n217[10]),
    .i1(1'b1),
    .sel(n139),
    .o(n218[10]));  // sources/rtl/camera_init.v(256)
  and mux37_b12_sel_is_2 (mux37_b12_sel_is_2_o, n139_neg, mux36_b12_sel_is_2_o);
  and mux37_b13_sel_is_2 (mux37_b13_sel_is_2_o, n139_neg, mux36_b13_sel_is_0_o);
  not mux37_b13_sel_is_2_o_inv (mux37_b13_sel_is_2_o_neg, mux37_b13_sel_is_2_o);
  AL_MUX mux37_b14 (
    .i0(1'b0),
    .i1(n216[14]),
    .sel(mux37_b0_sel_is_0_o),
    .o(n218[14]));
  and mux37_b15_sel_is_2 (mux37_b15_sel_is_2_o, n139_neg, mux36_b15_sel_is_2_o);
  and mux37_b1_sel_is_2 (mux37_b1_sel_is_2_o, n139_neg, mux36_b1_sel_is_2_o);
  AL_MUX mux37_b2 (
    .i0(1'b0),
    .i1(n212[2]),
    .sel(mux37_b1_sel_is_2_o),
    .o(n218[2]));
  AL_MUX mux37_b3 (
    .i0(1'b0),
    .i1(n209[3]),
    .sel(mux37_b3_sel_is_2_o),
    .o(n218[3]));
  and mux37_b3_sel_is_2 (mux37_b3_sel_is_2_o, n139_neg, mux36_b3_sel_is_2_o);
  AL_MUX mux37_b5 (
    .i0(1'b0),
    .i1(n212[5]),
    .sel(mux37_b1_sel_is_2_o),
    .o(n218[5]));
  AL_MUX mux37_b6 (
    .i0(1'b0),
    .i1(n215[6]),
    .sel(mux37_b6_sel_is_2_o),
    .o(n218[6]));
  and mux37_b6_sel_is_2 (mux37_b6_sel_is_2_o, n139_neg, mux36_b6_sel_is_0_o);
  AL_MUX mux37_b7 (
    .i0(1'b0),
    .i1(n214[7]),
    .sel(mux37_b12_sel_is_2_o),
    .o(n218[7]));
  AL_MUX mux37_b8 (
    .i0(1'b0),
    .i1(n216[8]),
    .sel(mux37_b0_sel_is_0_o),
    .o(n218[8]));
  and mux37_b9_sel_is_2 (mux37_b9_sel_is_2_o, n139_neg, mux36_b9_sel_is_2_o);
  not mux37_b9_sel_is_2_o_inv (mux37_b9_sel_is_2_o_neg, mux37_b9_sel_is_2_o);
  binary_mux_s1_w1 mux38_b0 (
    .i0(n218[0]),
    .i1(1'b1),
    .sel(n138),
    .o(n219[0]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux38_b10 (
    .i0(n218[10]),
    .i1(1'b0),
    .sel(n138),
    .o(n219[10]));  // sources/rtl/camera_init.v(256)
  and mux38_b11_sel_is_0 (mux38_b11_sel_is_0_o, n138_neg, n139_neg);
  AL_MUX mux38_b12 (
    .i0(1'b0),
    .i1(n214[12]),
    .sel(mux38_b12_sel_is_2_o),
    .o(n219[12]));
  and mux38_b12_sel_is_2 (mux38_b12_sel_is_2_o, n138_neg, mux37_b12_sel_is_2_o);
  and mux38_b13_sel_is_0 (mux38_b13_sel_is_0_o, n138_neg, mux37_b13_sel_is_2_o_neg);
  binary_mux_s1_w1 mux38_b14 (
    .i0(n218[14]),
    .i1(1'b1),
    .sel(n138),
    .o(n219[14]));  // sources/rtl/camera_init.v(256)
  and mux38_b15_sel_is_2 (mux38_b15_sel_is_2_o, n138_neg, mux37_b15_sel_is_2_o);
  and mux38_b1_sel_is_2 (mux38_b1_sel_is_2_o, n138_neg, mux37_b1_sel_is_2_o);
  binary_mux_s1_w1 mux38_b2 (
    .i0(n218[2]),
    .i1(1'b1),
    .sel(n138),
    .o(n219[2]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux38_b3 (
    .i0(n218[3]),
    .i1(1'b1),
    .sel(n138),
    .o(n219[3]));  // sources/rtl/camera_init.v(256)
  and mux38_b4_sel_is_2 (mux38_b4_sel_is_2_o, n138_neg, mux37_b0_sel_is_0_o);
  binary_mux_s1_w1 mux38_b5 (
    .i0(n218[5]),
    .i1(1'b1),
    .sel(n138),
    .o(n219[5]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux38_b6 (
    .i0(n218[6]),
    .i1(1'b1),
    .sel(n138),
    .o(n219[6]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux38_b7 (
    .i0(n218[7]),
    .i1(1'b1),
    .sel(n138),
    .o(n219[7]));  // sources/rtl/camera_init.v(256)
  and mux38_b9_sel_is_0 (mux38_b9_sel_is_0_o, n138_neg, mux37_b9_sel_is_2_o_neg);
  and mux39_b11_sel_is_2 (mux39_b11_sel_is_2_o, n137_neg, mux38_b11_sel_is_0_o);
  and mux39_b13_sel_is_2 (mux39_b13_sel_is_2_o, n137_neg, mux38_b13_sel_is_0_o);
  and mux39_b15_sel_is_2 (mux39_b15_sel_is_2_o, n137_neg, mux38_b15_sel_is_2_o);
  and mux39_b1_sel_is_2 (mux39_b1_sel_is_2_o, n137_neg, mux38_b1_sel_is_2_o);
  and mux39_b4_sel_is_2 (mux39_b4_sel_is_2_o, n137_neg, mux38_b4_sel_is_2_o);
  and mux39_b8_sel_is_0 (mux39_b8_sel_is_0_o, n137_neg, n138_neg);
  and mux39_b9_sel_is_2 (mux39_b9_sel_is_2_o, n137_neg, mux38_b9_sel_is_0_o);
  binary_mux_s1_w1 mux3_b0 (
    .i0(n183[0]),
    .i1(1'b1),
    .sel(n173),
    .o(n184[0]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux3_b10 (
    .i0(n183[10]),
    .i1(1'b1),
    .sel(n173),
    .o(n184[10]));  // sources/rtl/camera_init.v(256)
  AL_MUX mux3_b11 (
    .i0(1'b0),
    .i1(n181[11]),
    .sel(mux3_b11_sel_is_2_o),
    .o(n184[11]));
  and mux3_b11_sel_is_2 (mux3_b11_sel_is_2_o, n173_neg, mux2_b11_sel_is_0_o);
  not mux3_b13_sel_is_2_o_inv (mux3_b13_sel_is_2_o_neg, mux3_b11_sel_is_2_o);
  binary_mux_s1_w1 mux3_b3 (
    .i0(n183[3]),
    .i1(1'b1),
    .sel(n173),
    .o(n184[3]));  // sources/rtl/camera_init.v(256)
  and mux3_b7_sel_is_2 (mux3_b7_sel_is_2_o, n173_neg, mux2_b7_sel_is_2_o);
  AL_MUX mux3_b8 (
    .i0(1'b1),
    .i1(n182[10]),
    .sel(mux3_b8_sel_is_0_o),
    .o(n184[8]));
  and mux3_b8_sel_is_0 (mux3_b8_sel_is_0_o, n173_neg, n174_neg);
  and mux40_b0_sel_is_0 (mux40_b0_sel_is_0_o, n136_neg, n137_neg);
  and mux40_b11_sel_is_2 (mux40_b11_sel_is_2_o, n136_neg, mux39_b11_sel_is_2_o);
  and mux40_b13_sel_is_2 (mux40_b13_sel_is_2_o, n136_neg, mux39_b13_sel_is_2_o);
  and mux40_b15_sel_is_2 (mux40_b15_sel_is_2_o, n136_neg, mux39_b15_sel_is_2_o);
  and mux40_b1_sel_is_2 (mux40_b1_sel_is_2_o, n136_neg, mux39_b1_sel_is_2_o);
  and mux40_b4_sel_is_2 (mux40_b4_sel_is_2_o, n136_neg, mux39_b4_sel_is_2_o);
  AL_MUX mux40_b7 (
    .i0(1'b0),
    .i1(n219[7]),
    .sel(mux40_b0_sel_is_0_o),
    .o(n221[7]));
  and mux40_b8_sel_is_2 (mux40_b8_sel_is_2_o, n136_neg, mux39_b8_sel_is_0_o);
  and mux40_b9_sel_is_2 (mux40_b9_sel_is_2_o, n136_neg, mux39_b9_sel_is_2_o);
  and mux41_b0_sel_is_2 (mux41_b0_sel_is_2_o, n135_neg, mux40_b0_sel_is_0_o);
  and mux41_b11_sel_is_2 (mux41_b11_sel_is_2_o, n135_neg, mux40_b11_sel_is_2_o);
  and mux41_b13_sel_is_2 (mux41_b13_sel_is_2_o, n135_neg, mux40_b13_sel_is_2_o);
  and mux41_b15_sel_is_2 (mux41_b15_sel_is_2_o, n135_neg, mux40_b15_sel_is_2_o);
  and mux41_b1_sel_is_2 (mux41_b1_sel_is_2_o, n135_neg, mux40_b1_sel_is_2_o);
  AL_MUX mux41_b3 (
    .i0(1'b0),
    .i1(n219[3]),
    .sel(mux41_b0_sel_is_2_o),
    .o(n222[3]));
  AL_MUX mux41_b4 (
    .i0(1'b0),
    .i1(n216[4]),
    .sel(mux41_b4_sel_is_2_o),
    .o(n222[4]));
  and mux41_b4_sel_is_2 (mux41_b4_sel_is_2_o, n135_neg, mux40_b4_sel_is_2_o);
  and mux41_b8_sel_is_2 (mux41_b8_sel_is_2_o, n135_neg, mux40_b8_sel_is_2_o);
  and mux41_b9_sel_is_2 (mux41_b9_sel_is_2_o, n135_neg, mux40_b9_sel_is_2_o);
  and mux42_b0_sel_is_2 (mux42_b0_sel_is_2_o, n134_neg, mux41_b0_sel_is_2_o);
  AL_MUX mux42_b1 (
    .i0(1'b0),
    .i1(n212[1]),
    .sel(mux42_b1_sel_is_2_o),
    .o(n223[1]));
  and mux42_b11_sel_is_2 (mux42_b11_sel_is_2_o, n134_neg, mux41_b11_sel_is_2_o);
  and mux42_b13_sel_is_2 (mux42_b13_sel_is_2_o, n134_neg, mux41_b13_sel_is_2_o);
  and mux42_b15_sel_is_2 (mux42_b15_sel_is_2_o, n134_neg, mux41_b15_sel_is_2_o);
  and mux42_b1_sel_is_2 (mux42_b1_sel_is_2_o, n134_neg, mux41_b1_sel_is_2_o);
  binary_mux_s1_w1 mux42_b3 (
    .i0(n222[3]),
    .i1(1'b1),
    .sel(n134),
    .o(n223[3]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux42_b4 (
    .i0(n222[4]),
    .i1(1'b1),
    .sel(n134),
    .o(n223[4]));  // sources/rtl/camera_init.v(256)
  AL_MUX mux42_b7 (
    .i0(1'b1),
    .i1(n221[7]),
    .sel(mux42_b7_sel_is_0_o),
    .o(n223[7]));
  and mux42_b7_sel_is_0 (mux42_b7_sel_is_0_o, n134_neg, n135_neg);
  and mux42_b8_sel_is_2 (mux42_b8_sel_is_2_o, n134_neg, mux41_b8_sel_is_2_o);
  and mux42_b9_sel_is_2 (mux42_b9_sel_is_2_o, n134_neg, mux41_b9_sel_is_2_o);
  and mux43_b0_sel_is_2 (mux43_b0_sel_is_2_o, n133_neg, mux42_b0_sel_is_2_o);
  and mux43_b11_sel_is_2 (mux43_b11_sel_is_2_o, n133_neg, mux42_b11_sel_is_2_o);
  and mux43_b13_sel_is_2 (mux43_b13_sel_is_2_o, n133_neg, mux42_b13_sel_is_2_o);
  and mux43_b15_sel_is_2 (mux43_b15_sel_is_2_o, n133_neg, mux42_b15_sel_is_2_o);
  AL_MUX mux43_b2 (
    .i0(1'b0),
    .i1(n219[2]),
    .sel(mux43_b0_sel_is_2_o),
    .o(n224[2]));
  AL_MUX mux43_b5 (
    .i0(1'b0),
    .i1(n219[5]),
    .sel(mux43_b0_sel_is_2_o),
    .o(n224[5]));
  and mux43_b8_sel_is_2 (mux43_b8_sel_is_2_o, n133_neg, mux42_b8_sel_is_2_o);
  and mux43_b9_sel_is_2 (mux43_b9_sel_is_2_o, n133_neg, mux42_b9_sel_is_2_o);
  and mux44_b0_sel_is_2 (mux44_b0_sel_is_2_o, n132_neg, mux43_b0_sel_is_2_o);
  AL_MUX mux44_b1 (
    .i0(1'b1),
    .i1(n223[1]),
    .sel(mux44_b1_sel_is_0_o),
    .o(n225[1]));
  and mux44_b11_sel_is_2 (mux44_b11_sel_is_2_o, n132_neg, mux43_b11_sel_is_2_o);
  and mux44_b13_sel_is_2 (mux44_b13_sel_is_2_o, n132_neg, mux43_b13_sel_is_2_o);
  and mux44_b15_sel_is_2 (mux44_b15_sel_is_2_o, n132_neg, mux43_b15_sel_is_2_o);
  and mux44_b1_sel_is_0 (mux44_b1_sel_is_0_o, n132_neg, n133_neg);
  binary_mux_s1_w1 mux44_b2 (
    .i0(n224[2]),
    .i1(1'b1),
    .sel(n132),
    .o(n225[2]));  // sources/rtl/camera_init.v(256)
  AL_MUX mux44_b3 (
    .i0(1'b0),
    .i1(n223[3]),
    .sel(mux44_b1_sel_is_0_o),
    .o(n225[3]));
  and mux44_b8_sel_is_2 (mux44_b8_sel_is_2_o, n132_neg, mux43_b8_sel_is_2_o);
  and mux44_b9_sel_is_2 (mux44_b9_sel_is_2_o, n132_neg, mux43_b9_sel_is_2_o);
  and mux45_b0_sel_is_2 (mux45_b0_sel_is_2_o, n131_neg, mux44_b0_sel_is_2_o);
  and mux45_b11_sel_is_2 (mux45_b11_sel_is_2_o, n131_neg, mux44_b11_sel_is_2_o);
  and mux45_b13_sel_is_2 (mux45_b13_sel_is_2_o, n131_neg, mux44_b13_sel_is_2_o);
  and mux45_b15_sel_is_2 (mux45_b15_sel_is_2_o, n131_neg, mux44_b15_sel_is_2_o);
  binary_mux_s1_w1 mux45_b3 (
    .i0(n225[3]),
    .i1(1'b1),
    .sel(n131),
    .o(n226[3]));  // sources/rtl/camera_init.v(256)
  AL_MUX mux45_b4 (
    .i0(1'b0),
    .i1(n223[4]),
    .sel(mux45_b4_sel_is_2_o),
    .o(n226[4]));
  and mux45_b4_sel_is_2 (mux45_b4_sel_is_2_o, n131_neg, mux44_b1_sel_is_0_o);
  and mux45_b5_sel_is_0 (mux45_b5_sel_is_0_o, n131_neg, n132_neg);
  and mux45_b8_sel_is_2 (mux45_b8_sel_is_2_o, n131_neg, mux44_b8_sel_is_2_o);
  and mux45_b9_sel_is_2 (mux45_b9_sel_is_2_o, n131_neg, mux44_b9_sel_is_2_o);
  and mux46_b0_sel_is_2 (mux46_b0_sel_is_2_o, n130_neg, mux45_b0_sel_is_2_o);
  and mux46_b11_sel_is_2 (mux46_b11_sel_is_2_o, n130_neg, mux45_b11_sel_is_2_o);
  and mux46_b13_sel_is_2 (mux46_b13_sel_is_2_o, n130_neg, mux45_b13_sel_is_2_o);
  and mux46_b15_sel_is_2 (mux46_b15_sel_is_2_o, n130_neg, mux45_b15_sel_is_2_o);
  and mux46_b1_sel_is_0 (mux46_b1_sel_is_0_o, n130_neg, n131_neg);
  AL_MUX mux46_b2 (
    .i0(1'b0),
    .i1(n225[2]),
    .sel(mux46_b1_sel_is_0_o),
    .o(n227[2]));
  binary_mux_s1_w1 mux46_b4 (
    .i0(n226[4]),
    .i1(1'b1),
    .sel(n130),
    .o(n227[4]));  // sources/rtl/camera_init.v(256)
  and mux46_b5_sel_is_2 (mux46_b5_sel_is_2_o, n130_neg, mux45_b5_sel_is_0_o);
  and mux46_b7_sel_is_2 (mux46_b7_sel_is_2_o, n130_neg, mux45_b4_sel_is_2_o);
  and mux46_b8_sel_is_2 (mux46_b8_sel_is_2_o, n130_neg, mux45_b8_sel_is_2_o);
  and mux46_b9_sel_is_2 (mux46_b9_sel_is_2_o, n130_neg, mux45_b9_sel_is_2_o);
  and mux47_b0_sel_is_2 (mux47_b0_sel_is_2_o, n129_neg, mux46_b0_sel_is_2_o);
  and mux47_b11_sel_is_2 (mux47_b11_sel_is_2_o, n129_neg, mux46_b11_sel_is_2_o);
  and mux47_b13_sel_is_2 (mux47_b13_sel_is_2_o, n129_neg, mux46_b13_sel_is_2_o);
  and mux47_b15_sel_is_2 (mux47_b15_sel_is_2_o, n129_neg, mux46_b15_sel_is_2_o);
  and mux47_b1_sel_is_2 (mux47_b1_sel_is_2_o, n129_neg, mux46_b1_sel_is_0_o);
  AL_MUX mux47_b3 (
    .i0(1'b0),
    .i1(n226[3]),
    .sel(mux47_b3_sel_is_0_o),
    .o(n228[3]));
  and mux47_b3_sel_is_0 (mux47_b3_sel_is_0_o, n129_neg, n130_neg);
  AL_MUX mux47_b5 (
    .i0(1'b1),
    .i1(n224[5]),
    .sel(mux47_b5_sel_is_2_o),
    .o(n228[5]));
  and mux47_b5_sel_is_2 (mux47_b5_sel_is_2_o, n129_neg, mux46_b5_sel_is_2_o);
  and mux47_b7_sel_is_2 (mux47_b7_sel_is_2_o, n129_neg, mux46_b7_sel_is_2_o);
  and mux47_b8_sel_is_2 (mux47_b8_sel_is_2_o, n129_neg, mux46_b8_sel_is_2_o);
  and mux47_b9_sel_is_2 (mux47_b9_sel_is_2_o, n129_neg, mux46_b9_sel_is_2_o);
  and mux48_b0_sel_is_2 (mux48_b0_sel_is_2_o, n128_neg, mux47_b0_sel_is_2_o);
  AL_MUX mux48_b1 (
    .i0(1'b0),
    .i1(n225[1]),
    .sel(mux48_b1_sel_is_2_o),
    .o(n229[1]));
  and mux48_b11_sel_is_2 (mux48_b11_sel_is_2_o, n128_neg, mux47_b11_sel_is_2_o);
  and mux48_b13_sel_is_2 (mux48_b13_sel_is_2_o, n128_neg, mux47_b13_sel_is_2_o);
  and mux48_b15_sel_is_2 (mux48_b15_sel_is_2_o, n128_neg, mux47_b15_sel_is_2_o);
  and mux48_b1_sel_is_2 (mux48_b1_sel_is_2_o, n128_neg, mux47_b1_sel_is_2_o);
  AL_MUX mux48_b2 (
    .i0(1'b1),
    .i1(n227[2]),
    .sel(mux48_b2_sel_is_0_o),
    .o(n229[2]));
  and mux48_b2_sel_is_0 (mux48_b2_sel_is_0_o, n128_neg, n129_neg);
  binary_mux_s1_w1 mux48_b3 (
    .i0(n228[3]),
    .i1(1'b1),
    .sel(n128),
    .o(n229[3]));  // sources/rtl/camera_init.v(256)
  and mux48_b7_sel_is_2 (mux48_b7_sel_is_2_o, n128_neg, mux47_b7_sel_is_2_o);
  and mux48_b8_sel_is_2 (mux48_b8_sel_is_2_o, n128_neg, mux47_b8_sel_is_2_o);
  and mux48_b9_sel_is_2 (mux48_b9_sel_is_2_o, n128_neg, mux47_b9_sel_is_2_o);
  AL_MUX mux49_b0 (
    .i0(1'b0),
    .i1(n219[0]),
    .sel(mux49_b0_sel_is_2_o),
    .o(n230[0]));
  and mux49_b0_sel_is_2 (mux49_b0_sel_is_2_o, n127_neg, mux48_b0_sel_is_2_o);
  binary_mux_s1_w1 mux49_b1 (
    .i0(n229[1]),
    .i1(1'b1),
    .sel(n127),
    .o(n230[1]));  // sources/rtl/camera_init.v(256)
  and mux49_b11_sel_is_2 (mux49_b11_sel_is_2_o, n127_neg, mux48_b11_sel_is_2_o);
  and mux49_b13_sel_is_2 (mux49_b13_sel_is_2_o, n127_neg, mux48_b13_sel_is_2_o);
  and mux49_b15_sel_is_2 (mux49_b15_sel_is_2_o, n127_neg, mux48_b15_sel_is_2_o);
  binary_mux_s1_w1 mux49_b3 (
    .i0(n229[3]),
    .i1(1'b0),
    .sel(n127),
    .o(n230[3]));  // sources/rtl/camera_init.v(256)
  AL_MUX mux49_b4 (
    .i0(1'b0),
    .i1(n227[4]),
    .sel(mux49_b4_sel_is_2_o),
    .o(n230[4]));
  and mux49_b4_sel_is_2 (mux49_b4_sel_is_2_o, n127_neg, mux48_b2_sel_is_0_o);
  and mux49_b5_sel_is_0 (mux49_b5_sel_is_0_o, n127_neg, n128_neg);
  and mux49_b7_sel_is_2 (mux49_b7_sel_is_2_o, n127_neg, mux48_b7_sel_is_2_o);
  and mux49_b8_sel_is_2 (mux49_b8_sel_is_2_o, n127_neg, mux48_b8_sel_is_2_o);
  and mux49_b9_sel_is_2 (mux49_b9_sel_is_2_o, n127_neg, mux48_b9_sel_is_2_o);
  binary_mux_s1_w1 mux4_b10 (
    .i0(n184[10]),
    .i1(1'b0),
    .sel(n172),
    .o(n185[10]));  // sources/rtl/camera_init.v(256)
  and mux4_b13_sel_is_0 (mux4_b13_sel_is_0_o, n172_neg, mux3_b13_sel_is_2_o_neg);
  not mux4_b13_sel_is_0_o_inv (mux4_b13_sel_is_0_o_neg, mux4_b13_sel_is_0_o);
  AL_MUX mux4_b14 (
    .i0(1'b1),
    .i1(n181[11]),
    .sel(mux4_b14_sel_is_2_o),
    .o(n185[14]));
  and mux4_b14_sel_is_2 (mux4_b14_sel_is_2_o, n172_neg, mux3_b11_sel_is_2_o);
  binary_mux_s1_w1 mux4_b3 (
    .i0(n184[3]),
    .i1(1'b1),
    .sel(n172),
    .o(n185[3]));  // sources/rtl/camera_init.v(256)
  and mux4_b5_sel_is_0 (mux4_b5_sel_is_0_o, n172_neg, n173_neg);
  and mux4_b7_sel_is_2 (mux4_b7_sel_is_2_o, n172_neg, mux3_b7_sel_is_2_o);
  binary_mux_s1_w1 mux4_b8 (
    .i0(n184[8]),
    .i1(1'b0),
    .sel(n172),
    .o(n185[8]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux50_b0 (
    .i0(n230[0]),
    .i1(1'b1),
    .sel(n126),
    .o(n231[0]));  // sources/rtl/camera_init.v(256)
  and mux50_b10_sel_is_2 (mux50_b10_sel_is_2_o, n126_neg, mux49_b0_sel_is_2_o);
  and mux50_b11_sel_is_2 (mux50_b11_sel_is_2_o, n126_neg, mux49_b11_sel_is_2_o);
  and mux50_b13_sel_is_2 (mux50_b13_sel_is_2_o, n126_neg, mux49_b13_sel_is_2_o);
  and mux50_b15_sel_is_2 (mux50_b15_sel_is_2_o, n126_neg, mux49_b15_sel_is_2_o);
  and mux50_b2_sel_is_0 (mux50_b2_sel_is_0_o, n126_neg, n127_neg);
  binary_mux_s1_w1 mux50_b4 (
    .i0(n230[4]),
    .i1(1'b1),
    .sel(n126),
    .o(n231[4]));  // sources/rtl/camera_init.v(256)
  and mux50_b5_sel_is_2 (mux50_b5_sel_is_2_o, n126_neg, mux49_b5_sel_is_0_o);
  and mux50_b7_sel_is_2 (mux50_b7_sel_is_2_o, n126_neg, mux49_b7_sel_is_2_o);
  and mux50_b8_sel_is_2 (mux50_b8_sel_is_2_o, n126_neg, mux49_b8_sel_is_2_o);
  and mux50_b9_sel_is_2 (mux50_b9_sel_is_2_o, n126_neg, mux49_b9_sel_is_2_o);
  and mux51_b10_sel_is_2 (mux51_b10_sel_is_2_o, n125_neg, mux50_b10_sel_is_2_o);
  and mux51_b11_sel_is_2 (mux51_b11_sel_is_2_o, n125_neg, mux50_b11_sel_is_2_o);
  and mux51_b13_sel_is_2 (mux51_b13_sel_is_2_o, n125_neg, mux50_b13_sel_is_2_o);
  and mux51_b15_sel_is_2 (mux51_b15_sel_is_2_o, n125_neg, mux50_b15_sel_is_2_o);
  and mux51_b1_sel_is_0 (mux51_b1_sel_is_0_o, n125_neg, n126_neg);
  and mux51_b2_sel_is_2 (mux51_b2_sel_is_2_o, n125_neg, mux50_b2_sel_is_0_o);
  AL_MUX mux51_b3 (
    .i0(1'b1),
    .i1(n230[3]),
    .sel(mux51_b1_sel_is_0_o),
    .o(n232[3]));
  and mux51_b5_sel_is_2 (mux51_b5_sel_is_2_o, n125_neg, mux50_b5_sel_is_2_o);
  and mux51_b7_sel_is_2 (mux51_b7_sel_is_2_o, n125_neg, mux50_b7_sel_is_2_o);
  AL_MUX mux51_b8 (
    .i0(1'b1),
    .i1(n218[8]),
    .sel(mux51_b8_sel_is_2_o),
    .o(n232[8]));
  and mux51_b8_sel_is_2 (mux51_b8_sel_is_2_o, n125_neg, mux50_b8_sel_is_2_o);
  and mux51_b9_sel_is_2 (mux51_b9_sel_is_2_o, n125_neg, mux50_b9_sel_is_2_o);
  and mux52_b0_sel_is_0 (mux52_b0_sel_is_0_o, n124_neg, n125_neg);
  AL_MUX mux52_b10 (
    .i0(1'b1),
    .i1(n219[10]),
    .sel(mux52_b10_sel_is_2_o),
    .o(n233[10]));
  and mux52_b10_sel_is_2 (mux52_b10_sel_is_2_o, n124_neg, mux51_b10_sel_is_2_o);
  and mux52_b11_sel_is_2 (mux52_b11_sel_is_2_o, n124_neg, mux51_b11_sel_is_2_o);
  and mux52_b13_sel_is_2 (mux52_b13_sel_is_2_o, n124_neg, mux51_b13_sel_is_2_o);
  and mux52_b15_sel_is_2 (mux52_b15_sel_is_2_o, n124_neg, mux51_b15_sel_is_2_o);
  and mux52_b1_sel_is_2 (mux52_b1_sel_is_2_o, n124_neg, mux51_b1_sel_is_0_o);
  and mux52_b2_sel_is_2 (mux52_b2_sel_is_2_o, n124_neg, mux51_b2_sel_is_2_o);
  and mux52_b5_sel_is_2 (mux52_b5_sel_is_2_o, n124_neg, mux51_b5_sel_is_2_o);
  and mux52_b7_sel_is_2 (mux52_b7_sel_is_2_o, n124_neg, mux51_b7_sel_is_2_o);
  binary_mux_s1_w1 mux52_b8 (
    .i0(n232[8]),
    .i1(1'b0),
    .sel(n124),
    .o(n233[8]));  // sources/rtl/camera_init.v(256)
  and mux52_b9_sel_is_2 (mux52_b9_sel_is_2_o, n124_neg, mux51_b9_sel_is_2_o);
  and mux53_b0_sel_is_2 (mux53_b0_sel_is_2_o, n123_neg, mux52_b0_sel_is_0_o);
  and mux53_b11_sel_is_2 (mux53_b11_sel_is_2_o, n123_neg, mux52_b11_sel_is_2_o);
  and mux53_b12_sel_is_2 (mux53_b12_sel_is_2_o, n123_neg, mux52_b10_sel_is_2_o);
  and mux53_b13_sel_is_2 (mux53_b13_sel_is_2_o, n123_neg, mux52_b13_sel_is_2_o);
  and mux53_b15_sel_is_2 (mux53_b15_sel_is_2_o, n123_neg, mux52_b15_sel_is_2_o);
  and mux53_b1_sel_is_2 (mux53_b1_sel_is_2_o, n123_neg, mux52_b1_sel_is_2_o);
  and mux53_b2_sel_is_2 (mux53_b2_sel_is_2_o, n123_neg, mux52_b2_sel_is_2_o);
  and mux53_b3_sel_is_0 (mux53_b3_sel_is_0_o, n123_neg, n124_neg);
  and mux53_b5_sel_is_2 (mux53_b5_sel_is_2_o, n123_neg, mux52_b5_sel_is_2_o);
  and mux53_b7_sel_is_2 (mux53_b7_sel_is_2_o, n123_neg, mux52_b7_sel_is_2_o);
  and mux53_b9_sel_is_2 (mux53_b9_sel_is_2_o, n123_neg, mux52_b9_sel_is_2_o);
  and mux54_b0_sel_is_2 (mux54_b0_sel_is_2_o, n122_neg, mux53_b0_sel_is_2_o);
  and mux54_b10_sel_is_0 (mux54_b10_sel_is_0_o, n122_neg, n123_neg);
  and mux54_b11_sel_is_2 (mux54_b11_sel_is_2_o, n122_neg, mux53_b11_sel_is_2_o);
  and mux54_b12_sel_is_2 (mux54_b12_sel_is_2_o, n122_neg, mux53_b12_sel_is_2_o);
  and mux54_b13_sel_is_2 (mux54_b13_sel_is_2_o, n122_neg, mux53_b13_sel_is_2_o);
  and mux54_b15_sel_is_2 (mux54_b15_sel_is_2_o, n122_neg, mux53_b15_sel_is_2_o);
  and mux54_b1_sel_is_2 (mux54_b1_sel_is_2_o, n122_neg, mux53_b1_sel_is_2_o);
  and mux54_b2_sel_is_2 (mux54_b2_sel_is_2_o, n122_neg, mux53_b2_sel_is_2_o);
  and mux54_b3_sel_is_2 (mux54_b3_sel_is_2_o, n122_neg, mux53_b3_sel_is_0_o);
  and mux54_b5_sel_is_2 (mux54_b5_sel_is_2_o, n122_neg, mux53_b5_sel_is_2_o);
  and mux54_b7_sel_is_2 (mux54_b7_sel_is_2_o, n122_neg, mux53_b7_sel_is_2_o);
  and mux54_b9_sel_is_2 (mux54_b9_sel_is_2_o, n122_neg, mux53_b9_sel_is_2_o);
  and mux55_b0_sel_is_2 (mux55_b0_sel_is_2_o, n121_neg, mux54_b0_sel_is_2_o);
  and mux55_b10_sel_is_2 (mux55_b10_sel_is_2_o, n121_neg, mux54_b10_sel_is_0_o);
  and mux55_b11_sel_is_2 (mux55_b11_sel_is_2_o, n121_neg, mux54_b11_sel_is_2_o);
  and mux55_b12_sel_is_2 (mux55_b12_sel_is_2_o, n121_neg, mux54_b12_sel_is_2_o);
  and mux55_b13_sel_is_2 (mux55_b13_sel_is_2_o, n121_neg, mux54_b13_sel_is_2_o);
  and mux55_b15_sel_is_2 (mux55_b15_sel_is_2_o, n121_neg, mux54_b15_sel_is_2_o);
  and mux55_b1_sel_is_2 (mux55_b1_sel_is_2_o, n121_neg, mux54_b1_sel_is_2_o);
  and mux55_b2_sel_is_2 (mux55_b2_sel_is_2_o, n121_neg, mux54_b2_sel_is_2_o);
  and mux55_b3_sel_is_2 (mux55_b3_sel_is_2_o, n121_neg, mux54_b3_sel_is_2_o);
  and mux55_b5_sel_is_2 (mux55_b5_sel_is_2_o, n121_neg, mux54_b5_sel_is_2_o);
  and mux55_b7_sel_is_2 (mux55_b7_sel_is_2_o, n121_neg, mux54_b7_sel_is_2_o);
  and mux55_b9_sel_is_2 (mux55_b9_sel_is_2_o, n121_neg, mux54_b9_sel_is_2_o);
  and mux56_b0_sel_is_2 (mux56_b0_sel_is_2_o, n120_neg, mux55_b0_sel_is_2_o);
  and mux56_b10_sel_is_2 (mux56_b10_sel_is_2_o, n120_neg, mux55_b10_sel_is_2_o);
  and mux56_b11_sel_is_2 (mux56_b11_sel_is_2_o, n120_neg, mux55_b11_sel_is_2_o);
  and mux56_b12_sel_is_2 (mux56_b12_sel_is_2_o, n120_neg, mux55_b12_sel_is_2_o);
  and mux56_b13_sel_is_2 (mux56_b13_sel_is_2_o, n120_neg, mux55_b13_sel_is_2_o);
  and mux56_b15_sel_is_2 (mux56_b15_sel_is_2_o, n120_neg, mux55_b15_sel_is_2_o);
  and mux56_b1_sel_is_2 (mux56_b1_sel_is_2_o, n120_neg, mux55_b1_sel_is_2_o);
  and mux56_b2_sel_is_2 (mux56_b2_sel_is_2_o, n120_neg, mux55_b2_sel_is_2_o);
  and mux56_b3_sel_is_2 (mux56_b3_sel_is_2_o, n120_neg, mux55_b3_sel_is_2_o);
  and mux56_b5_sel_is_2 (mux56_b5_sel_is_2_o, n120_neg, mux55_b5_sel_is_2_o);
  and mux56_b7_sel_is_2 (mux56_b7_sel_is_2_o, n120_neg, mux55_b7_sel_is_2_o);
  and mux56_b9_sel_is_2 (mux56_b9_sel_is_2_o, n120_neg, mux55_b9_sel_is_2_o);
  and mux57_b0_sel_is_2 (mux57_b0_sel_is_2_o, n119_neg, mux56_b0_sel_is_2_o);
  and mux57_b10_sel_is_2 (mux57_b10_sel_is_2_o, n119_neg, mux56_b10_sel_is_2_o);
  and mux57_b11_sel_is_2 (mux57_b11_sel_is_2_o, n119_neg, mux56_b11_sel_is_2_o);
  and mux57_b12_sel_is_2 (mux57_b12_sel_is_2_o, n119_neg, mux56_b12_sel_is_2_o);
  and mux57_b13_sel_is_2 (mux57_b13_sel_is_2_o, n119_neg, mux56_b13_sel_is_2_o);
  and mux57_b15_sel_is_2 (mux57_b15_sel_is_2_o, n119_neg, mux56_b15_sel_is_2_o);
  and mux57_b1_sel_is_2 (mux57_b1_sel_is_2_o, n119_neg, mux56_b1_sel_is_2_o);
  and mux57_b2_sel_is_2 (mux57_b2_sel_is_2_o, n119_neg, mux56_b2_sel_is_2_o);
  and mux57_b3_sel_is_2 (mux57_b3_sel_is_2_o, n119_neg, mux56_b3_sel_is_2_o);
  and mux57_b5_sel_is_2 (mux57_b5_sel_is_2_o, n119_neg, mux56_b5_sel_is_2_o);
  and mux57_b7_sel_is_2 (mux57_b7_sel_is_2_o, n119_neg, mux56_b7_sel_is_2_o);
  and mux57_b9_sel_is_2 (mux57_b9_sel_is_2_o, n119_neg, mux56_b9_sel_is_2_o);
  and mux58_b0_sel_is_2 (mux58_b0_sel_is_2_o, n118_neg, mux57_b0_sel_is_2_o);
  and mux58_b10_sel_is_2 (mux58_b10_sel_is_2_o, n118_neg, mux57_b10_sel_is_2_o);
  and mux58_b11_sel_is_2 (mux58_b11_sel_is_2_o, n118_neg, mux57_b11_sel_is_2_o);
  and mux58_b12_sel_is_2 (mux58_b12_sel_is_2_o, n118_neg, mux57_b12_sel_is_2_o);
  and mux58_b13_sel_is_2 (mux58_b13_sel_is_2_o, n118_neg, mux57_b13_sel_is_2_o);
  and mux58_b15_sel_is_2 (mux58_b15_sel_is_2_o, n118_neg, mux57_b15_sel_is_2_o);
  and mux58_b1_sel_is_2 (mux58_b1_sel_is_2_o, n118_neg, mux57_b1_sel_is_2_o);
  and mux58_b2_sel_is_2 (mux58_b2_sel_is_2_o, n118_neg, mux57_b2_sel_is_2_o);
  and mux58_b3_sel_is_2 (mux58_b3_sel_is_2_o, n118_neg, mux57_b3_sel_is_2_o);
  and mux58_b5_sel_is_2 (mux58_b5_sel_is_2_o, n118_neg, mux57_b5_sel_is_2_o);
  and mux58_b7_sel_is_2 (mux58_b7_sel_is_2_o, n118_neg, mux57_b7_sel_is_2_o);
  and mux58_b9_sel_is_2 (mux58_b9_sel_is_2_o, n118_neg, mux57_b9_sel_is_2_o);
  and mux59_b0_sel_is_2 (mux59_b0_sel_is_2_o, n117_neg, mux58_b0_sel_is_2_o);
  and mux59_b10_sel_is_2 (mux59_b10_sel_is_2_o, n117_neg, mux58_b10_sel_is_2_o);
  and mux59_b11_sel_is_2 (mux59_b11_sel_is_2_o, n117_neg, mux58_b11_sel_is_2_o);
  and mux59_b12_sel_is_2 (mux59_b12_sel_is_2_o, n117_neg, mux58_b12_sel_is_2_o);
  and mux59_b13_sel_is_2 (mux59_b13_sel_is_2_o, n117_neg, mux58_b13_sel_is_2_o);
  and mux59_b15_sel_is_2 (mux59_b15_sel_is_2_o, n117_neg, mux58_b15_sel_is_2_o);
  and mux59_b1_sel_is_2 (mux59_b1_sel_is_2_o, n117_neg, mux58_b1_sel_is_2_o);
  AL_MUX mux59_b2 (
    .i0(1'b0),
    .i1(n229[2]),
    .sel(mux59_b2_sel_is_2_o),
    .o(n240[2]));
  and mux59_b2_sel_is_2 (mux59_b2_sel_is_2_o, n117_neg, mux58_b2_sel_is_2_o);
  and mux59_b3_sel_is_2 (mux59_b3_sel_is_2_o, n117_neg, mux58_b3_sel_is_2_o);
  and mux59_b5_sel_is_2 (mux59_b5_sel_is_2_o, n117_neg, mux58_b5_sel_is_2_o);
  and mux59_b7_sel_is_2 (mux59_b7_sel_is_2_o, n117_neg, mux58_b7_sel_is_2_o);
  and mux59_b9_sel_is_2 (mux59_b9_sel_is_2_o, n117_neg, mux58_b9_sel_is_2_o);
  AL_MUX mux5_b0 (
    .i0(1'b0),
    .i1(n184[0]),
    .sel(mux5_b0_sel_is_0_o),
    .o(n186[0]));
  and mux5_b0_sel_is_0 (mux5_b0_sel_is_0_o, n171_neg, n172_neg);
  binary_mux_s1_w1 mux5_b10 (
    .i0(n185[10]),
    .i1(1'b1),
    .sel(n171),
    .o(n186[10]));  // sources/rtl/camera_init.v(256)
  AL_MUX mux5_b11 (
    .i0(1'b1),
    .i1(n184[11]),
    .sel(mux5_b0_sel_is_0_o),
    .o(n186[11]));
  and mux5_b13_sel_is_0 (mux5_b13_sel_is_0_o, n171_neg, mux4_b13_sel_is_0_o_neg);
  not mux5_b13_sel_is_0_o_inv (mux5_b13_sel_is_0_o_neg, mux5_b13_sel_is_0_o);
  binary_mux_s1_w1 mux5_b15 (
    .i0(n185[14]),
    .i1(1'b0),
    .sel(n171),
    .o(n186[15]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux5_b3 (
    .i0(n185[3]),
    .i1(1'b0),
    .sel(n171),
    .o(n186[3]));  // sources/rtl/camera_init.v(256)
  AL_MUX mux5_b5 (
    .i0(1'b0),
    .i1(n183[0]),
    .sel(mux5_b5_sel_is_2_o),
    .o(n186[5]));
  and mux5_b5_sel_is_2 (mux5_b5_sel_is_2_o, n171_neg, mux4_b5_sel_is_0_o);
  AL_MUX mux5_b7 (
    .i0(1'b0),
    .i1(n178[2]),
    .sel(mux5_b7_sel_is_2_o),
    .o(n186[7]));
  and mux5_b7_sel_is_2 (mux5_b7_sel_is_2_o, n171_neg, mux4_b7_sel_is_2_o);
  and mux60_b0_sel_is_2 (mux60_b0_sel_is_2_o, n116_neg, mux59_b0_sel_is_2_o);
  and mux60_b10_sel_is_2 (mux60_b10_sel_is_2_o, n116_neg, mux59_b10_sel_is_2_o);
  and mux60_b11_sel_is_2 (mux60_b11_sel_is_2_o, n116_neg, mux59_b11_sel_is_2_o);
  and mux60_b12_sel_is_2 (mux60_b12_sel_is_2_o, n116_neg, mux59_b12_sel_is_2_o);
  and mux60_b13_sel_is_2 (mux60_b13_sel_is_2_o, n116_neg, mux59_b13_sel_is_2_o);
  and mux60_b15_sel_is_2 (mux60_b15_sel_is_2_o, n116_neg, mux59_b15_sel_is_2_o);
  and mux60_b1_sel_is_2 (mux60_b1_sel_is_2_o, n116_neg, mux59_b1_sel_is_2_o);
  binary_mux_s1_w1 mux60_b2 (
    .i0(n240[2]),
    .i1(1'b1),
    .sel(n116),
    .o(n241[2]));  // sources/rtl/camera_init.v(256)
  and mux60_b3_sel_is_2 (mux60_b3_sel_is_2_o, n116_neg, mux59_b3_sel_is_2_o);
  and mux60_b5_sel_is_2 (mux60_b5_sel_is_2_o, n116_neg, mux59_b5_sel_is_2_o);
  and mux60_b7_sel_is_2 (mux60_b7_sel_is_2_o, n116_neg, mux59_b7_sel_is_2_o);
  and mux60_b9_sel_is_2 (mux60_b9_sel_is_2_o, n116_neg, mux59_b9_sel_is_2_o);
  AL_MUX mux61_b0 (
    .i0(1'b0),
    .i1(n231[0]),
    .sel(mux61_b0_sel_is_2_o),
    .o(n242[0]));
  and mux61_b0_sel_is_2 (mux61_b0_sel_is_2_o, n115_neg, mux60_b0_sel_is_2_o);
  and mux61_b10_sel_is_2 (mux61_b10_sel_is_2_o, n115_neg, mux60_b10_sel_is_2_o);
  and mux61_b11_sel_is_2 (mux61_b11_sel_is_2_o, n115_neg, mux60_b11_sel_is_2_o);
  and mux61_b12_sel_is_2 (mux61_b12_sel_is_2_o, n115_neg, mux60_b12_sel_is_2_o);
  and mux61_b13_sel_is_2 (mux61_b13_sel_is_2_o, n115_neg, mux60_b13_sel_is_2_o);
  and mux61_b15_sel_is_2 (mux61_b15_sel_is_2_o, n115_neg, mux60_b15_sel_is_2_o);
  and mux61_b1_sel_is_2 (mux61_b1_sel_is_2_o, n115_neg, mux60_b1_sel_is_2_o);
  binary_mux_s1_w1 mux61_b2 (
    .i0(n241[2]),
    .i1(1'b0),
    .sel(n115),
    .o(n242[2]));  // sources/rtl/camera_init.v(256)
  and mux61_b3_sel_is_2 (mux61_b3_sel_is_2_o, n115_neg, mux60_b3_sel_is_2_o);
  and mux61_b5_sel_is_2 (mux61_b5_sel_is_2_o, n115_neg, mux60_b5_sel_is_2_o);
  and mux61_b7_sel_is_2 (mux61_b7_sel_is_2_o, n115_neg, mux60_b7_sel_is_2_o);
  and mux61_b9_sel_is_2 (mux61_b9_sel_is_2_o, n115_neg, mux60_b9_sel_is_2_o);
  and mux62_b10_sel_is_2 (mux62_b10_sel_is_2_o, n114_neg, mux61_b10_sel_is_2_o);
  and mux62_b11_sel_is_2 (mux62_b11_sel_is_2_o, n114_neg, mux61_b11_sel_is_2_o);
  and mux62_b12_sel_is_2 (mux62_b12_sel_is_2_o, n114_neg, mux61_b12_sel_is_2_o);
  and mux62_b13_sel_is_2 (mux62_b13_sel_is_2_o, n114_neg, mux61_b13_sel_is_2_o);
  and mux62_b15_sel_is_2 (mux62_b15_sel_is_2_o, n114_neg, mux61_b15_sel_is_2_o);
  and mux62_b1_sel_is_2 (mux62_b1_sel_is_2_o, n114_neg, mux61_b1_sel_is_2_o);
  and mux62_b3_sel_is_2 (mux62_b3_sel_is_2_o, n114_neg, mux61_b3_sel_is_2_o);
  and mux62_b4_sel_is_2 (mux62_b4_sel_is_2_o, n114_neg, mux61_b0_sel_is_2_o);
  and mux62_b5_sel_is_2 (mux62_b5_sel_is_2_o, n114_neg, mux61_b5_sel_is_2_o);
  and mux62_b7_sel_is_2 (mux62_b7_sel_is_2_o, n114_neg, mux61_b7_sel_is_2_o);
  and mux62_b9_sel_is_2 (mux62_b9_sel_is_2_o, n114_neg, mux61_b9_sel_is_2_o);
  and mux63_b0_sel_is_0 (mux63_b0_sel_is_0_o, n113_neg, n114_neg);
  AL_MUX mux63_b1 (
    .i0(1'b0),
    .i1(n230[1]),
    .sel(mux63_b1_sel_is_2_o),
    .o(n244[1]));
  and mux63_b10_sel_is_2 (mux63_b10_sel_is_2_o, n113_neg, mux62_b10_sel_is_2_o);
  and mux63_b11_sel_is_2 (mux63_b11_sel_is_2_o, n113_neg, mux62_b11_sel_is_2_o);
  and mux63_b12_sel_is_2 (mux63_b12_sel_is_2_o, n113_neg, mux62_b12_sel_is_2_o);
  and mux63_b13_sel_is_2 (mux63_b13_sel_is_2_o, n113_neg, mux62_b13_sel_is_2_o);
  and mux63_b15_sel_is_2 (mux63_b15_sel_is_2_o, n113_neg, mux62_b15_sel_is_2_o);
  and mux63_b1_sel_is_2 (mux63_b1_sel_is_2_o, n113_neg, mux62_b1_sel_is_2_o);
  AL_MUX mux63_b2 (
    .i0(1'b1),
    .i1(n242[2]),
    .sel(mux63_b0_sel_is_0_o),
    .o(n244[2]));
  and mux63_b3_sel_is_2 (mux63_b3_sel_is_2_o, n113_neg, mux62_b3_sel_is_2_o);
  and mux63_b4_sel_is_2 (mux63_b4_sel_is_2_o, n113_neg, mux62_b4_sel_is_2_o);
  AL_MUX mux63_b5 (
    .i0(1'b0),
    .i1(n228[5]),
    .sel(mux63_b5_sel_is_2_o),
    .o(n244[5]));
  and mux63_b5_sel_is_2 (mux63_b5_sel_is_2_o, n113_neg, mux62_b5_sel_is_2_o);
  AL_MUX mux63_b6 (
    .i0(1'b0),
    .i1(n219[6]),
    .sel(mux63_b12_sel_is_2_o),
    .o(n244[6]));
  AL_MUX mux63_b7 (
    .i0(1'b0),
    .i1(n223[7]),
    .sel(mux63_b7_sel_is_2_o),
    .o(n244[7]));
  and mux63_b7_sel_is_2 (mux63_b7_sel_is_2_o, n113_neg, mux62_b7_sel_is_2_o);
  and mux63_b9_sel_is_2 (mux63_b9_sel_is_2_o, n113_neg, mux62_b9_sel_is_2_o);
  AL_MUX mux64_b0 (
    .i0(1'b1),
    .i1(n242[0]),
    .sel(mux64_b0_sel_is_2_o),
    .o(n245[0]));
  and mux64_b0_sel_is_2 (mux64_b0_sel_is_2_o, n112_neg, mux63_b0_sel_is_0_o);
  and mux64_b10_sel_is_2 (mux64_b10_sel_is_2_o, n112_neg, mux63_b10_sel_is_2_o);
  and mux64_b11_sel_is_2 (mux64_b11_sel_is_2_o, n112_neg, mux63_b11_sel_is_2_o);
  and mux64_b12_sel_is_2 (mux64_b12_sel_is_2_o, n112_neg, mux63_b12_sel_is_2_o);
  and mux64_b13_sel_is_2 (mux64_b13_sel_is_2_o, n112_neg, mux63_b13_sel_is_2_o);
  and mux64_b15_sel_is_2 (mux64_b15_sel_is_2_o, n112_neg, mux63_b15_sel_is_2_o);
  binary_mux_s1_w1 mux64_b2 (
    .i0(n244[2]),
    .i1(1'b0),
    .sel(n112),
    .o(n245[2]));  // sources/rtl/camera_init.v(256)
  and mux64_b3_sel_is_2 (mux64_b3_sel_is_2_o, n112_neg, mux63_b3_sel_is_2_o);
  and mux64_b4_sel_is_2 (mux64_b4_sel_is_2_o, n112_neg, mux63_b4_sel_is_2_o);
  binary_mux_s1_w1 mux64_b5 (
    .i0(n244[5]),
    .i1(1'b1),
    .sel(n112),
    .o(n245[5]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux64_b6 (
    .i0(n244[6]),
    .i1(1'b1),
    .sel(n112),
    .o(n245[6]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux64_b7 (
    .i0(n244[7]),
    .i1(1'b1),
    .sel(n112),
    .o(n245[7]));  // sources/rtl/camera_init.v(256)
  and mux64_b9_sel_is_2 (mux64_b9_sel_is_2_o, n112_neg, mux63_b9_sel_is_2_o);
  AL_MUX mux65_b1 (
    .i0(1'b1),
    .i1(n244[1]),
    .sel(mux65_b1_sel_is_0_o),
    .o(n246[1]));
  and mux65_b10_sel_is_2 (mux65_b10_sel_is_2_o, n111_neg, mux64_b10_sel_is_2_o);
  and mux65_b11_sel_is_2 (mux65_b11_sel_is_2_o, n111_neg, mux64_b11_sel_is_2_o);
  and mux65_b12_sel_is_2 (mux65_b12_sel_is_2_o, n111_neg, mux64_b12_sel_is_2_o);
  and mux65_b13_sel_is_2 (mux65_b13_sel_is_2_o, n111_neg, mux64_b13_sel_is_2_o);
  and mux65_b15_sel_is_2 (mux65_b15_sel_is_2_o, n111_neg, mux64_b15_sel_is_2_o);
  and mux65_b1_sel_is_0 (mux65_b1_sel_is_0_o, n111_neg, n112_neg);
  binary_mux_s1_w1 mux65_b2 (
    .i0(n245[2]),
    .i1(1'b1),
    .sel(n111),
    .o(n246[2]));  // sources/rtl/camera_init.v(256)
  and mux65_b3_sel_is_2 (mux65_b3_sel_is_2_o, n111_neg, mux64_b3_sel_is_2_o);
  and mux65_b4_sel_is_2 (mux65_b4_sel_is_2_o, n111_neg, mux64_b4_sel_is_2_o);
  AL_MUX mux65_b8 (
    .i0(1'b1),
    .i1(n233[8]),
    .sel(mux65_b10_sel_is_2_o),
    .o(n246[8]));
  and mux65_b9_sel_is_2 (mux65_b9_sel_is_2_o, n111_neg, mux64_b9_sel_is_2_o);
  and mux66_b0_sel_is_0 (mux66_b0_sel_is_0_o, n110_neg, n111_neg);
  and mux66_b10_sel_is_2 (mux66_b10_sel_is_2_o, n110_neg, mux65_b10_sel_is_2_o);
  and mux66_b11_sel_is_2 (mux66_b11_sel_is_2_o, n110_neg, mux65_b11_sel_is_2_o);
  and mux66_b12_sel_is_2 (mux66_b12_sel_is_2_o, n110_neg, mux65_b12_sel_is_2_o);
  and mux66_b13_sel_is_2 (mux66_b13_sel_is_2_o, n110_neg, mux65_b13_sel_is_2_o);
  and mux66_b15_sel_is_2 (mux66_b15_sel_is_2_o, n110_neg, mux65_b15_sel_is_2_o);
  and mux66_b3_sel_is_2 (mux66_b3_sel_is_2_o, n110_neg, mux65_b3_sel_is_2_o);
  and mux66_b4_sel_is_2 (mux66_b4_sel_is_2_o, n110_neg, mux65_b4_sel_is_2_o);
  AL_MUX mux66_b5 (
    .i0(1'b0),
    .i1(n245[5]),
    .sel(mux66_b0_sel_is_0_o),
    .o(n247[5]));
  binary_mux_s1_w1 mux66_b8 (
    .i0(n246[8]),
    .i1(1'b0),
    .sel(n110),
    .o(n247[8]));  // sources/rtl/camera_init.v(256)
  and mux66_b9_sel_is_2 (mux66_b9_sel_is_2_o, n110_neg, mux65_b9_sel_is_2_o);
  not mux66_b9_sel_is_2_o_inv (mux66_b9_sel_is_2_o_neg, mux66_b9_sel_is_2_o);
  and mux67_b0_sel_is_2 (mux67_b0_sel_is_2_o, n109_neg, mux66_b0_sel_is_0_o);
  and mux67_b10_sel_is_2 (mux67_b10_sel_is_2_o, n109_neg, mux66_b10_sel_is_2_o);
  and mux67_b11_sel_is_2 (mux67_b11_sel_is_2_o, n109_neg, mux66_b11_sel_is_2_o);
  and mux67_b12_sel_is_2 (mux67_b12_sel_is_2_o, n109_neg, mux66_b12_sel_is_2_o);
  and mux67_b13_sel_is_2 (mux67_b13_sel_is_2_o, n109_neg, mux66_b13_sel_is_2_o);
  and mux67_b15_sel_is_2 (mux67_b15_sel_is_2_o, n109_neg, mux66_b15_sel_is_2_o);
  and mux67_b1_sel_is_0 (mux67_b1_sel_is_0_o, n109_neg, n110_neg);
  AL_MUX mux67_b3 (
    .i0(1'b0),
    .i1(n232[3]),
    .sel(mux67_b3_sel_is_2_o),
    .o(n248[3]));
  and mux67_b3_sel_is_2 (mux67_b3_sel_is_2_o, n109_neg, mux66_b3_sel_is_2_o);
  and mux67_b4_sel_is_2 (mux67_b4_sel_is_2_o, n109_neg, mux66_b4_sel_is_2_o);
  AL_MUX mux67_b6 (
    .i0(1'b0),
    .i1(n245[6]),
    .sel(mux67_b0_sel_is_2_o),
    .o(n248[6]));
  AL_MUX mux67_b7 (
    .i0(1'b0),
    .i1(n245[7]),
    .sel(mux67_b0_sel_is_2_o),
    .o(n248[7]));
  and mux67_b9_sel_is_0 (mux67_b9_sel_is_0_o, n109_neg, mux66_b9_sel_is_2_o_neg);
  AL_MUX mux68_b0 (
    .i0(1'b0),
    .i1(n245[0]),
    .sel(mux68_b0_sel_is_2_o),
    .o(n249[0]));
  and mux68_b0_sel_is_2 (mux68_b0_sel_is_2_o, n108_neg, mux67_b0_sel_is_2_o);
  AL_MUX mux68_b1 (
    .i0(1'b0),
    .i1(n246[1]),
    .sel(mux68_b1_sel_is_2_o),
    .o(n249[1]));
  and mux68_b10_sel_is_2 (mux68_b10_sel_is_2_o, n108_neg, mux67_b10_sel_is_2_o);
  and mux68_b11_sel_is_2 (mux68_b11_sel_is_2_o, n108_neg, mux67_b11_sel_is_2_o);
  and mux68_b12_sel_is_2 (mux68_b12_sel_is_2_o, n108_neg, mux67_b12_sel_is_2_o);
  and mux68_b13_sel_is_2 (mux68_b13_sel_is_2_o, n108_neg, mux67_b13_sel_is_2_o);
  and mux68_b15_sel_is_2 (mux68_b15_sel_is_2_o, n108_neg, mux67_b15_sel_is_2_o);
  and mux68_b1_sel_is_2 (mux68_b1_sel_is_2_o, n108_neg, mux67_b1_sel_is_0_o);
  AL_MUX mux68_b2 (
    .i0(1'b0),
    .i1(n246[2]),
    .sel(mux68_b1_sel_is_2_o),
    .o(n249[2]));
  binary_mux_s1_w1 mux68_b3 (
    .i0(n248[3]),
    .i1(1'b1),
    .sel(n108),
    .o(n249[3]));  // sources/rtl/camera_init.v(256)
  AL_MUX mux68_b4 (
    .i0(1'b0),
    .i1(n231[4]),
    .sel(mux68_b4_sel_is_2_o),
    .o(n249[4]));
  and mux68_b4_sel_is_2 (mux68_b4_sel_is_2_o, n108_neg, mux67_b4_sel_is_2_o);
  AL_MUX mux68_b5 (
    .i0(1'b1),
    .i1(n247[5]),
    .sel(mux68_b5_sel_is_0_o),
    .o(n249[5]));
  and mux68_b5_sel_is_0 (mux68_b5_sel_is_0_o, n108_neg, n109_neg);
  and mux68_b9_sel_is_2 (mux68_b9_sel_is_2_o, n108_neg, mux67_b9_sel_is_0_o);
  binary_mux_s1_w1 mux69_b0 (
    .i0(n249[0]),
    .i1(1'b1),
    .sel(n107),
    .o(n250[0]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux69_b1 (
    .i0(n249[1]),
    .i1(1'b1),
    .sel(n107),
    .o(n250[1]));  // sources/rtl/camera_init.v(256)
  and mux69_b10_sel_is_2 (mux69_b10_sel_is_2_o, n107_neg, mux68_b10_sel_is_2_o);
  and mux69_b11_sel_is_2 (mux69_b11_sel_is_2_o, n107_neg, mux68_b11_sel_is_2_o);
  and mux69_b12_sel_is_2 (mux69_b12_sel_is_2_o, n107_neg, mux68_b12_sel_is_2_o);
  and mux69_b13_sel_is_2 (mux69_b13_sel_is_2_o, n107_neg, mux68_b13_sel_is_2_o);
  and mux69_b15_sel_is_2 (mux69_b15_sel_is_2_o, n107_neg, mux68_b15_sel_is_2_o);
  binary_mux_s1_w1 mux69_b4 (
    .i0(n249[4]),
    .i1(1'b1),
    .sel(n107),
    .o(n250[4]));  // sources/rtl/camera_init.v(256)
  and mux69_b6_sel_is_0 (mux69_b6_sel_is_0_o, n107_neg, n108_neg);
  and mux69_b8_sel_is_2 (mux69_b8_sel_is_2_o, n107_neg, mux68_b5_sel_is_0_o);
  and mux69_b9_sel_is_2 (mux69_b9_sel_is_2_o, n107_neg, mux68_b9_sel_is_2_o);
  binary_mux_s1_w1 mux6_b0 (
    .i0(n186[0]),
    .i1(1'b1),
    .sel(n170),
    .o(n187[0]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux6_b1 (
    .i0(n186[0]),
    .i1(1'b0),
    .sel(n170),
    .o(n187[1]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux6_b11 (
    .i0(n186[11]),
    .i1(1'b0),
    .sel(n170),
    .o(n187[11]));  // sources/rtl/camera_init.v(256)
  and mux6_b13_sel_is_0 (mux6_b13_sel_is_0_o, n170_neg, mux5_b13_sel_is_0_o_neg);
  and mux6_b14_sel_is_0 (mux6_b14_sel_is_0_o, n170_neg, n171_neg);
  binary_mux_s1_w1 mux6_b3 (
    .i0(n186[3]),
    .i1(1'b1),
    .sel(n170),
    .o(n187[3]));  // sources/rtl/camera_init.v(256)
  and mux6_b4_sel_is_2 (mux6_b4_sel_is_2_o, n170_neg, mux5_b0_sel_is_0_o);
  binary_mux_s1_w1 mux6_b5 (
    .i0(n186[5]),
    .i1(1'b1),
    .sel(n170),
    .o(n187[5]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux70_b0 (
    .i0(n250[0]),
    .i1(1'b0),
    .sel(n106),
    .o(n251[0]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux70_b1 (
    .i0(n250[1]),
    .i1(1'b0),
    .sel(n106),
    .o(n251[1]));  // sources/rtl/camera_init.v(256)
  and mux70_b10_sel_is_2 (mux70_b10_sel_is_2_o, n106_neg, mux69_b10_sel_is_2_o);
  and mux70_b11_sel_is_2 (mux70_b11_sel_is_2_o, n106_neg, mux69_b11_sel_is_2_o);
  and mux70_b12_sel_is_2 (mux70_b12_sel_is_2_o, n106_neg, mux69_b12_sel_is_2_o);
  and mux70_b13_sel_is_2 (mux70_b13_sel_is_2_o, n106_neg, mux69_b13_sel_is_2_o);
  and mux70_b15_sel_is_2 (mux70_b15_sel_is_2_o, n106_neg, mux69_b15_sel_is_2_o);
  and mux70_b2_sel_is_0 (mux70_b2_sel_is_0_o, n106_neg, n107_neg);
  AL_MUX mux70_b3 (
    .i0(1'b0),
    .i1(n249[3]),
    .sel(mux70_b2_sel_is_0_o),
    .o(n251[3]));
  AL_MUX mux70_b5 (
    .i0(1'b0),
    .i1(n249[5]),
    .sel(mux70_b2_sel_is_0_o),
    .o(n251[5]));
  AL_MUX mux70_b6 (
    .i0(1'b1),
    .i1(n248[6]),
    .sel(mux70_b6_sel_is_2_o),
    .o(n251[6]));
  and mux70_b6_sel_is_2 (mux70_b6_sel_is_2_o, n106_neg, mux69_b6_sel_is_0_o);
  and mux70_b8_sel_is_2 (mux70_b8_sel_is_2_o, n106_neg, mux69_b8_sel_is_2_o);
  and mux70_b9_sel_is_2 (mux70_b9_sel_is_2_o, n106_neg, mux69_b9_sel_is_2_o);
  and mux71_b10_sel_is_2 (mux71_b10_sel_is_2_o, n105_neg, mux70_b10_sel_is_2_o);
  and mux71_b11_sel_is_2 (mux71_b11_sel_is_2_o, n105_neg, mux70_b11_sel_is_2_o);
  and mux71_b12_sel_is_2 (mux71_b12_sel_is_2_o, n105_neg, mux70_b12_sel_is_2_o);
  and mux71_b13_sel_is_2 (mux71_b13_sel_is_2_o, n105_neg, mux70_b13_sel_is_2_o);
  and mux71_b15_sel_is_2 (mux71_b15_sel_is_2_o, n105_neg, mux70_b15_sel_is_2_o);
  AL_MUX mux71_b2 (
    .i0(1'b1),
    .i1(n249[2]),
    .sel(mux71_b2_sel_is_2_o),
    .o(n252[2]));
  and mux71_b2_sel_is_2 (mux71_b2_sel_is_2_o, n105_neg, mux70_b2_sel_is_0_o);
  binary_mux_s1_w1 mux71_b3 (
    .i0(n251[3]),
    .i1(1'b1),
    .sel(n105),
    .o(n252[3]));  // sources/rtl/camera_init.v(256)
  and mux71_b4_sel_is_0 (mux71_b4_sel_is_0_o, n105_neg, n106_neg);
  and mux71_b7_sel_is_2 (mux71_b7_sel_is_2_o, n105_neg, mux70_b6_sel_is_2_o);
  and mux71_b8_sel_is_2 (mux71_b8_sel_is_2_o, n105_neg, mux70_b8_sel_is_2_o);
  and mux71_b9_sel_is_2 (mux71_b9_sel_is_2_o, n105_neg, mux70_b9_sel_is_2_o);
  AL_MUX mux72_b0 (
    .i0(1'b1),
    .i1(n251[0]),
    .sel(mux72_b0_sel_is_0_o),
    .o(n253[0]));
  and mux72_b0_sel_is_0 (mux72_b0_sel_is_0_o, n104_neg, n105_neg);
  and mux72_b10_sel_is_2 (mux72_b10_sel_is_2_o, n104_neg, mux71_b10_sel_is_2_o);
  and mux72_b11_sel_is_2 (mux72_b11_sel_is_2_o, n104_neg, mux71_b11_sel_is_2_o);
  and mux72_b12_sel_is_2 (mux72_b12_sel_is_2_o, n104_neg, mux71_b12_sel_is_2_o);
  and mux72_b13_sel_is_2 (mux72_b13_sel_is_2_o, n104_neg, mux71_b13_sel_is_2_o);
  and mux72_b15_sel_is_2 (mux72_b15_sel_is_2_o, n104_neg, mux71_b15_sel_is_2_o);
  binary_mux_s1_w1 mux72_b2 (
    .i0(n252[2]),
    .i1(1'b0),
    .sel(n104),
    .o(n253[2]));  // sources/rtl/camera_init.v(256)
  AL_MUX mux72_b4 (
    .i0(1'b0),
    .i1(n250[4]),
    .sel(mux72_b4_sel_is_2_o),
    .o(n253[4]));
  and mux72_b4_sel_is_2 (mux72_b4_sel_is_2_o, n104_neg, mux71_b4_sel_is_0_o);
  AL_MUX mux72_b5 (
    .i0(1'b1),
    .i1(n251[5]),
    .sel(mux72_b0_sel_is_0_o),
    .o(n253[5]));
  and mux72_b7_sel_is_2 (mux72_b7_sel_is_2_o, n104_neg, mux71_b7_sel_is_2_o);
  and mux72_b8_sel_is_2 (mux72_b8_sel_is_2_o, n104_neg, mux71_b8_sel_is_2_o);
  and mux72_b9_sel_is_2 (mux72_b9_sel_is_2_o, n104_neg, mux71_b9_sel_is_2_o);
  binary_mux_s1_w1 mux73_b0 (
    .i0(n253[0]),
    .i1(1'b0),
    .sel(n103),
    .o(n254[0]));  // sources/rtl/camera_init.v(256)
  and mux73_b10_sel_is_2 (mux73_b10_sel_is_2_o, n103_neg, mux72_b10_sel_is_2_o);
  and mux73_b11_sel_is_2 (mux73_b11_sel_is_2_o, n103_neg, mux72_b11_sel_is_2_o);
  and mux73_b12_sel_is_2 (mux73_b12_sel_is_2_o, n103_neg, mux72_b12_sel_is_2_o);
  and mux73_b13_sel_is_2 (mux73_b13_sel_is_2_o, n103_neg, mux72_b13_sel_is_2_o);
  and mux73_b15_sel_is_2 (mux73_b15_sel_is_2_o, n103_neg, mux72_b15_sel_is_2_o);
  and mux73_b1_sel_is_2 (mux73_b1_sel_is_2_o, n103_neg, mux72_b0_sel_is_0_o);
  AL_MUX mux73_b3 (
    .i0(1'b0),
    .i1(n252[3]),
    .sel(mux73_b3_sel_is_0_o),
    .o(n254[3]));
  and mux73_b3_sel_is_0 (mux73_b3_sel_is_0_o, n103_neg, n104_neg);
  binary_mux_s1_w1 mux73_b4 (
    .i0(n253[4]),
    .i1(1'b1),
    .sel(n103),
    .o(n254[4]));  // sources/rtl/camera_init.v(256)
  and mux73_b7_sel_is_2 (mux73_b7_sel_is_2_o, n103_neg, mux72_b7_sel_is_2_o);
  and mux73_b8_sel_is_2 (mux73_b8_sel_is_2_o, n103_neg, mux72_b8_sel_is_2_o);
  and mux73_b9_sel_is_2 (mux73_b9_sel_is_2_o, n103_neg, mux72_b9_sel_is_2_o);
  binary_mux_s1_w1 mux74_b0 (
    .i0(n254[0]),
    .i1(1'b1),
    .sel(n102),
    .o(n255[0]));  // sources/rtl/camera_init.v(256)
  AL_MUX mux74_b1 (
    .i0(1'b1),
    .i1(n251[1]),
    .sel(mux74_b1_sel_is_2_o),
    .o(n255[1]));
  and mux74_b10_sel_is_2 (mux74_b10_sel_is_2_o, n102_neg, mux73_b10_sel_is_2_o);
  and mux74_b11_sel_is_2 (mux74_b11_sel_is_2_o, n102_neg, mux73_b11_sel_is_2_o);
  and mux74_b12_sel_is_2 (mux74_b12_sel_is_2_o, n102_neg, mux73_b12_sel_is_2_o);
  and mux74_b13_sel_is_2 (mux74_b13_sel_is_2_o, n102_neg, mux73_b13_sel_is_2_o);
  and mux74_b15_sel_is_2 (mux74_b15_sel_is_2_o, n102_neg, mux73_b15_sel_is_2_o);
  and mux74_b1_sel_is_2 (mux74_b1_sel_is_2_o, n102_neg, mux73_b1_sel_is_2_o);
  AL_MUX mux74_b2 (
    .i0(1'b1),
    .i1(n253[2]),
    .sel(mux74_b2_sel_is_0_o),
    .o(n255[2]));
  and mux74_b2_sel_is_0 (mux74_b2_sel_is_0_o, n102_neg, n103_neg);
  and mux74_b7_sel_is_2 (mux74_b7_sel_is_2_o, n102_neg, mux73_b7_sel_is_2_o);
  and mux74_b8_sel_is_2 (mux74_b8_sel_is_2_o, n102_neg, mux73_b8_sel_is_2_o);
  and mux74_b9_sel_is_2 (mux74_b9_sel_is_2_o, n102_neg, mux73_b9_sel_is_2_o);
  binary_mux_s1_w1 mux75_b1 (
    .i0(n255[1]),
    .i1(1'b0),
    .sel(n101),
    .o(n256[1]));  // sources/rtl/camera_init.v(256)
  and mux75_b10_sel_is_2 (mux75_b10_sel_is_2_o, n101_neg, mux74_b10_sel_is_2_o);
  and mux75_b11_sel_is_2 (mux75_b11_sel_is_2_o, n101_neg, mux74_b11_sel_is_2_o);
  and mux75_b12_sel_is_2 (mux75_b12_sel_is_2_o, n101_neg, mux74_b12_sel_is_2_o);
  and mux75_b13_sel_is_2 (mux75_b13_sel_is_2_o, n101_neg, mux74_b13_sel_is_2_o);
  and mux75_b15_sel_is_2 (mux75_b15_sel_is_2_o, n101_neg, mux74_b15_sel_is_2_o);
  binary_mux_s1_w1 mux75_b2 (
    .i0(n255[2]),
    .i1(1'b0),
    .sel(n101),
    .o(n256[2]));  // sources/rtl/camera_init.v(256)
  and mux75_b3_sel_is_0 (mux75_b3_sel_is_0_o, n101_neg, n102_neg);
  AL_MUX mux75_b4 (
    .i0(1'b0),
    .i1(n254[4]),
    .sel(mux75_b3_sel_is_0_o),
    .o(n256[4]));
  AL_MUX mux75_b5 (
    .i0(1'b0),
    .i1(n253[5]),
    .sel(mux75_b5_sel_is_2_o),
    .o(n256[5]));
  and mux75_b5_sel_is_2 (mux75_b5_sel_is_2_o, n101_neg, mux74_b2_sel_is_0_o);
  AL_MUX mux75_b6 (
    .i0(1'b0),
    .i1(n251[6]),
    .sel(mux75_b6_sel_is_2_o),
    .o(n256[6]));
  and mux75_b6_sel_is_2 (mux75_b6_sel_is_2_o, n101_neg, mux74_b1_sel_is_2_o);
  AL_MUX mux75_b7 (
    .i0(1'b1),
    .i1(n248[7]),
    .sel(mux75_b7_sel_is_2_o),
    .o(n256[7]));
  and mux75_b7_sel_is_2 (mux75_b7_sel_is_2_o, n101_neg, mux74_b7_sel_is_2_o);
  and mux75_b8_sel_is_2 (mux75_b8_sel_is_2_o, n101_neg, mux74_b8_sel_is_2_o);
  and mux75_b9_sel_is_2 (mux75_b9_sel_is_2_o, n101_neg, mux74_b9_sel_is_2_o);
  AL_MUX mux76_b0 (
    .i0(1'b0),
    .i1(n255[0]),
    .sel(mux76_b0_sel_is_0_o),
    .o(n257[0]));
  and mux76_b0_sel_is_0 (mux76_b0_sel_is_0_o, n100_neg, n101_neg);
  binary_mux_s1_w1 mux76_b1 (
    .i0(n256[1]),
    .i1(1'b1),
    .sel(n100),
    .o(n257[1]));  // sources/rtl/camera_init.v(256)
  and mux76_b10_sel_is_2 (mux76_b10_sel_is_2_o, n100_neg, mux75_b10_sel_is_2_o);
  and mux76_b11_sel_is_2 (mux76_b11_sel_is_2_o, n100_neg, mux75_b11_sel_is_2_o);
  and mux76_b12_sel_is_2 (mux76_b12_sel_is_2_o, n100_neg, mux75_b12_sel_is_2_o);
  and mux76_b13_sel_is_2 (mux76_b13_sel_is_2_o, n100_neg, mux75_b13_sel_is_2_o);
  and mux76_b15_sel_is_2 (mux76_b15_sel_is_2_o, n100_neg, mux75_b15_sel_is_2_o);
  AL_MUX mux76_b3 (
    .i0(1'b1),
    .i1(n254[3]),
    .sel(mux76_b3_sel_is_2_o),
    .o(n257[3]));
  and mux76_b3_sel_is_2 (mux76_b3_sel_is_2_o, n100_neg, mux75_b3_sel_is_0_o);
  and mux76_b8_sel_is_2 (mux76_b8_sel_is_2_o, n100_neg, mux75_b8_sel_is_2_o);
  and mux76_b9_sel_is_2 (mux76_b9_sel_is_2_o, n100_neg, mux75_b9_sel_is_2_o);
  and mux77_b10_sel_is_2 (mux77_b10_sel_is_2_o, n99_neg, mux76_b10_sel_is_2_o);
  and mux77_b11_sel_is_2 (mux77_b11_sel_is_2_o, n99_neg, mux76_b11_sel_is_2_o);
  and mux77_b12_sel_is_2 (mux77_b12_sel_is_2_o, n99_neg, mux76_b12_sel_is_2_o);
  and mux77_b13_sel_is_2 (mux77_b13_sel_is_2_o, n99_neg, mux76_b13_sel_is_2_o);
  and mux77_b15_sel_is_2 (mux77_b15_sel_is_2_o, n99_neg, mux76_b15_sel_is_2_o);
  AL_MUX mux77_b2 (
    .i0(1'b1),
    .i1(n256[2]),
    .sel(mux77_b2_sel_is_0_o),
    .o(n258[2]));
  and mux77_b2_sel_is_0 (mux77_b2_sel_is_0_o, n99_neg, n100_neg);
  binary_mux_s1_w1 mux77_b3 (
    .i0(n257[3]),
    .i1(1'b0),
    .sel(n99),
    .o(n258[3]));  // sources/rtl/camera_init.v(256)
  AL_MUX mux77_b4 (
    .i0(1'b1),
    .i1(n256[4]),
    .sel(mux77_b2_sel_is_0_o),
    .o(n258[4]));
  and mux77_b8_sel_is_2 (mux77_b8_sel_is_2_o, n99_neg, mux76_b8_sel_is_2_o);
  and mux77_b9_sel_is_2 (mux77_b9_sel_is_2_o, n99_neg, mux76_b9_sel_is_2_o);
  AL_MUX mux78_b0 (
    .i0(1'b1),
    .i1(n257[0]),
    .sel(mux78_b0_sel_is_0_o),
    .o(n259[0]));
  and mux78_b0_sel_is_0 (mux78_b0_sel_is_0_o, n98_neg, n99_neg);
  AL_MUX mux78_b1 (
    .i0(1'b0),
    .i1(n257[1]),
    .sel(mux78_b0_sel_is_0_o),
    .o(n259[1]));
  and mux78_b10_sel_is_2 (mux78_b10_sel_is_2_o, n98_neg, mux77_b10_sel_is_2_o);
  and mux78_b11_sel_is_2 (mux78_b11_sel_is_2_o, n98_neg, mux77_b11_sel_is_2_o);
  and mux78_b12_sel_is_2 (mux78_b12_sel_is_2_o, n98_neg, mux77_b12_sel_is_2_o);
  and mux78_b13_sel_is_2 (mux78_b13_sel_is_2_o, n98_neg, mux77_b13_sel_is_2_o);
  and mux78_b15_sel_is_2 (mux78_b15_sel_is_2_o, n98_neg, mux77_b15_sel_is_2_o);
  binary_mux_s1_w1 mux78_b4 (
    .i0(n258[4]),
    .i1(1'b0),
    .sel(n98),
    .o(n259[4]));  // sources/rtl/camera_init.v(256)
  AL_MUX mux78_b5 (
    .i0(1'b1),
    .i1(n256[5]),
    .sel(mux78_b5_sel_is_2_o),
    .o(n259[5]));
  and mux78_b5_sel_is_2 (mux78_b5_sel_is_2_o, n98_neg, mux77_b2_sel_is_0_o);
  and mux78_b8_sel_is_2 (mux78_b8_sel_is_2_o, n98_neg, mux77_b8_sel_is_2_o);
  and mux78_b9_sel_is_2 (mux78_b9_sel_is_2_o, n98_neg, mux77_b9_sel_is_2_o);
  binary_mux_s1_w1 mux79_b0 (
    .i0(n259[0]),
    .i1(1'b0),
    .sel(n97),
    .o(n260[0]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux79_b1 (
    .i0(n259[1]),
    .i1(1'b1),
    .sel(n97),
    .o(n260[1]));  // sources/rtl/camera_init.v(256)
  and mux79_b10_sel_is_2 (mux79_b10_sel_is_2_o, n97_neg, mux78_b10_sel_is_2_o);
  and mux79_b11_sel_is_2 (mux79_b11_sel_is_2_o, n97_neg, mux78_b11_sel_is_2_o);
  and mux79_b12_sel_is_2 (mux79_b12_sel_is_2_o, n97_neg, mux78_b12_sel_is_2_o);
  and mux79_b13_sel_is_2 (mux79_b13_sel_is_2_o, n97_neg, mux78_b13_sel_is_2_o);
  and mux79_b15_sel_is_2 (mux79_b15_sel_is_2_o, n97_neg, mux78_b15_sel_is_2_o);
  and mux79_b2_sel_is_0 (mux79_b2_sel_is_0_o, n97_neg, n98_neg);
  AL_MUX mux79_b3 (
    .i0(1'b1),
    .i1(n258[3]),
    .sel(mux79_b2_sel_is_0_o),
    .o(n260[3]));
  binary_mux_s1_w1 mux79_b5 (
    .i0(n259[5]),
    .i1(1'b0),
    .sel(n97),
    .o(n260[5]));  // sources/rtl/camera_init.v(256)
  AL_MUX mux79_b6 (
    .i0(1'b1),
    .i1(n256[6]),
    .sel(mux79_b6_sel_is_2_o),
    .o(n260[6]));
  and mux79_b6_sel_is_2 (mux79_b6_sel_is_2_o, n97_neg, mux78_b5_sel_is_2_o);
  and mux79_b8_sel_is_2 (mux79_b8_sel_is_2_o, n97_neg, mux78_b8_sel_is_2_o);
  and mux79_b9_sel_is_2 (mux79_b9_sel_is_2_o, n97_neg, mux78_b9_sel_is_2_o);
  binary_mux_s1_w1 mux7_b1 (
    .i0(n187[1]),
    .i1(1'b1),
    .sel(n169),
    .o(n188[1]));  // sources/rtl/camera_init.v(256)
  AL_MUX mux7_b10 (
    .i0(1'b0),
    .i1(n186[10]),
    .sel(mux7_b10_sel_is_0_o),
    .o(n188[10]));
  and mux7_b10_sel_is_0 (mux7_b10_sel_is_0_o, n169_neg, n170_neg);
  binary_mux_s1_w1 mux7_b11 (
    .i0(n187[11]),
    .i1(1'b0),
    .sel(n169),
    .o(n188[11]));  // sources/rtl/camera_init.v(256)
  and mux7_b13_sel_is_2 (mux7_b13_sel_is_2_o, n169_neg, mux6_b13_sel_is_0_o);
  and mux7_b14_sel_is_2 (mux7_b14_sel_is_2_o, n169_neg, mux6_b14_sel_is_0_o);
  AL_MUX mux7_b15 (
    .i0(1'b1),
    .i1(n186[15]),
    .sel(mux7_b10_sel_is_0_o),
    .o(n188[15]));
  and mux7_b4_sel_is_2 (mux7_b4_sel_is_2_o, n169_neg, mux6_b4_sel_is_2_o);
  AL_MUX mux7_b7 (
    .i0(1'b1),
    .i1(n186[7]),
    .sel(mux7_b10_sel_is_0_o),
    .o(n188[7]));
  AL_MUX mux7_b8 (
    .i0(1'b1),
    .i1(n185[8]),
    .sel(mux7_b14_sel_is_2_o),
    .o(n188[8]));
  not mux7_b9_sel_is_2_o_inv (mux7_b9_sel_is_2_o_neg, mux7_b4_sel_is_2_o);
  binary_mux_s1_w1 mux80_b0 (
    .i0(n260[0]),
    .i1(1'b1),
    .sel(n96),
    .o(n261[0]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux80_b1 (
    .i0(n260[1]),
    .i1(1'b0),
    .sel(n96),
    .o(n261[1]));  // sources/rtl/camera_init.v(256)
  and mux80_b10_sel_is_2 (mux80_b10_sel_is_2_o, n96_neg, mux79_b10_sel_is_2_o);
  and mux80_b11_sel_is_2 (mux80_b11_sel_is_2_o, n96_neg, mux79_b11_sel_is_2_o);
  and mux80_b12_sel_is_2 (mux80_b12_sel_is_2_o, n96_neg, mux79_b12_sel_is_2_o);
  and mux80_b13_sel_is_2 (mux80_b13_sel_is_2_o, n96_neg, mux79_b13_sel_is_2_o);
  and mux80_b15_sel_is_2 (mux80_b15_sel_is_2_o, n96_neg, mux79_b15_sel_is_2_o);
  and mux80_b2_sel_is_2 (mux80_b2_sel_is_2_o, n96_neg, mux79_b2_sel_is_0_o);
  binary_mux_s1_w1 mux80_b3 (
    .i0(n260[3]),
    .i1(1'b0),
    .sel(n96),
    .o(n261[3]));  // sources/rtl/camera_init.v(256)
  and mux80_b4_sel_is_0 (mux80_b4_sel_is_0_o, n96_neg, n97_neg);
  binary_mux_s1_w1 mux80_b5 (
    .i0(n260[5]),
    .i1(1'b1),
    .sel(n96),
    .o(n261[5]));  // sources/rtl/camera_init.v(256)
  and mux80_b7_sel_is_2 (mux80_b7_sel_is_2_o, n96_neg, mux79_b6_sel_is_2_o);
  and mux80_b8_sel_is_2 (mux80_b8_sel_is_2_o, n96_neg, mux79_b8_sel_is_2_o);
  and mux80_b9_sel_is_2 (mux80_b9_sel_is_2_o, n96_neg, mux79_b9_sel_is_2_o);
  and mux81_b10_sel_is_2 (mux81_b10_sel_is_2_o, n95_neg, mux80_b10_sel_is_2_o);
  and mux81_b11_sel_is_2 (mux81_b11_sel_is_2_o, n95_neg, mux80_b11_sel_is_2_o);
  and mux81_b12_sel_is_2 (mux81_b12_sel_is_2_o, n95_neg, mux80_b12_sel_is_2_o);
  and mux81_b13_sel_is_2 (mux81_b13_sel_is_2_o, n95_neg, mux80_b13_sel_is_2_o);
  and mux81_b15_sel_is_2 (mux81_b15_sel_is_2_o, n95_neg, mux80_b15_sel_is_2_o);
  AL_MUX mux81_b2 (
    .i0(1'b0),
    .i1(n258[2]),
    .sel(mux81_b2_sel_is_2_o),
    .o(n262[2]));
  and mux81_b2_sel_is_2 (mux81_b2_sel_is_2_o, n95_neg, mux80_b2_sel_is_2_o);
  AL_MUX mux81_b4 (
    .i0(1'b1),
    .i1(n259[4]),
    .sel(mux81_b4_sel_is_2_o),
    .o(n262[4]));
  and mux81_b4_sel_is_2 (mux81_b4_sel_is_2_o, n95_neg, mux80_b4_sel_is_0_o);
  and mux81_b6_sel_is_0 (mux81_b6_sel_is_0_o, n95_neg, n96_neg);
  and mux81_b7_sel_is_2 (mux81_b7_sel_is_2_o, n95_neg, mux80_b7_sel_is_2_o);
  and mux81_b8_sel_is_2 (mux81_b8_sel_is_2_o, n95_neg, mux80_b8_sel_is_2_o);
  and mux81_b9_sel_is_2 (mux81_b9_sel_is_2_o, n95_neg, mux80_b9_sel_is_2_o);
  and mux82_b0_sel_is_0 (mux82_b0_sel_is_0_o, n94_neg, n95_neg);
  AL_MUX mux82_b1 (
    .i0(1'b1),
    .i1(n261[1]),
    .sel(mux82_b0_sel_is_0_o),
    .o(n263[1]));
  and mux82_b10_sel_is_2 (mux82_b10_sel_is_2_o, n94_neg, mux81_b10_sel_is_2_o);
  and mux82_b11_sel_is_2 (mux82_b11_sel_is_2_o, n94_neg, mux81_b11_sel_is_2_o);
  and mux82_b12_sel_is_2 (mux82_b12_sel_is_2_o, n94_neg, mux81_b12_sel_is_2_o);
  and mux82_b13_sel_is_2 (mux82_b13_sel_is_2_o, n94_neg, mux81_b13_sel_is_2_o);
  and mux82_b15_sel_is_2 (mux82_b15_sel_is_2_o, n94_neg, mux81_b15_sel_is_2_o);
  binary_mux_s1_w1 mux82_b2 (
    .i0(n262[2]),
    .i1(1'b1),
    .sel(n94),
    .o(n263[2]));  // sources/rtl/camera_init.v(256)
  AL_MUX mux82_b3 (
    .i0(1'b1),
    .i1(n261[3]),
    .sel(mux82_b0_sel_is_0_o),
    .o(n263[3]));
  and mux82_b6_sel_is_2 (mux82_b6_sel_is_2_o, n94_neg, mux81_b6_sel_is_0_o);
  and mux82_b7_sel_is_2 (mux82_b7_sel_is_2_o, n94_neg, mux81_b7_sel_is_2_o);
  AL_MUX mux82_b8 (
    .i0(1'b1),
    .i1(n247[8]),
    .sel(mux82_b8_sel_is_2_o),
    .o(n263[8]));
  and mux82_b8_sel_is_2 (mux82_b8_sel_is_2_o, n94_neg, mux81_b8_sel_is_2_o);
  and mux82_b9_sel_is_2 (mux82_b9_sel_is_2_o, n94_neg, mux81_b9_sel_is_2_o);
  and mux83_b0_sel_is_2 (mux83_b0_sel_is_2_o, n93_neg, mux82_b0_sel_is_0_o);
  binary_mux_s1_w1 mux83_b1 (
    .i0(n263[1]),
    .i1(1'b0),
    .sel(n93),
    .o(n264[1]));  // sources/rtl/camera_init.v(256)
  AL_MUX mux83_b10 (
    .i0(1'b0),
    .i1(n233[10]),
    .sel(mux83_b10_sel_is_2_o),
    .o(n264[10]));
  and mux83_b10_sel_is_2 (mux83_b10_sel_is_2_o, n93_neg, mux82_b10_sel_is_2_o);
  AL_MUX mux83_b11 (
    .i0(1'b0),
    .i1(n217[11]),
    .sel(mux83_b11_sel_is_2_o),
    .o(n264[11]));
  and mux83_b11_sel_is_2 (mux83_b11_sel_is_2_o, n93_neg, mux82_b11_sel_is_2_o);
  and mux83_b12_sel_is_2 (mux83_b12_sel_is_2_o, n93_neg, mux82_b12_sel_is_2_o);
  and mux83_b13_sel_is_2 (mux83_b13_sel_is_2_o, n93_neg, mux82_b13_sel_is_2_o);
  not mux83_b13_sel_is_2_o_inv (mux83_b13_sel_is_2_o_neg, mux83_b13_sel_is_2_o);
  AL_MUX mux83_b14 (
    .i0(1'b0),
    .i1(n219[14]),
    .sel(mux83_b12_sel_is_2_o),
    .o(n264[14]));
  AL_MUX mux83_b15 (
    .i0(1'b1),
    .i1(n197[15]),
    .sel(mux83_b15_sel_is_2_o),
    .o(n264[15]));
  and mux83_b15_sel_is_2 (mux83_b15_sel_is_2_o, n93_neg, mux82_b15_sel_is_2_o);
  binary_mux_s1_w1 mux83_b2 (
    .i0(n263[2]),
    .i1(1'b0),
    .sel(n93),
    .o(n264[2]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux83_b3 (
    .i0(n263[3]),
    .i1(1'b0),
    .sel(n93),
    .o(n264[3]));  // sources/rtl/camera_init.v(256)
  and mux83_b4_sel_is_0 (mux83_b4_sel_is_0_o, n93_neg, n94_neg);
  and mux83_b6_sel_is_2 (mux83_b6_sel_is_2_o, n93_neg, mux82_b6_sel_is_2_o);
  and mux83_b7_sel_is_2 (mux83_b7_sel_is_2_o, n93_neg, mux82_b7_sel_is_2_o);
  binary_mux_s1_w1 mux83_b8 (
    .i0(n263[8]),
    .i1(1'b0),
    .sel(n93),
    .o(n264[8]));  // sources/rtl/camera_init.v(256)
  and mux83_b9_sel_is_2 (mux83_b9_sel_is_2_o, n93_neg, mux82_b9_sel_is_2_o);
  and mux84_b0_sel_is_2 (mux84_b0_sel_is_2_o, n92_neg, mux83_b0_sel_is_2_o);
  binary_mux_s1_w1 mux84_b1 (
    .i0(n264[1]),
    .i1(1'b1),
    .sel(n92),
    .o(n265[1]));  // sources/rtl/camera_init.v(256)
  and mux84_b12_sel_is_2 (mux84_b12_sel_is_2_o, n92_neg, mux83_b12_sel_is_2_o);
  and mux84_b13_sel_is_0 (mux84_b13_sel_is_0_o, n92_neg, mux83_b13_sel_is_2_o_neg);
  binary_mux_s1_w1 mux84_b2 (
    .i0(n264[2]),
    .i1(1'b1),
    .sel(n92),
    .o(n265[2]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux84_b3 (
    .i0(n264[3]),
    .i1(1'b1),
    .sel(n92),
    .o(n265[3]));  // sources/rtl/camera_init.v(256)
  AL_MUX mux84_b4 (
    .i0(1'b0),
    .i1(n262[4]),
    .sel(mux84_b4_sel_is_2_o),
    .o(n265[4]));
  and mux84_b4_sel_is_2 (mux84_b4_sel_is_2_o, n92_neg, mux83_b4_sel_is_0_o);
  and mux84_b6_sel_is_2 (mux84_b6_sel_is_2_o, n92_neg, mux83_b6_sel_is_2_o);
  and mux84_b7_sel_is_2 (mux84_b7_sel_is_2_o, n92_neg, mux83_b7_sel_is_2_o);
  and mux84_b9_sel_is_2 (mux84_b9_sel_is_2_o, n92_neg, mux83_b9_sel_is_2_o);
  and mux85_b0_sel_is_2 (mux85_b0_sel_is_2_o, n91_neg, mux84_b0_sel_is_2_o);
  and mux85_b10_sel_is_0 (mux85_b10_sel_is_0_o, n91_neg, n92_neg);
  and mux85_b12_sel_is_2 (mux85_b12_sel_is_2_o, n91_neg, mux84_b12_sel_is_2_o);
  and mux85_b13_sel_is_2 (mux85_b13_sel_is_2_o, n91_neg, mux84_b13_sel_is_0_o);
  binary_mux_s1_w1 mux85_b4 (
    .i0(n265[4]),
    .i1(1'b1),
    .sel(n91),
    .o(n266[4]));  // sources/rtl/camera_init.v(256)
  AL_MUX mux85_b5 (
    .i0(1'b0),
    .i1(n261[5]),
    .sel(mux85_b0_sel_is_2_o),
    .o(n266[5]));
  and mux85_b6_sel_is_2 (mux85_b6_sel_is_2_o, n91_neg, mux84_b6_sel_is_2_o);
  and mux85_b7_sel_is_2 (mux85_b7_sel_is_2_o, n91_neg, mux84_b7_sel_is_2_o);
  and mux85_b9_sel_is_2 (mux85_b9_sel_is_2_o, n91_neg, mux84_b9_sel_is_2_o);
  and mux86_b0_sel_is_2 (mux86_b0_sel_is_2_o, n90_neg, mux85_b0_sel_is_2_o);
  and mux86_b10_sel_is_2 (mux86_b10_sel_is_2_o, n90_neg, mux85_b10_sel_is_0_o);
  and mux86_b12_sel_is_2 (mux86_b12_sel_is_2_o, n90_neg, mux85_b12_sel_is_2_o);
  and mux86_b13_sel_is_2 (mux86_b13_sel_is_2_o, n90_neg, mux85_b13_sel_is_2_o);
  and mux86_b1_sel_is_0 (mux86_b1_sel_is_0_o, n90_neg, n91_neg);
  AL_MUX mux86_b3 (
    .i0(1'b0),
    .i1(n265[3]),
    .sel(mux86_b1_sel_is_0_o),
    .o(n267[3]));
  binary_mux_s1_w1 mux86_b5 (
    .i0(n266[5]),
    .i1(1'b1),
    .sel(n90),
    .o(n267[5]));  // sources/rtl/camera_init.v(256)
  and mux86_b6_sel_is_2 (mux86_b6_sel_is_2_o, n90_neg, mux85_b6_sel_is_2_o);
  and mux86_b7_sel_is_2 (mux86_b7_sel_is_2_o, n90_neg, mux85_b7_sel_is_2_o);
  AL_MUX mux86_b8 (
    .i0(1'b1),
    .i1(n264[8]),
    .sel(mux86_b10_sel_is_2_o),
    .o(n267[8]));
  and mux86_b9_sel_is_2 (mux86_b9_sel_is_2_o, n90_neg, mux85_b9_sel_is_2_o);
  and mux87_b0_sel_is_2 (mux87_b0_sel_is_2_o, n89_neg, mux86_b0_sel_is_2_o);
  and mux87_b10_sel_is_2 (mux87_b10_sel_is_2_o, n89_neg, mux86_b10_sel_is_2_o);
  and mux87_b12_sel_is_2 (mux87_b12_sel_is_2_o, n89_neg, mux86_b12_sel_is_2_o);
  and mux87_b13_sel_is_2 (mux87_b13_sel_is_2_o, n89_neg, mux86_b13_sel_is_2_o);
  and mux87_b1_sel_is_2 (mux87_b1_sel_is_2_o, n89_neg, mux86_b1_sel_is_0_o);
  and mux87_b4_sel_is_0 (mux87_b4_sel_is_0_o, n89_neg, n90_neg);
  AL_MUX mux87_b6 (
    .i0(1'b0),
    .i1(n260[6]),
    .sel(mux87_b6_sel_is_2_o),
    .o(n268[6]));
  and mux87_b6_sel_is_2 (mux87_b6_sel_is_2_o, n89_neg, mux86_b6_sel_is_2_o);
  and mux87_b7_sel_is_2 (mux87_b7_sel_is_2_o, n89_neg, mux86_b7_sel_is_2_o);
  binary_mux_s1_w1 mux87_b8 (
    .i0(n267[8]),
    .i1(1'b0),
    .sel(n89),
    .o(n268[8]));  // sources/rtl/camera_init.v(256)
  and mux87_b9_sel_is_2 (mux87_b9_sel_is_2_o, n89_neg, mux86_b9_sel_is_2_o);
  and mux88_b0_sel_is_2 (mux88_b0_sel_is_2_o, n88_neg, mux87_b0_sel_is_2_o);
  and mux88_b10_sel_is_2 (mux88_b10_sel_is_2_o, n88_neg, mux87_b10_sel_is_2_o);
  and mux88_b12_sel_is_2 (mux88_b12_sel_is_2_o, n88_neg, mux87_b12_sel_is_2_o);
  and mux88_b13_sel_is_2 (mux88_b13_sel_is_2_o, n88_neg, mux87_b13_sel_is_2_o);
  and mux88_b1_sel_is_2 (mux88_b1_sel_is_2_o, n88_neg, mux87_b1_sel_is_2_o);
  and mux88_b3_sel_is_0 (mux88_b3_sel_is_0_o, n88_neg, n89_neg);
  and mux88_b4_sel_is_2 (mux88_b4_sel_is_2_o, n88_neg, mux87_b4_sel_is_0_o);
  and mux88_b7_sel_is_2 (mux88_b7_sel_is_2_o, n88_neg, mux87_b7_sel_is_2_o);
  and mux88_b9_sel_is_2 (mux88_b9_sel_is_2_o, n88_neg, mux87_b9_sel_is_2_o);
  AL_MUX mux89_b0 (
    .i0(1'b0),
    .i1(n261[0]),
    .sel(mux89_b0_sel_is_2_o),
    .o(n270[0]));
  and mux89_b0_sel_is_2 (mux89_b0_sel_is_2_o, n87_neg, mux88_b0_sel_is_2_o);
  AL_MUX mux89_b1 (
    .i0(1'b0),
    .i1(n265[1]),
    .sel(mux89_b1_sel_is_2_o),
    .o(n270[1]));
  and mux89_b10_sel_is_2 (mux89_b10_sel_is_2_o, n87_neg, mux88_b10_sel_is_2_o);
  and mux89_b12_sel_is_2 (mux89_b12_sel_is_2_o, n87_neg, mux88_b12_sel_is_2_o);
  and mux89_b13_sel_is_2 (mux89_b13_sel_is_2_o, n87_neg, mux88_b13_sel_is_2_o);
  and mux89_b1_sel_is_2 (mux89_b1_sel_is_2_o, n87_neg, mux88_b1_sel_is_2_o);
  AL_MUX mux89_b3 (
    .i0(1'b1),
    .i1(n267[3]),
    .sel(mux89_b3_sel_is_2_o),
    .o(n270[3]));
  and mux89_b3_sel_is_2 (mux89_b3_sel_is_2_o, n87_neg, mux88_b3_sel_is_0_o);
  and mux89_b4_sel_is_2 (mux89_b4_sel_is_2_o, n87_neg, mux88_b4_sel_is_2_o);
  AL_MUX mux89_b6 (
    .i0(1'b1),
    .i1(n268[6]),
    .sel(mux89_b6_sel_is_0_o),
    .o(n270[6]));
  and mux89_b6_sel_is_0 (mux89_b6_sel_is_0_o, n87_neg, n88_neg);
  and mux89_b7_sel_is_2 (mux89_b7_sel_is_2_o, n87_neg, mux88_b7_sel_is_2_o);
  AL_MUX mux89_b8 (
    .i0(1'b1),
    .i1(n268[8]),
    .sel(mux89_b6_sel_is_0_o),
    .o(n270[8]));
  and mux89_b9_sel_is_2 (mux89_b9_sel_is_2_o, n87_neg, mux88_b9_sel_is_2_o);
  AL_MUX mux8_b0 (
    .i0(1'b0),
    .i1(n187[0]),
    .sel(mux8_b0_sel_is_0_o),
    .o(n189[0]));
  and mux8_b0_sel_is_0 (mux8_b0_sel_is_0_o, n168_neg, n169_neg);
  binary_mux_s1_w1 mux8_b10 (
    .i0(n188[10]),
    .i1(1'b1),
    .sel(n168),
    .o(n189[10]));  // sources/rtl/camera_init.v(256)
  and mux8_b13_sel_is_2 (mux8_b13_sel_is_2_o, n168_neg, mux7_b13_sel_is_2_o);
  and mux8_b14_sel_is_2 (mux8_b14_sel_is_2_o, n168_neg, mux7_b14_sel_is_2_o);
  AL_MUX mux8_b3 (
    .i0(1'b0),
    .i1(n187[3]),
    .sel(mux8_b0_sel_is_0_o),
    .o(n189[3]));
  and mux8_b4_sel_is_2 (mux8_b4_sel_is_2_o, n168_neg, mux7_b4_sel_is_2_o);
  AL_MUX mux8_b5 (
    .i0(1'b0),
    .i1(n187[5]),
    .sel(mux8_b0_sel_is_0_o),
    .o(n189[5]));
  binary_mux_s1_w1 mux8_b8 (
    .i0(n188[8]),
    .i1(1'b0),
    .sel(n168),
    .o(n189[8]));  // sources/rtl/camera_init.v(256)
  and mux8_b9_sel_is_0 (mux8_b9_sel_is_0_o, n168_neg, mux7_b9_sel_is_2_o_neg);
  not mux8_b9_sel_is_0_o_inv (mux8_b9_sel_is_0_o_neg, mux8_b9_sel_is_0_o);
  binary_mux_s1_w1 mux90_b0 (
    .i0(n270[0]),
    .i1(1'b1),
    .sel(n86),
    .o(n271[0]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux90_b1 (
    .i0(n270[1]),
    .i1(1'b1),
    .sel(n86),
    .o(n271[1]));  // sources/rtl/camera_init.v(256)
  and mux90_b10_sel_is_2 (mux90_b10_sel_is_2_o, n86_neg, mux89_b10_sel_is_2_o);
  and mux90_b12_sel_is_2 (mux90_b12_sel_is_2_o, n86_neg, mux89_b12_sel_is_2_o);
  and mux90_b13_sel_is_2 (mux90_b13_sel_is_2_o, n86_neg, mux89_b13_sel_is_2_o);
  and mux90_b2_sel_is_2 (mux90_b2_sel_is_2_o, n86_neg, mux89_b1_sel_is_2_o);
  and mux90_b4_sel_is_2 (mux90_b4_sel_is_2_o, n86_neg, mux89_b4_sel_is_2_o);
  and mux90_b5_sel_is_2 (mux90_b5_sel_is_2_o, n86_neg, mux89_b3_sel_is_2_o);
  and mux90_b7_sel_is_2 (mux90_b7_sel_is_2_o, n86_neg, mux89_b7_sel_is_2_o);
  binary_mux_s1_w1 mux90_b8 (
    .i0(n270[8]),
    .i1(1'b0),
    .sel(n86),
    .o(n271[8]));  // sources/rtl/camera_init.v(256)
  and mux90_b9_sel_is_2 (mux90_b9_sel_is_2_o, n86_neg, mux89_b9_sel_is_2_o);
  and mux91_b10_sel_is_2 (mux91_b10_sel_is_2_o, n85_neg, mux90_b10_sel_is_2_o);
  and mux91_b12_sel_is_2 (mux91_b12_sel_is_2_o, n85_neg, mux90_b12_sel_is_2_o);
  and mux91_b13_sel_is_2 (mux91_b13_sel_is_2_o, n85_neg, mux90_b13_sel_is_2_o);
  and mux91_b2_sel_is_2 (mux91_b2_sel_is_2_o, n85_neg, mux90_b2_sel_is_2_o);
  and mux91_b3_sel_is_0 (mux91_b3_sel_is_0_o, n85_neg, n86_neg);
  and mux91_b4_sel_is_2 (mux91_b4_sel_is_2_o, n85_neg, mux90_b4_sel_is_2_o);
  and mux91_b5_sel_is_2 (mux91_b5_sel_is_2_o, n85_neg, mux90_b5_sel_is_2_o);
  and mux91_b7_sel_is_2 (mux91_b7_sel_is_2_o, n85_neg, mux90_b7_sel_is_2_o);
  binary_mux_s1_w1 mux91_b8 (
    .i0(n271[8]),
    .i1(1'b1),
    .sel(n85),
    .o(n272[8]));  // sources/rtl/camera_init.v(256)
  and mux91_b9_sel_is_2 (mux91_b9_sel_is_2_o, n85_neg, mux90_b9_sel_is_2_o);
  and mux92_b0_sel_is_0 (mux92_b0_sel_is_0_o, n84_neg, n85_neg);
  AL_MUX mux92_b10 (
    .i0(1'b1),
    .i1(n264[10]),
    .sel(mux92_b10_sel_is_2_o),
    .o(n273[10]));
  and mux92_b10_sel_is_2 (mux92_b10_sel_is_2_o, n84_neg, mux91_b10_sel_is_2_o);
  AL_MUX mux92_b12 (
    .i0(1'b1),
    .i1(n219[12]),
    .sel(mux92_b12_sel_is_2_o),
    .o(n273[12]));
  and mux92_b12_sel_is_2 (mux92_b12_sel_is_2_o, n84_neg, mux91_b12_sel_is_2_o);
  and mux92_b13_sel_is_2 (mux92_b13_sel_is_2_o, n84_neg, mux91_b13_sel_is_2_o);
  not mux92_b13_sel_is_2_o_inv (mux92_b13_sel_is_2_o_neg, mux92_b13_sel_is_2_o);
  AL_MUX mux92_b15 (
    .i0(1'b0),
    .i1(n264[15]),
    .sel(mux92_b10_sel_is_2_o),
    .o(n273[15]));
  and mux92_b2_sel_is_2 (mux92_b2_sel_is_2_o, n84_neg, mux91_b2_sel_is_2_o);
  and mux92_b3_sel_is_2 (mux92_b3_sel_is_2_o, n84_neg, mux91_b3_sel_is_0_o);
  and mux92_b4_sel_is_2 (mux92_b4_sel_is_2_o, n84_neg, mux91_b4_sel_is_2_o);
  and mux92_b5_sel_is_2 (mux92_b5_sel_is_2_o, n84_neg, mux91_b5_sel_is_2_o);
  AL_MUX mux92_b7 (
    .i0(1'b0),
    .i1(n256[7]),
    .sel(mux92_b7_sel_is_2_o),
    .o(n273[7]));
  and mux92_b7_sel_is_2 (mux92_b7_sel_is_2_o, n84_neg, mux91_b7_sel_is_2_o);
  binary_mux_s1_w1 mux92_b8 (
    .i0(n272[8]),
    .i1(1'b0),
    .sel(n84),
    .o(n273[8]));  // sources/rtl/camera_init.v(256)
  and mux92_b9_sel_is_2 (mux92_b9_sel_is_2_o, n84_neg, mux91_b9_sel_is_2_o);
  and mux93_b0_sel_is_2 (mux93_b0_sel_is_2_o, n83_neg, mux92_b0_sel_is_0_o);
  and mux93_b11_sel_is_2 (mux93_b11_sel_is_2_o, n83_neg, mux92_b10_sel_is_2_o);
  and mux93_b13_sel_is_0 (mux93_b13_sel_is_0_o, n83_neg, mux92_b13_sel_is_2_o_neg);
  and mux93_b2_sel_is_2 (mux93_b2_sel_is_2_o, n83_neg, mux92_b2_sel_is_2_o);
  AL_MUX mux93_b3 (
    .i0(1'b0),
    .i1(n270[3]),
    .sel(mux93_b3_sel_is_2_o),
    .o(n274[3]));
  and mux93_b3_sel_is_2 (mux93_b3_sel_is_2_o, n83_neg, mux92_b3_sel_is_2_o);
  and mux93_b4_sel_is_2 (mux93_b4_sel_is_2_o, n83_neg, mux92_b4_sel_is_2_o);
  and mux93_b5_sel_is_2 (mux93_b5_sel_is_2_o, n83_neg, mux92_b5_sel_is_2_o);
  binary_mux_s1_w1 mux93_b7 (
    .i0(n273[7]),
    .i1(1'b1),
    .sel(n83),
    .o(n274[7]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux93_b8 (
    .i0(n273[8]),
    .i1(1'b1),
    .sel(n83),
    .o(n274[8]));  // sources/rtl/camera_init.v(256)
  and mux93_b9_sel_is_2 (mux93_b9_sel_is_2_o, n83_neg, mux92_b9_sel_is_2_o);
  and mux94_b0_sel_is_2 (mux94_b0_sel_is_2_o, n82_neg, mux93_b0_sel_is_2_o);
  AL_MUX mux94_b1 (
    .i0(1'b0),
    .i1(n271[1]),
    .sel(mux94_b0_sel_is_2_o),
    .o(n275[1]));
  and mux94_b10_sel_is_0 (mux94_b10_sel_is_0_o, n82_neg, n83_neg);
  AL_MUX mux94_b11 (
    .i0(1'b1),
    .i1(n264[11]),
    .sel(mux94_b11_sel_is_2_o),
    .o(n275[11]));
  and mux94_b11_sel_is_2 (mux94_b11_sel_is_2_o, n82_neg, mux93_b11_sel_is_2_o);
  AL_MUX mux94_b12 (
    .i0(1'b0),
    .i1(n273[12]),
    .sel(mux94_b10_sel_is_0_o),
    .o(n275[12]));
  and mux94_b13_sel_is_2 (mux94_b13_sel_is_2_o, n82_neg, mux93_b13_sel_is_0_o);
  and mux94_b2_sel_is_2 (mux94_b2_sel_is_2_o, n82_neg, mux93_b2_sel_is_2_o);
  binary_mux_s1_w1 mux94_b3 (
    .i0(n274[3]),
    .i1(1'b1),
    .sel(n82),
    .o(n275[3]));  // sources/rtl/camera_init.v(256)
  and mux94_b4_sel_is_2 (mux94_b4_sel_is_2_o, n82_neg, mux93_b4_sel_is_2_o);
  and mux94_b5_sel_is_2 (mux94_b5_sel_is_2_o, n82_neg, mux93_b5_sel_is_2_o);
  and mux94_b6_sel_is_2 (mux94_b6_sel_is_2_o, n82_neg, mux93_b3_sel_is_2_o);
  binary_mux_s1_w1 mux94_b7 (
    .i0(n274[7]),
    .i1(1'b0),
    .sel(n82),
    .o(n275[7]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux94_b8 (
    .i0(n274[8]),
    .i1(1'b0),
    .sel(n82),
    .o(n275[8]));  // sources/rtl/camera_init.v(256)
  and mux94_b9_sel_is_2 (mux94_b9_sel_is_2_o, n82_neg, mux93_b9_sel_is_2_o);
  not mux94_b9_sel_is_2_o_inv (mux94_b9_sel_is_2_o_neg, mux94_b9_sel_is_2_o);
  and mux95_b0_sel_is_2 (mux95_b0_sel_is_2_o, n81_neg, mux94_b0_sel_is_2_o);
  binary_mux_s1_w1 mux95_b1 (
    .i0(n275[1]),
    .i1(1'b1),
    .sel(n81),
    .o(n276[1]));  // sources/rtl/camera_init.v(256)
  and mux95_b10_sel_is_2 (mux95_b10_sel_is_2_o, n81_neg, mux94_b10_sel_is_0_o);
  binary_mux_s1_w1 mux95_b11 (
    .i0(n275[11]),
    .i1(1'b0),
    .sel(n81),
    .o(n276[11]));  // sources/rtl/camera_init.v(256)
  and mux95_b13_sel_is_2 (mux95_b13_sel_is_2_o, n81_neg, mux94_b13_sel_is_2_o);
  and mux95_b14_sel_is_2 (mux95_b14_sel_is_2_o, n81_neg, mux94_b11_sel_is_2_o);
  and mux95_b2_sel_is_2 (mux95_b2_sel_is_2_o, n81_neg, mux94_b2_sel_is_2_o);
  AL_MUX mux95_b4 (
    .i0(1'b0),
    .i1(n266[4]),
    .sel(mux95_b4_sel_is_2_o),
    .o(n276[4]));
  and mux95_b4_sel_is_2 (mux95_b4_sel_is_2_o, n81_neg, mux94_b4_sel_is_2_o);
  and mux95_b5_sel_is_2 (mux95_b5_sel_is_2_o, n81_neg, mux94_b5_sel_is_2_o);
  and mux95_b6_sel_is_2 (mux95_b6_sel_is_2_o, n81_neg, mux94_b6_sel_is_2_o);
  binary_mux_s1_w1 mux95_b7 (
    .i0(n275[7]),
    .i1(1'b1),
    .sel(n81),
    .o(n276[7]));  // sources/rtl/camera_init.v(256)
  and mux95_b9_sel_is_0 (mux95_b9_sel_is_0_o, n81_neg, mux94_b9_sel_is_2_o_neg);
  not mux95_b9_sel_is_0_o_inv (mux95_b9_sel_is_0_o_neg, mux95_b9_sel_is_0_o);
  AL_MUX mux96_b0 (
    .i0(1'b0),
    .i1(n271[0]),
    .sel(mux96_b0_sel_is_2_o),
    .o(n277[0]));
  and mux96_b0_sel_is_2 (mux96_b0_sel_is_2_o, n80_neg, mux95_b0_sel_is_2_o);
  binary_mux_s1_w1 mux96_b1 (
    .i0(n276[1]),
    .i1(1'b0),
    .sel(n80),
    .o(n277[1]));  // sources/rtl/camera_init.v(256)
  AL_MUX mux96_b10 (
    .i0(1'b0),
    .i1(n273[10]),
    .sel(mux96_b10_sel_is_2_o),
    .o(n277[10]));
  and mux96_b10_sel_is_2 (mux96_b10_sel_is_2_o, n80_neg, mux95_b10_sel_is_2_o);
  binary_mux_s1_w1 mux96_b11 (
    .i0(n276[11]),
    .i1(1'b1),
    .sel(n80),
    .o(n277[11]));  // sources/rtl/camera_init.v(256)
  and mux96_b12_sel_is_0 (mux96_b12_sel_is_0_o, n80_neg, n81_neg);
  and mux96_b13_sel_is_2 (mux96_b13_sel_is_2_o, n80_neg, mux95_b13_sel_is_2_o);
  and mux96_b14_sel_is_2 (mux96_b14_sel_is_2_o, n80_neg, mux95_b14_sel_is_2_o);
  and mux96_b2_sel_is_2 (mux96_b2_sel_is_2_o, n80_neg, mux95_b2_sel_is_2_o);
  binary_mux_s1_w1 mux96_b4 (
    .i0(n276[4]),
    .i1(1'b1),
    .sel(n80),
    .o(n277[4]));  // sources/rtl/camera_init.v(256)
  and mux96_b5_sel_is_2 (mux96_b5_sel_is_2_o, n80_neg, mux95_b5_sel_is_2_o);
  and mux96_b6_sel_is_2 (mux96_b6_sel_is_2_o, n80_neg, mux95_b6_sel_is_2_o);
  and mux96_b9_sel_is_0 (mux96_b9_sel_is_0_o, n80_neg, mux95_b9_sel_is_0_o_neg);
  not mux96_b9_sel_is_0_o_inv (mux96_b9_sel_is_0_o_neg, mux96_b9_sel_is_0_o);
  binary_mux_s1_w1 mux97_b10 (
    .i0(n277[10]),
    .i1(1'b1),
    .sel(n79),
    .o(n278[10]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux97_b11 (
    .i0(n277[11]),
    .i1(1'b0),
    .sel(n79),
    .o(n278[11]));  // sources/rtl/camera_init.v(256)
  AL_MUX mux97_b12 (
    .i0(1'b1),
    .i1(n275[12]),
    .sel(mux97_b12_sel_is_2_o),
    .o(n278[12]));
  and mux97_b12_sel_is_2 (mux97_b12_sel_is_2_o, n79_neg, mux96_b12_sel_is_0_o);
  and mux97_b13_sel_is_2 (mux97_b13_sel_is_2_o, n79_neg, mux96_b13_sel_is_2_o);
  AL_MUX mux97_b14 (
    .i0(1'b1),
    .i1(n264[14]),
    .sel(mux97_b14_sel_is_2_o),
    .o(n278[14]));
  and mux97_b14_sel_is_2 (mux97_b14_sel_is_2_o, n79_neg, mux96_b14_sel_is_2_o);
  and mux97_b15_sel_is_2 (mux97_b15_sel_is_2_o, n79_neg, mux96_b10_sel_is_2_o);
  AL_MUX mux97_b2 (
    .i0(1'b0),
    .i1(n265[2]),
    .sel(mux97_b2_sel_is_2_o),
    .o(n278[2]));
  and mux97_b2_sel_is_2 (mux97_b2_sel_is_2_o, n79_neg, mux96_b2_sel_is_2_o);
  AL_MUX mux97_b3 (
    .i0(1'b0),
    .i1(n275[3]),
    .sel(mux97_b12_sel_is_2_o),
    .o(n278[3]));
  binary_mux_s1_w1 mux97_b4 (
    .i0(n277[4]),
    .i1(1'b0),
    .sel(n79),
    .o(n278[4]));  // sources/rtl/camera_init.v(256)
  AL_MUX mux97_b5 (
    .i0(1'b0),
    .i1(n267[5]),
    .sel(mux97_b5_sel_is_2_o),
    .o(n278[5]));
  and mux97_b5_sel_is_2 (mux97_b5_sel_is_2_o, n79_neg, mux96_b5_sel_is_2_o);
  and mux97_b6_sel_is_2 (mux97_b6_sel_is_2_o, n79_neg, mux96_b6_sel_is_2_o);
  and mux97_b7_sel_is_0 (mux97_b7_sel_is_0_o, n79_neg, n80_neg);
  AL_MUX mux97_b8 (
    .i0(1'b1),
    .i1(n275[8]),
    .sel(mux97_b12_sel_is_2_o),
    .o(n278[8]));
  and mux97_b9_sel_is_0 (mux97_b9_sel_is_0_o, n79_neg, mux96_b9_sel_is_0_o_neg);
  not mux97_b9_sel_is_0_o_inv (mux97_b9_sel_is_0_o_neg, mux97_b9_sel_is_0_o);
  and mux98_b0_sel_is_0 (mux98_b0_sel_is_0_o, n78_neg, n79_neg);
  AL_MUX mux98_b1 (
    .i0(1'b1),
    .i1(n277[1]),
    .sel(mux98_b0_sel_is_0_o),
    .o(n279[1]));
  binary_mux_s1_w1 mux98_b10 (
    .i0(n278[10]),
    .i1(1'b0),
    .sel(n78),
    .o(n279[10]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux98_b11 (
    .i0(n278[11]),
    .i1(1'b1),
    .sel(n78),
    .o(n279[11]));  // sources/rtl/camera_init.v(256)
  and mux98_b13_sel_is_2 (mux98_b13_sel_is_2_o, n78_neg, mux97_b13_sel_is_2_o);
  and mux98_b15_sel_is_2 (mux98_b15_sel_is_2_o, n78_neg, mux97_b15_sel_is_2_o);
  binary_mux_s1_w1 mux98_b3 (
    .i0(n278[3]),
    .i1(1'b1),
    .sel(n78),
    .o(n279[3]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux98_b5 (
    .i0(n278[5]),
    .i1(1'b1),
    .sel(n78),
    .o(n279[5]));  // sources/rtl/camera_init.v(256)
  AL_MUX mux98_b6 (
    .i0(1'b0),
    .i1(n270[6]),
    .sel(mux98_b6_sel_is_2_o),
    .o(n279[6]));
  and mux98_b6_sel_is_2 (mux98_b6_sel_is_2_o, n78_neg, mux97_b6_sel_is_2_o);
  AL_MUX mux98_b7 (
    .i0(1'b0),
    .i1(n276[7]),
    .sel(mux98_b7_sel_is_2_o),
    .o(n279[7]));
  and mux98_b7_sel_is_2 (mux98_b7_sel_is_2_o, n78_neg, mux97_b7_sel_is_0_o);
  binary_mux_s1_w1 mux98_b8 (
    .i0(n278[8]),
    .i1(1'b0),
    .sel(n78),
    .o(n279[8]));  // sources/rtl/camera_init.v(256)
  and mux98_b9_sel_is_0 (mux98_b9_sel_is_0_o, n78_neg, mux97_b9_sel_is_0_o_neg);
  not mux98_b9_sel_is_0_o_inv (mux98_b9_sel_is_0_o_neg, mux98_b9_sel_is_0_o);
  AL_MUX mux99_b0 (
    .i0(1'b1),
    .i1(n277[0]),
    .sel(mux99_b0_sel_is_2_o),
    .o(n280[0]));
  and mux99_b0_sel_is_2 (mux99_b0_sel_is_2_o, n77_neg, mux98_b0_sel_is_0_o);
  binary_mux_s1_w1 mux99_b11 (
    .i0(n279[11]),
    .i1(1'b0),
    .sel(n77),
    .o(n280[11]));  // sources/rtl/camera_init.v(256)
  and mux99_b12_sel_is_0 (mux99_b12_sel_is_0_o, n77_neg, n78_neg);
  and mux99_b13_sel_is_2 (mux99_b13_sel_is_2_o, n77_neg, mux98_b13_sel_is_2_o);
  AL_MUX mux99_b14 (
    .i0(1'b0),
    .i1(n278[14]),
    .sel(mux99_b12_sel_is_0_o),
    .o(n280[14]));
  AL_MUX mux99_b15 (
    .i0(1'b1),
    .i1(n273[15]),
    .sel(mux99_b15_sel_is_2_o),
    .o(n280[15]));
  and mux99_b15_sel_is_2 (mux99_b15_sel_is_2_o, n77_neg, mux98_b15_sel_is_2_o);
  AL_MUX mux99_b2 (
    .i0(1'b1),
    .i1(n278[2]),
    .sel(mux99_b12_sel_is_0_o),
    .o(n280[2]));
  AL_MUX mux99_b4 (
    .i0(1'b1),
    .i1(n278[4]),
    .sel(mux99_b12_sel_is_0_o),
    .o(n280[4]));
  binary_mux_s1_w1 mux99_b6 (
    .i0(n279[6]),
    .i1(1'b1),
    .sel(n77),
    .o(n280[6]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux99_b7 (
    .i0(n279[7]),
    .i1(1'b1),
    .sel(n77),
    .o(n280[7]));  // sources/rtl/camera_init.v(256)
  binary_mux_s1_w1 mux99_b8 (
    .i0(n279[8]),
    .i1(1'b1),
    .sel(n77),
    .o(n280[8]));  // sources/rtl/camera_init.v(256)
  and mux99_b9_sel_is_0 (mux99_b9_sel_is_0_o, n77_neg, mux98_b9_sel_is_0_o_neg);
  not mux99_b9_sel_is_0_o_inv (mux99_b9_sel_is_0_o_neg, mux99_b9_sel_is_0_o);
  binary_mux_s1_w1 mux9_b0 (
    .i0(n189[0]),
    .i1(1'b1),
    .sel(n167),
    .o(n190[0]));  // sources/rtl/camera_init.v(256)
  AL_MUX mux9_b1 (
    .i0(1'b0),
    .i1(n188[1]),
    .sel(mux9_b11_sel_is_0_o),
    .o(n190[1]));
  and mux9_b11_sel_is_0 (mux9_b11_sel_is_0_o, n167_neg, n168_neg);
  and mux9_b12_sel_is_2 (mux9_b12_sel_is_2_o, n167_neg, mux8_b0_sel_is_0_o);
  and mux9_b13_sel_is_2 (mux9_b13_sel_is_2_o, n167_neg, mux8_b13_sel_is_2_o);
  and mux9_b14_sel_is_2 (mux9_b14_sel_is_2_o, n167_neg, mux8_b14_sel_is_2_o);
  binary_mux_s1_w1 mux9_b3 (
    .i0(n189[3]),
    .i1(1'b1),
    .sel(n167),
    .o(n190[3]));  // sources/rtl/camera_init.v(256)
  AL_MUX mux9_b4 (
    .i0(1'b0),
    .i1(n184[3]),
    .sel(mux9_b4_sel_is_2_o),
    .o(n190[4]));
  and mux9_b4_sel_is_2 (mux9_b4_sel_is_2_o, n167_neg, mux8_b4_sel_is_2_o);
  binary_mux_s1_w1 mux9_b8 (
    .i0(n189[8]),
    .i1(1'b1),
    .sel(n167),
    .o(n190[8]));  // sources/rtl/camera_init.v(256)
  and mux9_b9_sel_is_0 (mux9_b9_sel_is_0_o, n167_neg, mux8_b9_sel_is_0_o_neg);
  not n100_inv (n100_neg, n100);
  not n101_inv (n101_neg, n101);
  not n102_inv (n102_neg, n102);
  not n103_inv (n103_neg, n103);
  not n104_inv (n104_neg, n104);
  not n105_inv (n105_neg, n105);
  not n106_inv (n106_neg, n106);
  not n107_inv (n107_neg, n107);
  not n108_inv (n108_neg, n108);
  not n109_inv (n109_neg, n109);
  not n10_inv (n10_neg, n10);
  not n110_inv (n110_neg, n110);
  not n111_inv (n111_neg, n111);
  not n112_inv (n112_neg, n112);
  not n113_inv (n113_neg, n113);
  not n114_inv (n114_neg, n114);
  not n115_inv (n115_neg, n115);
  not n116_inv (n116_neg, n116);
  not n117_inv (n117_neg, n117);
  not n118_inv (n118_neg, n118);
  not n119_inv (n119_neg, n119);
  not n11_inv (n11_neg, n11);
  not n120_inv (n120_neg, n120);
  not n121_inv (n121_neg, n121);
  not n122_inv (n122_neg, n122);
  not n123_inv (n123_neg, n123);
  not n124_inv (n124_neg, n124);
  not n125_inv (n125_neg, n125);
  not n126_inv (n126_neg, n126);
  not n127_inv (n127_neg, n127);
  not n128_inv (n128_neg, n128);
  not n129_inv (n129_neg, n129);
  not n12_inv (n12_neg, n12);
  not n130_inv (n130_neg, n130);
  not n131_inv (n131_neg, n131);
  not n132_inv (n132_neg, n132);
  not n133_inv (n133_neg, n133);
  not n134_inv (n134_neg, n134);
  not n135_inv (n135_neg, n135);
  not n136_inv (n136_neg, n136);
  not n137_inv (n137_neg, n137);
  not n138_inv (n138_neg, n138);
  not n139_inv (n139_neg, n139);
  not n13_inv (n13_neg, n13);
  not n140_inv (n140_neg, n140);
  not n141_inv (n141_neg, n141);
  not n142_inv (n142_neg, n142);
  not n143_inv (n143_neg, n143);
  not n144_inv (n144_neg, n144);
  not n145_inv (n145_neg, n145);
  not n146_inv (n146_neg, n146);
  not n147_inv (n147_neg, n147);
  not n148_inv (n148_neg, n148);
  not n149_inv (n149_neg, n149);
  not n14_inv (n14_neg, n14);
  not n150_inv (n150_neg, n150);
  not n151_inv (n151_neg, n151);
  not n152_inv (n152_neg, n152);
  not n153_inv (n153_neg, n153);
  not n154_inv (n154_neg, n154);
  not n155_inv (n155_neg, n155);
  not n156_inv (n156_neg, n156);
  not n157_inv (n157_neg, n157);
  not n158_inv (n158_neg, n158);
  not n159_inv (n159_neg, n159);
  not n15_inv (n15_neg, n15);
  not n160_inv (n160_neg, n160);
  not n161_inv (n161_neg, n161);
  not n162_inv (n162_neg, n162);
  not n163_inv (n163_neg, n163);
  not n164_inv (n164_neg, n164);
  not n165_inv (n165_neg, n165);
  not n166_inv (n166_neg, n166);
  not n167_inv (n167_neg, n167);
  not n168_inv (n168_neg, n168);
  not n169_inv (n169_neg, n169);
  not n16_inv (n16_neg, n16);
  not n170_inv (n170_neg, n170);
  not n171_inv (n171_neg, n171);
  not n172_inv (n172_neg, n172);
  not n173_inv (n173_neg, n173);
  not n174_inv (n174_neg, n174);
  not n175_inv (n175_neg, n175);
  not n176_inv (n176_neg, n176);
  not n17_inv (n17_neg, n17);
  not n18_inv (n18_neg, n18);
  not n19_inv (n19_neg, n19);
  not n1_inv (n1_neg, n1);
  not n20_inv (n20_neg, n20);
  not n21_inv (n21_neg, n21);
  not n22_inv (n22_neg, n22);
  not n23_inv (n23_neg, n23);
  not n24_inv (n24_neg, n24);
  not n25_inv (n25_neg, n25);
  not n26_inv (n26_neg, n26);
  not n27_inv (n27_neg, n27);
  not n28_inv (n28_neg, n28);
  not n29_inv (n29_neg, n29);
  not n2_inv (n2_neg, n2);
  not n30_inv (n30_neg, n30);
  not n31_inv (n31_neg, n31);
  not n32_inv (n32_neg, n32);
  not n33_inv (n33_neg, n33);
  not n34_inv (n34_neg, n34);
  not n35_inv (n35_neg, n35);
  not n36_inv (n36_neg, n36);
  not n37_inv (n37_neg, n37);
  not n38_inv (n38_neg, n38);
  not n39_inv (n39_neg, n39);
  not n3_inv (n3_neg, n3);
  not n40_inv (n40_neg, n40);
  not n41_inv (n41_neg, n41);
  not n42_inv (n42_neg, n42);
  not n43_inv (n43_neg, n43);
  not n44_inv (n44_neg, n44);
  not n45_inv (n45_neg, n45);
  not n46_inv (n46_neg, n46);
  not n47_inv (n47_neg, n47);
  not n48_inv (n48_neg, n48);
  not n49_inv (n49_neg, n49);
  not n4_inv (n4_neg, n4);
  not n50_inv (n50_neg, n50);
  not n51_inv (n51_neg, n51);
  not n52_inv (n52_neg, n52);
  not n53_inv (n53_neg, n53);
  not n54_inv (n54_neg, n54);
  not n55_inv (n55_neg, n55);
  not n56_inv (n56_neg, n56);
  not n57_inv (n57_neg, n57);
  not n58_inv (n58_neg, n58);
  not n59_inv (n59_neg, n59);
  not n5_inv (n5_neg, n5);
  not n60_inv (n60_neg, n60);
  not n61_inv (n61_neg, n61);
  not n62_inv (n62_neg, n62);
  not n63_inv (n63_neg, n63);
  not n64_inv (n64_neg, n64);
  not n65_inv (n65_neg, n65);
  not n66_inv (n66_neg, n66);
  not n67_inv (n67_neg, n67);
  not n68_inv (n68_neg, n68);
  not n69_inv (n69_neg, n69);
  not n6_inv (n6_neg, n6);
  not n70_inv (n70_neg, n70);
  not n71_inv (n71_neg, n71);
  not n72_inv (n72_neg, n72);
  not n73_inv (n73_neg, n73);
  not n74_inv (n74_neg, n74);
  not n75_inv (n75_neg, n75);
  not n76_inv (n76_neg, n76);
  not n77_inv (n77_neg, n77);
  not n78_inv (n78_neg, n78);
  not n79_inv (n79_neg, n79);
  not n7_inv (n7_neg, n7);
  not n80_inv (n80_neg, n80);
  not n81_inv (n81_neg, n81);
  not n82_inv (n82_neg, n82);
  not n83_inv (n83_neg, n83);
  not n84_inv (n84_neg, n84);
  not n85_inv (n85_neg, n85);
  not n86_inv (n86_neg, n86);
  not n87_inv (n87_neg, n87);
  not n88_inv (n88_neg, n88);
  not n89_inv (n89_neg, n89);
  not n8_inv (n8_neg, n8);
  not n90_inv (n90_neg, n90);
  not n91_inv (n91_neg, n91);
  not n92_inv (n92_neg, n92);
  not n93_inv (n93_neg, n93);
  not n94_inv (n94_neg, n94);
  not n95_inv (n95_neg, n95);
  not n96_inv (n96_neg, n96);
  not n97_inv (n97_neg, n97);
  not n98_inv (n98_neg, n98);
  not n99_inv (n99_neg, n99);
  not n9_inv (n9_neg, n9);
  reg_ar_as_w1 ready_reg (
    .clk(clk),
    .d(n382),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(ready));  // sources/rtl/camera_init.v(265)
  reg_ar_as_w1 reg0_b0 (
    .clk(divider2[8]),
    .d(sel1_b0_sel_o),
    .en(1'b1),
    .reset(~reset_n),
    .set(1'b0),
    .q(reg_address[0]));  // sources/rtl/camera_init.v(389)
  reg_ar_as_w1 reg0_b1 (
    .clk(divider2[8]),
    .d(sel1_b1_sel_o),
    .en(1'b1),
    .reset(~reset_n),
    .set(1'b0),
    .q(reg_address[1]));  // sources/rtl/camera_init.v(389)
  reg_ar_as_w1 reg1_b0 (
    .clk(divider2[8]),
    .d(\sel2_b0/or_or_B4_B5_o_or_B6__o ),
    .en(1'b1),
    .reset(~reset_n),
    .set(1'b0),
    .q(data_in_bus[0]));  // sources/rtl/camera_init.v(389)
  reg_ar_as_w1 reg1_b1 (
    .clk(divider2[8]),
    .d(\sel2_b1/or_B6_or_B7_B8_o_o ),
    .en(1'b1),
    .reset(~reset_n),
    .set(1'b0),
    .q(data_in_bus[1]));  // sources/rtl/camera_init.v(389)
  reg_ar_as_w1 reg1_b2 (
    .clk(divider2[8]),
    .d(\sel2_b2/or_B6_or_B7_B8_o_o ),
    .en(1'b1),
    .reset(~reset_n),
    .set(1'b0),
    .q(data_in_bus[2]));  // sources/rtl/camera_init.v(389)
  reg_ar_as_w1 reg1_b3 (
    .clk(divider2[8]),
    .d(\sel2_b3/or_B6_or_B7_B8_o_o ),
    .en(1'b1),
    .reset(~reset_n),
    .set(1'b0),
    .q(data_in_bus[3]));  // sources/rtl/camera_init.v(389)
  reg_ar_as_w1 reg1_b4 (
    .clk(divider2[8]),
    .d(\sel2_b4/or_B6_or_B7_B8_o_o ),
    .en(1'b1),
    .reset(~reset_n),
    .set(1'b0),
    .q(data_in_bus[4]));  // sources/rtl/camera_init.v(389)
  reg_ar_as_w1 reg1_b5 (
    .clk(divider2[8]),
    .d(\sel2_b5/or_B6_or_B7_B8_o_o ),
    .en(1'b1),
    .reset(~reset_n),
    .set(1'b0),
    .q(data_in_bus[5]));  // sources/rtl/camera_init.v(389)
  reg_ar_as_w1 reg1_b6 (
    .clk(divider2[8]),
    .d(\sel2_b6/or_B6_or_B7_B8_o_o ),
    .en(1'b1),
    .reset(~reset_n),
    .set(1'b0),
    .q(data_in_bus[6]));  // sources/rtl/camera_init.v(389)
  reg_ar_as_w1 reg1_b7 (
    .clk(divider2[8]),
    .d(\sel2_b7/or_B6_or_B7_B8_o_o ),
    .en(1'b1),
    .reset(~reset_n),
    .set(1'b0),
    .q(data_in_bus[7]));  // sources/rtl/camera_init.v(389)
  reg_ar_as_w1 reg2_b0 (
    .clk(divider2[8]),
    .d(n374[0]),
    .en(n380),
    .reset(~reset_n),
    .set(1'b0),
    .q(counter[0]));  // sources/rtl/camera_init.v(389)
  reg_ar_as_w1 reg2_b1 (
    .clk(divider2[8]),
    .d(n374[1]),
    .en(n380),
    .reset(~reset_n),
    .set(1'b0),
    .q(counter[1]));  // sources/rtl/camera_init.v(389)
  reg_ar_as_w1 reg2_b2 (
    .clk(divider2[8]),
    .d(n374[2]),
    .en(n380),
    .reset(~reset_n),
    .set(1'b0),
    .q(counter[2]));  // sources/rtl/camera_init.v(389)
  reg_ar_as_w1 reg2_b3 (
    .clk(divider2[8]),
    .d(n374[3]),
    .en(n380),
    .reset(~reset_n),
    .set(1'b0),
    .q(counter[3]));  // sources/rtl/camera_init.v(389)
  reg_ar_as_w1 reg2_b4 (
    .clk(divider2[8]),
    .d(n374[4]),
    .en(n380),
    .reset(~reset_n),
    .set(1'b0),
    .q(counter[4]));  // sources/rtl/camera_init.v(389)
  reg_ar_as_w1 reg2_b5 (
    .clk(divider2[8]),
    .d(n374[5]),
    .en(n380),
    .reset(~reset_n),
    .set(1'b0),
    .q(counter[5]));  // sources/rtl/camera_init.v(389)
  reg_ar_as_w1 reg2_b6 (
    .clk(divider2[8]),
    .d(n374[6]),
    .en(n380),
    .reset(~reset_n),
    .set(1'b0),
    .q(counter[6]));  // sources/rtl/camera_init.v(389)
  reg_ar_as_w1 reg2_b7 (
    .clk(divider2[8]),
    .d(n374[7]),
    .en(n380),
    .reset(~reset_n),
    .set(1'b0),
    .q(counter[7]));  // sources/rtl/camera_init.v(389)
  reg_ar_as_w1 reg3_b0 (
    .clk(divider2[8]),
    .d(n371[0]),
    .en(mux181_b0_sel_is_2_o),
    .reset(1'b0),
    .set(1'b0),
    .q(cnt[0]));  // sources/rtl/camera_init.v(389)
  reg_ar_as_w1 reg3_b1 (
    .clk(divider2[8]),
    .d(n371[1]),
    .en(mux181_b0_sel_is_2_o),
    .reset(1'b0),
    .set(1'b0),
    .q(cnt[1]));  // sources/rtl/camera_init.v(389)
  reg_ar_as_w1 reg3_b2 (
    .clk(divider2[8]),
    .d(n371[2]),
    .en(mux181_b0_sel_is_2_o),
    .reset(1'b0),
    .set(1'b0),
    .q(cnt[2]));  // sources/rtl/camera_init.v(389)
  reg_ar_as_w1 reg3_b3 (
    .clk(divider2[8]),
    .d(n371[3]),
    .en(mux181_b0_sel_is_2_o),
    .reset(1'b0),
    .set(1'b0),
    .q(cnt[3]));  // sources/rtl/camera_init.v(389)
  reg_ar_as_w1 reg3_b4 (
    .clk(divider2[8]),
    .d(n371[4]),
    .en(mux181_b0_sel_is_2_o),
    .reset(1'b0),
    .set(1'b0),
    .q(cnt[4]));  // sources/rtl/camera_init.v(389)
  reg_ar_as_w1 reg3_b5 (
    .clk(divider2[8]),
    .d(n371[5]),
    .en(mux181_b0_sel_is_2_o),
    .reset(1'b0),
    .set(1'b0),
    .q(cnt[5]));  // sources/rtl/camera_init.v(389)
  reg_ar_as_w1 reg3_b6 (
    .clk(divider2[8]),
    .d(n371[6]),
    .en(mux181_b0_sel_is_2_o),
    .reset(1'b0),
    .set(1'b0),
    .q(cnt[6]));  // sources/rtl/camera_init.v(389)
  reg_ar_as_w1 reg3_b7 (
    .clk(divider2[8]),
    .d(n371[7]),
    .en(mux181_b0_sel_is_2_o),
    .reset(1'b0),
    .set(1'b0),
    .q(cnt[7]));  // sources/rtl/camera_init.v(389)
  reg_ar_as_w1 reg4_b0 (
    .clk(clk),
    .d(n0[0]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(divider2[0]));  // sources/rtl/camera_init.v(72)
  reg_ar_as_w1 reg4_b1 (
    .clk(clk),
    .d(n0[1]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(divider2[1]));  // sources/rtl/camera_init.v(72)
  reg_ar_as_w1 reg4_b2 (
    .clk(clk),
    .d(n0[2]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(divider2[2]));  // sources/rtl/camera_init.v(72)
  reg_ar_as_w1 reg4_b3 (
    .clk(clk),
    .d(n0[3]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(divider2[3]));  // sources/rtl/camera_init.v(72)
  reg_ar_as_w1 reg4_b4 (
    .clk(clk),
    .d(n0[4]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(divider2[4]));  // sources/rtl/camera_init.v(72)
  reg_ar_as_w1 reg4_b5 (
    .clk(clk),
    .d(n0[5]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(divider2[5]));  // sources/rtl/camera_init.v(72)
  reg_ar_as_w1 reg4_b6 (
    .clk(clk),
    .d(n0[6]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(divider2[6]));  // sources/rtl/camera_init.v(72)
  reg_ar_as_w1 reg4_b7 (
    .clk(clk),
    .d(n0[7]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(divider2[7]));  // sources/rtl/camera_init.v(72)
  reg_ar_as_w1 reg4_b8 (
    .clk(clk),
    .d(n0[8]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(divider2[8]));  // sources/rtl/camera_init.v(72)
  reg_ar_as_w1 reg5_b0 (
    .clk(divider2[8]),
    .d(n369[0]),
    .en(1'b1),
    .reset(1'b0),
    .set(~reset_n),
    .q(state_next[0]));  // sources/rtl/camera_init.v(311)
  reg_ar_as_w1 reg5_b1 (
    .clk(divider2[8]),
    .d(n369[1]),
    .en(1'b1),
    .reset(1'b0),
    .set(~reset_n),
    .q(state_next[1]));  // sources/rtl/camera_init.v(311)
  reg_ar_as_w1 reg5_b2 (
    .clk(divider2[8]),
    .d(n369[2]),
    .en(1'b1),
    .reset(~reset_n),
    .set(1'b0),
    .q(state_next[2]));  // sources/rtl/camera_init.v(311)
  reg_ar_as_w1 reg5_b3 (
    .clk(divider2[8]),
    .d(n369[3]),
    .en(1'b1),
    .reset(1'b0),
    .set(~reset_n),
    .q(state_next[3]));  // sources/rtl/camera_init.v(311)
  reg_ar_as_w1 reg5_b4 (
    .clk(divider2[8]),
    .d(n369[4]),
    .en(1'b1),
    .reset(~reset_n),
    .set(1'b0),
    .q(state_next[4]));  // sources/rtl/camera_init.v(311)
  reg_ar_as_w1 reg5_b5 (
    .clk(divider2[8]),
    .d(n369[5]),
    .en(1'b1),
    .reset(~reset_n),
    .set(1'b0),
    .q(state_next[5]));  // sources/rtl/camera_init.v(311)
  reg_ar_as_w1 reg5_b6 (
    .clk(divider2[8]),
    .d(n369[6]),
    .en(1'b1),
    .reset(~reset_n),
    .set(1'b0),
    .q(state_next[6]));  // sources/rtl/camera_init.v(311)
  reg_ar_as_w1 reg5_b7 (
    .clk(divider2[8]),
    .d(n369[7]),
    .en(1'b1),
    .reset(~reset_n),
    .set(1'b0),
    .q(state_next[7]));  // sources/rtl/camera_init.v(311)
  and \sel0_b0/and_b0_0  (\sel0_b0/B0 , state_next[0], n383);
  and \sel0_b0/and_b0_3  (\sel0_b0/B3 , n363[0], n379);
  and \sel0_b0/and_b0_4  (\sel0_b0/B4 , n357[0], n381);
  or \sel0_b0/or_B4_B5  (\sel0_b0/or_B4_B5_o , \sel0_b0/B4 , n378);
  or \sel0_b0/or_or_B0_B1_o_or_B2_  (\sel0_b0/or_or_B0_B1_o_or_B2__o , \sel0_b0/B0 , \sel0_b0/B3 );
  or \sel0_b0/or_or_B4_B5_o_or_B6_  (\sel0_b0/or_or_B4_B5_o_or_B6__o , \sel0_b0/or_B4_B5_o , n376);
  or \sel0_b0/or_or_or_B0_B1_o_or_  (n369[0], \sel0_b0/or_or_B0_B1_o_or_B2__o , \sel0_b0/or_or_B4_B5_o_or_B6__o );
  and \sel0_b1/and_b0_0  (\sel0_b1/B0 , state_next[1], n383);
  and \sel0_b1/and_b0_3  (\sel0_b1/B3 , n363[1], n379);
  and \sel0_b1/and_b0_4  (\sel0_b1/B4 , n357[1], n381);
  or \sel0_b1/or_B0_B1  (\sel0_b1/or_B0_B1_o , \sel0_b1/B0 , n382);
  or \sel0_b1/or_or_B0_B1_o_or_B2_  (\sel0_b1/or_or_B0_B1_o_or_B2__o , \sel0_b1/or_B0_B1_o , \sel0_b1/B3 );
  or \sel0_b1/or_or_B4_B5_o_or_B6_  (\sel0_b1/or_or_B4_B5_o_or_B6__o , \sel0_b1/B4 , n377);
  or \sel0_b1/or_or_or_B0_B1_o_or_  (n369[1], \sel0_b1/or_or_B0_B1_o_or_B2__o , \sel0_b1/or_or_B4_B5_o_or_B6__o );
  and \sel0_b2/and_b0_0  (\sel0_b2/B0 , state_next[2], n383);
  and \sel0_b2/and_b0_3  (\sel0_b2/B3 , n363[2], n379);
  and \sel0_b2/and_b0_4  (\sel0_b2/B4 , n357[2], n381);
  or \sel0_b2/or_B2_B3  (\sel0_b2/or_B2_B3_o , n380, \sel0_b2/B3 );
  or \sel0_b2/or_B6_or_B7_B8_o  (\sel0_b2/or_B6_or_B7_B8_o_o , n377, \sel0_b2/or_B7_B8_o );
  or \sel0_b2/or_B7_B8  (\sel0_b2/or_B7_B8_o , n376, n375);
  or \sel0_b2/or_or_B0_B1_o_or_B2_  (\sel0_b2/or_or_B0_B1_o_or_B2__o , \sel0_b2/B0 , \sel0_b2/or_B2_B3_o );
  or \sel0_b2/or_or_B4_B5_o_or_B6_  (\sel0_b2/or_or_B4_B5_o_or_B6__o , \sel0_b2/B4 , \sel0_b2/or_B6_or_B7_B8_o_o );
  or \sel0_b2/or_or_or_B0_B1_o_or_  (n369[2], \sel0_b2/or_or_B0_B1_o_or_B2__o , \sel0_b2/or_or_B4_B5_o_or_B6__o );
  and \sel0_b3/and_b0_0  (\sel0_b3/B0 , state_next[3], n383);
  and \sel0_b3/and_b0_3  (\sel0_b3/B3 , n363[3], n379);
  and \sel0_b3/and_b0_4  (\sel0_b3/B4 , n357[3], n381);
  or \sel0_b3/or_B2_B3  (\sel0_b3/or_B2_B3_o , n380, \sel0_b3/B3 );
  or \sel0_b3/or_or_B0_B1_o_or_B2_  (\sel0_b3/or_or_B0_B1_o_or_B2__o , \sel0_b3/B0 , \sel0_b3/or_B2_B3_o );
  or \sel0_b3/or_or_B4_B5_o_or_B6_  (\sel0_b3/or_or_B4_B5_o_or_B6__o , \sel0_b3/B4 , \sel0_b2/or_B6_or_B7_B8_o_o );
  or \sel0_b3/or_or_or_B0_B1_o_or_  (n369[3], \sel0_b3/or_or_B0_B1_o_or_B2__o , \sel0_b3/or_or_B4_B5_o_or_B6__o );
  and \sel0_b4/and_b0_0  (\sel0_b4/B0 , state_next[4], n383);
  and \sel0_b4/and_b0_3  (\sel0_b4/B3 , n363[4], n379);
  and \sel0_b4/and_b0_4  (\sel0_b4/B4 , n357[4], n381);
  or \sel0_b4/or_B0_B1  (\sel0_b4/or_B0_B1_o , \sel0_b4/B0 , n382);
  or \sel0_b4/or_B4_B5  (\sel0_b4/or_B4_B5_o , \sel0_b4/B4 , n378);
  or \sel0_b4/or_or_B0_B1_o_or_B2_  (\sel0_b4/or_or_B0_B1_o_or_B2__o , \sel0_b4/or_B0_B1_o , \sel0_b4/B3 );
  or \sel0_b4/or_or_or_B0_B1_o_or_  (n369[4], \sel0_b4/or_or_B0_B1_o_or_B2__o , \sel0_b4/or_B4_B5_o );
  and \sel0_b5/and_b0_0  (\sel0_b5/B0 , state_next[5], n383);
  and \sel0_b5/and_b0_3  (\sel0_b5/B3 , n363[5], n379);
  and \sel0_b5/and_b0_4  (\sel0_b5/B4 , n357[5], n381);
  or \sel0_b5/or_or_B0_B1_o_or_B2_  (\sel0_b5/or_or_B0_B1_o_or_B2__o , \sel0_b5/B0 , \sel0_b5/B3 );
  or \sel0_b5/or_or_or_B0_B1_o_or_  (n369[5], \sel0_b5/or_or_B0_B1_o_or_B2__o , \sel0_b5/B4 );
  and \sel0_b6/and_b0_0  (\sel0_b6/B0 , state_next[6], n383);
  and \sel0_b6/and_b0_3  (\sel0_b6/B3 , n363[6], n379);
  and \sel0_b6/and_b0_4  (\sel0_b6/B4 , n357[6], n381);
  or \sel0_b6/or_or_B0_B1_o_or_B2_  (\sel0_b6/or_or_B0_B1_o_or_B2__o , \sel0_b6/B0 , \sel0_b6/B3 );
  or \sel0_b6/or_or_or_B0_B1_o_or_  (n369[6], \sel0_b6/or_or_B0_B1_o_or_B2__o , \sel0_b6/B4 );
  and \sel0_b7/and_b0_0  (\sel0_b7/B0 , state_next[7], n383);
  and \sel0_b7/and_b0_3  (\sel0_b7/B3 , n363[7], n379);
  and \sel0_b7/and_b0_4  (\sel0_b7/B4 , n357[7], n381);
  or \sel0_b7/or_or_B0_B1_o_or_B2_  (\sel0_b7/or_or_B0_B1_o_or_B2__o , \sel0_b7/B0 , \sel0_b7/B3 );
  or \sel0_b7/or_or_or_B0_B1_o_or_  (n369[7], \sel0_b7/or_or_B0_B1_o_or_B2__o , \sel0_b7/B4 );
  or sel1_b0_sel (sel1_b0_sel_o, n377, n375);  // sources/rtl/camera_init.v(388)
  or sel1_b1_sel (sel1_b1_sel_o, n377, n376);  // sources/rtl/camera_init.v(388)
  and \sel2_b0/and_b0_6  (\sel2_b0/B6 , regs_data[0], n377);
  and \sel2_b0/and_b0_7  (\sel2_b0/B7 , regs_data[8], n376);
  or \sel2_b0/or_B6_or_B7_B8_o  (\sel2_b0/or_B6_or_B7_B8_o_o , \sel2_b0/B6 , \sel2_b0/B7 );
  or \sel2_b0/or_or_B4_B5_o_or_B6_  (\sel2_b0/or_or_B4_B5_o_or_B6__o , n378, \sel2_b0/or_B6_or_B7_B8_o_o );
  and \sel2_b1/and_b0_6  (\sel2_b1/B6 , regs_data[1], n377);
  and \sel2_b1/and_b0_7  (\sel2_b1/B7 , regs_data[9], n376);
  or \sel2_b1/or_B6_or_B7_B8_o  (\sel2_b1/or_B6_or_B7_B8_o_o , \sel2_b1/B6 , \sel2_b1/B7 );
  and \sel2_b2/and_b0_6  (\sel2_b2/B6 , regs_data[2], n377);
  and \sel2_b2/and_b0_7  (\sel2_b2/B7 , regs_data[10], n376);
  or \sel2_b2/or_B6_or_B7_B8_o  (\sel2_b2/or_B6_or_B7_B8_o_o , \sel2_b2/B6 , \sel2_b2/B7 );
  and \sel2_b3/and_b0_6  (\sel2_b3/B6 , regs_data[3], n377);
  and \sel2_b3/and_b0_7  (\sel2_b3/B7 , regs_data[11], n376);
  or \sel2_b3/or_B6_or_B7_B8_o  (\sel2_b3/or_B6_or_B7_B8_o_o , \sel2_b3/B6 , \sel2_b3/B7 );
  and \sel2_b4/and_b0_6  (\sel2_b4/B6 , regs_data[4], n377);
  and \sel2_b4/and_b0_7  (\sel2_b4/B7 , regs_data[12], n376);
  or \sel2_b4/or_B6_or_B7_B8_o  (\sel2_b4/or_B6_or_B7_B8_o_o , \sel2_b4/B6 , \sel2_b4/B7 );
  and \sel2_b5/and_b0_6  (\sel2_b5/B6 , regs_data[5], n377);
  and \sel2_b5/and_b0_7  (\sel2_b5/B7 , regs_data[13], n376);
  or \sel2_b5/or_B6_or_B7_B8_o  (\sel2_b5/or_B6_or_B7_B8_o_o , \sel2_b5/B6 , \sel2_b5/or_B7_B8_o );
  or \sel2_b5/or_B7_B8  (\sel2_b5/or_B7_B8_o , \sel2_b5/B7 , n375);
  and \sel2_b6/and_b0_6  (\sel2_b6/B6 , regs_data[6], n377);
  and \sel2_b6/and_b0_7  (\sel2_b6/B7 , regs_data[14], n376);
  or \sel2_b6/or_B6_or_B7_B8_o  (\sel2_b6/or_B6_or_B7_B8_o_o , \sel2_b6/B6 , \sel2_b6/or_B7_B8_o );
  or \sel2_b6/or_B7_B8  (\sel2_b6/or_B7_B8_o , \sel2_b6/B7 , n375);
  and \sel2_b7/and_b0_6  (\sel2_b7/B6 , regs_data[7], n377);
  and \sel2_b7/and_b0_7  (\sel2_b7/B7 , regs_data[15], n376);
  or \sel2_b7/or_B6_or_B7_B8_o  (\sel2_b7/or_B6_or_B7_B8_o_o , \sel2_b7/B6 , \sel2_b7/B7 );
  and sel3_b0_sel_is_3 (sel3_b0_sel_is_3_o, n380, n177);
  or u10 (n366, n365, \sel0_b2/or_B7_B8_o );  // sources/rtl/camera_init.v(388)
  or u12 (n365, n378, n377);  // sources/rtl/camera_init.v(388)
  or u13 (n180, n382, n381);  // sources/rtl/camera_init.v(388)
  or u14 (n356, n180, n179);  // sources/rtl/camera_init.v(388)
  or u15 (n179, n380, n379);  // sources/rtl/camera_init.v(388)
  not u2 (n178[2], n177);  // sources/rtl/camera_init.v(256)
  not u4 (n359[3], n358);  // sources/rtl/camera_init.v(299)
  not u8 (n383, n364);  // sources/rtl/camera_init.v(388)
  or u9 (n364, n356, n366);  // sources/rtl/camera_init.v(388)
  i2c_module u_i2c_write (
    .address({1'b0,reg_address[1:0]}),
    .clk(clk),
    .reset_n(reset_n),
    .sda_in(sda_in),
    .write(bus_write),
    .writedata(data_in_bus),
    .ready(ready_out),
    .scl_out(scl),
    .sda(sda),
    .sda_oe(sda_oe),
    .success_out(success_out));  // sources/rtl/camera_init.v(48)

endmodule 

module add_pu20_pu20_o20
  (
  i0,
  i1,
  o
  );

  input [19:0] i0;
  input [19:0] i1;
  output [19:0] o;

  wire net_a0;
  wire net_a1;
  wire net_a10;
  wire net_a11;
  wire net_a12;
  wire net_a13;
  wire net_a14;
  wire net_a15;
  wire net_a16;
  wire net_a17;
  wire net_a18;
  wire net_a19;
  wire net_a2;
  wire net_a3;
  wire net_a4;
  wire net_a5;
  wire net_a6;
  wire net_a7;
  wire net_a8;
  wire net_a9;
  wire net_b0;
  wire net_b1;
  wire net_b10;
  wire net_b11;
  wire net_b12;
  wire net_b13;
  wire net_b14;
  wire net_b15;
  wire net_b16;
  wire net_b17;
  wire net_b18;
  wire net_b19;
  wire net_b2;
  wire net_b3;
  wire net_b4;
  wire net_b5;
  wire net_b6;
  wire net_b7;
  wire net_b8;
  wire net_b9;
  wire net_cout0;
  wire net_cout1;
  wire net_cout10;
  wire net_cout11;
  wire net_cout12;
  wire net_cout13;
  wire net_cout14;
  wire net_cout15;
  wire net_cout16;
  wire net_cout17;
  wire net_cout18;
  wire net_cout19;
  wire net_cout2;
  wire net_cout3;
  wire net_cout4;
  wire net_cout5;
  wire net_cout6;
  wire net_cout7;
  wire net_cout8;
  wire net_cout9;
  wire net_sum0;
  wire net_sum1;
  wire net_sum10;
  wire net_sum11;
  wire net_sum12;
  wire net_sum13;
  wire net_sum14;
  wire net_sum15;
  wire net_sum16;
  wire net_sum17;
  wire net_sum18;
  wire net_sum19;
  wire net_sum2;
  wire net_sum3;
  wire net_sum4;
  wire net_sum5;
  wire net_sum6;
  wire net_sum7;
  wire net_sum8;
  wire net_sum9;

  assign net_a19 = i0[19];
  assign net_a18 = i0[18];
  assign net_a17 = i0[17];
  assign net_a16 = i0[16];
  assign net_a15 = i0[15];
  assign net_a14 = i0[14];
  assign net_a13 = i0[13];
  assign net_a12 = i0[12];
  assign net_a11 = i0[11];
  assign net_a10 = i0[10];
  assign net_a9 = i0[9];
  assign net_a8 = i0[8];
  assign net_a7 = i0[7];
  assign net_a6 = i0[6];
  assign net_a5 = i0[5];
  assign net_a4 = i0[4];
  assign net_a3 = i0[3];
  assign net_a2 = i0[2];
  assign net_a1 = i0[1];
  assign net_a0 = i0[0];
  assign net_b19 = i1[19];
  assign net_b18 = i1[18];
  assign net_b17 = i1[17];
  assign net_b16 = i1[16];
  assign net_b15 = i1[15];
  assign net_b14 = i1[14];
  assign net_b13 = i1[13];
  assign net_b12 = i1[12];
  assign net_b11 = i1[11];
  assign net_b10 = i1[10];
  assign net_b9 = i1[9];
  assign net_b8 = i1[8];
  assign net_b7 = i1[7];
  assign net_b6 = i1[6];
  assign net_b5 = i1[5];
  assign net_b4 = i1[4];
  assign net_b3 = i1[3];
  assign net_b2 = i1[2];
  assign net_b1 = i1[1];
  assign net_b0 = i1[0];
  assign o[19] = net_sum19;
  assign o[18] = net_sum18;
  assign o[17] = net_sum17;
  assign o[16] = net_sum16;
  assign o[15] = net_sum15;
  assign o[14] = net_sum14;
  assign o[13] = net_sum13;
  assign o[12] = net_sum12;
  assign o[11] = net_sum11;
  assign o[10] = net_sum10;
  assign o[9] = net_sum9;
  assign o[8] = net_sum8;
  assign o[7] = net_sum7;
  assign o[6] = net_sum6;
  assign o[5] = net_sum5;
  assign o[4] = net_sum4;
  assign o[3] = net_sum3;
  assign o[2] = net_sum2;
  assign o[1] = net_sum1;
  assign o[0] = net_sum0;
  AL_FADD comp_0 (
    .a(net_a0),
    .b(net_b0),
    .c(1'b0),
    .cout(net_cout0),
    .sum(net_sum0));
  AL_FADD comp_1 (
    .a(net_a1),
    .b(net_b1),
    .c(net_cout0),
    .cout(net_cout1),
    .sum(net_sum1));
  AL_FADD comp_10 (
    .a(net_a10),
    .b(net_b10),
    .c(net_cout9),
    .cout(net_cout10),
    .sum(net_sum10));
  AL_FADD comp_11 (
    .a(net_a11),
    .b(net_b11),
    .c(net_cout10),
    .cout(net_cout11),
    .sum(net_sum11));
  AL_FADD comp_12 (
    .a(net_a12),
    .b(net_b12),
    .c(net_cout11),
    .cout(net_cout12),
    .sum(net_sum12));
  AL_FADD comp_13 (
    .a(net_a13),
    .b(net_b13),
    .c(net_cout12),
    .cout(net_cout13),
    .sum(net_sum13));
  AL_FADD comp_14 (
    .a(net_a14),
    .b(net_b14),
    .c(net_cout13),
    .cout(net_cout14),
    .sum(net_sum14));
  AL_FADD comp_15 (
    .a(net_a15),
    .b(net_b15),
    .c(net_cout14),
    .cout(net_cout15),
    .sum(net_sum15));
  AL_FADD comp_16 (
    .a(net_a16),
    .b(net_b16),
    .c(net_cout15),
    .cout(net_cout16),
    .sum(net_sum16));
  AL_FADD comp_17 (
    .a(net_a17),
    .b(net_b17),
    .c(net_cout16),
    .cout(net_cout17),
    .sum(net_sum17));
  AL_FADD comp_18 (
    .a(net_a18),
    .b(net_b18),
    .c(net_cout17),
    .cout(net_cout18),
    .sum(net_sum18));
  AL_FADD comp_19 (
    .a(net_a19),
    .b(net_b19),
    .c(net_cout18),
    .cout(net_cout19),
    .sum(net_sum19));
  AL_FADD comp_2 (
    .a(net_a2),
    .b(net_b2),
    .c(net_cout1),
    .cout(net_cout2),
    .sum(net_sum2));
  AL_FADD comp_3 (
    .a(net_a3),
    .b(net_b3),
    .c(net_cout2),
    .cout(net_cout3),
    .sum(net_sum3));
  AL_FADD comp_4 (
    .a(net_a4),
    .b(net_b4),
    .c(net_cout3),
    .cout(net_cout4),
    .sum(net_sum4));
  AL_FADD comp_5 (
    .a(net_a5),
    .b(net_b5),
    .c(net_cout4),
    .cout(net_cout5),
    .sum(net_sum5));
  AL_FADD comp_6 (
    .a(net_a6),
    .b(net_b6),
    .c(net_cout5),
    .cout(net_cout6),
    .sum(net_sum6));
  AL_FADD comp_7 (
    .a(net_a7),
    .b(net_b7),
    .c(net_cout6),
    .cout(net_cout7),
    .sum(net_sum7));
  AL_FADD comp_8 (
    .a(net_a8),
    .b(net_b8),
    .c(net_cout7),
    .cout(net_cout8),
    .sum(net_sum8));
  AL_FADD comp_9 (
    .a(net_a9),
    .b(net_b9),
    .c(net_cout8),
    .cout(net_cout9),
    .sum(net_sum9));

endmodule 

module add_pu16_pu16_o16
  (
  i0,
  i1,
  o
  );

  input [15:0] i0;
  input [15:0] i1;
  output [15:0] o;

  wire net_a0;
  wire net_a1;
  wire net_a10;
  wire net_a11;
  wire net_a12;
  wire net_a13;
  wire net_a14;
  wire net_a15;
  wire net_a2;
  wire net_a3;
  wire net_a4;
  wire net_a5;
  wire net_a6;
  wire net_a7;
  wire net_a8;
  wire net_a9;
  wire net_b0;
  wire net_b1;
  wire net_b10;
  wire net_b11;
  wire net_b12;
  wire net_b13;
  wire net_b14;
  wire net_b15;
  wire net_b2;
  wire net_b3;
  wire net_b4;
  wire net_b5;
  wire net_b6;
  wire net_b7;
  wire net_b8;
  wire net_b9;
  wire net_cout0;
  wire net_cout1;
  wire net_cout10;
  wire net_cout11;
  wire net_cout12;
  wire net_cout13;
  wire net_cout14;
  wire net_cout15;
  wire net_cout2;
  wire net_cout3;
  wire net_cout4;
  wire net_cout5;
  wire net_cout6;
  wire net_cout7;
  wire net_cout8;
  wire net_cout9;
  wire net_sum0;
  wire net_sum1;
  wire net_sum10;
  wire net_sum11;
  wire net_sum12;
  wire net_sum13;
  wire net_sum14;
  wire net_sum15;
  wire net_sum2;
  wire net_sum3;
  wire net_sum4;
  wire net_sum5;
  wire net_sum6;
  wire net_sum7;
  wire net_sum8;
  wire net_sum9;

  assign net_a15 = i0[15];
  assign net_a14 = i0[14];
  assign net_a13 = i0[13];
  assign net_a12 = i0[12];
  assign net_a11 = i0[11];
  assign net_a10 = i0[10];
  assign net_a9 = i0[9];
  assign net_a8 = i0[8];
  assign net_a7 = i0[7];
  assign net_a6 = i0[6];
  assign net_a5 = i0[5];
  assign net_a4 = i0[4];
  assign net_a3 = i0[3];
  assign net_a2 = i0[2];
  assign net_a1 = i0[1];
  assign net_a0 = i0[0];
  assign net_b15 = i1[15];
  assign net_b14 = i1[14];
  assign net_b13 = i1[13];
  assign net_b12 = i1[12];
  assign net_b11 = i1[11];
  assign net_b10 = i1[10];
  assign net_b9 = i1[9];
  assign net_b8 = i1[8];
  assign net_b7 = i1[7];
  assign net_b6 = i1[6];
  assign net_b5 = i1[5];
  assign net_b4 = i1[4];
  assign net_b3 = i1[3];
  assign net_b2 = i1[2];
  assign net_b1 = i1[1];
  assign net_b0 = i1[0];
  assign o[15] = net_sum15;
  assign o[14] = net_sum14;
  assign o[13] = net_sum13;
  assign o[12] = net_sum12;
  assign o[11] = net_sum11;
  assign o[10] = net_sum10;
  assign o[9] = net_sum9;
  assign o[8] = net_sum8;
  assign o[7] = net_sum7;
  assign o[6] = net_sum6;
  assign o[5] = net_sum5;
  assign o[4] = net_sum4;
  assign o[3] = net_sum3;
  assign o[2] = net_sum2;
  assign o[1] = net_sum1;
  assign o[0] = net_sum0;
  AL_FADD comp_0 (
    .a(net_a0),
    .b(net_b0),
    .c(1'b0),
    .cout(net_cout0),
    .sum(net_sum0));
  AL_FADD comp_1 (
    .a(net_a1),
    .b(net_b1),
    .c(net_cout0),
    .cout(net_cout1),
    .sum(net_sum1));
  AL_FADD comp_10 (
    .a(net_a10),
    .b(net_b10),
    .c(net_cout9),
    .cout(net_cout10),
    .sum(net_sum10));
  AL_FADD comp_11 (
    .a(net_a11),
    .b(net_b11),
    .c(net_cout10),
    .cout(net_cout11),
    .sum(net_sum11));
  AL_FADD comp_12 (
    .a(net_a12),
    .b(net_b12),
    .c(net_cout11),
    .cout(net_cout12),
    .sum(net_sum12));
  AL_FADD comp_13 (
    .a(net_a13),
    .b(net_b13),
    .c(net_cout12),
    .cout(net_cout13),
    .sum(net_sum13));
  AL_FADD comp_14 (
    .a(net_a14),
    .b(net_b14),
    .c(net_cout13),
    .cout(net_cout14),
    .sum(net_sum14));
  AL_FADD comp_15 (
    .a(net_a15),
    .b(net_b15),
    .c(net_cout14),
    .cout(net_cout15),
    .sum(net_sum15));
  AL_FADD comp_2 (
    .a(net_a2),
    .b(net_b2),
    .c(net_cout1),
    .cout(net_cout2),
    .sum(net_sum2));
  AL_FADD comp_3 (
    .a(net_a3),
    .b(net_b3),
    .c(net_cout2),
    .cout(net_cout3),
    .sum(net_sum3));
  AL_FADD comp_4 (
    .a(net_a4),
    .b(net_b4),
    .c(net_cout3),
    .cout(net_cout4),
    .sum(net_sum4));
  AL_FADD comp_5 (
    .a(net_a5),
    .b(net_b5),
    .c(net_cout4),
    .cout(net_cout5),
    .sum(net_sum5));
  AL_FADD comp_6 (
    .a(net_a6),
    .b(net_b6),
    .c(net_cout5),
    .cout(net_cout6),
    .sum(net_sum6));
  AL_FADD comp_7 (
    .a(net_a7),
    .b(net_b7),
    .c(net_cout6),
    .cout(net_cout7),
    .sum(net_sum7));
  AL_FADD comp_8 (
    .a(net_a8),
    .b(net_b8),
    .c(net_cout7),
    .cout(net_cout8),
    .sum(net_sum8));
  AL_FADD comp_9 (
    .a(net_a9),
    .b(net_b9),
    .c(net_cout8),
    .cout(net_cout9),
    .sum(net_sum9));

endmodule 

module eq_w1
  (
  i0,
  i1,
  o
  );

  input i0;
  input i1;
  output o;

  wire xor_i0_i1_o;

  not none_diff (o, xor_i0_i1_o);
  xor xor_i0_i1 (xor_i0_i1_o, i0, i1);

endmodule 

module lt_u20_u20
  (
  ci,
  i0,
  i1,
  o
  );

  input ci;
  input [19:0] i0;
  input [19:0] i1;
  output o;

  wire [19:0] diff;
  wire diff_12_18;
  wire diff_6_11;
  wire less_12_18;
  wire \less_12_18_inst/diff_0 ;
  wire \less_12_18_inst/diff_1 ;
  wire \less_12_18_inst/diff_2 ;
  wire \less_12_18_inst/diff_3 ;
  wire \less_12_18_inst/diff_4 ;
  wire \less_12_18_inst/diff_5 ;
  wire \less_12_18_inst/diff_6 ;
  wire \less_12_18_inst/o_0 ;
  wire \less_12_18_inst/o_1 ;
  wire \less_12_18_inst/o_2 ;
  wire \less_12_18_inst/o_3 ;
  wire \less_12_18_inst/o_4 ;
  wire \less_12_18_inst/o_5 ;
  wire less_6_11;
  wire \less_6_11_inst/diff_0 ;
  wire \less_6_11_inst/diff_1 ;
  wire \less_6_11_inst/diff_2 ;
  wire \less_6_11_inst/diff_3 ;
  wire \less_6_11_inst/diff_4 ;
  wire \less_6_11_inst/diff_5 ;
  wire \less_6_11_inst/o_0 ;
  wire \less_6_11_inst/o_1 ;
  wire \less_6_11_inst/o_2 ;
  wire \less_6_11_inst/o_3 ;
  wire \less_6_11_inst/o_4 ;
  wire o_0;
  wire o_1;
  wire o_2;
  wire o_3;
  wire o_4;
  wire o_5;
  wire o_6;
  wire o_7;

  or any_diff_12_18 (diff_12_18, diff[12], diff[13], diff[14], diff[15], diff[16], diff[17], diff[18]);
  or any_diff_6_11 (diff_6_11, diff[6], diff[7], diff[8], diff[9], diff[10], diff[11]);
  xor diff_0 (diff[0], i0[0], i1[0]);
  xor diff_1 (diff[1], i0[1], i1[1]);
  xor diff_10 (diff[10], i0[10], i1[10]);
  xor diff_11 (diff[11], i0[11], i1[11]);
  xor diff_12 (diff[12], i0[12], i1[12]);
  xor diff_13 (diff[13], i0[13], i1[13]);
  xor diff_14 (diff[14], i0[14], i1[14]);
  xor diff_15 (diff[15], i0[15], i1[15]);
  xor diff_16 (diff[16], i0[16], i1[16]);
  xor diff_17 (diff[17], i0[17], i1[17]);
  xor diff_18 (diff[18], i0[18], i1[18]);
  xor diff_19 (diff[19], i0[19], i1[19]);
  xor diff_2 (diff[2], i0[2], i1[2]);
  xor diff_3 (diff[3], i0[3], i1[3]);
  xor diff_4 (diff[4], i0[4], i1[4]);
  xor diff_5 (diff[5], i0[5], i1[5]);
  xor diff_6 (diff[6], i0[6], i1[6]);
  xor diff_7 (diff[7], i0[7], i1[7]);
  xor diff_8 (diff[8], i0[8], i1[8]);
  xor diff_9 (diff[9], i0[9], i1[9]);
  AL_MUX \less_12_18_inst/mux_0  (
    .i0(1'b0),
    .i1(i1[12]),
    .sel(\less_12_18_inst/diff_0 ),
    .o(\less_12_18_inst/o_0 ));
  AL_MUX \less_12_18_inst/mux_1  (
    .i0(\less_12_18_inst/o_0 ),
    .i1(i1[13]),
    .sel(\less_12_18_inst/diff_1 ),
    .o(\less_12_18_inst/o_1 ));
  AL_MUX \less_12_18_inst/mux_2  (
    .i0(\less_12_18_inst/o_1 ),
    .i1(i1[14]),
    .sel(\less_12_18_inst/diff_2 ),
    .o(\less_12_18_inst/o_2 ));
  AL_MUX \less_12_18_inst/mux_3  (
    .i0(\less_12_18_inst/o_2 ),
    .i1(i1[15]),
    .sel(\less_12_18_inst/diff_3 ),
    .o(\less_12_18_inst/o_3 ));
  AL_MUX \less_12_18_inst/mux_4  (
    .i0(\less_12_18_inst/o_3 ),
    .i1(i1[16]),
    .sel(\less_12_18_inst/diff_4 ),
    .o(\less_12_18_inst/o_4 ));
  AL_MUX \less_12_18_inst/mux_5  (
    .i0(\less_12_18_inst/o_4 ),
    .i1(i1[17]),
    .sel(\less_12_18_inst/diff_5 ),
    .o(\less_12_18_inst/o_5 ));
  AL_MUX \less_12_18_inst/mux_6  (
    .i0(\less_12_18_inst/o_5 ),
    .i1(i1[18]),
    .sel(\less_12_18_inst/diff_6 ),
    .o(less_12_18));
  xor \less_12_18_inst/xor_0  (\less_12_18_inst/diff_0 , i0[12], i1[12]);
  xor \less_12_18_inst/xor_1  (\less_12_18_inst/diff_1 , i0[13], i1[13]);
  xor \less_12_18_inst/xor_2  (\less_12_18_inst/diff_2 , i0[14], i1[14]);
  xor \less_12_18_inst/xor_3  (\less_12_18_inst/diff_3 , i0[15], i1[15]);
  xor \less_12_18_inst/xor_4  (\less_12_18_inst/diff_4 , i0[16], i1[16]);
  xor \less_12_18_inst/xor_5  (\less_12_18_inst/diff_5 , i0[17], i1[17]);
  xor \less_12_18_inst/xor_6  (\less_12_18_inst/diff_6 , i0[18], i1[18]);
  AL_MUX \less_6_11_inst/mux_0  (
    .i0(1'b0),
    .i1(i1[6]),
    .sel(\less_6_11_inst/diff_0 ),
    .o(\less_6_11_inst/o_0 ));
  AL_MUX \less_6_11_inst/mux_1  (
    .i0(\less_6_11_inst/o_0 ),
    .i1(i1[7]),
    .sel(\less_6_11_inst/diff_1 ),
    .o(\less_6_11_inst/o_1 ));
  AL_MUX \less_6_11_inst/mux_2  (
    .i0(\less_6_11_inst/o_1 ),
    .i1(i1[8]),
    .sel(\less_6_11_inst/diff_2 ),
    .o(\less_6_11_inst/o_2 ));
  AL_MUX \less_6_11_inst/mux_3  (
    .i0(\less_6_11_inst/o_2 ),
    .i1(i1[9]),
    .sel(\less_6_11_inst/diff_3 ),
    .o(\less_6_11_inst/o_3 ));
  AL_MUX \less_6_11_inst/mux_4  (
    .i0(\less_6_11_inst/o_3 ),
    .i1(i1[10]),
    .sel(\less_6_11_inst/diff_4 ),
    .o(\less_6_11_inst/o_4 ));
  AL_MUX \less_6_11_inst/mux_5  (
    .i0(\less_6_11_inst/o_4 ),
    .i1(i1[11]),
    .sel(\less_6_11_inst/diff_5 ),
    .o(less_6_11));
  xor \less_6_11_inst/xor_0  (\less_6_11_inst/diff_0 , i0[6], i1[6]);
  xor \less_6_11_inst/xor_1  (\less_6_11_inst/diff_1 , i0[7], i1[7]);
  xor \less_6_11_inst/xor_2  (\less_6_11_inst/diff_2 , i0[8], i1[8]);
  xor \less_6_11_inst/xor_3  (\less_6_11_inst/diff_3 , i0[9], i1[9]);
  xor \less_6_11_inst/xor_4  (\less_6_11_inst/diff_4 , i0[10], i1[10]);
  xor \less_6_11_inst/xor_5  (\less_6_11_inst/diff_5 , i0[11], i1[11]);
  AL_MUX mux_0 (
    .i0(ci),
    .i1(i1[0]),
    .sel(diff[0]),
    .o(o_0));
  AL_MUX mux_1 (
    .i0(o_0),
    .i1(i1[1]),
    .sel(diff[1]),
    .o(o_1));
  AL_MUX mux_2 (
    .i0(o_1),
    .i1(i1[2]),
    .sel(diff[2]),
    .o(o_2));
  AL_MUX mux_3 (
    .i0(o_2),
    .i1(i1[3]),
    .sel(diff[3]),
    .o(o_3));
  AL_MUX mux_4 (
    .i0(o_3),
    .i1(i1[4]),
    .sel(diff[4]),
    .o(o_4));
  AL_MUX mux_5 (
    .i0(o_4),
    .i1(i1[5]),
    .sel(diff[5]),
    .o(o_5));
  AL_MUX mux_6 (
    .i0(o_5),
    .i1(less_6_11),
    .sel(diff_6_11),
    .o(o_6));
  AL_MUX mux_7 (
    .i0(o_6),
    .i1(less_12_18),
    .sel(diff_12_18),
    .o(o_7));
  AL_MUX mux_8 (
    .i0(o_7),
    .i1(i1[19]),
    .sel(diff[19]),
    .o(o));

endmodule 

module reg_ar_as_w1
  (
  clk,
  d,
  en,
  reset,
  set,
  q
  );

  input clk;
  input d;
  input en;
  input reset;
  input set;
  output q;

  parameter REGSET = "RESET";
  wire enout;

  AL_MUX u_en0 (
    .i0(q),
    .i1(d),
    .sel(en),
    .o(enout));
  AL_DFF #(
    .INI((REGSET == "SET") ? 1'b1 : 1'b0))
    u_seq0 (
    .clk(clk),
    .d(enout),
    .reset(reset),
    .set(set),
    .q(q));

endmodule 

module reg_ar_ss_w1
  (
  clk,
  d,
  en,
  reset,
  set,
  q
  );

  input clk;
  input d;
  input en;
  input reset;
  input set;
  output q;

  parameter REGSET = "RESET";
  wire enout;
  wire setout;

  AL_MUX u_en0 (
    .i0(q),
    .i1(d),
    .sel(en),
    .o(enout));
  AL_DFF #(
    .INI((REGSET == "SET") ? 1'b1 : 1'b0))
    u_seq0 (
    .clk(clk),
    .d(setout),
    .reset(reset),
    .set(1'b0),
    .q(q));
  AL_MUX u_set0 (
    .i0(enout),
    .i1(1'b1),
    .sel(set),
    .o(setout));

endmodule 

module \lcd_sync(IMG_Y=1)   // sources/rtl/lcd_sync.v(14)
  (
  clk,
  rest_n,
  addr,
  hsync_cnt,
  img_ack,
  lcd_clk,
  lcd_de,
  lcd_hsync,
  lcd_pwm,
  lcd_vsync,
  vsync_cnt
  );

  input clk;  // sources/rtl/lcd_sync.v(23)
  input rest_n;  // sources/rtl/lcd_sync.v(24)
  output [15:0] addr;  // sources/rtl/lcd_sync.v(33)
  output [10:0] hsync_cnt;  // sources/rtl/lcd_sync.v(30)
  output img_ack;  // sources/rtl/lcd_sync.v(32)
  output lcd_clk;  // sources/rtl/lcd_sync.v(25)
  output lcd_de;  // sources/rtl/lcd_sync.v(29)
  output lcd_hsync;  // sources/rtl/lcd_sync.v(27)
  output lcd_pwm;  // sources/rtl/lcd_sync.v(26)
  output lcd_vsync;  // sources/rtl/lcd_sync.v(28)
  output [10:0] vsync_cnt;  // sources/rtl/lcd_sync.v(31)

  parameter IMG_H = 164;
  parameter IMG_W = 200;
  parameter IMG_X = 0;
  parameter IMG_Y = 1;
  // localparam TFT_H = 640;
  // localparam TFT_V = 480;
  // localparam TH = 800;
  // localparam THB = 160;
  // localparam TV = 525;
  // localparam TVB = 45;
  wire [10:0] n10;
  wire [10:0] n2;
  wire [11:0] n21;
  wire [11:0] n24;
  wire [11:0] n28;
  wire [31:0] n29;
  wire [10:0] n3;
  wire [11:0] n30;
  wire [31:0] n31;
  wire [39:0] n32;
  wire [31:0] n33;
  wire [15:0] n34;
  wire [10:0] n8;
  wire [10:0] n9;
  wire n1;
  wire n11;
  wire n12;
  wire n13;
  wire n14;
  wire n15;
  wire n16;
  wire n17;
  wire n18;
  wire n19;
  wire n20;
  wire n22;
  wire n23;
  wire n25;
  wire n26;
  wire n27;
  wire n4;
  wire n5;
  wire n6;
  wire n7;

  add_pu11_pu11_o11 add0 (
    .i0(hsync_cnt),
    .i1(11'b00000000001),
    .o(n2));  // sources/rtl/lcd_sync.v(61)
  add_pu11_pu11_o11 add1 (
    .i0(vsync_cnt),
    .i1(11'b00000000001),
    .o(n8));  // sources/rtl/lcd_sync.v(71)
  add_pu16_pu16_o16 add2 (
    .i0(n29[15:0]),
    .i1({n32[15:3],3'b000}),
    .o(n33[15:0]));  // sources/rtl/lcd_sync.v(93)
  eq_w11 eq0 (
    .i0(hsync_cnt),
    .i1(11'b01100100000),
    .o(n1));  // sources/rtl/lcd_sync.v(58)
  eq_w11 eq1 (
    .i0(vsync_cnt),
    .i1(11'b01000001101),
    .o(n4));  // sources/rtl/lcd_sync.v(68)
  eq_w1 eq2 (
    .i0(rest_n),
    .i1(1'b1),
    .o(lcd_pwm));  // sources/rtl/lcd_sync.v(74)
  lt_u11_u11 lt0 (
    .ci(1'b1),
    .i0(11'b00000010000),
    .i1(hsync_cnt),
    .o(n11));  // sources/rtl/lcd_sync.v(76)
  lt_u11_u11 lt1 (
    .ci(1'b0),
    .i0(hsync_cnt),
    .i1(11'b00001110000),
    .o(n12));  // sources/rtl/lcd_sync.v(76)
  lt_u12_u12 lt10_2 (
    .ci(1'b0),
    .i0(n24),
    .i1(12'b000010100101),
    .o(n26));  // sources/rtl/lcd_sync.v(84)
  lt_u11_u11 lt2 (
    .ci(1'b1),
    .i0(11'b00000001010),
    .i1(vsync_cnt),
    .o(n13));  // sources/rtl/lcd_sync.v(77)
  lt_u11_u11 lt3 (
    .ci(1'b0),
    .i0(vsync_cnt),
    .i1(11'b00000001100),
    .o(n14));  // sources/rtl/lcd_sync.v(77)
  lt_u11_u11 lt4 (
    .ci(1'b1),
    .i0(11'b00010100000),
    .i1(hsync_cnt),
    .o(n15));  // sources/rtl/lcd_sync.v(78)
  lt_u11_u11 lt5 (
    .ci(1'b1),
    .i0(hsync_cnt),
    .i1(11'b01100100000),
    .o(n16));  // sources/rtl/lcd_sync.v(78)
  lt_u11_u11 lt6 (
    .ci(1'b1),
    .i0(11'b00000101101),
    .i1(vsync_cnt),
    .o(n18));  // sources/rtl/lcd_sync.v(78)
  lt_u11_u11 lt7 (
    .ci(1'b0),
    .i0(vsync_cnt),
    .i1(11'b01000001101),
    .o(n20));  // sources/rtl/lcd_sync.v(78)
  lt_u12_u12 lt8_2 (
    .ci(1'b0),
    .i0(n21),
    .i1(12'b000011001000),
    .o(n22));  // sources/rtl/lcd_sync.v(83)
  lt_u12_u12 lt9_2 (
    .ci(1'b1),
    .i0(12'b000000000001),
    .i1(n24),
    .o(n25));  // sources/rtl/lcd_sync.v(84)
  mult_u13_u5_o13 mult0 (
    .i0(n31[12:0]),
    .i1(5'b11001),
    .o(n32[15:3]));  // sources/rtl/lcd_sync.v(93)
  binary_mux_s1_w1 mux0_b0 (
    .i0(n2[0]),
    .i1(1'b0),
    .sel(n1),
    .o(n3[0]));  // sources/rtl/lcd_sync.v(61)
  binary_mux_s1_w1 mux0_b1 (
    .i0(n2[1]),
    .i1(1'b0),
    .sel(n1),
    .o(n3[1]));  // sources/rtl/lcd_sync.v(61)
  binary_mux_s1_w1 mux0_b10 (
    .i0(n2[10]),
    .i1(1'b0),
    .sel(n1),
    .o(n3[10]));  // sources/rtl/lcd_sync.v(61)
  binary_mux_s1_w1 mux0_b2 (
    .i0(n2[2]),
    .i1(1'b0),
    .sel(n1),
    .o(n3[2]));  // sources/rtl/lcd_sync.v(61)
  binary_mux_s1_w1 mux0_b3 (
    .i0(n2[3]),
    .i1(1'b0),
    .sel(n1),
    .o(n3[3]));  // sources/rtl/lcd_sync.v(61)
  binary_mux_s1_w1 mux0_b4 (
    .i0(n2[4]),
    .i1(1'b0),
    .sel(n1),
    .o(n3[4]));  // sources/rtl/lcd_sync.v(61)
  binary_mux_s1_w1 mux0_b5 (
    .i0(n2[5]),
    .i1(1'b0),
    .sel(n1),
    .o(n3[5]));  // sources/rtl/lcd_sync.v(61)
  binary_mux_s1_w1 mux0_b6 (
    .i0(n2[6]),
    .i1(1'b0),
    .sel(n1),
    .o(n3[6]));  // sources/rtl/lcd_sync.v(61)
  binary_mux_s1_w1 mux0_b7 (
    .i0(n2[7]),
    .i1(1'b0),
    .sel(n1),
    .o(n3[7]));  // sources/rtl/lcd_sync.v(61)
  binary_mux_s1_w1 mux0_b8 (
    .i0(n2[8]),
    .i1(1'b0),
    .sel(n1),
    .o(n3[8]));  // sources/rtl/lcd_sync.v(61)
  binary_mux_s1_w1 mux0_b9 (
    .i0(n2[9]),
    .i1(1'b0),
    .sel(n1),
    .o(n3[9]));  // sources/rtl/lcd_sync.v(61)
  binary_mux_s1_w1 mux1_b0 (
    .i0(vsync_cnt[0]),
    .i1(n8[0]),
    .sel(n7),
    .o(n9[0]));  // sources/rtl/lcd_sync.v(71)
  binary_mux_s1_w1 mux1_b1 (
    .i0(vsync_cnt[1]),
    .i1(n8[1]),
    .sel(n7),
    .o(n9[1]));  // sources/rtl/lcd_sync.v(71)
  binary_mux_s1_w1 mux1_b10 (
    .i0(vsync_cnt[10]),
    .i1(n8[10]),
    .sel(n7),
    .o(n9[10]));  // sources/rtl/lcd_sync.v(71)
  binary_mux_s1_w1 mux1_b2 (
    .i0(vsync_cnt[2]),
    .i1(n8[2]),
    .sel(n7),
    .o(n9[2]));  // sources/rtl/lcd_sync.v(71)
  binary_mux_s1_w1 mux1_b3 (
    .i0(vsync_cnt[3]),
    .i1(n8[3]),
    .sel(n7),
    .o(n9[3]));  // sources/rtl/lcd_sync.v(71)
  binary_mux_s1_w1 mux1_b4 (
    .i0(vsync_cnt[4]),
    .i1(n8[4]),
    .sel(n7),
    .o(n9[4]));  // sources/rtl/lcd_sync.v(71)
  binary_mux_s1_w1 mux1_b5 (
    .i0(vsync_cnt[5]),
    .i1(n8[5]),
    .sel(n7),
    .o(n9[5]));  // sources/rtl/lcd_sync.v(71)
  binary_mux_s1_w1 mux1_b6 (
    .i0(vsync_cnt[6]),
    .i1(n8[6]),
    .sel(n7),
    .o(n9[6]));  // sources/rtl/lcd_sync.v(71)
  binary_mux_s1_w1 mux1_b7 (
    .i0(vsync_cnt[7]),
    .i1(n8[7]),
    .sel(n7),
    .o(n9[7]));  // sources/rtl/lcd_sync.v(71)
  binary_mux_s1_w1 mux1_b8 (
    .i0(vsync_cnt[8]),
    .i1(n8[8]),
    .sel(n7),
    .o(n9[8]));  // sources/rtl/lcd_sync.v(71)
  binary_mux_s1_w1 mux1_b9 (
    .i0(vsync_cnt[9]),
    .i1(n8[9]),
    .sel(n7),
    .o(n9[9]));  // sources/rtl/lcd_sync.v(71)
  binary_mux_s1_w1 mux2_b0 (
    .i0(n9[0]),
    .i1(1'b0),
    .sel(n5),
    .o(n10[0]));  // sources/rtl/lcd_sync.v(71)
  binary_mux_s1_w1 mux2_b1 (
    .i0(n9[1]),
    .i1(1'b0),
    .sel(n5),
    .o(n10[1]));  // sources/rtl/lcd_sync.v(71)
  binary_mux_s1_w1 mux2_b10 (
    .i0(n9[10]),
    .i1(1'b0),
    .sel(n5),
    .o(n10[10]));  // sources/rtl/lcd_sync.v(71)
  binary_mux_s1_w1 mux2_b2 (
    .i0(n9[2]),
    .i1(1'b0),
    .sel(n5),
    .o(n10[2]));  // sources/rtl/lcd_sync.v(71)
  binary_mux_s1_w1 mux2_b3 (
    .i0(n9[3]),
    .i1(1'b0),
    .sel(n5),
    .o(n10[3]));  // sources/rtl/lcd_sync.v(71)
  binary_mux_s1_w1 mux2_b4 (
    .i0(n9[4]),
    .i1(1'b0),
    .sel(n5),
    .o(n10[4]));  // sources/rtl/lcd_sync.v(71)
  binary_mux_s1_w1 mux2_b5 (
    .i0(n9[5]),
    .i1(1'b0),
    .sel(n5),
    .o(n10[5]));  // sources/rtl/lcd_sync.v(71)
  binary_mux_s1_w1 mux2_b6 (
    .i0(n9[6]),
    .i1(1'b0),
    .sel(n5),
    .o(n10[6]));  // sources/rtl/lcd_sync.v(71)
  binary_mux_s1_w1 mux2_b7 (
    .i0(n9[7]),
    .i1(1'b0),
    .sel(n5),
    .o(n10[7]));  // sources/rtl/lcd_sync.v(71)
  binary_mux_s1_w1 mux2_b8 (
    .i0(n9[8]),
    .i1(1'b0),
    .sel(n5),
    .o(n10[8]));  // sources/rtl/lcd_sync.v(71)
  binary_mux_s1_w1 mux2_b9 (
    .i0(n9[9]),
    .i1(1'b0),
    .sel(n5),
    .o(n10[9]));  // sources/rtl/lcd_sync.v(71)
  binary_mux_s1_w1 mux3_b0 (
    .i0(1'b0),
    .i1(n33[0]),
    .sel(img_ack),
    .o(n34[0]));  // sources/rtl/lcd_sync.v(95)
  binary_mux_s1_w1 mux3_b1 (
    .i0(1'b0),
    .i1(n33[1]),
    .sel(img_ack),
    .o(n34[1]));  // sources/rtl/lcd_sync.v(95)
  binary_mux_s1_w1 mux3_b10 (
    .i0(1'b0),
    .i1(n33[10]),
    .sel(img_ack),
    .o(n34[10]));  // sources/rtl/lcd_sync.v(95)
  binary_mux_s1_w1 mux3_b11 (
    .i0(1'b0),
    .i1(n33[11]),
    .sel(img_ack),
    .o(n34[11]));  // sources/rtl/lcd_sync.v(95)
  binary_mux_s1_w1 mux3_b12 (
    .i0(1'b0),
    .i1(n33[12]),
    .sel(img_ack),
    .o(n34[12]));  // sources/rtl/lcd_sync.v(95)
  binary_mux_s1_w1 mux3_b13 (
    .i0(1'b0),
    .i1(n33[13]),
    .sel(img_ack),
    .o(n34[13]));  // sources/rtl/lcd_sync.v(95)
  binary_mux_s1_w1 mux3_b14 (
    .i0(1'b0),
    .i1(n33[14]),
    .sel(img_ack),
    .o(n34[14]));  // sources/rtl/lcd_sync.v(95)
  binary_mux_s1_w1 mux3_b15 (
    .i0(1'b0),
    .i1(n33[15]),
    .sel(img_ack),
    .o(n34[15]));  // sources/rtl/lcd_sync.v(95)
  binary_mux_s1_w1 mux3_b2 (
    .i0(1'b0),
    .i1(n33[2]),
    .sel(img_ack),
    .o(n34[2]));  // sources/rtl/lcd_sync.v(95)
  binary_mux_s1_w1 mux3_b3 (
    .i0(1'b0),
    .i1(n33[3]),
    .sel(img_ack),
    .o(n34[3]));  // sources/rtl/lcd_sync.v(95)
  binary_mux_s1_w1 mux3_b4 (
    .i0(1'b0),
    .i1(n33[4]),
    .sel(img_ack),
    .o(n34[4]));  // sources/rtl/lcd_sync.v(95)
  binary_mux_s1_w1 mux3_b5 (
    .i0(1'b0),
    .i1(n33[5]),
    .sel(img_ack),
    .o(n34[5]));  // sources/rtl/lcd_sync.v(95)
  binary_mux_s1_w1 mux3_b6 (
    .i0(1'b0),
    .i1(n33[6]),
    .sel(img_ack),
    .o(n34[6]));  // sources/rtl/lcd_sync.v(95)
  binary_mux_s1_w1 mux3_b7 (
    .i0(1'b0),
    .i1(n33[7]),
    .sel(img_ack),
    .o(n34[7]));  // sources/rtl/lcd_sync.v(95)
  binary_mux_s1_w1 mux3_b8 (
    .i0(1'b0),
    .i1(n33[8]),
    .sel(img_ack),
    .o(n34[8]));  // sources/rtl/lcd_sync.v(95)
  binary_mux_s1_w1 mux3_b9 (
    .i0(1'b0),
    .i1(n33[9]),
    .sel(img_ack),
    .o(n34[9]));  // sources/rtl/lcd_sync.v(95)
  ne_w11 neq0 (
    .i0(vsync_cnt),
    .i1(11'b01000001101),
    .o(n6));  // sources/rtl/lcd_sync.v(70)
  reg_ar_as_w1 reg0_b0 (
    .clk(clk),
    .d(n10[0]),
    .en(1'b1),
    .reset(~rest_n),
    .set(1'b0),
    .q(vsync_cnt[0]));  // sources/rtl/lcd_sync.v(71)
  reg_ar_as_w1 reg0_b1 (
    .clk(clk),
    .d(n10[1]),
    .en(1'b1),
    .reset(~rest_n),
    .set(1'b0),
    .q(vsync_cnt[1]));  // sources/rtl/lcd_sync.v(71)
  reg_ar_as_w1 reg0_b10 (
    .clk(clk),
    .d(n10[10]),
    .en(1'b1),
    .reset(~rest_n),
    .set(1'b0),
    .q(vsync_cnt[10]));  // sources/rtl/lcd_sync.v(71)
  reg_ar_as_w1 reg0_b2 (
    .clk(clk),
    .d(n10[2]),
    .en(1'b1),
    .reset(~rest_n),
    .set(1'b0),
    .q(vsync_cnt[2]));  // sources/rtl/lcd_sync.v(71)
  reg_ar_as_w1 reg0_b3 (
    .clk(clk),
    .d(n10[3]),
    .en(1'b1),
    .reset(~rest_n),
    .set(1'b0),
    .q(vsync_cnt[3]));  // sources/rtl/lcd_sync.v(71)
  reg_ar_as_w1 reg0_b4 (
    .clk(clk),
    .d(n10[4]),
    .en(1'b1),
    .reset(~rest_n),
    .set(1'b0),
    .q(vsync_cnt[4]));  // sources/rtl/lcd_sync.v(71)
  reg_ar_as_w1 reg0_b5 (
    .clk(clk),
    .d(n10[5]),
    .en(1'b1),
    .reset(~rest_n),
    .set(1'b0),
    .q(vsync_cnt[5]));  // sources/rtl/lcd_sync.v(71)
  reg_ar_as_w1 reg0_b6 (
    .clk(clk),
    .d(n10[6]),
    .en(1'b1),
    .reset(~rest_n),
    .set(1'b0),
    .q(vsync_cnt[6]));  // sources/rtl/lcd_sync.v(71)
  reg_ar_as_w1 reg0_b7 (
    .clk(clk),
    .d(n10[7]),
    .en(1'b1),
    .reset(~rest_n),
    .set(1'b0),
    .q(vsync_cnt[7]));  // sources/rtl/lcd_sync.v(71)
  reg_ar_as_w1 reg0_b8 (
    .clk(clk),
    .d(n10[8]),
    .en(1'b1),
    .reset(~rest_n),
    .set(1'b0),
    .q(vsync_cnt[8]));  // sources/rtl/lcd_sync.v(71)
  reg_ar_as_w1 reg0_b9 (
    .clk(clk),
    .d(n10[9]),
    .en(1'b1),
    .reset(~rest_n),
    .set(1'b0),
    .q(vsync_cnt[9]));  // sources/rtl/lcd_sync.v(71)
  reg_ar_as_w1 reg1_b0 (
    .clk(clk),
    .d(n34[0]),
    .en(1'b1),
    .reset(~rest_n),
    .set(1'b0),
    .q(addr[0]));  // sources/rtl/lcd_sync.v(95)
  reg_ar_as_w1 reg1_b1 (
    .clk(clk),
    .d(n34[1]),
    .en(1'b1),
    .reset(~rest_n),
    .set(1'b0),
    .q(addr[1]));  // sources/rtl/lcd_sync.v(95)
  reg_ar_as_w1 reg1_b10 (
    .clk(clk),
    .d(n34[10]),
    .en(1'b1),
    .reset(~rest_n),
    .set(1'b0),
    .q(addr[10]));  // sources/rtl/lcd_sync.v(95)
  reg_ar_as_w1 reg1_b11 (
    .clk(clk),
    .d(n34[11]),
    .en(1'b1),
    .reset(~rest_n),
    .set(1'b0),
    .q(addr[11]));  // sources/rtl/lcd_sync.v(95)
  reg_ar_as_w1 reg1_b12 (
    .clk(clk),
    .d(n34[12]),
    .en(1'b1),
    .reset(~rest_n),
    .set(1'b0),
    .q(addr[12]));  // sources/rtl/lcd_sync.v(95)
  reg_ar_as_w1 reg1_b13 (
    .clk(clk),
    .d(n34[13]),
    .en(1'b1),
    .reset(~rest_n),
    .set(1'b0),
    .q(addr[13]));  // sources/rtl/lcd_sync.v(95)
  reg_ar_as_w1 reg1_b14 (
    .clk(clk),
    .d(n34[14]),
    .en(1'b1),
    .reset(~rest_n),
    .set(1'b0),
    .q(addr[14]));  // sources/rtl/lcd_sync.v(95)
  reg_ar_as_w1 reg1_b15 (
    .clk(clk),
    .d(n34[15]),
    .en(1'b1),
    .reset(~rest_n),
    .set(1'b0),
    .q(addr[15]));  // sources/rtl/lcd_sync.v(95)
  reg_ar_as_w1 reg1_b2 (
    .clk(clk),
    .d(n34[2]),
    .en(1'b1),
    .reset(~rest_n),
    .set(1'b0),
    .q(addr[2]));  // sources/rtl/lcd_sync.v(95)
  reg_ar_as_w1 reg1_b3 (
    .clk(clk),
    .d(n34[3]),
    .en(1'b1),
    .reset(~rest_n),
    .set(1'b0),
    .q(addr[3]));  // sources/rtl/lcd_sync.v(95)
  reg_ar_as_w1 reg1_b4 (
    .clk(clk),
    .d(n34[4]),
    .en(1'b1),
    .reset(~rest_n),
    .set(1'b0),
    .q(addr[4]));  // sources/rtl/lcd_sync.v(95)
  reg_ar_as_w1 reg1_b5 (
    .clk(clk),
    .d(n34[5]),
    .en(1'b1),
    .reset(~rest_n),
    .set(1'b0),
    .q(addr[5]));  // sources/rtl/lcd_sync.v(95)
  reg_ar_as_w1 reg1_b6 (
    .clk(clk),
    .d(n34[6]),
    .en(1'b1),
    .reset(~rest_n),
    .set(1'b0),
    .q(addr[6]));  // sources/rtl/lcd_sync.v(95)
  reg_ar_as_w1 reg1_b7 (
    .clk(clk),
    .d(n34[7]),
    .en(1'b1),
    .reset(~rest_n),
    .set(1'b0),
    .q(addr[7]));  // sources/rtl/lcd_sync.v(95)
  reg_ar_as_w1 reg1_b8 (
    .clk(clk),
    .d(n34[8]),
    .en(1'b1),
    .reset(~rest_n),
    .set(1'b0),
    .q(addr[8]));  // sources/rtl/lcd_sync.v(95)
  reg_ar_as_w1 reg1_b9 (
    .clk(clk),
    .d(n34[9]),
    .en(1'b1),
    .reset(~rest_n),
    .set(1'b0),
    .q(addr[9]));  // sources/rtl/lcd_sync.v(95)
  reg_ar_as_w1 reg2_b0 (
    .clk(clk),
    .d(n3[0]),
    .en(1'b1),
    .reset(~rest_n),
    .set(1'b0),
    .q(hsync_cnt[0]));  // sources/rtl/lcd_sync.v(61)
  reg_ar_as_w1 reg2_b1 (
    .clk(clk),
    .d(n3[1]),
    .en(1'b1),
    .reset(~rest_n),
    .set(1'b0),
    .q(hsync_cnt[1]));  // sources/rtl/lcd_sync.v(61)
  reg_ar_as_w1 reg2_b10 (
    .clk(clk),
    .d(n3[10]),
    .en(1'b1),
    .reset(~rest_n),
    .set(1'b0),
    .q(hsync_cnt[10]));  // sources/rtl/lcd_sync.v(61)
  reg_ar_as_w1 reg2_b2 (
    .clk(clk),
    .d(n3[2]),
    .en(1'b1),
    .reset(~rest_n),
    .set(1'b0),
    .q(hsync_cnt[2]));  // sources/rtl/lcd_sync.v(61)
  reg_ar_as_w1 reg2_b3 (
    .clk(clk),
    .d(n3[3]),
    .en(1'b1),
    .reset(~rest_n),
    .set(1'b0),
    .q(hsync_cnt[3]));  // sources/rtl/lcd_sync.v(61)
  reg_ar_as_w1 reg2_b4 (
    .clk(clk),
    .d(n3[4]),
    .en(1'b1),
    .reset(~rest_n),
    .set(1'b0),
    .q(hsync_cnt[4]));  // sources/rtl/lcd_sync.v(61)
  reg_ar_as_w1 reg2_b5 (
    .clk(clk),
    .d(n3[5]),
    .en(1'b1),
    .reset(~rest_n),
    .set(1'b0),
    .q(hsync_cnt[5]));  // sources/rtl/lcd_sync.v(61)
  reg_ar_as_w1 reg2_b6 (
    .clk(clk),
    .d(n3[6]),
    .en(1'b1),
    .reset(~rest_n),
    .set(1'b0),
    .q(hsync_cnt[6]));  // sources/rtl/lcd_sync.v(61)
  reg_ar_as_w1 reg2_b7 (
    .clk(clk),
    .d(n3[7]),
    .en(1'b1),
    .reset(~rest_n),
    .set(1'b0),
    .q(hsync_cnt[7]));  // sources/rtl/lcd_sync.v(61)
  reg_ar_as_w1 reg2_b8 (
    .clk(clk),
    .d(n3[8]),
    .en(1'b1),
    .reset(~rest_n),
    .set(1'b0),
    .q(hsync_cnt[8]));  // sources/rtl/lcd_sync.v(61)
  reg_ar_as_w1 reg2_b9 (
    .clk(clk),
    .d(n3[9]),
    .en(1'b1),
    .reset(~rest_n),
    .set(1'b0),
    .q(hsync_cnt[9]));  // sources/rtl/lcd_sync.v(61)
  add_pu11_mu11_o12 sub0 (
    .i0(hsync_cnt),
    .i1(11'b00010100000),
    .o(n21));  // sources/rtl/lcd_sync.v(83)
  add_pu11_mu11_o12 sub1 (
    .i0(vsync_cnt),
    .i1(11'b00000101101),
    .o(n24));  // sources/rtl/lcd_sync.v(84)
  add_pu11_mu11_o12 sub2 (
    .i0(hsync_cnt),
    .i1(11'b00000000000),
    .o(n28));  // sources/rtl/lcd_sync.v(93)
  add_pu16_mu16_o16 sub3 (
    .i0({n28[11],n28[11],n28[11],n28[11],n28}),
    .i1(16'b0000000010100000),
    .o(n29[15:0]));  // sources/rtl/lcd_sync.v(93)
  add_pu11_mu11_o12 sub4 (
    .i0(vsync_cnt),
    .i1(11'b00000000001),
    .o(n30));  // sources/rtl/lcd_sync.v(93)
  add_pu13_mu13_o13 sub5 (
    .i0({n30[11],n30}),
    .i1(13'b0000000101101),
    .o(n31[12:0]));  // sources/rtl/lcd_sync.v(93)
  and u11 (n7, n1, n6);  // sources/rtl/lcd_sync.v(70)
  AL_MUX u12 (
    .i0(1'b0),
    .i1(clk),
    .sel(lcd_pwm),
    .o(lcd_clk));  // sources/rtl/lcd_sync.v(74)
  and u14 (lcd_hsync, n11, n12);  // sources/rtl/lcd_sync.v(76)
  and u15 (lcd_vsync, n13, n14);  // sources/rtl/lcd_sync.v(77)
  and u16 (n17, n15, n16);  // sources/rtl/lcd_sync.v(78)
  and u17 (n19, n17, n18);  // sources/rtl/lcd_sync.v(78)
  and u18 (lcd_de, n19, n20);  // sources/rtl/lcd_sync.v(78)
  and u21 (n23, lcd_de, n22);  // sources/rtl/lcd_sync.v(83)
  and u23 (n27, n25, n26);  // sources/rtl/lcd_sync.v(84)
  and u24 (img_ack, n23, n27);  // sources/rtl/lcd_sync.v(84)
  and u9 (n5, n1, n4);  // sources/rtl/lcd_sync.v(68)

endmodule 

module add_pu9_pu9_o9
  (
  i0,
  i1,
  o
  );

  input [8:0] i0;
  input [8:0] i1;
  output [8:0] o;

  wire net_a0;
  wire net_a1;
  wire net_a2;
  wire net_a3;
  wire net_a4;
  wire net_a5;
  wire net_a6;
  wire net_a7;
  wire net_a8;
  wire net_b0;
  wire net_b1;
  wire net_b2;
  wire net_b3;
  wire net_b4;
  wire net_b5;
  wire net_b6;
  wire net_b7;
  wire net_b8;
  wire net_cout0;
  wire net_cout1;
  wire net_cout2;
  wire net_cout3;
  wire net_cout4;
  wire net_cout5;
  wire net_cout6;
  wire net_cout7;
  wire net_cout8;
  wire net_sum0;
  wire net_sum1;
  wire net_sum2;
  wire net_sum3;
  wire net_sum4;
  wire net_sum5;
  wire net_sum6;
  wire net_sum7;
  wire net_sum8;

  assign net_a8 = i0[8];
  assign net_a7 = i0[7];
  assign net_a6 = i0[6];
  assign net_a5 = i0[5];
  assign net_a4 = i0[4];
  assign net_a3 = i0[3];
  assign net_a2 = i0[2];
  assign net_a1 = i0[1];
  assign net_a0 = i0[0];
  assign net_b8 = i1[8];
  assign net_b7 = i1[7];
  assign net_b6 = i1[6];
  assign net_b5 = i1[5];
  assign net_b4 = i1[4];
  assign net_b3 = i1[3];
  assign net_b2 = i1[2];
  assign net_b1 = i1[1];
  assign net_b0 = i1[0];
  assign o[8] = net_sum8;
  assign o[7] = net_sum7;
  assign o[6] = net_sum6;
  assign o[5] = net_sum5;
  assign o[4] = net_sum4;
  assign o[3] = net_sum3;
  assign o[2] = net_sum2;
  assign o[1] = net_sum1;
  assign o[0] = net_sum0;
  AL_FADD comp_0 (
    .a(net_a0),
    .b(net_b0),
    .c(1'b0),
    .cout(net_cout0),
    .sum(net_sum0));
  AL_FADD comp_1 (
    .a(net_a1),
    .b(net_b1),
    .c(net_cout0),
    .cout(net_cout1),
    .sum(net_sum1));
  AL_FADD comp_2 (
    .a(net_a2),
    .b(net_b2),
    .c(net_cout1),
    .cout(net_cout2),
    .sum(net_sum2));
  AL_FADD comp_3 (
    .a(net_a3),
    .b(net_b3),
    .c(net_cout2),
    .cout(net_cout3),
    .sum(net_sum3));
  AL_FADD comp_4 (
    .a(net_a4),
    .b(net_b4),
    .c(net_cout3),
    .cout(net_cout4),
    .sum(net_sum4));
  AL_FADD comp_5 (
    .a(net_a5),
    .b(net_b5),
    .c(net_cout4),
    .cout(net_cout5),
    .sum(net_sum5));
  AL_FADD comp_6 (
    .a(net_a6),
    .b(net_b6),
    .c(net_cout5),
    .cout(net_cout6),
    .sum(net_sum6));
  AL_FADD comp_7 (
    .a(net_a7),
    .b(net_b7),
    .c(net_cout6),
    .cout(net_cout7),
    .sum(net_sum7));
  AL_FADD comp_8 (
    .a(net_a8),
    .b(net_b8),
    .c(net_cout7),
    .cout(net_cout8),
    .sum(net_sum8));

endmodule 

module add_pu8_pu8_o8
  (
  i0,
  i1,
  o
  );

  input [7:0] i0;
  input [7:0] i1;
  output [7:0] o;

  wire net_a0;
  wire net_a1;
  wire net_a2;
  wire net_a3;
  wire net_a4;
  wire net_a5;
  wire net_a6;
  wire net_a7;
  wire net_b0;
  wire net_b1;
  wire net_b2;
  wire net_b3;
  wire net_b4;
  wire net_b5;
  wire net_b6;
  wire net_b7;
  wire net_cout0;
  wire net_cout1;
  wire net_cout2;
  wire net_cout3;
  wire net_cout4;
  wire net_cout5;
  wire net_cout6;
  wire net_cout7;
  wire net_sum0;
  wire net_sum1;
  wire net_sum2;
  wire net_sum3;
  wire net_sum4;
  wire net_sum5;
  wire net_sum6;
  wire net_sum7;

  assign net_a7 = i0[7];
  assign net_a6 = i0[6];
  assign net_a5 = i0[5];
  assign net_a4 = i0[4];
  assign net_a3 = i0[3];
  assign net_a2 = i0[2];
  assign net_a1 = i0[1];
  assign net_a0 = i0[0];
  assign net_b7 = i1[7];
  assign net_b6 = i1[6];
  assign net_b5 = i1[5];
  assign net_b4 = i1[4];
  assign net_b3 = i1[3];
  assign net_b2 = i1[2];
  assign net_b1 = i1[1];
  assign net_b0 = i1[0];
  assign o[7] = net_sum7;
  assign o[6] = net_sum6;
  assign o[5] = net_sum5;
  assign o[4] = net_sum4;
  assign o[3] = net_sum3;
  assign o[2] = net_sum2;
  assign o[1] = net_sum1;
  assign o[0] = net_sum0;
  AL_FADD comp_0 (
    .a(net_a0),
    .b(net_b0),
    .c(1'b0),
    .cout(net_cout0),
    .sum(net_sum0));
  AL_FADD comp_1 (
    .a(net_a1),
    .b(net_b1),
    .c(net_cout0),
    .cout(net_cout1),
    .sum(net_sum1));
  AL_FADD comp_2 (
    .a(net_a2),
    .b(net_b2),
    .c(net_cout1),
    .cout(net_cout2),
    .sum(net_sum2));
  AL_FADD comp_3 (
    .a(net_a3),
    .b(net_b3),
    .c(net_cout2),
    .cout(net_cout3),
    .sum(net_sum3));
  AL_FADD comp_4 (
    .a(net_a4),
    .b(net_b4),
    .c(net_cout3),
    .cout(net_cout4),
    .sum(net_sum4));
  AL_FADD comp_5 (
    .a(net_a5),
    .b(net_b5),
    .c(net_cout4),
    .cout(net_cout5),
    .sum(net_sum5));
  AL_FADD comp_6 (
    .a(net_a6),
    .b(net_b6),
    .c(net_cout5),
    .cout(net_cout6),
    .sum(net_sum6));
  AL_FADD comp_7 (
    .a(net_a7),
    .b(net_b7),
    .c(net_cout6),
    .cout(net_cout7),
    .sum(net_sum7));

endmodule 

module eq_w8
  (
  i0,
  i1,
  o
  );

  input [7:0] i0;
  input [7:0] i1;
  output o;

  wire \or_or_or_xor_i0[0]_i_o ;
  wire \or_or_xor_i0[0]_i1[0_o ;
  wire \or_or_xor_i0[4]_i1[4_o ;
  wire \or_xor_i0[0]_i1[0]_o_o ;
  wire \or_xor_i0[2]_i1[2]_o_o ;
  wire \or_xor_i0[4]_i1[4]_o_o ;
  wire \or_xor_i0[6]_i1[6]_o_o ;
  wire \xor_i0[0]_i1[0]_o ;
  wire \xor_i0[1]_i1[1]_o ;
  wire \xor_i0[2]_i1[2]_o ;
  wire \xor_i0[3]_i1[3]_o ;
  wire \xor_i0[4]_i1[4]_o ;
  wire \xor_i0[5]_i1[5]_o ;
  wire \xor_i0[6]_i1[6]_o ;
  wire \xor_i0[7]_i1[7]_o ;

  not none_diff (o, \or_or_or_xor_i0[0]_i_o );
  or \or_or_or_xor_i0[0]_i  (\or_or_or_xor_i0[0]_i_o , \or_or_xor_i0[0]_i1[0_o , \or_or_xor_i0[4]_i1[4_o );
  or \or_or_xor_i0[0]_i1[0  (\or_or_xor_i0[0]_i1[0_o , \or_xor_i0[0]_i1[0]_o_o , \or_xor_i0[2]_i1[2]_o_o );
  or \or_or_xor_i0[4]_i1[4  (\or_or_xor_i0[4]_i1[4_o , \or_xor_i0[4]_i1[4]_o_o , \or_xor_i0[6]_i1[6]_o_o );
  or \or_xor_i0[0]_i1[0]_o  (\or_xor_i0[0]_i1[0]_o_o , \xor_i0[0]_i1[0]_o , \xor_i0[1]_i1[1]_o );
  or \or_xor_i0[2]_i1[2]_o  (\or_xor_i0[2]_i1[2]_o_o , \xor_i0[2]_i1[2]_o , \xor_i0[3]_i1[3]_o );
  or \or_xor_i0[4]_i1[4]_o  (\or_xor_i0[4]_i1[4]_o_o , \xor_i0[4]_i1[4]_o , \xor_i0[5]_i1[5]_o );
  or \or_xor_i0[6]_i1[6]_o  (\or_xor_i0[6]_i1[6]_o_o , \xor_i0[6]_i1[6]_o , \xor_i0[7]_i1[7]_o );
  xor \xor_i0[0]_i1[0]  (\xor_i0[0]_i1[0]_o , i0[0], i1[0]);
  xor \xor_i0[1]_i1[1]  (\xor_i0[1]_i1[1]_o , i0[1], i1[1]);
  xor \xor_i0[2]_i1[2]  (\xor_i0[2]_i1[2]_o , i0[2], i1[2]);
  xor \xor_i0[3]_i1[3]  (\xor_i0[3]_i1[3]_o , i0[3], i1[3]);
  xor \xor_i0[4]_i1[4]  (\xor_i0[4]_i1[4]_o , i0[4], i1[4]);
  xor \xor_i0[5]_i1[5]  (\xor_i0[5]_i1[5]_o , i0[5], i1[5]);
  xor \xor_i0[6]_i1[6]  (\xor_i0[6]_i1[6]_o , i0[6], i1[6]);
  xor \xor_i0[7]_i1[7]  (\xor_i0[7]_i1[7]_o , i0[7], i1[7]);

endmodule 

module i2c_module  // sources/rtl/i2c_module.v(2)
  (
  address,
  clk,
  reset_n,
  sda_in,
  write,
  writedata,
  ready,
  scl_out,
  sda,
  sda_oe,
  success_out
  );

  input [2:0] address;  // sources/rtl/i2c_module.v(14)
  input clk;  // sources/rtl/i2c_module.v(3)
  input reset_n;  // sources/rtl/i2c_module.v(4)
  input sda_in;  // sources/rtl/i2c_module.v(7)
  input write;  // sources/rtl/i2c_module.v(13)
  input [7:0] writedata;  // sources/rtl/i2c_module.v(12)
  output ready;  // sources/rtl/i2c_module.v(16)
  output scl_out;  // sources/rtl/i2c_module.v(10)
  output sda;  // sources/rtl/i2c_module.v(8)
  output sda_oe;  // sources/rtl/i2c_module.v(6)
  output success_out;  // sources/rtl/i2c_module.v(17)

  // localparam STATE_ADDRESS_ACK = 10;
  // localparam STATE_ADDRESS_BIT_1 = 2;
  // localparam STATE_ADDRESS_BIT_2 = 3;
  // localparam STATE_ADDRESS_BIT_3 = 4;
  // localparam STATE_ADDRESS_BIT_4 = 5;
  // localparam STATE_ADDRESS_BIT_5 = 6;
  // localparam STATE_ADDRESS_BIT_6 = 7;
  // localparam STATE_ADDRESS_BIT_7 = 8;
  // localparam STATE_ADDRESS_BIT_8 = 9;
  // localparam STATE_ADDRESS_START = 1;
  // localparam STATE_ADDRESS_START_2 = 111;
  // localparam STATE_ADDRESS_START_3 = 112;
  // localparam STATE_DATA_ACK = 28;
  // localparam STATE_DATA_BIT_1 = 20;
  // localparam STATE_DATA_BIT_2 = 21;
  // localparam STATE_DATA_BIT_3 = 22;
  // localparam STATE_DATA_BIT_4 = 23;
  // localparam STATE_DATA_BIT_5 = 24;
  // localparam STATE_DATA_BIT_6 = 25;
  // localparam STATE_DATA_BIT_7 = 26;
  // localparam STATE_DATA_BIT_8 = 27;
  // localparam STATE_IDLE = 0;
  // localparam STATE_REG_ACK = 19;
  // localparam STATE_REG_BIT_1 = 11;
  // localparam STATE_REG_BIT_2 = 12;
  // localparam STATE_REG_BIT_3 = 13;
  // localparam STATE_REG_BIT_4 = 14;
  // localparam STATE_REG_BIT_5 = 15;
  // localparam STATE_REG_BIT_6 = 16;
  // localparam STATE_REG_BIT_7 = 17;
  // localparam STATE_REG_BIT_8 = 18;
  // localparam STATE_STOP = 29;
  // localparam STATE_STOP_1 = 30;
  // localparam STATE_STOP_2 = 31;
  // localparam STATE_TRANSIT_1 = 102;
  // localparam STATE_TRANSIT_2 = 192;
  wire [7:0] control_reg;  // sources/rtl/i2c_module.v(85)
  wire [7:0] divider2;  // sources/rtl/i2c_module.v(71)
  wire [7:0] n1;
  wire [7:0] n35;
  wire [7:0] n37;
  wire [7:0] n38;
  wire [7:0] n48;
  wire [7:0] n53;
  wire [7:0] n55;
  wire [7:0] n56;
  wire [7:0] n57;
  wire [7:0] n58;
  wire [7:0] n59;
  wire [7:0] n69;
  wire [7:0] n70;
  wire [7:0] n71;
  wire [7:0] n72;
  wire [7:0] n99;
  wire  \sel0_b0/B0 ;
  wire  \sel0_b0/B1 ;
  wire  \sel0_b0/B10 ;
  wire  \sel0_b0/B11 ;
  wire  \sel0_b0/B12 ;
  wire  \sel0_b0/B13 ;
  wire  \sel0_b0/B14 ;
  wire  \sel0_b0/B15 ;
  wire  \sel0_b0/B16 ;
  wire  \sel0_b0/B17 ;
  wire  \sel0_b0/B18 ;
  wire  \sel0_b0/B19 ;
  wire  \sel0_b0/B2 ;
  wire  \sel0_b0/B20 ;
  wire  \sel0_b0/B21 ;
  wire  \sel0_b0/B22 ;
  wire  \sel0_b0/B23 ;
  wire  \sel0_b0/B24 ;
  wire  \sel0_b0/B25 ;
  wire  \sel0_b0/B26 ;
  wire  \sel0_b0/B27 ;
  wire  \sel0_b0/B28 ;
  wire  \sel0_b0/B29 ;
  wire  \sel0_b0/B3 ;
  wire  \sel0_b0/B30 ;
  wire  \sel0_b0/B31 ;
  wire  \sel0_b0/B32 ;
  wire  \sel0_b0/B33 ;
  wire  \sel0_b0/B34 ;
  wire  \sel0_b0/B35 ;
  wire  \sel0_b0/B36 ;
  wire  \sel0_b0/B4 ;
  wire  \sel0_b0/B5 ;
  wire  \sel0_b0/B6 ;
  wire  \sel0_b0/B7 ;
  wire  \sel0_b0/B8 ;
  wire  \sel0_b0/B9 ;
  wire  \sel0_b1/B0 ;
  wire  \sel0_b1/B1 ;
  wire  \sel0_b1/B10 ;
  wire  \sel0_b1/B11 ;
  wire  \sel0_b1/B12 ;
  wire  \sel0_b1/B13 ;
  wire  \sel0_b1/B14 ;
  wire  \sel0_b1/B15 ;
  wire  \sel0_b1/B16 ;
  wire  \sel0_b1/B17 ;
  wire  \sel0_b1/B18 ;
  wire  \sel0_b1/B19 ;
  wire  \sel0_b1/B2 ;
  wire  \sel0_b1/B20 ;
  wire  \sel0_b1/B21 ;
  wire  \sel0_b1/B22 ;
  wire  \sel0_b1/B23 ;
  wire  \sel0_b1/B24 ;
  wire  \sel0_b1/B25 ;
  wire  \sel0_b1/B26 ;
  wire  \sel0_b1/B27 ;
  wire  \sel0_b1/B28 ;
  wire  \sel0_b1/B29 ;
  wire  \sel0_b1/B3 ;
  wire  \sel0_b1/B30 ;
  wire  \sel0_b1/B31 ;
  wire  \sel0_b1/B32 ;
  wire  \sel0_b1/B33 ;
  wire  \sel0_b1/B34 ;
  wire  \sel0_b1/B35 ;
  wire  \sel0_b1/B36 ;
  wire  \sel0_b1/B4 ;
  wire  \sel0_b1/B5 ;
  wire  \sel0_b1/B6 ;
  wire  \sel0_b1/B7 ;
  wire  \sel0_b1/B8 ;
  wire  \sel0_b1/B9 ;
  wire  \sel0_b2/B0 ;
  wire  \sel0_b2/B1 ;
  wire  \sel0_b2/B10 ;
  wire  \sel0_b2/B11 ;
  wire  \sel0_b2/B12 ;
  wire  \sel0_b2/B13 ;
  wire  \sel0_b2/B14 ;
  wire  \sel0_b2/B15 ;
  wire  \sel0_b2/B16 ;
  wire  \sel0_b2/B17 ;
  wire  \sel0_b2/B18 ;
  wire  \sel0_b2/B19 ;
  wire  \sel0_b2/B2 ;
  wire  \sel0_b2/B20 ;
  wire  \sel0_b2/B21 ;
  wire  \sel0_b2/B22 ;
  wire  \sel0_b2/B23 ;
  wire  \sel0_b2/B24 ;
  wire  \sel0_b2/B25 ;
  wire  \sel0_b2/B26 ;
  wire  \sel0_b2/B27 ;
  wire  \sel0_b2/B28 ;
  wire  \sel0_b2/B29 ;
  wire  \sel0_b2/B3 ;
  wire  \sel0_b2/B30 ;
  wire  \sel0_b2/B31 ;
  wire  \sel0_b2/B32 ;
  wire  \sel0_b2/B33 ;
  wire  \sel0_b2/B34 ;
  wire  \sel0_b2/B35 ;
  wire  \sel0_b2/B36 ;
  wire  \sel0_b2/B4 ;
  wire  \sel0_b2/B5 ;
  wire  \sel0_b2/B6 ;
  wire  \sel0_b2/B7 ;
  wire  \sel0_b2/B8 ;
  wire  \sel0_b2/B9 ;
  wire  \sel0_b3/B0 ;
  wire  \sel0_b3/B1 ;
  wire  \sel0_b3/B10 ;
  wire  \sel0_b3/B11 ;
  wire  \sel0_b3/B12 ;
  wire  \sel0_b3/B13 ;
  wire  \sel0_b3/B14 ;
  wire  \sel0_b3/B15 ;
  wire  \sel0_b3/B16 ;
  wire  \sel0_b3/B17 ;
  wire  \sel0_b3/B18 ;
  wire  \sel0_b3/B19 ;
  wire  \sel0_b3/B2 ;
  wire  \sel0_b3/B20 ;
  wire  \sel0_b3/B21 ;
  wire  \sel0_b3/B22 ;
  wire  \sel0_b3/B23 ;
  wire  \sel0_b3/B24 ;
  wire  \sel0_b3/B25 ;
  wire  \sel0_b3/B26 ;
  wire  \sel0_b3/B27 ;
  wire  \sel0_b3/B28 ;
  wire  \sel0_b3/B29 ;
  wire  \sel0_b3/B3 ;
  wire  \sel0_b3/B30 ;
  wire  \sel0_b3/B31 ;
  wire  \sel0_b3/B32 ;
  wire  \sel0_b3/B33 ;
  wire  \sel0_b3/B34 ;
  wire  \sel0_b3/B35 ;
  wire  \sel0_b3/B36 ;
  wire  \sel0_b3/B4 ;
  wire  \sel0_b3/B5 ;
  wire  \sel0_b3/B6 ;
  wire  \sel0_b3/B7 ;
  wire  \sel0_b3/B8 ;
  wire  \sel0_b3/B9 ;
  wire  \sel0_b4/B0 ;
  wire  \sel0_b4/B1 ;
  wire  \sel0_b4/B10 ;
  wire  \sel0_b4/B11 ;
  wire  \sel0_b4/B12 ;
  wire  \sel0_b4/B13 ;
  wire  \sel0_b4/B14 ;
  wire  \sel0_b4/B15 ;
  wire  \sel0_b4/B16 ;
  wire  \sel0_b4/B17 ;
  wire  \sel0_b4/B18 ;
  wire  \sel0_b4/B19 ;
  wire  \sel0_b4/B2 ;
  wire  \sel0_b4/B20 ;
  wire  \sel0_b4/B21 ;
  wire  \sel0_b4/B22 ;
  wire  \sel0_b4/B23 ;
  wire  \sel0_b4/B24 ;
  wire  \sel0_b4/B25 ;
  wire  \sel0_b4/B26 ;
  wire  \sel0_b4/B27 ;
  wire  \sel0_b4/B28 ;
  wire  \sel0_b4/B29 ;
  wire  \sel0_b4/B3 ;
  wire  \sel0_b4/B30 ;
  wire  \sel0_b4/B31 ;
  wire  \sel0_b4/B32 ;
  wire  \sel0_b4/B33 ;
  wire  \sel0_b4/B34 ;
  wire  \sel0_b4/B35 ;
  wire  \sel0_b4/B36 ;
  wire  \sel0_b4/B4 ;
  wire  \sel0_b4/B5 ;
  wire  \sel0_b4/B6 ;
  wire  \sel0_b4/B7 ;
  wire  \sel0_b4/B8 ;
  wire  \sel0_b4/B9 ;
  wire  \sel0_b5/B0 ;
  wire  \sel0_b5/B1 ;
  wire  \sel0_b5/B10 ;
  wire  \sel0_b5/B11 ;
  wire  \sel0_b5/B12 ;
  wire  \sel0_b5/B13 ;
  wire  \sel0_b5/B14 ;
  wire  \sel0_b5/B15 ;
  wire  \sel0_b5/B16 ;
  wire  \sel0_b5/B17 ;
  wire  \sel0_b5/B18 ;
  wire  \sel0_b5/B19 ;
  wire  \sel0_b5/B2 ;
  wire  \sel0_b5/B20 ;
  wire  \sel0_b5/B21 ;
  wire  \sel0_b5/B22 ;
  wire  \sel0_b5/B23 ;
  wire  \sel0_b5/B24 ;
  wire  \sel0_b5/B25 ;
  wire  \sel0_b5/B26 ;
  wire  \sel0_b5/B27 ;
  wire  \sel0_b5/B28 ;
  wire  \sel0_b5/B29 ;
  wire  \sel0_b5/B3 ;
  wire  \sel0_b5/B30 ;
  wire  \sel0_b5/B31 ;
  wire  \sel0_b5/B32 ;
  wire  \sel0_b5/B33 ;
  wire  \sel0_b5/B34 ;
  wire  \sel0_b5/B35 ;
  wire  \sel0_b5/B36 ;
  wire  \sel0_b5/B4 ;
  wire  \sel0_b5/B5 ;
  wire  \sel0_b5/B6 ;
  wire  \sel0_b5/B7 ;
  wire  \sel0_b5/B8 ;
  wire  \sel0_b5/B9 ;
  wire  \sel0_b6/B0 ;
  wire  \sel0_b6/B1 ;
  wire  \sel0_b6/B10 ;
  wire  \sel0_b6/B11 ;
  wire  \sel0_b6/B12 ;
  wire  \sel0_b6/B13 ;
  wire  \sel0_b6/B14 ;
  wire  \sel0_b6/B15 ;
  wire  \sel0_b6/B16 ;
  wire  \sel0_b6/B17 ;
  wire  \sel0_b6/B18 ;
  wire  \sel0_b6/B19 ;
  wire  \sel0_b6/B2 ;
  wire  \sel0_b6/B20 ;
  wire  \sel0_b6/B21 ;
  wire  \sel0_b6/B22 ;
  wire  \sel0_b6/B23 ;
  wire  \sel0_b6/B24 ;
  wire  \sel0_b6/B25 ;
  wire  \sel0_b6/B26 ;
  wire  \sel0_b6/B27 ;
  wire  \sel0_b6/B28 ;
  wire  \sel0_b6/B29 ;
  wire  \sel0_b6/B3 ;
  wire  \sel0_b6/B30 ;
  wire  \sel0_b6/B31 ;
  wire  \sel0_b6/B32 ;
  wire  \sel0_b6/B33 ;
  wire  \sel0_b6/B34 ;
  wire  \sel0_b6/B35 ;
  wire  \sel0_b6/B36 ;
  wire  \sel0_b6/B4 ;
  wire  \sel0_b6/B5 ;
  wire  \sel0_b6/B6 ;
  wire  \sel0_b6/B7 ;
  wire  \sel0_b6/B8 ;
  wire  \sel0_b6/B9 ;
  wire  \sel0_b7/B0 ;
  wire  \sel0_b7/B1 ;
  wire  \sel0_b7/B10 ;
  wire  \sel0_b7/B11 ;
  wire  \sel0_b7/B12 ;
  wire  \sel0_b7/B13 ;
  wire  \sel0_b7/B14 ;
  wire  \sel0_b7/B15 ;
  wire  \sel0_b7/B16 ;
  wire  \sel0_b7/B17 ;
  wire  \sel0_b7/B18 ;
  wire  \sel0_b7/B19 ;
  wire  \sel0_b7/B2 ;
  wire  \sel0_b7/B20 ;
  wire  \sel0_b7/B21 ;
  wire  \sel0_b7/B22 ;
  wire  \sel0_b7/B23 ;
  wire  \sel0_b7/B24 ;
  wire  \sel0_b7/B25 ;
  wire  \sel0_b7/B26 ;
  wire  \sel0_b7/B27 ;
  wire  \sel0_b7/B28 ;
  wire  \sel0_b7/B29 ;
  wire  \sel0_b7/B3 ;
  wire  \sel0_b7/B30 ;
  wire  \sel0_b7/B31 ;
  wire  \sel0_b7/B32 ;
  wire  \sel0_b7/B33 ;
  wire  \sel0_b7/B34 ;
  wire  \sel0_b7/B35 ;
  wire  \sel0_b7/B36 ;
  wire  \sel0_b7/B4 ;
  wire  \sel0_b7/B5 ;
  wire  \sel0_b7/B6 ;
  wire  \sel0_b7/B7 ;
  wire  \sel0_b7/B8 ;
  wire  \sel0_b7/B9 ;
  wire  \sel1/B0 ;
  wire  \sel1/B1 ;
  wire  \sel1/B10 ;
  wire  \sel1/B11 ;
  wire  \sel1/B12 ;
  wire  \sel1/B13 ;
  wire  \sel1/B14 ;
  wire  \sel1/B15 ;
  wire  \sel1/B16 ;
  wire  \sel1/B17 ;
  wire  \sel1/B18 ;
  wire  \sel1/B19 ;
  wire  \sel1/B2 ;
  wire  \sel1/B20 ;
  wire  \sel1/B21 ;
  wire  \sel1/B22 ;
  wire  \sel1/B23 ;
  wire  \sel1/B24 ;
  wire  \sel1/B25 ;
  wire  \sel1/B26 ;
  wire  \sel1/B27 ;
  wire  \sel1/B28 ;
  wire  \sel1/B29 ;
  wire  \sel1/B3 ;
  wire  \sel1/B30 ;
  wire  \sel1/B31 ;
  wire  \sel1/B32 ;
  wire  \sel1/B33 ;
  wire  \sel1/B34 ;
  wire  \sel1/B4 ;
  wire  \sel1/B5 ;
  wire  \sel1/B6 ;
  wire  \sel1/B7 ;
  wire  \sel1/B8 ;
  wire  \sel1/B9 ;
  wire  \sel2/B0 ;
  wire  \sel2/B1 ;
  wire  \sel2/B10 ;
  wire  \sel2/B11 ;
  wire  \sel2/B12 ;
  wire  \sel2/B13 ;
  wire  \sel2/B14 ;
  wire  \sel2/B15 ;
  wire  \sel2/B16 ;
  wire  \sel2/B17 ;
  wire  \sel2/B18 ;
  wire  \sel2/B19 ;
  wire  \sel2/B2 ;
  wire  \sel2/B20 ;
  wire  \sel2/B21 ;
  wire  \sel2/B22 ;
  wire  \sel2/B23 ;
  wire  \sel2/B24 ;
  wire  \sel2/B25 ;
  wire  \sel2/B26 ;
  wire  \sel2/B27 ;
  wire  \sel2/B28 ;
  wire  \sel2/B29 ;
  wire  \sel2/B3 ;
  wire  \sel2/B30 ;
  wire  \sel2/B31 ;
  wire  \sel2/B32 ;
  wire  \sel2/B33 ;
  wire  \sel2/B34 ;
  wire  \sel2/B4 ;
  wire  \sel2/B5 ;
  wire  \sel2/B6 ;
  wire  \sel2/B7 ;
  wire  \sel2/B8 ;
  wire  \sel2/B9 ;
  wire  \sel3/B0 ;
  wire  \sel3/B1 ;
  wire  \sel3/B10 ;
  wire  \sel3/B11 ;
  wire  \sel3/B12 ;
  wire  \sel3/B13 ;
  wire  \sel3/B14 ;
  wire  \sel3/B15 ;
  wire  \sel3/B16 ;
  wire  \sel3/B17 ;
  wire  \sel3/B18 ;
  wire  \sel3/B19 ;
  wire  \sel3/B2 ;
  wire  \sel3/B20 ;
  wire  \sel3/B21 ;
  wire  \sel3/B22 ;
  wire  \sel3/B23 ;
  wire  \sel3/B24 ;
  wire  \sel3/B25 ;
  wire  \sel3/B26 ;
  wire  \sel3/B27 ;
  wire  \sel3/B28 ;
  wire  \sel3/B29 ;
  wire  \sel3/B3 ;
  wire  \sel3/B30 ;
  wire  \sel3/B31 ;
  wire  \sel3/B32 ;
  wire  \sel3/B33 ;
  wire  \sel3/B34 ;
  wire  \sel3/B4 ;
  wire  \sel3/B5 ;
  wire  \sel3/B6 ;
  wire  \sel3/B7 ;
  wire  \sel3/B8 ;
  wire  \sel3/B9 ;
  wire  \sel4/B0 ;
  wire  \sel4/B1 ;
  wire  \sel4/B10 ;
  wire  \sel4/B11 ;
  wire  \sel4/B12 ;
  wire  \sel4/B13 ;
  wire  \sel4/B14 ;
  wire  \sel4/B15 ;
  wire  \sel4/B16 ;
  wire  \sel4/B17 ;
  wire  \sel4/B18 ;
  wire  \sel4/B19 ;
  wire  \sel4/B2 ;
  wire  \sel4/B20 ;
  wire  \sel4/B21 ;
  wire  \sel4/B22 ;
  wire  \sel4/B23 ;
  wire  \sel4/B24 ;
  wire  \sel4/B25 ;
  wire  \sel4/B26 ;
  wire  \sel4/B27 ;
  wire  \sel4/B28 ;
  wire  \sel4/B29 ;
  wire  \sel4/B3 ;
  wire  \sel4/B30 ;
  wire  \sel4/B31 ;
  wire  \sel4/B32 ;
  wire  \sel4/B33 ;
  wire  \sel4/B34 ;
  wire  \sel4/B4 ;
  wire  \sel4/B5 ;
  wire  \sel4/B6 ;
  wire  \sel4/B7 ;
  wire  \sel4/B8 ;
  wire  \sel4/B9 ;
  wire  \sel5/B0 ;
  wire  \sel5/B1 ;
  wire  \sel5/B10 ;
  wire  \sel5/B11 ;
  wire  \sel5/B12 ;
  wire  \sel5/B13 ;
  wire  \sel5/B14 ;
  wire  \sel5/B15 ;
  wire  \sel5/B16 ;
  wire  \sel5/B17 ;
  wire  \sel5/B18 ;
  wire  \sel5/B19 ;
  wire  \sel5/B2 ;
  wire  \sel5/B20 ;
  wire  \sel5/B21 ;
  wire  \sel5/B22 ;
  wire  \sel5/B23 ;
  wire  \sel5/B24 ;
  wire  \sel5/B25 ;
  wire  \sel5/B26 ;
  wire  \sel5/B27 ;
  wire  \sel5/B28 ;
  wire  \sel5/B29 ;
  wire  \sel5/B3 ;
  wire  \sel5/B30 ;
  wire  \sel5/B31 ;
  wire  \sel5/B32 ;
  wire  \sel5/B33 ;
  wire  \sel5/B34 ;
  wire  \sel5/B4 ;
  wire  \sel5/B5 ;
  wire  \sel5/B6 ;
  wire  \sel5/B7 ;
  wire  \sel5/B8 ;
  wire  \sel5/B9 ;
  wire  \sel6/B0 ;
  wire  \sel6/B1 ;
  wire  \sel6/B10 ;
  wire  \sel6/B11 ;
  wire  \sel6/B12 ;
  wire  \sel6/B13 ;
  wire  \sel6/B14 ;
  wire  \sel6/B15 ;
  wire  \sel6/B16 ;
  wire  \sel6/B17 ;
  wire  \sel6/B18 ;
  wire  \sel6/B19 ;
  wire  \sel6/B2 ;
  wire  \sel6/B20 ;
  wire  \sel6/B21 ;
  wire  \sel6/B22 ;
  wire  \sel6/B23 ;
  wire  \sel6/B24 ;
  wire  \sel6/B25 ;
  wire  \sel6/B26 ;
  wire  \sel6/B27 ;
  wire  \sel6/B28 ;
  wire  \sel6/B29 ;
  wire  \sel6/B3 ;
  wire  \sel6/B30 ;
  wire  \sel6/B31 ;
  wire  \sel6/B32 ;
  wire  \sel6/B33 ;
  wire  \sel6/B34 ;
  wire  \sel6/B4 ;
  wire  \sel6/B5 ;
  wire  \sel6/B6 ;
  wire  \sel6/B7 ;
  wire  \sel6/B8 ;
  wire  \sel6/B9 ;
  wire [7:0] slave_address;  // sources/rtl/i2c_module.v(86)
  wire [7:0] slave_data_1;  // sources/rtl/i2c_module.v(88)
  wire [7:0] slave_reg_address;  // sources/rtl/i2c_module.v(87)
  wire [7:0] state_next;  // sources/rtl/i2c_module.v(21)
  wire ack_ok;  // sources/rtl/i2c_module.v(143)
  wire \address[0]_neg ;
  wire \address[1]_neg ;
  wire clk_div;  // sources/rtl/i2c_module.v(69)
  wire mux0_b0_sel_is_3_o;
  wire mux1_b0_sel_is_2_o;
  wire mux2_b0_sel_is_1_o;
  wire mux3_b0_sel_is_0_o;
  wire mux4_b0_sel_is_3_o;
  wire mux5_b0_sel_is_3_o;
  wire mux6_b0_sel_is_3_o;
  wire mux7_b0_sel_is_3_o;
  wire mux9_b0_sel_is_0_o;
  wire n0;
  wire n102;
  wire n103;
  wire n104;
  wire n105;
  wire n106;
  wire n107;
  wire n108;
  wire n109;
  wire n11;
  wire n110;
  wire n111;
  wire n112;
  wire n113;
  wire n114;
  wire n115;
  wire n116;
  wire n117;
  wire n118;
  wire n119;
  wire n11_neg;
  wire n120;
  wire n121;
  wire n122;
  wire n123;
  wire n124;
  wire n125;
  wire n126;
  wire n127;
  wire n128;
  wire n129;
  wire n130;
  wire n131;
  wire n132;
  wire n133;
  wire n134;
  wire n135;
  wire n136;
  wire n137;
  wire n138;
  wire n139;
  wire n140;
  wire n141;
  wire n142;
  wire n143;
  wire n144;
  wire n145;
  wire n146;
  wire n147;
  wire n148;
  wire n149;
  wire n150;
  wire n151;
  wire n152;
  wire n153;
  wire n154;
  wire n155;
  wire n156;
  wire n157;
  wire n158;
  wire n159;
  wire n160;
  wire n161;
  wire n162;
  wire n163;
  wire n164;
  wire n165;
  wire n166;
  wire n167;
  wire n168;
  wire n169;
  wire n17;
  wire n170;
  wire n171;
  wire n172;
  wire n173;
  wire n174;
  wire n175;
  wire n176;
  wire n177;
  wire n178;
  wire n179;
  wire n18;
  wire n180;
  wire n181;
  wire n182;
  wire n183;
  wire n184;
  wire n185;
  wire n186;
  wire n187;
  wire n188;
  wire n189;
  wire n19;
  wire n190;
  wire n191;
  wire n192;
  wire n193;
  wire n194;
  wire n2;
  wire n20;
  wire n21;
  wire n22;
  wire n23;
  wire n24;
  wire n25;
  wire n26;
  wire n27;
  wire n28;
  wire n29;
  wire n2_neg;
  wire n30;
  wire n31;
  wire n32;
  wire n33;
  wire n36;
  wire n73;
  wire n74;
  wire n75;
  wire n76;
  wire n77;
  wire n78;
  wire n79;
  wire n80;
  wire n81;
  wire n82;
  wire n83;
  wire n84;
  wire n85;
  wire n86;
  wire n87;
  wire n88;
  wire n89;
  wire n90;
  wire n91;
  wire n92;
  wire n93;
  wire n94;
  wire n95;
  wire n96;
  wire n97;
  wire n98;
  wire scl_output_enable;  // sources/rtl/i2c_module.v(120)
  wire scl_output_zero;  // sources/rtl/i2c_module.v(121)
  wire \sel0_b0/or_B0_B1_o ;
  wire \sel0_b0/or_B11_B12_o ;
  wire \sel0_b0/or_B13_B14_o ;
  wire \sel0_b0/or_B15_or_B16_B17_o_o ;
  wire \sel0_b0/or_B16_B17_o ;
  wire \sel0_b0/or_B18_B19_o ;
  wire \sel0_b0/or_B20_B21_o ;
  wire \sel0_b0/or_B22_B23_o ;
  wire \sel0_b0/or_B24_or_B25_B26_o_o ;
  wire \sel0_b0/or_B25_B26_o ;
  wire \sel0_b0/or_B27_B28_o ;
  wire \sel0_b0/or_B29_or_B30_B31_o_o ;
  wire \sel0_b0/or_B2_B3_o ;
  wire \sel0_b0/or_B30_B31_o ;
  wire \sel0_b0/or_B32_B33_o ;
  wire \sel0_b0/or_B34_or_B35_B36_o_o ;
  wire \sel0_b0/or_B35_B36_o ;
  wire \sel0_b0/or_B4_B5_o ;
  wire \sel0_b0/or_B6_or_B7_B8_o_o ;
  wire \sel0_b0/or_B7_B8_o ;
  wire \sel0_b0/or_B9_B10_o ;
  wire \sel0_b0/or_or_B0_B1_o_or_B2__o ;
  wire \sel0_b0/or_or_B13_B14_o_or_B_o ;
  wire \sel0_b0/or_or_B18_B19_o_or_B_o ;
  wire \sel0_b0/or_or_B22_B23_o_or_B_o ;
  wire \sel0_b0/or_or_B27_B28_o_or_B_o ;
  wire \sel0_b0/or_or_B32_B33_o_or_B_o ;
  wire \sel0_b0/or_or_B4_B5_o_or_B6__o ;
  wire \sel0_b0/or_or_B9_B10_o_or_B1_o ;
  wire \sel0_b0/or_or_or_B0_B1_o_or__o ;
  wire \sel0_b0/or_or_or_B18_B19_o_o_o ;
  wire \sel0_b0/or_or_or_B27_B28_o_o_o ;
  wire \sel0_b0/or_or_or_B9_B10_o_or_o ;
  wire \sel0_b0/or_or_or_or_B0_B1_o__o ;
  wire \sel0_b0/or_or_or_or_B18_B19__o ;
  wire \sel0_b1/or_B0_B1_o ;
  wire \sel0_b1/or_B11_B12_o ;
  wire \sel0_b1/or_B13_B14_o ;
  wire \sel0_b1/or_B15_or_B16_B17_o_o ;
  wire \sel0_b1/or_B16_B17_o ;
  wire \sel0_b1/or_B18_B19_o ;
  wire \sel0_b1/or_B20_B21_o ;
  wire \sel0_b1/or_B22_B23_o ;
  wire \sel0_b1/or_B24_or_B25_B26_o_o ;
  wire \sel0_b1/or_B25_B26_o ;
  wire \sel0_b1/or_B27_B28_o ;
  wire \sel0_b1/or_B29_or_B30_B31_o_o ;
  wire \sel0_b1/or_B2_B3_o ;
  wire \sel0_b1/or_B30_B31_o ;
  wire \sel0_b1/or_B32_B33_o ;
  wire \sel0_b1/or_B34_or_B35_B36_o_o ;
  wire \sel0_b1/or_B35_B36_o ;
  wire \sel0_b1/or_B4_B5_o ;
  wire \sel0_b1/or_B6_or_B7_B8_o_o ;
  wire \sel0_b1/or_B7_B8_o ;
  wire \sel0_b1/or_B9_B10_o ;
  wire \sel0_b1/or_or_B0_B1_o_or_B2__o ;
  wire \sel0_b1/or_or_B13_B14_o_or_B_o ;
  wire \sel0_b1/or_or_B18_B19_o_or_B_o ;
  wire \sel0_b1/or_or_B22_B23_o_or_B_o ;
  wire \sel0_b1/or_or_B27_B28_o_or_B_o ;
  wire \sel0_b1/or_or_B32_B33_o_or_B_o ;
  wire \sel0_b1/or_or_B4_B5_o_or_B6__o ;
  wire \sel0_b1/or_or_B9_B10_o_or_B1_o ;
  wire \sel0_b1/or_or_or_B0_B1_o_or__o ;
  wire \sel0_b1/or_or_or_B18_B19_o_o_o ;
  wire \sel0_b1/or_or_or_B27_B28_o_o_o ;
  wire \sel0_b1/or_or_or_B9_B10_o_or_o ;
  wire \sel0_b1/or_or_or_or_B0_B1_o__o ;
  wire \sel0_b1/or_or_or_or_B18_B19__o ;
  wire \sel0_b2/or_B0_B1_o ;
  wire \sel0_b2/or_B11_B12_o ;
  wire \sel0_b2/or_B13_B14_o ;
  wire \sel0_b2/or_B15_or_B16_B17_o_o ;
  wire \sel0_b2/or_B16_B17_o ;
  wire \sel0_b2/or_B18_B19_o ;
  wire \sel0_b2/or_B20_B21_o ;
  wire \sel0_b2/or_B22_B23_o ;
  wire \sel0_b2/or_B24_or_B25_B26_o_o ;
  wire \sel0_b2/or_B25_B26_o ;
  wire \sel0_b2/or_B27_B28_o ;
  wire \sel0_b2/or_B29_or_B30_B31_o_o ;
  wire \sel0_b2/or_B2_B3_o ;
  wire \sel0_b2/or_B30_B31_o ;
  wire \sel0_b2/or_B32_B33_o ;
  wire \sel0_b2/or_B34_or_B35_B36_o_o ;
  wire \sel0_b2/or_B35_B36_o ;
  wire \sel0_b2/or_B4_B5_o ;
  wire \sel0_b2/or_B6_or_B7_B8_o_o ;
  wire \sel0_b2/or_B7_B8_o ;
  wire \sel0_b2/or_B9_B10_o ;
  wire \sel0_b2/or_or_B0_B1_o_or_B2__o ;
  wire \sel0_b2/or_or_B13_B14_o_or_B_o ;
  wire \sel0_b2/or_or_B18_B19_o_or_B_o ;
  wire \sel0_b2/or_or_B22_B23_o_or_B_o ;
  wire \sel0_b2/or_or_B27_B28_o_or_B_o ;
  wire \sel0_b2/or_or_B32_B33_o_or_B_o ;
  wire \sel0_b2/or_or_B4_B5_o_or_B6__o ;
  wire \sel0_b2/or_or_B9_B10_o_or_B1_o ;
  wire \sel0_b2/or_or_or_B0_B1_o_or__o ;
  wire \sel0_b2/or_or_or_B18_B19_o_o_o ;
  wire \sel0_b2/or_or_or_B27_B28_o_o_o ;
  wire \sel0_b2/or_or_or_B9_B10_o_or_o ;
  wire \sel0_b2/or_or_or_or_B0_B1_o__o ;
  wire \sel0_b2/or_or_or_or_B18_B19__o ;
  wire \sel0_b3/or_B0_B1_o ;
  wire \sel0_b3/or_B11_B12_o ;
  wire \sel0_b3/or_B13_B14_o ;
  wire \sel0_b3/or_B15_or_B16_B17_o_o ;
  wire \sel0_b3/or_B16_B17_o ;
  wire \sel0_b3/or_B18_B19_o ;
  wire \sel0_b3/or_B20_B21_o ;
  wire \sel0_b3/or_B22_B23_o ;
  wire \sel0_b3/or_B24_or_B25_B26_o_o ;
  wire \sel0_b3/or_B25_B26_o ;
  wire \sel0_b3/or_B27_B28_o ;
  wire \sel0_b3/or_B29_or_B30_B31_o_o ;
  wire \sel0_b3/or_B2_B3_o ;
  wire \sel0_b3/or_B30_B31_o ;
  wire \sel0_b3/or_B32_B33_o ;
  wire \sel0_b3/or_B34_or_B35_B36_o_o ;
  wire \sel0_b3/or_B35_B36_o ;
  wire \sel0_b3/or_B4_B5_o ;
  wire \sel0_b3/or_B6_or_B7_B8_o_o ;
  wire \sel0_b3/or_B7_B8_o ;
  wire \sel0_b3/or_B9_B10_o ;
  wire \sel0_b3/or_or_B0_B1_o_or_B2__o ;
  wire \sel0_b3/or_or_B13_B14_o_or_B_o ;
  wire \sel0_b3/or_or_B18_B19_o_or_B_o ;
  wire \sel0_b3/or_or_B22_B23_o_or_B_o ;
  wire \sel0_b3/or_or_B27_B28_o_or_B_o ;
  wire \sel0_b3/or_or_B32_B33_o_or_B_o ;
  wire \sel0_b3/or_or_B4_B5_o_or_B6__o ;
  wire \sel0_b3/or_or_B9_B10_o_or_B1_o ;
  wire \sel0_b3/or_or_or_B0_B1_o_or__o ;
  wire \sel0_b3/or_or_or_B18_B19_o_o_o ;
  wire \sel0_b3/or_or_or_B27_B28_o_o_o ;
  wire \sel0_b3/or_or_or_B9_B10_o_or_o ;
  wire \sel0_b3/or_or_or_or_B0_B1_o__o ;
  wire \sel0_b3/or_or_or_or_B18_B19__o ;
  wire \sel0_b4/or_B0_B1_o ;
  wire \sel0_b4/or_B11_B12_o ;
  wire \sel0_b4/or_B13_B14_o ;
  wire \sel0_b4/or_B15_or_B16_B17_o_o ;
  wire \sel0_b4/or_B16_B17_o ;
  wire \sel0_b4/or_B18_B19_o ;
  wire \sel0_b4/or_B20_B21_o ;
  wire \sel0_b4/or_B22_B23_o ;
  wire \sel0_b4/or_B24_or_B25_B26_o_o ;
  wire \sel0_b4/or_B25_B26_o ;
  wire \sel0_b4/or_B27_B28_o ;
  wire \sel0_b4/or_B29_or_B30_B31_o_o ;
  wire \sel0_b4/or_B2_B3_o ;
  wire \sel0_b4/or_B30_B31_o ;
  wire \sel0_b4/or_B32_B33_o ;
  wire \sel0_b4/or_B34_or_B35_B36_o_o ;
  wire \sel0_b4/or_B35_B36_o ;
  wire \sel0_b4/or_B4_B5_o ;
  wire \sel0_b4/or_B6_or_B7_B8_o_o ;
  wire \sel0_b4/or_B7_B8_o ;
  wire \sel0_b4/or_B9_B10_o ;
  wire \sel0_b4/or_or_B0_B1_o_or_B2__o ;
  wire \sel0_b4/or_or_B13_B14_o_or_B_o ;
  wire \sel0_b4/or_or_B18_B19_o_or_B_o ;
  wire \sel0_b4/or_or_B22_B23_o_or_B_o ;
  wire \sel0_b4/or_or_B27_B28_o_or_B_o ;
  wire \sel0_b4/or_or_B32_B33_o_or_B_o ;
  wire \sel0_b4/or_or_B4_B5_o_or_B6__o ;
  wire \sel0_b4/or_or_B9_B10_o_or_B1_o ;
  wire \sel0_b4/or_or_or_B0_B1_o_or__o ;
  wire \sel0_b4/or_or_or_B18_B19_o_o_o ;
  wire \sel0_b4/or_or_or_B27_B28_o_o_o ;
  wire \sel0_b4/or_or_or_B9_B10_o_or_o ;
  wire \sel0_b4/or_or_or_or_B0_B1_o__o ;
  wire \sel0_b4/or_or_or_or_B18_B19__o ;
  wire \sel0_b5/or_B0_B1_o ;
  wire \sel0_b5/or_B11_B12_o ;
  wire \sel0_b5/or_B13_B14_o ;
  wire \sel0_b5/or_B15_or_B16_B17_o_o ;
  wire \sel0_b5/or_B16_B17_o ;
  wire \sel0_b5/or_B18_B19_o ;
  wire \sel0_b5/or_B20_B21_o ;
  wire \sel0_b5/or_B22_B23_o ;
  wire \sel0_b5/or_B24_or_B25_B26_o_o ;
  wire \sel0_b5/or_B25_B26_o ;
  wire \sel0_b5/or_B27_B28_o ;
  wire \sel0_b5/or_B29_or_B30_B31_o_o ;
  wire \sel0_b5/or_B2_B3_o ;
  wire \sel0_b5/or_B30_B31_o ;
  wire \sel0_b5/or_B32_B33_o ;
  wire \sel0_b5/or_B34_or_B35_B36_o_o ;
  wire \sel0_b5/or_B35_B36_o ;
  wire \sel0_b5/or_B4_B5_o ;
  wire \sel0_b5/or_B6_or_B7_B8_o_o ;
  wire \sel0_b5/or_B7_B8_o ;
  wire \sel0_b5/or_B9_B10_o ;
  wire \sel0_b5/or_or_B0_B1_o_or_B2__o ;
  wire \sel0_b5/or_or_B13_B14_o_or_B_o ;
  wire \sel0_b5/or_or_B18_B19_o_or_B_o ;
  wire \sel0_b5/or_or_B22_B23_o_or_B_o ;
  wire \sel0_b5/or_or_B27_B28_o_or_B_o ;
  wire \sel0_b5/or_or_B32_B33_o_or_B_o ;
  wire \sel0_b5/or_or_B4_B5_o_or_B6__o ;
  wire \sel0_b5/or_or_B9_B10_o_or_B1_o ;
  wire \sel0_b5/or_or_or_B0_B1_o_or__o ;
  wire \sel0_b5/or_or_or_B18_B19_o_o_o ;
  wire \sel0_b5/or_or_or_B27_B28_o_o_o ;
  wire \sel0_b5/or_or_or_B9_B10_o_or_o ;
  wire \sel0_b5/or_or_or_or_B0_B1_o__o ;
  wire \sel0_b5/or_or_or_or_B18_B19__o ;
  wire \sel0_b6/or_B0_B1_o ;
  wire \sel0_b6/or_B11_B12_o ;
  wire \sel0_b6/or_B13_B14_o ;
  wire \sel0_b6/or_B15_or_B16_B17_o_o ;
  wire \sel0_b6/or_B16_B17_o ;
  wire \sel0_b6/or_B18_B19_o ;
  wire \sel0_b6/or_B20_B21_o ;
  wire \sel0_b6/or_B22_B23_o ;
  wire \sel0_b6/or_B24_or_B25_B26_o_o ;
  wire \sel0_b6/or_B25_B26_o ;
  wire \sel0_b6/or_B27_B28_o ;
  wire \sel0_b6/or_B29_or_B30_B31_o_o ;
  wire \sel0_b6/or_B2_B3_o ;
  wire \sel0_b6/or_B30_B31_o ;
  wire \sel0_b6/or_B32_B33_o ;
  wire \sel0_b6/or_B34_or_B35_B36_o_o ;
  wire \sel0_b6/or_B35_B36_o ;
  wire \sel0_b6/or_B4_B5_o ;
  wire \sel0_b6/or_B6_or_B7_B8_o_o ;
  wire \sel0_b6/or_B7_B8_o ;
  wire \sel0_b6/or_B9_B10_o ;
  wire \sel0_b6/or_or_B0_B1_o_or_B2__o ;
  wire \sel0_b6/or_or_B13_B14_o_or_B_o ;
  wire \sel0_b6/or_or_B18_B19_o_or_B_o ;
  wire \sel0_b6/or_or_B22_B23_o_or_B_o ;
  wire \sel0_b6/or_or_B27_B28_o_or_B_o ;
  wire \sel0_b6/or_or_B32_B33_o_or_B_o ;
  wire \sel0_b6/or_or_B4_B5_o_or_B6__o ;
  wire \sel0_b6/or_or_B9_B10_o_or_B1_o ;
  wire \sel0_b6/or_or_or_B0_B1_o_or__o ;
  wire \sel0_b6/or_or_or_B18_B19_o_o_o ;
  wire \sel0_b6/or_or_or_B27_B28_o_o_o ;
  wire \sel0_b6/or_or_or_B9_B10_o_or_o ;
  wire \sel0_b6/or_or_or_or_B0_B1_o__o ;
  wire \sel0_b6/or_or_or_or_B18_B19__o ;
  wire \sel0_b7/or_B0_B1_o ;
  wire \sel0_b7/or_B11_B12_o ;
  wire \sel0_b7/or_B13_B14_o ;
  wire \sel0_b7/or_B15_or_B16_B17_o_o ;
  wire \sel0_b7/or_B16_B17_o ;
  wire \sel0_b7/or_B18_B19_o ;
  wire \sel0_b7/or_B20_B21_o ;
  wire \sel0_b7/or_B22_B23_o ;
  wire \sel0_b7/or_B24_or_B25_B26_o_o ;
  wire \sel0_b7/or_B25_B26_o ;
  wire \sel0_b7/or_B27_B28_o ;
  wire \sel0_b7/or_B29_or_B30_B31_o_o ;
  wire \sel0_b7/or_B2_B3_o ;
  wire \sel0_b7/or_B30_B31_o ;
  wire \sel0_b7/or_B32_B33_o ;
  wire \sel0_b7/or_B34_or_B35_B36_o_o ;
  wire \sel0_b7/or_B35_B36_o ;
  wire \sel0_b7/or_B4_B5_o ;
  wire \sel0_b7/or_B6_or_B7_B8_o_o ;
  wire \sel0_b7/or_B7_B8_o ;
  wire \sel0_b7/or_B9_B10_o ;
  wire \sel0_b7/or_or_B0_B1_o_or_B2__o ;
  wire \sel0_b7/or_or_B13_B14_o_or_B_o ;
  wire \sel0_b7/or_or_B18_B19_o_or_B_o ;
  wire \sel0_b7/or_or_B22_B23_o_or_B_o ;
  wire \sel0_b7/or_or_B27_B28_o_or_B_o ;
  wire \sel0_b7/or_or_B32_B33_o_or_B_o ;
  wire \sel0_b7/or_or_B4_B5_o_or_B6__o ;
  wire \sel0_b7/or_or_B9_B10_o_or_B1_o ;
  wire \sel0_b7/or_or_or_B0_B1_o_or__o ;
  wire \sel0_b7/or_or_or_B18_B19_o_o_o ;
  wire \sel0_b7/or_or_or_B27_B28_o_o_o ;
  wire \sel0_b7/or_or_or_B9_B10_o_or_o ;
  wire \sel0_b7/or_or_or_or_B0_B1_o__o ;
  wire \sel0_b7/or_or_or_or_B18_B19__o ;
  wire \sel1/or_B0_B1_o ;
  wire \sel1/or_B11_B12_o ;
  wire \sel1/or_B13_B14_o ;
  wire \sel1/or_B15_or_B16_B17_o_o ;
  wire \sel1/or_B16_B17_o ;
  wire \sel1/or_B18_B19_o ;
  wire \sel1/or_B20_B21_o ;
  wire \sel1/or_B22_B23_o ;
  wire \sel1/or_B24_or_B25_B26_o_o ;
  wire \sel1/or_B25_B26_o ;
  wire \sel1/or_B27_B28_o ;
  wire \sel1/or_B29_B30_o ;
  wire \sel1/or_B2_B3_o ;
  wire \sel1/or_B31_B32_o ;
  wire \sel1/or_B33_or_B34_B35_o_o ;
  wire \sel1/or_B34_B35_o ;
  wire \sel1/or_B4_B5_o ;
  wire \sel1/or_B6_or_B7_B8_o_o ;
  wire \sel1/or_B7_B8_o ;
  wire \sel1/or_B9_B10_o ;
  wire \sel1/or_or_B0_B1_o_or_B2__o ;
  wire \sel1/or_or_B13_B14_o_or_B_o ;
  wire \sel1/or_or_B18_B19_o_or_B_o ;
  wire \sel1/or_or_B22_B23_o_or_B_o ;
  wire \sel1/or_or_B27_B28_o_or_B_o ;
  wire \sel1/or_or_B31_B32_o_or_B_o ;
  wire \sel1/or_or_B4_B5_o_or_B6__o ;
  wire \sel1/or_or_B9_B10_o_or_B1_o ;
  wire \sel1/or_or_or_B0_B1_o_or__o ;
  wire \sel1/or_or_or_B18_B19_o_o_o ;
  wire \sel1/or_or_or_B27_B28_o_o_o ;
  wire \sel1/or_or_or_B9_B10_o_or_o ;
  wire \sel1/or_or_or_or_B0_B1_o__o ;
  wire \sel1/or_or_or_or_B18_B19__o ;
  wire \sel2/or_B0_B1_o ;
  wire \sel2/or_B11_B12_o ;
  wire \sel2/or_B13_B14_o ;
  wire \sel2/or_B15_or_B16_B17_o_o ;
  wire \sel2/or_B16_B17_o ;
  wire \sel2/or_B18_B19_o ;
  wire \sel2/or_B20_B21_o ;
  wire \sel2/or_B22_B23_o ;
  wire \sel2/or_B24_or_B25_B26_o_o ;
  wire \sel2/or_B25_B26_o ;
  wire \sel2/or_B27_B28_o ;
  wire \sel2/or_B29_B30_o ;
  wire \sel2/or_B2_B3_o ;
  wire \sel2/or_B31_B32_o ;
  wire \sel2/or_B33_or_B34_B35_o_o ;
  wire \sel2/or_B34_B35_o ;
  wire \sel2/or_B4_B5_o ;
  wire \sel2/or_B6_or_B7_B8_o_o ;
  wire \sel2/or_B7_B8_o ;
  wire \sel2/or_B9_B10_o ;
  wire \sel2/or_or_B0_B1_o_or_B2__o ;
  wire \sel2/or_or_B13_B14_o_or_B_o ;
  wire \sel2/or_or_B18_B19_o_or_B_o ;
  wire \sel2/or_or_B22_B23_o_or_B_o ;
  wire \sel2/or_or_B27_B28_o_or_B_o ;
  wire \sel2/or_or_B31_B32_o_or_B_o ;
  wire \sel2/or_or_B4_B5_o_or_B6__o ;
  wire \sel2/or_or_B9_B10_o_or_B1_o ;
  wire \sel2/or_or_or_B0_B1_o_or__o ;
  wire \sel2/or_or_or_B18_B19_o_o_o ;
  wire \sel2/or_or_or_B27_B28_o_o_o ;
  wire \sel2/or_or_or_B9_B10_o_or_o ;
  wire \sel2/or_or_or_or_B0_B1_o__o ;
  wire \sel2/or_or_or_or_B18_B19__o ;
  wire \sel3/or_B0_B1_o ;
  wire \sel3/or_B11_B12_o ;
  wire \sel3/or_B13_B14_o ;
  wire \sel3/or_B15_or_B16_B17_o_o ;
  wire \sel3/or_B16_B17_o ;
  wire \sel3/or_B18_B19_o ;
  wire \sel3/or_B20_B21_o ;
  wire \sel3/or_B22_B23_o ;
  wire \sel3/or_B24_or_B25_B26_o_o ;
  wire \sel3/or_B25_B26_o ;
  wire \sel3/or_B27_B28_o ;
  wire \sel3/or_B29_B30_o ;
  wire \sel3/or_B2_B3_o ;
  wire \sel3/or_B31_B32_o ;
  wire \sel3/or_B33_or_B34_B35_o_o ;
  wire \sel3/or_B4_B5_o ;
  wire \sel3/or_B6_or_B7_B8_o_o ;
  wire \sel3/or_B7_B8_o ;
  wire \sel3/or_B9_B10_o ;
  wire \sel3/or_or_B0_B1_o_or_B2__o ;
  wire \sel3/or_or_B13_B14_o_or_B_o ;
  wire \sel3/or_or_B18_B19_o_or_B_o ;
  wire \sel3/or_or_B22_B23_o_or_B_o ;
  wire \sel3/or_or_B27_B28_o_or_B_o ;
  wire \sel3/or_or_B31_B32_o_or_B_o ;
  wire \sel3/or_or_B4_B5_o_or_B6__o ;
  wire \sel3/or_or_B9_B10_o_or_B1_o ;
  wire \sel3/or_or_or_B0_B1_o_or__o ;
  wire \sel3/or_or_or_B18_B19_o_o_o ;
  wire \sel3/or_or_or_B27_B28_o_o_o ;
  wire \sel3/or_or_or_B9_B10_o_or_o ;
  wire \sel3/or_or_or_or_B0_B1_o__o ;
  wire \sel3/or_or_or_or_B18_B19__o ;
  wire \sel4/or_B0_B1_o ;
  wire \sel4/or_B11_B12_o ;
  wire \sel4/or_B13_B14_o ;
  wire \sel4/or_B15_or_B16_B17_o_o ;
  wire \sel4/or_B16_B17_o ;
  wire \sel4/or_B18_B19_o ;
  wire \sel4/or_B20_B21_o ;
  wire \sel4/or_B22_B23_o ;
  wire \sel4/or_B24_or_B25_B26_o_o ;
  wire \sel4/or_B25_B26_o ;
  wire \sel4/or_B27_B28_o ;
  wire \sel4/or_B29_B30_o ;
  wire \sel4/or_B2_B3_o ;
  wire \sel4/or_B31_B32_o ;
  wire \sel4/or_B33_or_B34_B35_o_o ;
  wire \sel4/or_B34_B35_o ;
  wire \sel4/or_B4_B5_o ;
  wire \sel4/or_B6_or_B7_B8_o_o ;
  wire \sel4/or_B7_B8_o ;
  wire \sel4/or_B9_B10_o ;
  wire \sel4/or_or_B0_B1_o_or_B2__o ;
  wire \sel4/or_or_B13_B14_o_or_B_o ;
  wire \sel4/or_or_B18_B19_o_or_B_o ;
  wire \sel4/or_or_B22_B23_o_or_B_o ;
  wire \sel4/or_or_B27_B28_o_or_B_o ;
  wire \sel4/or_or_B31_B32_o_or_B_o ;
  wire \sel4/or_or_B4_B5_o_or_B6__o ;
  wire \sel4/or_or_B9_B10_o_or_B1_o ;
  wire \sel4/or_or_or_B0_B1_o_or__o ;
  wire \sel4/or_or_or_B18_B19_o_o_o ;
  wire \sel4/or_or_or_B27_B28_o_o_o ;
  wire \sel4/or_or_or_B9_B10_o_or_o ;
  wire \sel4/or_or_or_or_B0_B1_o__o ;
  wire \sel4/or_or_or_or_B18_B19__o ;
  wire \sel5/or_B0_B1_o ;
  wire \sel5/or_B11_B12_o ;
  wire \sel5/or_B13_B14_o ;
  wire \sel5/or_B15_or_B16_B17_o_o ;
  wire \sel5/or_B16_B17_o ;
  wire \sel5/or_B18_B19_o ;
  wire \sel5/or_B20_B21_o ;
  wire \sel5/or_B22_B23_o ;
  wire \sel5/or_B24_or_B25_B26_o_o ;
  wire \sel5/or_B25_B26_o ;
  wire \sel5/or_B27_B28_o ;
  wire \sel5/or_B29_B30_o ;
  wire \sel5/or_B2_B3_o ;
  wire \sel5/or_B31_B32_o ;
  wire \sel5/or_B33_or_B34_B35_o_o ;
  wire \sel5/or_B4_B5_o ;
  wire \sel5/or_B6_or_B7_B8_o_o ;
  wire \sel5/or_B7_B8_o ;
  wire \sel5/or_B9_B10_o ;
  wire \sel5/or_or_B0_B1_o_or_B2__o ;
  wire \sel5/or_or_B13_B14_o_or_B_o ;
  wire \sel5/or_or_B18_B19_o_or_B_o ;
  wire \sel5/or_or_B22_B23_o_or_B_o ;
  wire \sel5/or_or_B27_B28_o_or_B_o ;
  wire \sel5/or_or_B31_B32_o_or_B_o ;
  wire \sel5/or_or_B4_B5_o_or_B6__o ;
  wire \sel5/or_or_B9_B10_o_or_B1_o ;
  wire \sel5/or_or_or_B0_B1_o_or__o ;
  wire \sel5/or_or_or_B18_B19_o_o_o ;
  wire \sel5/or_or_or_B27_B28_o_o_o ;
  wire \sel5/or_or_or_B9_B10_o_or_o ;
  wire \sel5/or_or_or_or_B0_B1_o__o ;
  wire \sel5/or_or_or_or_B18_B19__o ;
  wire \sel6/or_B0_B1_o ;
  wire \sel6/or_B11_B12_o ;
  wire \sel6/or_B13_B14_o ;
  wire \sel6/or_B15_or_B16_B17_o_o ;
  wire \sel6/or_B16_B17_o ;
  wire \sel6/or_B18_B19_o ;
  wire \sel6/or_B20_B21_o ;
  wire \sel6/or_B22_B23_o ;
  wire \sel6/or_B24_or_B25_B26_o_o ;
  wire \sel6/or_B25_B26_o ;
  wire \sel6/or_B27_B28_o ;
  wire \sel6/or_B29_B30_o ;
  wire \sel6/or_B2_B3_o ;
  wire \sel6/or_B31_B32_o ;
  wire \sel6/or_B33_or_B34_B35_o_o ;
  wire \sel6/or_B4_B5_o ;
  wire \sel6/or_B6_or_B7_B8_o_o ;
  wire \sel6/or_B7_B8_o ;
  wire \sel6/or_B9_B10_o ;
  wire \sel6/or_or_B0_B1_o_or_B2__o ;
  wire \sel6/or_or_B13_B14_o_or_B_o ;
  wire \sel6/or_or_B18_B19_o_or_B_o ;
  wire \sel6/or_or_B22_B23_o_or_B_o ;
  wire \sel6/or_or_B27_B28_o_or_B_o ;
  wire \sel6/or_or_B31_B32_o_or_B_o ;
  wire \sel6/or_or_B4_B5_o_or_B6__o ;
  wire \sel6/or_or_B9_B10_o_or_B1_o ;
  wire \sel6/or_or_or_B0_B1_o_or__o ;
  wire \sel6/or_or_or_B18_B19_o_o_o ;
  wire \sel6/or_or_or_B27_B28_o_o_o ;
  wire \sel6/or_or_or_B9_B10_o_or_o ;
  wire \sel6/or_or_or_or_B0_B1_o__o ;
  wire \sel6/or_or_or_or_B18_B19__o ;
  wire success;  // sources/rtl/i2c_module.v(141)

  reg_ar_as_w1 ack_ok_reg (
    .clk(divider2[7]),
    .d(n29),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(ack_ok));  // sources/rtl/i2c_module.v(153)
  add_pu8_pu8_o8 add0 (
    .i0(divider2),
    .i1(8'b00000001),
    .o(n1));  // sources/rtl/i2c_module.v(80)
  not \address[0]_inv  (\address[0]_neg , address[0]);
  not \address[1]_inv  (\address[1]_neg , address[1]);
  reg_ar_as_w1 clk_div_reg (
    .clk(divider2[7]),
    .d(n0),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(clk_div));  // sources/rtl/i2c_module.v(76)
  eq_w1 eq0 (
    .i0(reset_n),
    .i1(1'b0),
    .o(n2));  // sources/rtl/i2c_module.v(93)
  eq_w1 eq1 (
    .i0(scl_output_enable),
    .i1(1'b1),
    .o(n17));  // sources/rtl/i2c_module.v(125)
  eq_w8 eq10 (
    .i0(state_next),
    .i1(8'b00000000),
    .o(n146));  // sources/rtl/i2c_module.v(179)
  eq_w8 eq11 (
    .i0(state_next),
    .i1(8'b01101111),
    .o(n148));  // sources/rtl/i2c_module.v(195)
  eq_w8 eq12 (
    .i0(state_next),
    .i1(8'b01110000),
    .o(n149));  // sources/rtl/i2c_module.v(203)
  eq_w8 eq13 (
    .i0(state_next),
    .i1(8'b00000010),
    .o(n150));  // sources/rtl/i2c_module.v(211)
  eq_w8 eq14 (
    .i0(state_next),
    .i1(8'b00000011),
    .o(n151));  // sources/rtl/i2c_module.v(219)
  eq_w8 eq15 (
    .i0(state_next),
    .i1(8'b00000100),
    .o(n152));  // sources/rtl/i2c_module.v(227)
  eq_w8 eq16 (
    .i0(state_next),
    .i1(8'b00000101),
    .o(n153));  // sources/rtl/i2c_module.v(235)
  eq_w8 eq17 (
    .i0(state_next),
    .i1(8'b00000110),
    .o(n154));  // sources/rtl/i2c_module.v(243)
  eq_w8 eq18 (
    .i0(state_next),
    .i1(8'b00000111),
    .o(n155));  // sources/rtl/i2c_module.v(251)
  eq_w8 eq19 (
    .i0(state_next),
    .i1(8'b00001000),
    .o(n156));  // sources/rtl/i2c_module.v(259)
  eq_w1 eq2 (
    .i0(scl_output_zero),
    .i1(1'b0),
    .o(n19));  // sources/rtl/i2c_module.v(131)
  eq_w8 eq20 (
    .i0(state_next),
    .i1(8'b00001001),
    .o(n157));  // sources/rtl/i2c_module.v(267)
  eq_w8 eq21 (
    .i0(state_next),
    .i1(8'b01100110),
    .o(n159));  // sources/rtl/i2c_module.v(290)
  eq_w8 eq22 (
    .i0(state_next),
    .i1(8'b00001011),
    .o(n160));  // sources/rtl/i2c_module.v(306)
  eq_w8 eq23 (
    .i0(state_next),
    .i1(8'b00001100),
    .o(n161));  // sources/rtl/i2c_module.v(314)
  eq_w8 eq24 (
    .i0(state_next),
    .i1(8'b00001101),
    .o(n162));  // sources/rtl/i2c_module.v(322)
  eq_w8 eq25 (
    .i0(state_next),
    .i1(8'b00001110),
    .o(n163));  // sources/rtl/i2c_module.v(330)
  eq_w8 eq26 (
    .i0(state_next),
    .i1(8'b00001111),
    .o(n164));  // sources/rtl/i2c_module.v(338)
  eq_w8 eq27 (
    .i0(state_next),
    .i1(8'b00010000),
    .o(n165));  // sources/rtl/i2c_module.v(346)
  eq_w8 eq28 (
    .i0(state_next),
    .i1(8'b00010001),
    .o(n166));  // sources/rtl/i2c_module.v(354)
  eq_w8 eq29 (
    .i0(state_next),
    .i1(8'b00010010),
    .o(n167));  // sources/rtl/i2c_module.v(362)
  eq_w8 eq3 (
    .i0(state_next),
    .i1(8'b00001010),
    .o(n158));  // sources/rtl/i2c_module.v(147)
  eq_w8 eq30 (
    .i0(state_next),
    .i1(8'b11000000),
    .o(n169));  // sources/rtl/i2c_module.v(393)
  eq_w8 eq31 (
    .i0(state_next),
    .i1(8'b00010100),
    .o(n170));  // sources/rtl/i2c_module.v(402)
  eq_w8 eq32 (
    .i0(state_next),
    .i1(8'b00010101),
    .o(n171));  // sources/rtl/i2c_module.v(410)
  eq_w8 eq33 (
    .i0(state_next),
    .i1(8'b00010110),
    .o(n172));  // sources/rtl/i2c_module.v(418)
  eq_w8 eq34 (
    .i0(state_next),
    .i1(8'b00010111),
    .o(n173));  // sources/rtl/i2c_module.v(426)
  eq_w8 eq35 (
    .i0(state_next),
    .i1(8'b00011000),
    .o(n174));  // sources/rtl/i2c_module.v(434)
  eq_w8 eq36 (
    .i0(state_next),
    .i1(8'b00011001),
    .o(n175));  // sources/rtl/i2c_module.v(442)
  eq_w8 eq37 (
    .i0(state_next),
    .i1(8'b00011010),
    .o(n176));  // sources/rtl/i2c_module.v(450)
  eq_w8 eq38 (
    .i0(state_next),
    .i1(8'b00011011),
    .o(n177));  // sources/rtl/i2c_module.v(458)
  eq_w8 eq39 (
    .i0(state_next),
    .i1(8'b00011110),
    .o(n180));  // sources/rtl/i2c_module.v(492)
  eq_w8 eq4 (
    .i0(state_next),
    .i1(8'b00010011),
    .o(n168));  // sources/rtl/i2c_module.v(147)
  eq_w8 eq40 (
    .i0(state_next),
    .i1(8'b00011111),
    .o(n181));  // sources/rtl/i2c_module.v(500)
  eq_w8 eq5 (
    .i0(state_next),
    .i1(8'b00011100),
    .o(n178));  // sources/rtl/i2c_module.v(147)
  eq_w1 eq6 (
    .i0(clk_div),
    .i1(1'b1),
    .o(n28));  // sources/rtl/i2c_module.v(147)
  eq_w8 eq7 (
    .i0(state_next),
    .i1(8'b00011101),
    .o(n179));  // sources/rtl/i2c_module.v(160)
  eq_w8 eq8 (
    .i0(state_next),
    .i1(8'b00000001),
    .o(n147));  // sources/rtl/i2c_module.v(163)
  eq_w1 eq9 (
    .i0(clk_div),
    .i1(1'b0),
    .o(n36));  // sources/rtl/i2c_module.v(189)
  and mux0_b0_sel_is_3 (mux0_b0_sel_is_3_o, address[0], address[1]);
  binary_mux_s1_w1 mux13_b0 (
    .i0(state_next[0]),
    .i1(1'b1),
    .sel(control_reg[0]),
    .o(n35[0]));  // sources/rtl/i2c_module.v(184)
  binary_mux_s1_w1 mux13_b1 (
    .i0(state_next[1]),
    .i1(1'b0),
    .sel(control_reg[0]),
    .o(n35[1]));  // sources/rtl/i2c_module.v(184)
  binary_mux_s1_w1 mux13_b2 (
    .i0(state_next[2]),
    .i1(1'b0),
    .sel(control_reg[0]),
    .o(n35[2]));  // sources/rtl/i2c_module.v(184)
  binary_mux_s1_w1 mux13_b3 (
    .i0(state_next[3]),
    .i1(1'b0),
    .sel(control_reg[0]),
    .o(n35[3]));  // sources/rtl/i2c_module.v(184)
  binary_mux_s1_w1 mux13_b4 (
    .i0(state_next[4]),
    .i1(1'b0),
    .sel(control_reg[0]),
    .o(n35[4]));  // sources/rtl/i2c_module.v(184)
  binary_mux_s1_w1 mux13_b5 (
    .i0(state_next[5]),
    .i1(1'b0),
    .sel(control_reg[0]),
    .o(n35[5]));  // sources/rtl/i2c_module.v(184)
  binary_mux_s1_w1 mux13_b6 (
    .i0(state_next[6]),
    .i1(1'b0),
    .sel(control_reg[0]),
    .o(n35[6]));  // sources/rtl/i2c_module.v(184)
  binary_mux_s1_w1 mux13_b7 (
    .i0(state_next[7]),
    .i1(1'b0),
    .sel(control_reg[0]),
    .o(n35[7]));  // sources/rtl/i2c_module.v(184)
  binary_mux_s1_w1 mux14_b0 (
    .i0(state_next[0]),
    .i1(1'b0),
    .sel(n28),
    .o(n72[0]));  // sources/rtl/i2c_module.v(200)
  binary_mux_s1_w1 mux14_b1 (
    .i0(state_next[1]),
    .i1(1'b0),
    .sel(n28),
    .o(n72[1]));  // sources/rtl/i2c_module.v(200)
  binary_mux_s1_w1 mux14_b10 (
    .i0(state_next[2]),
    .i1(1'b1),
    .sel(n28),
    .o(n70[2]));  // sources/rtl/i2c_module.v(200)
  binary_mux_s1_w1 mux14_b11 (
    .i0(state_next[3]),
    .i1(1'b1),
    .sel(n28),
    .o(n70[3]));  // sources/rtl/i2c_module.v(200)
  binary_mux_s1_w1 mux14_b12 (
    .i0(state_next[4]),
    .i1(1'b1),
    .sel(n28),
    .o(n70[4]));  // sources/rtl/i2c_module.v(200)
  binary_mux_s1_w1 mux14_b13 (
    .i0(state_next[5]),
    .i1(1'b0),
    .sel(n28),
    .o(n70[5]));  // sources/rtl/i2c_module.v(200)
  binary_mux_s1_w1 mux14_b14 (
    .i0(state_next[6]),
    .i1(1'b0),
    .sel(n28),
    .o(n70[6]));  // sources/rtl/i2c_module.v(200)
  binary_mux_s1_w1 mux14_b15 (
    .i0(state_next[7]),
    .i1(1'b0),
    .sel(n28),
    .o(n70[7]));  // sources/rtl/i2c_module.v(200)
  binary_mux_s1_w1 mux14_b18 (
    .i0(state_next[2]),
    .i1(1'b0),
    .sel(n28),
    .o(n38[2]));  // sources/rtl/i2c_module.v(200)
  binary_mux_s1_w1 mux14_b19 (
    .i0(state_next[3]),
    .i1(1'b0),
    .sel(n28),
    .o(n38[3]));  // sources/rtl/i2c_module.v(200)
  binary_mux_s1_w1 mux14_b21 (
    .i0(state_next[5]),
    .i1(1'b1),
    .sel(n28),
    .o(n38[5]));  // sources/rtl/i2c_module.v(200)
  binary_mux_s1_w1 mux14_b22 (
    .i0(state_next[6]),
    .i1(1'b1),
    .sel(n28),
    .o(n38[6]));  // sources/rtl/i2c_module.v(200)
  binary_mux_s1_w1 mux14_b4 (
    .i0(state_next[4]),
    .i1(1'b0),
    .sel(n28),
    .o(n72[4]));  // sources/rtl/i2c_module.v(200)
  binary_mux_s1_w1 mux14_b9 (
    .i0(state_next[1]),
    .i1(1'b1),
    .sel(n28),
    .o(n70[1]));  // sources/rtl/i2c_module.v(200)
  binary_mux_s1_w1 mux15_b0 (
    .i0(state_next[0]),
    .i1(1'b0),
    .sel(n36),
    .o(n71[0]));  // sources/rtl/i2c_module.v(192)
  binary_mux_s1_w1 mux15_b1 (
    .i0(state_next[1]),
    .i1(1'b0),
    .sel(n36),
    .o(n71[1]));  // sources/rtl/i2c_module.v(192)
  binary_mux_s1_w1 mux15_b10 (
    .i0(state_next[2]),
    .i1(1'b1),
    .sel(n36),
    .o(n69[2]));  // sources/rtl/i2c_module.v(192)
  binary_mux_s1_w1 mux15_b100 (
    .i0(state_next[4]),
    .i1(1'b1),
    .sel(n36),
    .o(n57[4]));  // sources/rtl/i2c_module.v(192)
  binary_mux_s1_w1 mux15_b101 (
    .i0(state_next[5]),
    .i1(1'b0),
    .sel(n36),
    .o(n57[5]));  // sources/rtl/i2c_module.v(192)
  binary_mux_s1_w1 mux15_b102 (
    .i0(state_next[6]),
    .i1(1'b0),
    .sel(n36),
    .o(n57[6]));  // sources/rtl/i2c_module.v(192)
  binary_mux_s1_w1 mux15_b103 (
    .i0(state_next[7]),
    .i1(1'b0),
    .sel(n36),
    .o(n57[7]));  // sources/rtl/i2c_module.v(192)
  binary_mux_s1_w1 mux15_b105 (
    .i0(state_next[1]),
    .i1(1'b1),
    .sel(n36),
    .o(n56[1]));  // sources/rtl/i2c_module.v(192)
  binary_mux_s1_w1 mux15_b106 (
    .i0(state_next[2]),
    .i1(1'b0),
    .sel(n36),
    .o(n56[2]));  // sources/rtl/i2c_module.v(192)
  binary_mux_s1_w1 mux15_b107 (
    .i0(state_next[3]),
    .i1(1'b0),
    .sel(n36),
    .o(n56[3]));  // sources/rtl/i2c_module.v(192)
  binary_mux_s1_w1 mux15_b11 (
    .i0(state_next[3]),
    .i1(1'b1),
    .sel(n36),
    .o(n69[3]));  // sources/rtl/i2c_module.v(192)
  binary_mux_s1_w1 mux15_b112 (
    .i0(state_next[0]),
    .i1(1'b1),
    .sel(n36),
    .o(n55[0]));  // sources/rtl/i2c_module.v(192)
  binary_mux_s1_w1 mux15_b132 (
    .i0(state_next[4]),
    .i1(1'b0),
    .sel(n36),
    .o(n53[4]));  // sources/rtl/i2c_module.v(192)
  binary_mux_s1_w1 mux15_b168 (
    .i0(state_next[0]),
    .i1(n58[0]),
    .sel(n36),
    .o(n48[0]));  // sources/rtl/i2c_module.v(192)
  binary_mux_s1_w1 mux15_b169 (
    .i0(state_next[1]),
    .i1(ack_ok),
    .sel(n36),
    .o(n48[1]));  // sources/rtl/i2c_module.v(192)
  binary_mux_s1_w1 mux15_b171 (
    .i0(state_next[3]),
    .i1(n58[0]),
    .sel(n36),
    .o(n48[3]));  // sources/rtl/i2c_module.v(192)
  binary_mux_s1_w1 mux15_b172 (
    .i0(state_next[4]),
    .i1(n58[0]),
    .sel(n36),
    .o(n48[4]));  // sources/rtl/i2c_module.v(192)
  binary_mux_s1_w1 mux15_b173 (
    .i0(state_next[5]),
    .i1(ack_ok),
    .sel(n36),
    .o(n48[5]));  // sources/rtl/i2c_module.v(192)
  binary_mux_s1_w1 mux15_b174 (
    .i0(state_next[6]),
    .i1(ack_ok),
    .sel(n36),
    .o(n48[6]));  // sources/rtl/i2c_module.v(192)
  binary_mux_s1_w1 mux15_b253 (
    .i0(state_next[5]),
    .i1(1'b1),
    .sel(n36),
    .o(n37[5]));  // sources/rtl/i2c_module.v(192)
  binary_mux_s1_w1 mux15_b254 (
    .i0(state_next[6]),
    .i1(1'b1),
    .sel(n36),
    .o(n37[6]));  // sources/rtl/i2c_module.v(192)
  binary_mux_s1_w1 mux15_b90 (
    .i0(state_next[2]),
    .i1(n58[0]),
    .sel(n36),
    .o(n59[2]));  // sources/rtl/i2c_module.v(192)
  binary_mux_s1_w1 mux15_b95 (
    .i0(state_next[7]),
    .i1(ack_ok),
    .sel(n36),
    .o(n59[7]));  // sources/rtl/i2c_module.v(192)
  and mux1_b0_sel_is_2 (mux1_b0_sel_is_2_o, \address[0]_neg , address[1]);
  and mux2_b0_sel_is_1 (mux2_b0_sel_is_1_o, address[0], \address[1]_neg );
  and mux3_b0_sel_is_0 (mux3_b0_sel_is_0_o, \address[0]_neg , \address[1]_neg );
  and mux4_b0_sel_is_3 (mux4_b0_sel_is_3_o, write, mux0_b0_sel_is_3_o);
  and mux5_b0_sel_is_3 (mux5_b0_sel_is_3_o, write, mux1_b0_sel_is_2_o);
  and mux6_b0_sel_is_3 (mux6_b0_sel_is_3_o, write, mux2_b0_sel_is_1_o);
  and mux7_b0_sel_is_3 (mux7_b0_sel_is_3_o, write, mux3_b0_sel_is_0_o);
  and mux9_b0_sel_is_0 (mux9_b0_sel_is_0_o, n2_neg, n11_neg);
  not n11_inv (n11_neg, n11);
  not n2_inv (n2_neg, n2);
  ne_w8 neq0 (
    .i0(state_next),
    .i1(8'b00000000),
    .o(n11));  // sources/rtl/i2c_module.v(114)
  reg_ar_ss_w1 ready_reg (
    .clk(~divider2[7]),
    .d(n190),
    .en(1'b1),
    .reset(1'b0),
    .set(~reset_n),
    .q(ready));  // sources/rtl/i2c_module.v(1066)
  reg_ar_as_w1 reg0_b0 (
    .clk(clk),
    .d(n1[0]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(divider2[0]));  // sources/rtl/i2c_module.v(81)
  reg_ar_as_w1 reg0_b1 (
    .clk(clk),
    .d(n1[1]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(divider2[1]));  // sources/rtl/i2c_module.v(81)
  reg_ar_as_w1 reg0_b2 (
    .clk(clk),
    .d(n1[2]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(divider2[2]));  // sources/rtl/i2c_module.v(81)
  reg_ar_as_w1 reg0_b3 (
    .clk(clk),
    .d(n1[3]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(divider2[3]));  // sources/rtl/i2c_module.v(81)
  reg_ar_as_w1 reg0_b4 (
    .clk(clk),
    .d(n1[4]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(divider2[4]));  // sources/rtl/i2c_module.v(81)
  reg_ar_as_w1 reg0_b5 (
    .clk(clk),
    .d(n1[5]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(divider2[5]));  // sources/rtl/i2c_module.v(81)
  reg_ar_as_w1 reg0_b6 (
    .clk(clk),
    .d(n1[6]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(divider2[6]));  // sources/rtl/i2c_module.v(81)
  reg_ar_as_w1 reg0_b7 (
    .clk(clk),
    .d(n1[7]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(divider2[7]));  // sources/rtl/i2c_module.v(81)
  reg_sr_as_w1 reg1_b0 (
    .clk(clk),
    .d(writedata[0]),
    .en(mux7_b0_sel_is_3_o),
    .reset(~mux9_b0_sel_is_0_o),
    .set(1'b0),
    .q(control_reg[0]));  // sources/rtl/i2c_module.v(117)
  reg_sr_as_w1 reg2_b0 (
    .clk(clk),
    .d(writedata[0]),
    .en(mux6_b0_sel_is_3_o),
    .reset(n2),
    .set(1'b0),
    .q(slave_address[0]));  // sources/rtl/i2c_module.v(117)
  reg_sr_as_w1 reg2_b1 (
    .clk(clk),
    .d(writedata[1]),
    .en(mux6_b0_sel_is_3_o),
    .reset(n2),
    .set(1'b0),
    .q(slave_address[1]));  // sources/rtl/i2c_module.v(117)
  reg_sr_as_w1 reg2_b2 (
    .clk(clk),
    .d(writedata[2]),
    .en(mux6_b0_sel_is_3_o),
    .reset(n2),
    .set(1'b0),
    .q(slave_address[2]));  // sources/rtl/i2c_module.v(117)
  reg_sr_as_w1 reg2_b3 (
    .clk(clk),
    .d(writedata[3]),
    .en(mux6_b0_sel_is_3_o),
    .reset(n2),
    .set(1'b0),
    .q(slave_address[3]));  // sources/rtl/i2c_module.v(117)
  reg_sr_as_w1 reg2_b4 (
    .clk(clk),
    .d(writedata[4]),
    .en(mux6_b0_sel_is_3_o),
    .reset(n2),
    .set(1'b0),
    .q(slave_address[4]));  // sources/rtl/i2c_module.v(117)
  reg_sr_as_w1 reg2_b5 (
    .clk(clk),
    .d(writedata[5]),
    .en(mux6_b0_sel_is_3_o),
    .reset(n2),
    .set(1'b0),
    .q(slave_address[5]));  // sources/rtl/i2c_module.v(117)
  reg_sr_as_w1 reg2_b6 (
    .clk(clk),
    .d(writedata[6]),
    .en(mux6_b0_sel_is_3_o),
    .reset(n2),
    .set(1'b0),
    .q(slave_address[6]));  // sources/rtl/i2c_module.v(117)
  reg_sr_as_w1 reg2_b7 (
    .clk(clk),
    .d(writedata[7]),
    .en(mux6_b0_sel_is_3_o),
    .reset(n2),
    .set(1'b0),
    .q(slave_address[7]));  // sources/rtl/i2c_module.v(117)
  reg_sr_as_w1 reg3_b0 (
    .clk(clk),
    .d(writedata[0]),
    .en(mux5_b0_sel_is_3_o),
    .reset(n2),
    .set(1'b0),
    .q(slave_reg_address[0]));  // sources/rtl/i2c_module.v(117)
  reg_sr_as_w1 reg3_b1 (
    .clk(clk),
    .d(writedata[1]),
    .en(mux5_b0_sel_is_3_o),
    .reset(n2),
    .set(1'b0),
    .q(slave_reg_address[1]));  // sources/rtl/i2c_module.v(117)
  reg_sr_as_w1 reg3_b2 (
    .clk(clk),
    .d(writedata[2]),
    .en(mux5_b0_sel_is_3_o),
    .reset(n2),
    .set(1'b0),
    .q(slave_reg_address[2]));  // sources/rtl/i2c_module.v(117)
  reg_sr_as_w1 reg3_b3 (
    .clk(clk),
    .d(writedata[3]),
    .en(mux5_b0_sel_is_3_o),
    .reset(n2),
    .set(1'b0),
    .q(slave_reg_address[3]));  // sources/rtl/i2c_module.v(117)
  reg_sr_as_w1 reg3_b4 (
    .clk(clk),
    .d(writedata[4]),
    .en(mux5_b0_sel_is_3_o),
    .reset(n2),
    .set(1'b0),
    .q(slave_reg_address[4]));  // sources/rtl/i2c_module.v(117)
  reg_sr_as_w1 reg3_b5 (
    .clk(clk),
    .d(writedata[5]),
    .en(mux5_b0_sel_is_3_o),
    .reset(n2),
    .set(1'b0),
    .q(slave_reg_address[5]));  // sources/rtl/i2c_module.v(117)
  reg_sr_as_w1 reg3_b6 (
    .clk(clk),
    .d(writedata[6]),
    .en(mux5_b0_sel_is_3_o),
    .reset(n2),
    .set(1'b0),
    .q(slave_reg_address[6]));  // sources/rtl/i2c_module.v(117)
  reg_sr_as_w1 reg3_b7 (
    .clk(clk),
    .d(writedata[7]),
    .en(mux5_b0_sel_is_3_o),
    .reset(n2),
    .set(1'b0),
    .q(slave_reg_address[7]));  // sources/rtl/i2c_module.v(117)
  reg_sr_as_w1 reg4_b0 (
    .clk(clk),
    .d(writedata[0]),
    .en(mux4_b0_sel_is_3_o),
    .reset(n2),
    .set(1'b0),
    .q(slave_data_1[0]));  // sources/rtl/i2c_module.v(117)
  reg_sr_as_w1 reg4_b1 (
    .clk(clk),
    .d(writedata[1]),
    .en(mux4_b0_sel_is_3_o),
    .reset(n2),
    .set(1'b0),
    .q(slave_data_1[1]));  // sources/rtl/i2c_module.v(117)
  reg_sr_as_w1 reg4_b2 (
    .clk(clk),
    .d(writedata[2]),
    .en(mux4_b0_sel_is_3_o),
    .reset(n2),
    .set(1'b0),
    .q(slave_data_1[2]));  // sources/rtl/i2c_module.v(117)
  reg_sr_as_w1 reg4_b3 (
    .clk(clk),
    .d(writedata[3]),
    .en(mux4_b0_sel_is_3_o),
    .reset(n2),
    .set(1'b0),
    .q(slave_data_1[3]));  // sources/rtl/i2c_module.v(117)
  reg_sr_as_w1 reg4_b4 (
    .clk(clk),
    .d(writedata[4]),
    .en(mux4_b0_sel_is_3_o),
    .reset(n2),
    .set(1'b0),
    .q(slave_data_1[4]));  // sources/rtl/i2c_module.v(117)
  reg_sr_as_w1 reg4_b5 (
    .clk(clk),
    .d(writedata[5]),
    .en(mux4_b0_sel_is_3_o),
    .reset(n2),
    .set(1'b0),
    .q(slave_data_1[5]));  // sources/rtl/i2c_module.v(117)
  reg_sr_as_w1 reg4_b6 (
    .clk(clk),
    .d(writedata[6]),
    .en(mux4_b0_sel_is_3_o),
    .reset(n2),
    .set(1'b0),
    .q(slave_data_1[6]));  // sources/rtl/i2c_module.v(117)
  reg_sr_as_w1 reg4_b7 (
    .clk(clk),
    .d(writedata[7]),
    .en(mux4_b0_sel_is_3_o),
    .reset(n2),
    .set(1'b0),
    .q(slave_data_1[7]));  // sources/rtl/i2c_module.v(117)
  reg_sr_as_w1 reg5_b0 (
    .clk(~divider2[7]),
    .d(n99[0]),
    .en(1'b1),
    .reset(n2),
    .set(1'b0),
    .q(state_next[0]));  // sources/rtl/i2c_module.v(510)
  reg_sr_as_w1 reg5_b1 (
    .clk(~divider2[7]),
    .d(n99[1]),
    .en(1'b1),
    .reset(n2),
    .set(1'b0),
    .q(state_next[1]));  // sources/rtl/i2c_module.v(510)
  reg_sr_as_w1 reg5_b2 (
    .clk(~divider2[7]),
    .d(n99[2]),
    .en(1'b1),
    .reset(n2),
    .set(1'b0),
    .q(state_next[2]));  // sources/rtl/i2c_module.v(510)
  reg_sr_as_w1 reg5_b3 (
    .clk(~divider2[7]),
    .d(n99[3]),
    .en(1'b1),
    .reset(n2),
    .set(1'b0),
    .q(state_next[3]));  // sources/rtl/i2c_module.v(510)
  reg_sr_as_w1 reg5_b4 (
    .clk(~divider2[7]),
    .d(n99[4]),
    .en(1'b1),
    .reset(n2),
    .set(1'b0),
    .q(state_next[4]));  // sources/rtl/i2c_module.v(510)
  reg_sr_as_w1 reg5_b5 (
    .clk(~divider2[7]),
    .d(n99[5]),
    .en(1'b1),
    .reset(n2),
    .set(1'b0),
    .q(state_next[5]));  // sources/rtl/i2c_module.v(510)
  reg_sr_as_w1 reg5_b6 (
    .clk(~divider2[7]),
    .d(n99[6]),
    .en(1'b1),
    .reset(n2),
    .set(1'b0),
    .q(state_next[6]));  // sources/rtl/i2c_module.v(510)
  reg_sr_as_w1 reg5_b7 (
    .clk(~divider2[7]),
    .d(n99[7]),
    .en(1'b1),
    .reset(n2),
    .set(1'b0),
    .q(state_next[7]));  // sources/rtl/i2c_module.v(510)
  reg_ar_as_w1 scl_out_reg (
    .clk(divider2[7]),
    .d(n20),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(scl_out));  // sources/rtl/i2c_module.v(137)
  reg_sr_as_w1 scl_output_enable_reg (
    .clk(~divider2[7]),
    .d(n188),
    .en(1'b1),
    .reset(~reset_n),
    .set(1'b0),
    .q(scl_output_enable));  // sources/rtl/i2c_module.v(1066)
  reg_ar_as_w1 scl_output_zero_reg (
    .clk(~divider2[7]),
    .d(n194),
    .en(~n102),
    .reset(1'b0),
    .set(1'b0),
    .q(scl_output_zero));  // sources/rtl/i2c_module.v(1066)
  reg_ar_ss_w1 sda_oe_reg (
    .clk(~divider2[7]),
    .d(n186),
    .en(1'b1),
    .reset(1'b0),
    .set(~reset_n),
    .q(sda_oe));  // sources/rtl/i2c_module.v(1066)
  reg_ar_ss_w1 sda_reg (
    .clk(~divider2[7]),
    .d(n184),
    .en(1'b1),
    .reset(1'b0),
    .set(~reset_n),
    .q(sda));  // sources/rtl/i2c_module.v(1066)
  and \sel0_b0/and_b0_0  (\sel0_b0/B0 , state_next[0], n182);
  and \sel0_b0/and_b0_1  (\sel0_b0/B1 , n72[0], n181);
  and \sel0_b0/and_b0_10  (\sel0_b0/B10 , n55[0], n172);
  and \sel0_b0/and_b0_11  (\sel0_b0/B11 , n71[0], n171);
  and \sel0_b0/and_b0_12  (\sel0_b0/B12 , n55[0], n170);
  and \sel0_b0/and_b0_13  (\sel0_b0/B13 , n71[0], n169);
  and \sel0_b0/and_b0_14  (\sel0_b0/B14 , n48[0], n168);
  and \sel0_b0/and_b0_15  (\sel0_b0/B15 , n55[0], n167);
  and \sel0_b0/and_b0_16  (\sel0_b0/B16 , n71[0], n166);
  and \sel0_b0/and_b0_17  (\sel0_b0/B17 , n55[0], n165);
  and \sel0_b0/and_b0_18  (\sel0_b0/B18 , n71[0], n164);
  and \sel0_b0/and_b0_19  (\sel0_b0/B19 , n55[0], n163);
  and \sel0_b0/and_b0_2  (\sel0_b0/B2 , n71[0], n180);
  and \sel0_b0/and_b0_20  (\sel0_b0/B20 , n71[0], n162);
  and \sel0_b0/and_b0_21  (\sel0_b0/B21 , n55[0], n161);
  and \sel0_b0/and_b0_22  (\sel0_b0/B22 , n71[0], n160);
  and \sel0_b0/and_b0_23  (\sel0_b0/B23 , n55[0], n159);
  and \sel0_b0/and_b0_24  (\sel0_b0/B24 , n48[0], n158);
  and \sel0_b0/and_b0_25  (\sel0_b0/B25 , n71[0], n157);
  and \sel0_b0/and_b0_26  (\sel0_b0/B26 , n55[0], n156);
  and \sel0_b0/and_b0_27  (\sel0_b0/B27 , n71[0], n155);
  and \sel0_b0/and_b0_28  (\sel0_b0/B28 , n55[0], n154);
  and \sel0_b0/and_b0_29  (\sel0_b0/B29 , n71[0], n153);
  and \sel0_b0/and_b0_3  (\sel0_b0/B3 , n72[0], n179);
  and \sel0_b0/and_b0_30  (\sel0_b0/B30 , n55[0], n152);
  and \sel0_b0/and_b0_31  (\sel0_b0/B31 , n71[0], n151);
  and \sel0_b0/and_b0_32  (\sel0_b0/B32 , n55[0], n150);
  and \sel0_b0/and_b0_33  (\sel0_b0/B33 , n71[0], n149);
  and \sel0_b0/and_b0_34  (\sel0_b0/B34 , n72[0], n148);
  and \sel0_b0/and_b0_35  (\sel0_b0/B35 , n55[0], n147);
  and \sel0_b0/and_b0_36  (\sel0_b0/B36 , n35[0], n146);
  and \sel0_b0/and_b0_4  (\sel0_b0/B4 , n55[0], n178);
  and \sel0_b0/and_b0_5  (\sel0_b0/B5 , n71[0], n177);
  and \sel0_b0/and_b0_6  (\sel0_b0/B6 , n55[0], n176);
  and \sel0_b0/and_b0_7  (\sel0_b0/B7 , n71[0], n175);
  and \sel0_b0/and_b0_8  (\sel0_b0/B8 , n55[0], n174);
  and \sel0_b0/and_b0_9  (\sel0_b0/B9 , n71[0], n173);
  or \sel0_b0/or_B0_B1  (\sel0_b0/or_B0_B1_o , \sel0_b0/B0 , \sel0_b0/B1 );
  or \sel0_b0/or_B11_B12  (\sel0_b0/or_B11_B12_o , \sel0_b0/B11 , \sel0_b0/B12 );
  or \sel0_b0/or_B13_B14  (\sel0_b0/or_B13_B14_o , \sel0_b0/B13 , \sel0_b0/B14 );
  or \sel0_b0/or_B15_or_B16_B17_o  (\sel0_b0/or_B15_or_B16_B17_o_o , \sel0_b0/B15 , \sel0_b0/or_B16_B17_o );
  or \sel0_b0/or_B16_B17  (\sel0_b0/or_B16_B17_o , \sel0_b0/B16 , \sel0_b0/B17 );
  or \sel0_b0/or_B18_B19  (\sel0_b0/or_B18_B19_o , \sel0_b0/B18 , \sel0_b0/B19 );
  or \sel0_b0/or_B20_B21  (\sel0_b0/or_B20_B21_o , \sel0_b0/B20 , \sel0_b0/B21 );
  or \sel0_b0/or_B22_B23  (\sel0_b0/or_B22_B23_o , \sel0_b0/B22 , \sel0_b0/B23 );
  or \sel0_b0/or_B24_or_B25_B26_o  (\sel0_b0/or_B24_or_B25_B26_o_o , \sel0_b0/B24 , \sel0_b0/or_B25_B26_o );
  or \sel0_b0/or_B25_B26  (\sel0_b0/or_B25_B26_o , \sel0_b0/B25 , \sel0_b0/B26 );
  or \sel0_b0/or_B27_B28  (\sel0_b0/or_B27_B28_o , \sel0_b0/B27 , \sel0_b0/B28 );
  or \sel0_b0/or_B29_or_B30_B31_o  (\sel0_b0/or_B29_or_B30_B31_o_o , \sel0_b0/B29 , \sel0_b0/or_B30_B31_o );
  or \sel0_b0/or_B2_B3  (\sel0_b0/or_B2_B3_o , \sel0_b0/B2 , \sel0_b0/B3 );
  or \sel0_b0/or_B30_B31  (\sel0_b0/or_B30_B31_o , \sel0_b0/B30 , \sel0_b0/B31 );
  or \sel0_b0/or_B32_B33  (\sel0_b0/or_B32_B33_o , \sel0_b0/B32 , \sel0_b0/B33 );
  or \sel0_b0/or_B34_or_B35_B36_o  (\sel0_b0/or_B34_or_B35_B36_o_o , \sel0_b0/B34 , \sel0_b0/or_B35_B36_o );
  or \sel0_b0/or_B35_B36  (\sel0_b0/or_B35_B36_o , \sel0_b0/B35 , \sel0_b0/B36 );
  or \sel0_b0/or_B4_B5  (\sel0_b0/or_B4_B5_o , \sel0_b0/B4 , \sel0_b0/B5 );
  or \sel0_b0/or_B6_or_B7_B8_o  (\sel0_b0/or_B6_or_B7_B8_o_o , \sel0_b0/B6 , \sel0_b0/or_B7_B8_o );
  or \sel0_b0/or_B7_B8  (\sel0_b0/or_B7_B8_o , \sel0_b0/B7 , \sel0_b0/B8 );
  or \sel0_b0/or_B9_B10  (\sel0_b0/or_B9_B10_o , \sel0_b0/B9 , \sel0_b0/B10 );
  or \sel0_b0/or_or_B0_B1_o_or_B2_  (\sel0_b0/or_or_B0_B1_o_or_B2__o , \sel0_b0/or_B0_B1_o , \sel0_b0/or_B2_B3_o );
  or \sel0_b0/or_or_B13_B14_o_or_B  (\sel0_b0/or_or_B13_B14_o_or_B_o , \sel0_b0/or_B13_B14_o , \sel0_b0/or_B15_or_B16_B17_o_o );
  or \sel0_b0/or_or_B18_B19_o_or_B  (\sel0_b0/or_or_B18_B19_o_or_B_o , \sel0_b0/or_B18_B19_o , \sel0_b0/or_B20_B21_o );
  or \sel0_b0/or_or_B22_B23_o_or_B  (\sel0_b0/or_or_B22_B23_o_or_B_o , \sel0_b0/or_B22_B23_o , \sel0_b0/or_B24_or_B25_B26_o_o );
  or \sel0_b0/or_or_B27_B28_o_or_B  (\sel0_b0/or_or_B27_B28_o_or_B_o , \sel0_b0/or_B27_B28_o , \sel0_b0/or_B29_or_B30_B31_o_o );
  or \sel0_b0/or_or_B32_B33_o_or_B  (\sel0_b0/or_or_B32_B33_o_or_B_o , \sel0_b0/or_B32_B33_o , \sel0_b0/or_B34_or_B35_B36_o_o );
  or \sel0_b0/or_or_B4_B5_o_or_B6_  (\sel0_b0/or_or_B4_B5_o_or_B6__o , \sel0_b0/or_B4_B5_o , \sel0_b0/or_B6_or_B7_B8_o_o );
  or \sel0_b0/or_or_B9_B10_o_or_B1  (\sel0_b0/or_or_B9_B10_o_or_B1_o , \sel0_b0/or_B9_B10_o , \sel0_b0/or_B11_B12_o );
  or \sel0_b0/or_or_or_B0_B1_o_or_  (\sel0_b0/or_or_or_B0_B1_o_or__o , \sel0_b0/or_or_B0_B1_o_or_B2__o , \sel0_b0/or_or_B4_B5_o_or_B6__o );
  or \sel0_b0/or_or_or_B18_B19_o_o  (\sel0_b0/or_or_or_B18_B19_o_o_o , \sel0_b0/or_or_B18_B19_o_or_B_o , \sel0_b0/or_or_B22_B23_o_or_B_o );
  or \sel0_b0/or_or_or_B27_B28_o_o  (\sel0_b0/or_or_or_B27_B28_o_o_o , \sel0_b0/or_or_B27_B28_o_or_B_o , \sel0_b0/or_or_B32_B33_o_or_B_o );
  or \sel0_b0/or_or_or_B9_B10_o_or  (\sel0_b0/or_or_or_B9_B10_o_or_o , \sel0_b0/or_or_B9_B10_o_or_B1_o , \sel0_b0/or_or_B13_B14_o_or_B_o );
  or \sel0_b0/or_or_or_or_B0_B1_o_  (\sel0_b0/or_or_or_or_B0_B1_o__o , \sel0_b0/or_or_or_B0_B1_o_or__o , \sel0_b0/or_or_or_B9_B10_o_or_o );
  or \sel0_b0/or_or_or_or_B18_B19_  (\sel0_b0/or_or_or_or_B18_B19__o , \sel0_b0/or_or_or_B18_B19_o_o_o , \sel0_b0/or_or_or_B27_B28_o_o_o );
  or \sel0_b0/or_or_or_or_or_B0_B1  (n99[0], \sel0_b0/or_or_or_or_B0_B1_o__o , \sel0_b0/or_or_or_or_B18_B19__o );
  and \sel0_b1/and_b0_0  (\sel0_b1/B0 , state_next[1], n182);
  and \sel0_b1/and_b0_1  (\sel0_b1/B1 , n72[1], n181);
  and \sel0_b1/and_b0_10  (\sel0_b1/B10 , n56[1], n172);
  and \sel0_b1/and_b0_11  (\sel0_b1/B11 , n56[1], n171);
  and \sel0_b1/and_b0_12  (\sel0_b1/B12 , n71[1], n170);
  and \sel0_b1/and_b0_13  (\sel0_b1/B13 , n71[1], n169);
  and \sel0_b1/and_b0_14  (\sel0_b1/B14 , n71[1], n168);
  and \sel0_b1/and_b0_15  (\sel0_b1/B15 , n56[1], n167);
  and \sel0_b1/and_b0_16  (\sel0_b1/B16 , n56[1], n166);
  and \sel0_b1/and_b0_17  (\sel0_b1/B17 , n71[1], n165);
  and \sel0_b1/and_b0_18  (\sel0_b1/B18 , n71[1], n164);
  and \sel0_b1/and_b0_19  (\sel0_b1/B19 , n56[1], n163);
  and \sel0_b1/and_b0_2  (\sel0_b1/B2 , n71[1], n180);
  and \sel0_b1/and_b0_20  (\sel0_b1/B20 , n56[1], n162);
  and \sel0_b1/and_b0_21  (\sel0_b1/B21 , n71[1], n161);
  and \sel0_b1/and_b0_22  (\sel0_b1/B22 , n71[1], n160);
  and \sel0_b1/and_b0_23  (\sel0_b1/B23 , n56[1], n159);
  and \sel0_b1/and_b0_24  (\sel0_b1/B24 , n48[1], n158);
  and \sel0_b1/and_b0_25  (\sel0_b1/B25 , n56[1], n157);
  and \sel0_b1/and_b0_26  (\sel0_b1/B26 , n71[1], n156);
  and \sel0_b1/and_b0_27  (\sel0_b1/B27 , n71[1], n155);
  and \sel0_b1/and_b0_28  (\sel0_b1/B28 , n56[1], n154);
  and \sel0_b1/and_b0_29  (\sel0_b1/B29 , n56[1], n153);
  and \sel0_b1/and_b0_3  (\sel0_b1/B3 , n70[1], n179);
  and \sel0_b1/and_b0_30  (\sel0_b1/B30 , n71[1], n152);
  and \sel0_b1/and_b0_31  (\sel0_b1/B31 , n71[1], n151);
  and \sel0_b1/and_b0_32  (\sel0_b1/B32 , n56[1], n150);
  and \sel0_b1/and_b0_33  (\sel0_b1/B33 , n56[1], n149);
  and \sel0_b1/and_b0_34  (\sel0_b1/B34 , n72[1], n148);
  and \sel0_b1/and_b0_35  (\sel0_b1/B35 , n56[1], n147);
  and \sel0_b1/and_b0_36  (\sel0_b1/B36 , n35[1], n146);
  and \sel0_b1/and_b0_4  (\sel0_b1/B4 , n71[1], n178);
  and \sel0_b1/and_b0_5  (\sel0_b1/B5 , n71[1], n177);
  and \sel0_b1/and_b0_6  (\sel0_b1/B6 , n56[1], n176);
  and \sel0_b1/and_b0_7  (\sel0_b1/B7 , n56[1], n175);
  and \sel0_b1/and_b0_8  (\sel0_b1/B8 , n71[1], n174);
  and \sel0_b1/and_b0_9  (\sel0_b1/B9 , n71[1], n173);
  or \sel0_b1/or_B0_B1  (\sel0_b1/or_B0_B1_o , \sel0_b1/B0 , \sel0_b1/B1 );
  or \sel0_b1/or_B11_B12  (\sel0_b1/or_B11_B12_o , \sel0_b1/B11 , \sel0_b1/B12 );
  or \sel0_b1/or_B13_B14  (\sel0_b1/or_B13_B14_o , \sel0_b1/B13 , \sel0_b1/B14 );
  or \sel0_b1/or_B15_or_B16_B17_o  (\sel0_b1/or_B15_or_B16_B17_o_o , \sel0_b1/B15 , \sel0_b1/or_B16_B17_o );
  or \sel0_b1/or_B16_B17  (\sel0_b1/or_B16_B17_o , \sel0_b1/B16 , \sel0_b1/B17 );
  or \sel0_b1/or_B18_B19  (\sel0_b1/or_B18_B19_o , \sel0_b1/B18 , \sel0_b1/B19 );
  or \sel0_b1/or_B20_B21  (\sel0_b1/or_B20_B21_o , \sel0_b1/B20 , \sel0_b1/B21 );
  or \sel0_b1/or_B22_B23  (\sel0_b1/or_B22_B23_o , \sel0_b1/B22 , \sel0_b1/B23 );
  or \sel0_b1/or_B24_or_B25_B26_o  (\sel0_b1/or_B24_or_B25_B26_o_o , \sel0_b1/B24 , \sel0_b1/or_B25_B26_o );
  or \sel0_b1/or_B25_B26  (\sel0_b1/or_B25_B26_o , \sel0_b1/B25 , \sel0_b1/B26 );
  or \sel0_b1/or_B27_B28  (\sel0_b1/or_B27_B28_o , \sel0_b1/B27 , \sel0_b1/B28 );
  or \sel0_b1/or_B29_or_B30_B31_o  (\sel0_b1/or_B29_or_B30_B31_o_o , \sel0_b1/B29 , \sel0_b1/or_B30_B31_o );
  or \sel0_b1/or_B2_B3  (\sel0_b1/or_B2_B3_o , \sel0_b1/B2 , \sel0_b1/B3 );
  or \sel0_b1/or_B30_B31  (\sel0_b1/or_B30_B31_o , \sel0_b1/B30 , \sel0_b1/B31 );
  or \sel0_b1/or_B32_B33  (\sel0_b1/or_B32_B33_o , \sel0_b1/B32 , \sel0_b1/B33 );
  or \sel0_b1/or_B34_or_B35_B36_o  (\sel0_b1/or_B34_or_B35_B36_o_o , \sel0_b1/B34 , \sel0_b1/or_B35_B36_o );
  or \sel0_b1/or_B35_B36  (\sel0_b1/or_B35_B36_o , \sel0_b1/B35 , \sel0_b1/B36 );
  or \sel0_b1/or_B4_B5  (\sel0_b1/or_B4_B5_o , \sel0_b1/B4 , \sel0_b1/B5 );
  or \sel0_b1/or_B6_or_B7_B8_o  (\sel0_b1/or_B6_or_B7_B8_o_o , \sel0_b1/B6 , \sel0_b1/or_B7_B8_o );
  or \sel0_b1/or_B7_B8  (\sel0_b1/or_B7_B8_o , \sel0_b1/B7 , \sel0_b1/B8 );
  or \sel0_b1/or_B9_B10  (\sel0_b1/or_B9_B10_o , \sel0_b1/B9 , \sel0_b1/B10 );
  or \sel0_b1/or_or_B0_B1_o_or_B2_  (\sel0_b1/or_or_B0_B1_o_or_B2__o , \sel0_b1/or_B0_B1_o , \sel0_b1/or_B2_B3_o );
  or \sel0_b1/or_or_B13_B14_o_or_B  (\sel0_b1/or_or_B13_B14_o_or_B_o , \sel0_b1/or_B13_B14_o , \sel0_b1/or_B15_or_B16_B17_o_o );
  or \sel0_b1/or_or_B18_B19_o_or_B  (\sel0_b1/or_or_B18_B19_o_or_B_o , \sel0_b1/or_B18_B19_o , \sel0_b1/or_B20_B21_o );
  or \sel0_b1/or_or_B22_B23_o_or_B  (\sel0_b1/or_or_B22_B23_o_or_B_o , \sel0_b1/or_B22_B23_o , \sel0_b1/or_B24_or_B25_B26_o_o );
  or \sel0_b1/or_or_B27_B28_o_or_B  (\sel0_b1/or_or_B27_B28_o_or_B_o , \sel0_b1/or_B27_B28_o , \sel0_b1/or_B29_or_B30_B31_o_o );
  or \sel0_b1/or_or_B32_B33_o_or_B  (\sel0_b1/or_or_B32_B33_o_or_B_o , \sel0_b1/or_B32_B33_o , \sel0_b1/or_B34_or_B35_B36_o_o );
  or \sel0_b1/or_or_B4_B5_o_or_B6_  (\sel0_b1/or_or_B4_B5_o_or_B6__o , \sel0_b1/or_B4_B5_o , \sel0_b1/or_B6_or_B7_B8_o_o );
  or \sel0_b1/or_or_B9_B10_o_or_B1  (\sel0_b1/or_or_B9_B10_o_or_B1_o , \sel0_b1/or_B9_B10_o , \sel0_b1/or_B11_B12_o );
  or \sel0_b1/or_or_or_B0_B1_o_or_  (\sel0_b1/or_or_or_B0_B1_o_or__o , \sel0_b1/or_or_B0_B1_o_or_B2__o , \sel0_b1/or_or_B4_B5_o_or_B6__o );
  or \sel0_b1/or_or_or_B18_B19_o_o  (\sel0_b1/or_or_or_B18_B19_o_o_o , \sel0_b1/or_or_B18_B19_o_or_B_o , \sel0_b1/or_or_B22_B23_o_or_B_o );
  or \sel0_b1/or_or_or_B27_B28_o_o  (\sel0_b1/or_or_or_B27_B28_o_o_o , \sel0_b1/or_or_B27_B28_o_or_B_o , \sel0_b1/or_or_B32_B33_o_or_B_o );
  or \sel0_b1/or_or_or_B9_B10_o_or  (\sel0_b1/or_or_or_B9_B10_o_or_o , \sel0_b1/or_or_B9_B10_o_or_B1_o , \sel0_b1/or_or_B13_B14_o_or_B_o );
  or \sel0_b1/or_or_or_or_B0_B1_o_  (\sel0_b1/or_or_or_or_B0_B1_o__o , \sel0_b1/or_or_or_B0_B1_o_or__o , \sel0_b1/or_or_or_B9_B10_o_or_o );
  or \sel0_b1/or_or_or_or_B18_B19_  (\sel0_b1/or_or_or_or_B18_B19__o , \sel0_b1/or_or_or_B18_B19_o_o_o , \sel0_b1/or_or_or_B27_B28_o_o_o );
  or \sel0_b1/or_or_or_or_or_B0_B1  (n99[1], \sel0_b1/or_or_or_or_B0_B1_o__o , \sel0_b1/or_or_or_or_B18_B19__o );
  and \sel0_b2/and_b0_0  (\sel0_b2/B0 , state_next[2], n182);
  and \sel0_b2/and_b0_1  (\sel0_b2/B1 , n38[2], n181);
  and \sel0_b2/and_b0_10  (\sel0_b2/B10 , n69[2], n172);
  and \sel0_b2/and_b0_11  (\sel0_b2/B11 , n69[2], n171);
  and \sel0_b2/and_b0_12  (\sel0_b2/B12 , n69[2], n170);
  and \sel0_b2/and_b0_13  (\sel0_b2/B13 , n69[2], n169);
  and \sel0_b2/and_b0_14  (\sel0_b2/B14 , n59[2], n168);
  and \sel0_b2/and_b0_15  (\sel0_b2/B15 , n56[2], n167);
  and \sel0_b2/and_b0_16  (\sel0_b2/B16 , n56[2], n166);
  and \sel0_b2/and_b0_17  (\sel0_b2/B17 , n56[2], n165);
  and \sel0_b2/and_b0_18  (\sel0_b2/B18 , n56[2], n164);
  and \sel0_b2/and_b0_19  (\sel0_b2/B19 , n69[2], n163);
  and \sel0_b2/and_b0_2  (\sel0_b2/B2 , n56[2], n180);
  and \sel0_b2/and_b0_20  (\sel0_b2/B20 , n69[2], n162);
  and \sel0_b2/and_b0_21  (\sel0_b2/B21 , n69[2], n161);
  and \sel0_b2/and_b0_22  (\sel0_b2/B22 , n69[2], n160);
  and \sel0_b2/and_b0_23  (\sel0_b2/B23 , n56[2], n159);
  and \sel0_b2/and_b0_24  (\sel0_b2/B24 , n69[2], n158);
  and \sel0_b2/and_b0_25  (\sel0_b2/B25 , n56[2], n157);
  and \sel0_b2/and_b0_26  (\sel0_b2/B26 , n56[2], n156);
  and \sel0_b2/and_b0_27  (\sel0_b2/B27 , n56[2], n155);
  and \sel0_b2/and_b0_28  (\sel0_b2/B28 , n69[2], n154);
  and \sel0_b2/and_b0_29  (\sel0_b2/B29 , n69[2], n153);
  and \sel0_b2/and_b0_3  (\sel0_b2/B3 , n70[2], n179);
  and \sel0_b2/and_b0_30  (\sel0_b2/B30 , n69[2], n152);
  and \sel0_b2/and_b0_31  (\sel0_b2/B31 , n69[2], n151);
  and \sel0_b2/and_b0_32  (\sel0_b2/B32 , n56[2], n150);
  and \sel0_b2/and_b0_33  (\sel0_b2/B33 , n56[2], n149);
  and \sel0_b2/and_b0_34  (\sel0_b2/B34 , n38[2], n148);
  and \sel0_b2/and_b0_35  (\sel0_b2/B35 , n69[2], n147);
  and \sel0_b2/and_b0_36  (\sel0_b2/B36 , n35[2], n146);
  and \sel0_b2/and_b0_4  (\sel0_b2/B4 , n69[2], n178);
  and \sel0_b2/and_b0_5  (\sel0_b2/B5 , n69[2], n177);
  and \sel0_b2/and_b0_6  (\sel0_b2/B6 , n56[2], n176);
  and \sel0_b2/and_b0_7  (\sel0_b2/B7 , n56[2], n175);
  and \sel0_b2/and_b0_8  (\sel0_b2/B8 , n56[2], n174);
  and \sel0_b2/and_b0_9  (\sel0_b2/B9 , n56[2], n173);
  or \sel0_b2/or_B0_B1  (\sel0_b2/or_B0_B1_o , \sel0_b2/B0 , \sel0_b2/B1 );
  or \sel0_b2/or_B11_B12  (\sel0_b2/or_B11_B12_o , \sel0_b2/B11 , \sel0_b2/B12 );
  or \sel0_b2/or_B13_B14  (\sel0_b2/or_B13_B14_o , \sel0_b2/B13 , \sel0_b2/B14 );
  or \sel0_b2/or_B15_or_B16_B17_o  (\sel0_b2/or_B15_or_B16_B17_o_o , \sel0_b2/B15 , \sel0_b2/or_B16_B17_o );
  or \sel0_b2/or_B16_B17  (\sel0_b2/or_B16_B17_o , \sel0_b2/B16 , \sel0_b2/B17 );
  or \sel0_b2/or_B18_B19  (\sel0_b2/or_B18_B19_o , \sel0_b2/B18 , \sel0_b2/B19 );
  or \sel0_b2/or_B20_B21  (\sel0_b2/or_B20_B21_o , \sel0_b2/B20 , \sel0_b2/B21 );
  or \sel0_b2/or_B22_B23  (\sel0_b2/or_B22_B23_o , \sel0_b2/B22 , \sel0_b2/B23 );
  or \sel0_b2/or_B24_or_B25_B26_o  (\sel0_b2/or_B24_or_B25_B26_o_o , \sel0_b2/B24 , \sel0_b2/or_B25_B26_o );
  or \sel0_b2/or_B25_B26  (\sel0_b2/or_B25_B26_o , \sel0_b2/B25 , \sel0_b2/B26 );
  or \sel0_b2/or_B27_B28  (\sel0_b2/or_B27_B28_o , \sel0_b2/B27 , \sel0_b2/B28 );
  or \sel0_b2/or_B29_or_B30_B31_o  (\sel0_b2/or_B29_or_B30_B31_o_o , \sel0_b2/B29 , \sel0_b2/or_B30_B31_o );
  or \sel0_b2/or_B2_B3  (\sel0_b2/or_B2_B3_o , \sel0_b2/B2 , \sel0_b2/B3 );
  or \sel0_b2/or_B30_B31  (\sel0_b2/or_B30_B31_o , \sel0_b2/B30 , \sel0_b2/B31 );
  or \sel0_b2/or_B32_B33  (\sel0_b2/or_B32_B33_o , \sel0_b2/B32 , \sel0_b2/B33 );
  or \sel0_b2/or_B34_or_B35_B36_o  (\sel0_b2/or_B34_or_B35_B36_o_o , \sel0_b2/B34 , \sel0_b2/or_B35_B36_o );
  or \sel0_b2/or_B35_B36  (\sel0_b2/or_B35_B36_o , \sel0_b2/B35 , \sel0_b2/B36 );
  or \sel0_b2/or_B4_B5  (\sel0_b2/or_B4_B5_o , \sel0_b2/B4 , \sel0_b2/B5 );
  or \sel0_b2/or_B6_or_B7_B8_o  (\sel0_b2/or_B6_or_B7_B8_o_o , \sel0_b2/B6 , \sel0_b2/or_B7_B8_o );
  or \sel0_b2/or_B7_B8  (\sel0_b2/or_B7_B8_o , \sel0_b2/B7 , \sel0_b2/B8 );
  or \sel0_b2/or_B9_B10  (\sel0_b2/or_B9_B10_o , \sel0_b2/B9 , \sel0_b2/B10 );
  or \sel0_b2/or_or_B0_B1_o_or_B2_  (\sel0_b2/or_or_B0_B1_o_or_B2__o , \sel0_b2/or_B0_B1_o , \sel0_b2/or_B2_B3_o );
  or \sel0_b2/or_or_B13_B14_o_or_B  (\sel0_b2/or_or_B13_B14_o_or_B_o , \sel0_b2/or_B13_B14_o , \sel0_b2/or_B15_or_B16_B17_o_o );
  or \sel0_b2/or_or_B18_B19_o_or_B  (\sel0_b2/or_or_B18_B19_o_or_B_o , \sel0_b2/or_B18_B19_o , \sel0_b2/or_B20_B21_o );
  or \sel0_b2/or_or_B22_B23_o_or_B  (\sel0_b2/or_or_B22_B23_o_or_B_o , \sel0_b2/or_B22_B23_o , \sel0_b2/or_B24_or_B25_B26_o_o );
  or \sel0_b2/or_or_B27_B28_o_or_B  (\sel0_b2/or_or_B27_B28_o_or_B_o , \sel0_b2/or_B27_B28_o , \sel0_b2/or_B29_or_B30_B31_o_o );
  or \sel0_b2/or_or_B32_B33_o_or_B  (\sel0_b2/or_or_B32_B33_o_or_B_o , \sel0_b2/or_B32_B33_o , \sel0_b2/or_B34_or_B35_B36_o_o );
  or \sel0_b2/or_or_B4_B5_o_or_B6_  (\sel0_b2/or_or_B4_B5_o_or_B6__o , \sel0_b2/or_B4_B5_o , \sel0_b2/or_B6_or_B7_B8_o_o );
  or \sel0_b2/or_or_B9_B10_o_or_B1  (\sel0_b2/or_or_B9_B10_o_or_B1_o , \sel0_b2/or_B9_B10_o , \sel0_b2/or_B11_B12_o );
  or \sel0_b2/or_or_or_B0_B1_o_or_  (\sel0_b2/or_or_or_B0_B1_o_or__o , \sel0_b2/or_or_B0_B1_o_or_B2__o , \sel0_b2/or_or_B4_B5_o_or_B6__o );
  or \sel0_b2/or_or_or_B18_B19_o_o  (\sel0_b2/or_or_or_B18_B19_o_o_o , \sel0_b2/or_or_B18_B19_o_or_B_o , \sel0_b2/or_or_B22_B23_o_or_B_o );
  or \sel0_b2/or_or_or_B27_B28_o_o  (\sel0_b2/or_or_or_B27_B28_o_o_o , \sel0_b2/or_or_B27_B28_o_or_B_o , \sel0_b2/or_or_B32_B33_o_or_B_o );
  or \sel0_b2/or_or_or_B9_B10_o_or  (\sel0_b2/or_or_or_B9_B10_o_or_o , \sel0_b2/or_or_B9_B10_o_or_B1_o , \sel0_b2/or_or_B13_B14_o_or_B_o );
  or \sel0_b2/or_or_or_or_B0_B1_o_  (\sel0_b2/or_or_or_or_B0_B1_o__o , \sel0_b2/or_or_or_B0_B1_o_or__o , \sel0_b2/or_or_or_B9_B10_o_or_o );
  or \sel0_b2/or_or_or_or_B18_B19_  (\sel0_b2/or_or_or_or_B18_B19__o , \sel0_b2/or_or_or_B18_B19_o_o_o , \sel0_b2/or_or_or_B27_B28_o_o_o );
  or \sel0_b2/or_or_or_or_or_B0_B1  (n99[2], \sel0_b2/or_or_or_or_B0_B1_o__o , \sel0_b2/or_or_or_or_B18_B19__o );
  and \sel0_b3/and_b0_0  (\sel0_b3/B0 , state_next[3], n182);
  and \sel0_b3/and_b0_1  (\sel0_b3/B1 , n38[3], n181);
  and \sel0_b3/and_b0_10  (\sel0_b3/B10 , n56[3], n172);
  and \sel0_b3/and_b0_11  (\sel0_b3/B11 , n56[3], n171);
  and \sel0_b3/and_b0_12  (\sel0_b3/B12 , n56[3], n170);
  and \sel0_b3/and_b0_13  (\sel0_b3/B13 , n56[3], n169);
  and \sel0_b3/and_b0_14  (\sel0_b3/B14 , n48[3], n168);
  and \sel0_b3/and_b0_15  (\sel0_b3/B15 , n56[3], n167);
  and \sel0_b3/and_b0_16  (\sel0_b3/B16 , n56[3], n166);
  and \sel0_b3/and_b0_17  (\sel0_b3/B17 , n56[3], n165);
  and \sel0_b3/and_b0_18  (\sel0_b3/B18 , n56[3], n164);
  and \sel0_b3/and_b0_19  (\sel0_b3/B19 , n69[3], n163);
  and \sel0_b3/and_b0_2  (\sel0_b3/B2 , n56[3], n180);
  and \sel0_b3/and_b0_20  (\sel0_b3/B20 , n69[3], n162);
  and \sel0_b3/and_b0_21  (\sel0_b3/B21 , n69[3], n161);
  and \sel0_b3/and_b0_22  (\sel0_b3/B22 , n69[3], n160);
  and \sel0_b3/and_b0_23  (\sel0_b3/B23 , n69[3], n159);
  and \sel0_b3/and_b0_24  (\sel0_b3/B24 , n48[3], n158);
  and \sel0_b3/and_b0_25  (\sel0_b3/B25 , n69[3], n157);
  and \sel0_b3/and_b0_26  (\sel0_b3/B26 , n69[3], n156);
  and \sel0_b3/and_b0_27  (\sel0_b3/B27 , n69[3], n155);
  and \sel0_b3/and_b0_28  (\sel0_b3/B28 , n56[3], n154);
  and \sel0_b3/and_b0_29  (\sel0_b3/B29 , n56[3], n153);
  and \sel0_b3/and_b0_3  (\sel0_b3/B3 , n70[3], n179);
  and \sel0_b3/and_b0_30  (\sel0_b3/B30 , n56[3], n152);
  and \sel0_b3/and_b0_31  (\sel0_b3/B31 , n56[3], n151);
  and \sel0_b3/and_b0_32  (\sel0_b3/B32 , n56[3], n150);
  and \sel0_b3/and_b0_33  (\sel0_b3/B33 , n56[3], n149);
  and \sel0_b3/and_b0_34  (\sel0_b3/B34 , n38[3], n148);
  and \sel0_b3/and_b0_35  (\sel0_b3/B35 , n69[3], n147);
  and \sel0_b3/and_b0_36  (\sel0_b3/B36 , n35[3], n146);
  and \sel0_b3/and_b0_4  (\sel0_b3/B4 , n69[3], n178);
  and \sel0_b3/and_b0_5  (\sel0_b3/B5 , n69[3], n177);
  and \sel0_b3/and_b0_6  (\sel0_b3/B6 , n69[3], n176);
  and \sel0_b3/and_b0_7  (\sel0_b3/B7 , n69[3], n175);
  and \sel0_b3/and_b0_8  (\sel0_b3/B8 , n69[3], n174);
  and \sel0_b3/and_b0_9  (\sel0_b3/B9 , n69[3], n173);
  or \sel0_b3/or_B0_B1  (\sel0_b3/or_B0_B1_o , \sel0_b3/B0 , \sel0_b3/B1 );
  or \sel0_b3/or_B11_B12  (\sel0_b3/or_B11_B12_o , \sel0_b3/B11 , \sel0_b3/B12 );
  or \sel0_b3/or_B13_B14  (\sel0_b3/or_B13_B14_o , \sel0_b3/B13 , \sel0_b3/B14 );
  or \sel0_b3/or_B15_or_B16_B17_o  (\sel0_b3/or_B15_or_B16_B17_o_o , \sel0_b3/B15 , \sel0_b3/or_B16_B17_o );
  or \sel0_b3/or_B16_B17  (\sel0_b3/or_B16_B17_o , \sel0_b3/B16 , \sel0_b3/B17 );
  or \sel0_b3/or_B18_B19  (\sel0_b3/or_B18_B19_o , \sel0_b3/B18 , \sel0_b3/B19 );
  or \sel0_b3/or_B20_B21  (\sel0_b3/or_B20_B21_o , \sel0_b3/B20 , \sel0_b3/B21 );
  or \sel0_b3/or_B22_B23  (\sel0_b3/or_B22_B23_o , \sel0_b3/B22 , \sel0_b3/B23 );
  or \sel0_b3/or_B24_or_B25_B26_o  (\sel0_b3/or_B24_or_B25_B26_o_o , \sel0_b3/B24 , \sel0_b3/or_B25_B26_o );
  or \sel0_b3/or_B25_B26  (\sel0_b3/or_B25_B26_o , \sel0_b3/B25 , \sel0_b3/B26 );
  or \sel0_b3/or_B27_B28  (\sel0_b3/or_B27_B28_o , \sel0_b3/B27 , \sel0_b3/B28 );
  or \sel0_b3/or_B29_or_B30_B31_o  (\sel0_b3/or_B29_or_B30_B31_o_o , \sel0_b3/B29 , \sel0_b3/or_B30_B31_o );
  or \sel0_b3/or_B2_B3  (\sel0_b3/or_B2_B3_o , \sel0_b3/B2 , \sel0_b3/B3 );
  or \sel0_b3/or_B30_B31  (\sel0_b3/or_B30_B31_o , \sel0_b3/B30 , \sel0_b3/B31 );
  or \sel0_b3/or_B32_B33  (\sel0_b3/or_B32_B33_o , \sel0_b3/B32 , \sel0_b3/B33 );
  or \sel0_b3/or_B34_or_B35_B36_o  (\sel0_b3/or_B34_or_B35_B36_o_o , \sel0_b3/B34 , \sel0_b3/or_B35_B36_o );
  or \sel0_b3/or_B35_B36  (\sel0_b3/or_B35_B36_o , \sel0_b3/B35 , \sel0_b3/B36 );
  or \sel0_b3/or_B4_B5  (\sel0_b3/or_B4_B5_o , \sel0_b3/B4 , \sel0_b3/B5 );
  or \sel0_b3/or_B6_or_B7_B8_o  (\sel0_b3/or_B6_or_B7_B8_o_o , \sel0_b3/B6 , \sel0_b3/or_B7_B8_o );
  or \sel0_b3/or_B7_B8  (\sel0_b3/or_B7_B8_o , \sel0_b3/B7 , \sel0_b3/B8 );
  or \sel0_b3/or_B9_B10  (\sel0_b3/or_B9_B10_o , \sel0_b3/B9 , \sel0_b3/B10 );
  or \sel0_b3/or_or_B0_B1_o_or_B2_  (\sel0_b3/or_or_B0_B1_o_or_B2__o , \sel0_b3/or_B0_B1_o , \sel0_b3/or_B2_B3_o );
  or \sel0_b3/or_or_B13_B14_o_or_B  (\sel0_b3/or_or_B13_B14_o_or_B_o , \sel0_b3/or_B13_B14_o , \sel0_b3/or_B15_or_B16_B17_o_o );
  or \sel0_b3/or_or_B18_B19_o_or_B  (\sel0_b3/or_or_B18_B19_o_or_B_o , \sel0_b3/or_B18_B19_o , \sel0_b3/or_B20_B21_o );
  or \sel0_b3/or_or_B22_B23_o_or_B  (\sel0_b3/or_or_B22_B23_o_or_B_o , \sel0_b3/or_B22_B23_o , \sel0_b3/or_B24_or_B25_B26_o_o );
  or \sel0_b3/or_or_B27_B28_o_or_B  (\sel0_b3/or_or_B27_B28_o_or_B_o , \sel0_b3/or_B27_B28_o , \sel0_b3/or_B29_or_B30_B31_o_o );
  or \sel0_b3/or_or_B32_B33_o_or_B  (\sel0_b3/or_or_B32_B33_o_or_B_o , \sel0_b3/or_B32_B33_o , \sel0_b3/or_B34_or_B35_B36_o_o );
  or \sel0_b3/or_or_B4_B5_o_or_B6_  (\sel0_b3/or_or_B4_B5_o_or_B6__o , \sel0_b3/or_B4_B5_o , \sel0_b3/or_B6_or_B7_B8_o_o );
  or \sel0_b3/or_or_B9_B10_o_or_B1  (\sel0_b3/or_or_B9_B10_o_or_B1_o , \sel0_b3/or_B9_B10_o , \sel0_b3/or_B11_B12_o );
  or \sel0_b3/or_or_or_B0_B1_o_or_  (\sel0_b3/or_or_or_B0_B1_o_or__o , \sel0_b3/or_or_B0_B1_o_or_B2__o , \sel0_b3/or_or_B4_B5_o_or_B6__o );
  or \sel0_b3/or_or_or_B18_B19_o_o  (\sel0_b3/or_or_or_B18_B19_o_o_o , \sel0_b3/or_or_B18_B19_o_or_B_o , \sel0_b3/or_or_B22_B23_o_or_B_o );
  or \sel0_b3/or_or_or_B27_B28_o_o  (\sel0_b3/or_or_or_B27_B28_o_o_o , \sel0_b3/or_or_B27_B28_o_or_B_o , \sel0_b3/or_or_B32_B33_o_or_B_o );
  or \sel0_b3/or_or_or_B9_B10_o_or  (\sel0_b3/or_or_or_B9_B10_o_or_o , \sel0_b3/or_or_B9_B10_o_or_B1_o , \sel0_b3/or_or_B13_B14_o_or_B_o );
  or \sel0_b3/or_or_or_or_B0_B1_o_  (\sel0_b3/or_or_or_or_B0_B1_o__o , \sel0_b3/or_or_or_B0_B1_o_or__o , \sel0_b3/or_or_or_B9_B10_o_or_o );
  or \sel0_b3/or_or_or_or_B18_B19_  (\sel0_b3/or_or_or_or_B18_B19__o , \sel0_b3/or_or_or_B18_B19_o_o_o , \sel0_b3/or_or_or_B27_B28_o_o_o );
  or \sel0_b3/or_or_or_or_or_B0_B1  (n99[3], \sel0_b3/or_or_or_or_B0_B1_o__o , \sel0_b3/or_or_or_or_B18_B19__o );
  and \sel0_b4/and_b0_0  (\sel0_b4/B0 , state_next[4], n182);
  and \sel0_b4/and_b0_1  (\sel0_b4/B1 , n72[4], n181);
  and \sel0_b4/and_b0_10  (\sel0_b4/B10 , n57[4], n172);
  and \sel0_b4/and_b0_11  (\sel0_b4/B11 , n57[4], n171);
  and \sel0_b4/and_b0_12  (\sel0_b4/B12 , n57[4], n170);
  and \sel0_b4/and_b0_13  (\sel0_b4/B13 , n57[4], n169);
  and \sel0_b4/and_b0_14  (\sel0_b4/B14 , n48[4], n168);
  and \sel0_b4/and_b0_15  (\sel0_b4/B15 , n57[4], n167);
  and \sel0_b4/and_b0_16  (\sel0_b4/B16 , n57[4], n166);
  and \sel0_b4/and_b0_17  (\sel0_b4/B17 , n57[4], n165);
  and \sel0_b4/and_b0_18  (\sel0_b4/B18 , n57[4], n164);
  and \sel0_b4/and_b0_19  (\sel0_b4/B19 , n53[4], n163);
  and \sel0_b4/and_b0_2  (\sel0_b4/B2 , n53[4], n180);
  and \sel0_b4/and_b0_20  (\sel0_b4/B20 , n53[4], n162);
  and \sel0_b4/and_b0_21  (\sel0_b4/B21 , n53[4], n161);
  and \sel0_b4/and_b0_22  (\sel0_b4/B22 , n53[4], n160);
  and \sel0_b4/and_b0_23  (\sel0_b4/B23 , n53[4], n159);
  and \sel0_b4/and_b0_24  (\sel0_b4/B24 , n48[4], n158);
  and \sel0_b4/and_b0_25  (\sel0_b4/B25 , n53[4], n157);
  and \sel0_b4/and_b0_26  (\sel0_b4/B26 , n53[4], n156);
  and \sel0_b4/and_b0_27  (\sel0_b4/B27 , n53[4], n155);
  and \sel0_b4/and_b0_28  (\sel0_b4/B28 , n53[4], n154);
  and \sel0_b4/and_b0_29  (\sel0_b4/B29 , n53[4], n153);
  and \sel0_b4/and_b0_3  (\sel0_b4/B3 , n70[4], n179);
  and \sel0_b4/and_b0_30  (\sel0_b4/B30 , n53[4], n152);
  and \sel0_b4/and_b0_31  (\sel0_b4/B31 , n53[4], n151);
  and \sel0_b4/and_b0_32  (\sel0_b4/B32 , n53[4], n150);
  and \sel0_b4/and_b0_33  (\sel0_b4/B33 , n53[4], n149);
  and \sel0_b4/and_b0_34  (\sel0_b4/B34 , n70[4], n148);
  and \sel0_b4/and_b0_35  (\sel0_b4/B35 , n53[4], n147);
  and \sel0_b4/and_b0_36  (\sel0_b4/B36 , n35[4], n146);
  and \sel0_b4/and_b0_4  (\sel0_b4/B4 , n57[4], n178);
  and \sel0_b4/and_b0_5  (\sel0_b4/B5 , n57[4], n177);
  and \sel0_b4/and_b0_6  (\sel0_b4/B6 , n57[4], n176);
  and \sel0_b4/and_b0_7  (\sel0_b4/B7 , n57[4], n175);
  and \sel0_b4/and_b0_8  (\sel0_b4/B8 , n57[4], n174);
  and \sel0_b4/and_b0_9  (\sel0_b4/B9 , n57[4], n173);
  or \sel0_b4/or_B0_B1  (\sel0_b4/or_B0_B1_o , \sel0_b4/B0 , \sel0_b4/B1 );
  or \sel0_b4/or_B11_B12  (\sel0_b4/or_B11_B12_o , \sel0_b4/B11 , \sel0_b4/B12 );
  or \sel0_b4/or_B13_B14  (\sel0_b4/or_B13_B14_o , \sel0_b4/B13 , \sel0_b4/B14 );
  or \sel0_b4/or_B15_or_B16_B17_o  (\sel0_b4/or_B15_or_B16_B17_o_o , \sel0_b4/B15 , \sel0_b4/or_B16_B17_o );
  or \sel0_b4/or_B16_B17  (\sel0_b4/or_B16_B17_o , \sel0_b4/B16 , \sel0_b4/B17 );
  or \sel0_b4/or_B18_B19  (\sel0_b4/or_B18_B19_o , \sel0_b4/B18 , \sel0_b4/B19 );
  or \sel0_b4/or_B20_B21  (\sel0_b4/or_B20_B21_o , \sel0_b4/B20 , \sel0_b4/B21 );
  or \sel0_b4/or_B22_B23  (\sel0_b4/or_B22_B23_o , \sel0_b4/B22 , \sel0_b4/B23 );
  or \sel0_b4/or_B24_or_B25_B26_o  (\sel0_b4/or_B24_or_B25_B26_o_o , \sel0_b4/B24 , \sel0_b4/or_B25_B26_o );
  or \sel0_b4/or_B25_B26  (\sel0_b4/or_B25_B26_o , \sel0_b4/B25 , \sel0_b4/B26 );
  or \sel0_b4/or_B27_B28  (\sel0_b4/or_B27_B28_o , \sel0_b4/B27 , \sel0_b4/B28 );
  or \sel0_b4/or_B29_or_B30_B31_o  (\sel0_b4/or_B29_or_B30_B31_o_o , \sel0_b4/B29 , \sel0_b4/or_B30_B31_o );
  or \sel0_b4/or_B2_B3  (\sel0_b4/or_B2_B3_o , \sel0_b4/B2 , \sel0_b4/B3 );
  or \sel0_b4/or_B30_B31  (\sel0_b4/or_B30_B31_o , \sel0_b4/B30 , \sel0_b4/B31 );
  or \sel0_b4/or_B32_B33  (\sel0_b4/or_B32_B33_o , \sel0_b4/B32 , \sel0_b4/B33 );
  or \sel0_b4/or_B34_or_B35_B36_o  (\sel0_b4/or_B34_or_B35_B36_o_o , \sel0_b4/B34 , \sel0_b4/or_B35_B36_o );
  or \sel0_b4/or_B35_B36  (\sel0_b4/or_B35_B36_o , \sel0_b4/B35 , \sel0_b4/B36 );
  or \sel0_b4/or_B4_B5  (\sel0_b4/or_B4_B5_o , \sel0_b4/B4 , \sel0_b4/B5 );
  or \sel0_b4/or_B6_or_B7_B8_o  (\sel0_b4/or_B6_or_B7_B8_o_o , \sel0_b4/B6 , \sel0_b4/or_B7_B8_o );
  or \sel0_b4/or_B7_B8  (\sel0_b4/or_B7_B8_o , \sel0_b4/B7 , \sel0_b4/B8 );
  or \sel0_b4/or_B9_B10  (\sel0_b4/or_B9_B10_o , \sel0_b4/B9 , \sel0_b4/B10 );
  or \sel0_b4/or_or_B0_B1_o_or_B2_  (\sel0_b4/or_or_B0_B1_o_or_B2__o , \sel0_b4/or_B0_B1_o , \sel0_b4/or_B2_B3_o );
  or \sel0_b4/or_or_B13_B14_o_or_B  (\sel0_b4/or_or_B13_B14_o_or_B_o , \sel0_b4/or_B13_B14_o , \sel0_b4/or_B15_or_B16_B17_o_o );
  or \sel0_b4/or_or_B18_B19_o_or_B  (\sel0_b4/or_or_B18_B19_o_or_B_o , \sel0_b4/or_B18_B19_o , \sel0_b4/or_B20_B21_o );
  or \sel0_b4/or_or_B22_B23_o_or_B  (\sel0_b4/or_or_B22_B23_o_or_B_o , \sel0_b4/or_B22_B23_o , \sel0_b4/or_B24_or_B25_B26_o_o );
  or \sel0_b4/or_or_B27_B28_o_or_B  (\sel0_b4/or_or_B27_B28_o_or_B_o , \sel0_b4/or_B27_B28_o , \sel0_b4/or_B29_or_B30_B31_o_o );
  or \sel0_b4/or_or_B32_B33_o_or_B  (\sel0_b4/or_or_B32_B33_o_or_B_o , \sel0_b4/or_B32_B33_o , \sel0_b4/or_B34_or_B35_B36_o_o );
  or \sel0_b4/or_or_B4_B5_o_or_B6_  (\sel0_b4/or_or_B4_B5_o_or_B6__o , \sel0_b4/or_B4_B5_o , \sel0_b4/or_B6_or_B7_B8_o_o );
  or \sel0_b4/or_or_B9_B10_o_or_B1  (\sel0_b4/or_or_B9_B10_o_or_B1_o , \sel0_b4/or_B9_B10_o , \sel0_b4/or_B11_B12_o );
  or \sel0_b4/or_or_or_B0_B1_o_or_  (\sel0_b4/or_or_or_B0_B1_o_or__o , \sel0_b4/or_or_B0_B1_o_or_B2__o , \sel0_b4/or_or_B4_B5_o_or_B6__o );
  or \sel0_b4/or_or_or_B18_B19_o_o  (\sel0_b4/or_or_or_B18_B19_o_o_o , \sel0_b4/or_or_B18_B19_o_or_B_o , \sel0_b4/or_or_B22_B23_o_or_B_o );
  or \sel0_b4/or_or_or_B27_B28_o_o  (\sel0_b4/or_or_or_B27_B28_o_o_o , \sel0_b4/or_or_B27_B28_o_or_B_o , \sel0_b4/or_or_B32_B33_o_or_B_o );
  or \sel0_b4/or_or_or_B9_B10_o_or  (\sel0_b4/or_or_or_B9_B10_o_or_o , \sel0_b4/or_or_B9_B10_o_or_B1_o , \sel0_b4/or_or_B13_B14_o_or_B_o );
  or \sel0_b4/or_or_or_or_B0_B1_o_  (\sel0_b4/or_or_or_or_B0_B1_o__o , \sel0_b4/or_or_or_B0_B1_o_or__o , \sel0_b4/or_or_or_B9_B10_o_or_o );
  or \sel0_b4/or_or_or_or_B18_B19_  (\sel0_b4/or_or_or_or_B18_B19__o , \sel0_b4/or_or_or_B18_B19_o_o_o , \sel0_b4/or_or_or_B27_B28_o_o_o );
  or \sel0_b4/or_or_or_or_or_B0_B1  (n99[4], \sel0_b4/or_or_or_or_B0_B1_o__o , \sel0_b4/or_or_or_or_B18_B19__o );
  and \sel0_b5/and_b0_0  (\sel0_b5/B0 , state_next[5], n182);
  and \sel0_b5/and_b0_1  (\sel0_b5/B1 , n70[5], n181);
  and \sel0_b5/and_b0_10  (\sel0_b5/B10 , n57[5], n172);
  and \sel0_b5/and_b0_11  (\sel0_b5/B11 , n57[5], n171);
  and \sel0_b5/and_b0_12  (\sel0_b5/B12 , n57[5], n170);
  and \sel0_b5/and_b0_13  (\sel0_b5/B13 , n57[5], n169);
  and \sel0_b5/and_b0_14  (\sel0_b5/B14 , n57[5], n168);
  and \sel0_b5/and_b0_15  (\sel0_b5/B15 , n57[5], n167);
  and \sel0_b5/and_b0_16  (\sel0_b5/B16 , n57[5], n166);
  and \sel0_b5/and_b0_17  (\sel0_b5/B17 , n57[5], n165);
  and \sel0_b5/and_b0_18  (\sel0_b5/B18 , n57[5], n164);
  and \sel0_b5/and_b0_19  (\sel0_b5/B19 , n57[5], n163);
  and \sel0_b5/and_b0_2  (\sel0_b5/B2 , n57[5], n180);
  and \sel0_b5/and_b0_20  (\sel0_b5/B20 , n57[5], n162);
  and \sel0_b5/and_b0_21  (\sel0_b5/B21 , n57[5], n161);
  and \sel0_b5/and_b0_22  (\sel0_b5/B22 , n57[5], n160);
  and \sel0_b5/and_b0_23  (\sel0_b5/B23 , n57[5], n159);
  and \sel0_b5/and_b0_24  (\sel0_b5/B24 , n48[5], n158);
  and \sel0_b5/and_b0_25  (\sel0_b5/B25 , n57[5], n157);
  and \sel0_b5/and_b0_26  (\sel0_b5/B26 , n57[5], n156);
  and \sel0_b5/and_b0_27  (\sel0_b5/B27 , n57[5], n155);
  and \sel0_b5/and_b0_28  (\sel0_b5/B28 , n57[5], n154);
  and \sel0_b5/and_b0_29  (\sel0_b5/B29 , n57[5], n153);
  and \sel0_b5/and_b0_3  (\sel0_b5/B3 , n70[5], n179);
  and \sel0_b5/and_b0_30  (\sel0_b5/B30 , n57[5], n152);
  and \sel0_b5/and_b0_31  (\sel0_b5/B31 , n57[5], n151);
  and \sel0_b5/and_b0_32  (\sel0_b5/B32 , n57[5], n150);
  and \sel0_b5/and_b0_33  (\sel0_b5/B33 , n57[5], n149);
  and \sel0_b5/and_b0_34  (\sel0_b5/B34 , n38[5], n148);
  and \sel0_b5/and_b0_35  (\sel0_b5/B35 , n37[5], n147);
  and \sel0_b5/and_b0_36  (\sel0_b5/B36 , n35[5], n146);
  and \sel0_b5/and_b0_4  (\sel0_b5/B4 , n57[5], n178);
  and \sel0_b5/and_b0_5  (\sel0_b5/B5 , n57[5], n177);
  and \sel0_b5/and_b0_6  (\sel0_b5/B6 , n57[5], n176);
  and \sel0_b5/and_b0_7  (\sel0_b5/B7 , n57[5], n175);
  and \sel0_b5/and_b0_8  (\sel0_b5/B8 , n57[5], n174);
  and \sel0_b5/and_b0_9  (\sel0_b5/B9 , n57[5], n173);
  or \sel0_b5/or_B0_B1  (\sel0_b5/or_B0_B1_o , \sel0_b5/B0 , \sel0_b5/B1 );
  or \sel0_b5/or_B11_B12  (\sel0_b5/or_B11_B12_o , \sel0_b5/B11 , \sel0_b5/B12 );
  or \sel0_b5/or_B13_B14  (\sel0_b5/or_B13_B14_o , \sel0_b5/B13 , \sel0_b5/B14 );
  or \sel0_b5/or_B15_or_B16_B17_o  (\sel0_b5/or_B15_or_B16_B17_o_o , \sel0_b5/B15 , \sel0_b5/or_B16_B17_o );
  or \sel0_b5/or_B16_B17  (\sel0_b5/or_B16_B17_o , \sel0_b5/B16 , \sel0_b5/B17 );
  or \sel0_b5/or_B18_B19  (\sel0_b5/or_B18_B19_o , \sel0_b5/B18 , \sel0_b5/B19 );
  or \sel0_b5/or_B20_B21  (\sel0_b5/or_B20_B21_o , \sel0_b5/B20 , \sel0_b5/B21 );
  or \sel0_b5/or_B22_B23  (\sel0_b5/or_B22_B23_o , \sel0_b5/B22 , \sel0_b5/B23 );
  or \sel0_b5/or_B24_or_B25_B26_o  (\sel0_b5/or_B24_or_B25_B26_o_o , \sel0_b5/B24 , \sel0_b5/or_B25_B26_o );
  or \sel0_b5/or_B25_B26  (\sel0_b5/or_B25_B26_o , \sel0_b5/B25 , \sel0_b5/B26 );
  or \sel0_b5/or_B27_B28  (\sel0_b5/or_B27_B28_o , \sel0_b5/B27 , \sel0_b5/B28 );
  or \sel0_b5/or_B29_or_B30_B31_o  (\sel0_b5/or_B29_or_B30_B31_o_o , \sel0_b5/B29 , \sel0_b5/or_B30_B31_o );
  or \sel0_b5/or_B2_B3  (\sel0_b5/or_B2_B3_o , \sel0_b5/B2 , \sel0_b5/B3 );
  or \sel0_b5/or_B30_B31  (\sel0_b5/or_B30_B31_o , \sel0_b5/B30 , \sel0_b5/B31 );
  or \sel0_b5/or_B32_B33  (\sel0_b5/or_B32_B33_o , \sel0_b5/B32 , \sel0_b5/B33 );
  or \sel0_b5/or_B34_or_B35_B36_o  (\sel0_b5/or_B34_or_B35_B36_o_o , \sel0_b5/B34 , \sel0_b5/or_B35_B36_o );
  or \sel0_b5/or_B35_B36  (\sel0_b5/or_B35_B36_o , \sel0_b5/B35 , \sel0_b5/B36 );
  or \sel0_b5/or_B4_B5  (\sel0_b5/or_B4_B5_o , \sel0_b5/B4 , \sel0_b5/B5 );
  or \sel0_b5/or_B6_or_B7_B8_o  (\sel0_b5/or_B6_or_B7_B8_o_o , \sel0_b5/B6 , \sel0_b5/or_B7_B8_o );
  or \sel0_b5/or_B7_B8  (\sel0_b5/or_B7_B8_o , \sel0_b5/B7 , \sel0_b5/B8 );
  or \sel0_b5/or_B9_B10  (\sel0_b5/or_B9_B10_o , \sel0_b5/B9 , \sel0_b5/B10 );
  or \sel0_b5/or_or_B0_B1_o_or_B2_  (\sel0_b5/or_or_B0_B1_o_or_B2__o , \sel0_b5/or_B0_B1_o , \sel0_b5/or_B2_B3_o );
  or \sel0_b5/or_or_B13_B14_o_or_B  (\sel0_b5/or_or_B13_B14_o_or_B_o , \sel0_b5/or_B13_B14_o , \sel0_b5/or_B15_or_B16_B17_o_o );
  or \sel0_b5/or_or_B18_B19_o_or_B  (\sel0_b5/or_or_B18_B19_o_or_B_o , \sel0_b5/or_B18_B19_o , \sel0_b5/or_B20_B21_o );
  or \sel0_b5/or_or_B22_B23_o_or_B  (\sel0_b5/or_or_B22_B23_o_or_B_o , \sel0_b5/or_B22_B23_o , \sel0_b5/or_B24_or_B25_B26_o_o );
  or \sel0_b5/or_or_B27_B28_o_or_B  (\sel0_b5/or_or_B27_B28_o_or_B_o , \sel0_b5/or_B27_B28_o , \sel0_b5/or_B29_or_B30_B31_o_o );
  or \sel0_b5/or_or_B32_B33_o_or_B  (\sel0_b5/or_or_B32_B33_o_or_B_o , \sel0_b5/or_B32_B33_o , \sel0_b5/or_B34_or_B35_B36_o_o );
  or \sel0_b5/or_or_B4_B5_o_or_B6_  (\sel0_b5/or_or_B4_B5_o_or_B6__o , \sel0_b5/or_B4_B5_o , \sel0_b5/or_B6_or_B7_B8_o_o );
  or \sel0_b5/or_or_B9_B10_o_or_B1  (\sel0_b5/or_or_B9_B10_o_or_B1_o , \sel0_b5/or_B9_B10_o , \sel0_b5/or_B11_B12_o );
  or \sel0_b5/or_or_or_B0_B1_o_or_  (\sel0_b5/or_or_or_B0_B1_o_or__o , \sel0_b5/or_or_B0_B1_o_or_B2__o , \sel0_b5/or_or_B4_B5_o_or_B6__o );
  or \sel0_b5/or_or_or_B18_B19_o_o  (\sel0_b5/or_or_or_B18_B19_o_o_o , \sel0_b5/or_or_B18_B19_o_or_B_o , \sel0_b5/or_or_B22_B23_o_or_B_o );
  or \sel0_b5/or_or_or_B27_B28_o_o  (\sel0_b5/or_or_or_B27_B28_o_o_o , \sel0_b5/or_or_B27_B28_o_or_B_o , \sel0_b5/or_or_B32_B33_o_or_B_o );
  or \sel0_b5/or_or_or_B9_B10_o_or  (\sel0_b5/or_or_or_B9_B10_o_or_o , \sel0_b5/or_or_B9_B10_o_or_B1_o , \sel0_b5/or_or_B13_B14_o_or_B_o );
  or \sel0_b5/or_or_or_or_B0_B1_o_  (\sel0_b5/or_or_or_or_B0_B1_o__o , \sel0_b5/or_or_or_B0_B1_o_or__o , \sel0_b5/or_or_or_B9_B10_o_or_o );
  or \sel0_b5/or_or_or_or_B18_B19_  (\sel0_b5/or_or_or_or_B18_B19__o , \sel0_b5/or_or_or_B18_B19_o_o_o , \sel0_b5/or_or_or_B27_B28_o_o_o );
  or \sel0_b5/or_or_or_or_or_B0_B1  (n99[5], \sel0_b5/or_or_or_or_B0_B1_o__o , \sel0_b5/or_or_or_or_B18_B19__o );
  and \sel0_b6/and_b0_0  (\sel0_b6/B0 , state_next[6], n182);
  and \sel0_b6/and_b0_1  (\sel0_b6/B1 , n70[6], n181);
  and \sel0_b6/and_b0_10  (\sel0_b6/B10 , n57[6], n172);
  and \sel0_b6/and_b0_11  (\sel0_b6/B11 , n57[6], n171);
  and \sel0_b6/and_b0_12  (\sel0_b6/B12 , n57[6], n170);
  and \sel0_b6/and_b0_13  (\sel0_b6/B13 , n57[6], n169);
  and \sel0_b6/and_b0_14  (\sel0_b6/B14 , n48[6], n168);
  and \sel0_b6/and_b0_15  (\sel0_b6/B15 , n57[6], n167);
  and \sel0_b6/and_b0_16  (\sel0_b6/B16 , n57[6], n166);
  and \sel0_b6/and_b0_17  (\sel0_b6/B17 , n57[6], n165);
  and \sel0_b6/and_b0_18  (\sel0_b6/B18 , n57[6], n164);
  and \sel0_b6/and_b0_19  (\sel0_b6/B19 , n57[6], n163);
  and \sel0_b6/and_b0_2  (\sel0_b6/B2 , n57[6], n180);
  and \sel0_b6/and_b0_20  (\sel0_b6/B20 , n57[6], n162);
  and \sel0_b6/and_b0_21  (\sel0_b6/B21 , n57[6], n161);
  and \sel0_b6/and_b0_22  (\sel0_b6/B22 , n57[6], n160);
  and \sel0_b6/and_b0_23  (\sel0_b6/B23 , n57[6], n159);
  and \sel0_b6/and_b0_24  (\sel0_b6/B24 , n48[6], n158);
  and \sel0_b6/and_b0_25  (\sel0_b6/B25 , n57[6], n157);
  and \sel0_b6/and_b0_26  (\sel0_b6/B26 , n57[6], n156);
  and \sel0_b6/and_b0_27  (\sel0_b6/B27 , n57[6], n155);
  and \sel0_b6/and_b0_28  (\sel0_b6/B28 , n57[6], n154);
  and \sel0_b6/and_b0_29  (\sel0_b6/B29 , n57[6], n153);
  and \sel0_b6/and_b0_3  (\sel0_b6/B3 , n70[6], n179);
  and \sel0_b6/and_b0_30  (\sel0_b6/B30 , n57[6], n152);
  and \sel0_b6/and_b0_31  (\sel0_b6/B31 , n57[6], n151);
  and \sel0_b6/and_b0_32  (\sel0_b6/B32 , n57[6], n150);
  and \sel0_b6/and_b0_33  (\sel0_b6/B33 , n57[6], n149);
  and \sel0_b6/and_b0_34  (\sel0_b6/B34 , n38[6], n148);
  and \sel0_b6/and_b0_35  (\sel0_b6/B35 , n37[6], n147);
  and \sel0_b6/and_b0_36  (\sel0_b6/B36 , n35[6], n146);
  and \sel0_b6/and_b0_4  (\sel0_b6/B4 , n57[6], n178);
  and \sel0_b6/and_b0_5  (\sel0_b6/B5 , n57[6], n177);
  and \sel0_b6/and_b0_6  (\sel0_b6/B6 , n57[6], n176);
  and \sel0_b6/and_b0_7  (\sel0_b6/B7 , n57[6], n175);
  and \sel0_b6/and_b0_8  (\sel0_b6/B8 , n57[6], n174);
  and \sel0_b6/and_b0_9  (\sel0_b6/B9 , n57[6], n173);
  or \sel0_b6/or_B0_B1  (\sel0_b6/or_B0_B1_o , \sel0_b6/B0 , \sel0_b6/B1 );
  or \sel0_b6/or_B11_B12  (\sel0_b6/or_B11_B12_o , \sel0_b6/B11 , \sel0_b6/B12 );
  or \sel0_b6/or_B13_B14  (\sel0_b6/or_B13_B14_o , \sel0_b6/B13 , \sel0_b6/B14 );
  or \sel0_b6/or_B15_or_B16_B17_o  (\sel0_b6/or_B15_or_B16_B17_o_o , \sel0_b6/B15 , \sel0_b6/or_B16_B17_o );
  or \sel0_b6/or_B16_B17  (\sel0_b6/or_B16_B17_o , \sel0_b6/B16 , \sel0_b6/B17 );
  or \sel0_b6/or_B18_B19  (\sel0_b6/or_B18_B19_o , \sel0_b6/B18 , \sel0_b6/B19 );
  or \sel0_b6/or_B20_B21  (\sel0_b6/or_B20_B21_o , \sel0_b6/B20 , \sel0_b6/B21 );
  or \sel0_b6/or_B22_B23  (\sel0_b6/or_B22_B23_o , \sel0_b6/B22 , \sel0_b6/B23 );
  or \sel0_b6/or_B24_or_B25_B26_o  (\sel0_b6/or_B24_or_B25_B26_o_o , \sel0_b6/B24 , \sel0_b6/or_B25_B26_o );
  or \sel0_b6/or_B25_B26  (\sel0_b6/or_B25_B26_o , \sel0_b6/B25 , \sel0_b6/B26 );
  or \sel0_b6/or_B27_B28  (\sel0_b6/or_B27_B28_o , \sel0_b6/B27 , \sel0_b6/B28 );
  or \sel0_b6/or_B29_or_B30_B31_o  (\sel0_b6/or_B29_or_B30_B31_o_o , \sel0_b6/B29 , \sel0_b6/or_B30_B31_o );
  or \sel0_b6/or_B2_B3  (\sel0_b6/or_B2_B3_o , \sel0_b6/B2 , \sel0_b6/B3 );
  or \sel0_b6/or_B30_B31  (\sel0_b6/or_B30_B31_o , \sel0_b6/B30 , \sel0_b6/B31 );
  or \sel0_b6/or_B32_B33  (\sel0_b6/or_B32_B33_o , \sel0_b6/B32 , \sel0_b6/B33 );
  or \sel0_b6/or_B34_or_B35_B36_o  (\sel0_b6/or_B34_or_B35_B36_o_o , \sel0_b6/B34 , \sel0_b6/or_B35_B36_o );
  or \sel0_b6/or_B35_B36  (\sel0_b6/or_B35_B36_o , \sel0_b6/B35 , \sel0_b6/B36 );
  or \sel0_b6/or_B4_B5  (\sel0_b6/or_B4_B5_o , \sel0_b6/B4 , \sel0_b6/B5 );
  or \sel0_b6/or_B6_or_B7_B8_o  (\sel0_b6/or_B6_or_B7_B8_o_o , \sel0_b6/B6 , \sel0_b6/or_B7_B8_o );
  or \sel0_b6/or_B7_B8  (\sel0_b6/or_B7_B8_o , \sel0_b6/B7 , \sel0_b6/B8 );
  or \sel0_b6/or_B9_B10  (\sel0_b6/or_B9_B10_o , \sel0_b6/B9 , \sel0_b6/B10 );
  or \sel0_b6/or_or_B0_B1_o_or_B2_  (\sel0_b6/or_or_B0_B1_o_or_B2__o , \sel0_b6/or_B0_B1_o , \sel0_b6/or_B2_B3_o );
  or \sel0_b6/or_or_B13_B14_o_or_B  (\sel0_b6/or_or_B13_B14_o_or_B_o , \sel0_b6/or_B13_B14_o , \sel0_b6/or_B15_or_B16_B17_o_o );
  or \sel0_b6/or_or_B18_B19_o_or_B  (\sel0_b6/or_or_B18_B19_o_or_B_o , \sel0_b6/or_B18_B19_o , \sel0_b6/or_B20_B21_o );
  or \sel0_b6/or_or_B22_B23_o_or_B  (\sel0_b6/or_or_B22_B23_o_or_B_o , \sel0_b6/or_B22_B23_o , \sel0_b6/or_B24_or_B25_B26_o_o );
  or \sel0_b6/or_or_B27_B28_o_or_B  (\sel0_b6/or_or_B27_B28_o_or_B_o , \sel0_b6/or_B27_B28_o , \sel0_b6/or_B29_or_B30_B31_o_o );
  or \sel0_b6/or_or_B32_B33_o_or_B  (\sel0_b6/or_or_B32_B33_o_or_B_o , \sel0_b6/or_B32_B33_o , \sel0_b6/or_B34_or_B35_B36_o_o );
  or \sel0_b6/or_or_B4_B5_o_or_B6_  (\sel0_b6/or_or_B4_B5_o_or_B6__o , \sel0_b6/or_B4_B5_o , \sel0_b6/or_B6_or_B7_B8_o_o );
  or \sel0_b6/or_or_B9_B10_o_or_B1  (\sel0_b6/or_or_B9_B10_o_or_B1_o , \sel0_b6/or_B9_B10_o , \sel0_b6/or_B11_B12_o );
  or \sel0_b6/or_or_or_B0_B1_o_or_  (\sel0_b6/or_or_or_B0_B1_o_or__o , \sel0_b6/or_or_B0_B1_o_or_B2__o , \sel0_b6/or_or_B4_B5_o_or_B6__o );
  or \sel0_b6/or_or_or_B18_B19_o_o  (\sel0_b6/or_or_or_B18_B19_o_o_o , \sel0_b6/or_or_B18_B19_o_or_B_o , \sel0_b6/or_or_B22_B23_o_or_B_o );
  or \sel0_b6/or_or_or_B27_B28_o_o  (\sel0_b6/or_or_or_B27_B28_o_o_o , \sel0_b6/or_or_B27_B28_o_or_B_o , \sel0_b6/or_or_B32_B33_o_or_B_o );
  or \sel0_b6/or_or_or_B9_B10_o_or  (\sel0_b6/or_or_or_B9_B10_o_or_o , \sel0_b6/or_or_B9_B10_o_or_B1_o , \sel0_b6/or_or_B13_B14_o_or_B_o );
  or \sel0_b6/or_or_or_or_B0_B1_o_  (\sel0_b6/or_or_or_or_B0_B1_o__o , \sel0_b6/or_or_or_B0_B1_o_or__o , \sel0_b6/or_or_or_B9_B10_o_or_o );
  or \sel0_b6/or_or_or_or_B18_B19_  (\sel0_b6/or_or_or_or_B18_B19__o , \sel0_b6/or_or_or_B18_B19_o_o_o , \sel0_b6/or_or_or_B27_B28_o_o_o );
  or \sel0_b6/or_or_or_or_or_B0_B1  (n99[6], \sel0_b6/or_or_or_or_B0_B1_o__o , \sel0_b6/or_or_or_or_B18_B19__o );
  and \sel0_b7/and_b0_0  (\sel0_b7/B0 , state_next[7], n182);
  and \sel0_b7/and_b0_1  (\sel0_b7/B1 , n70[7], n181);
  and \sel0_b7/and_b0_10  (\sel0_b7/B10 , n57[7], n172);
  and \sel0_b7/and_b0_11  (\sel0_b7/B11 , n57[7], n171);
  and \sel0_b7/and_b0_12  (\sel0_b7/B12 , n57[7], n170);
  and \sel0_b7/and_b0_13  (\sel0_b7/B13 , n57[7], n169);
  and \sel0_b7/and_b0_14  (\sel0_b7/B14 , n59[7], n168);
  and \sel0_b7/and_b0_15  (\sel0_b7/B15 , n57[7], n167);
  and \sel0_b7/and_b0_16  (\sel0_b7/B16 , n57[7], n166);
  and \sel0_b7/and_b0_17  (\sel0_b7/B17 , n57[7], n165);
  and \sel0_b7/and_b0_18  (\sel0_b7/B18 , n57[7], n164);
  and \sel0_b7/and_b0_19  (\sel0_b7/B19 , n57[7], n163);
  and \sel0_b7/and_b0_2  (\sel0_b7/B2 , n57[7], n180);
  and \sel0_b7/and_b0_20  (\sel0_b7/B20 , n57[7], n162);
  and \sel0_b7/and_b0_21  (\sel0_b7/B21 , n57[7], n161);
  and \sel0_b7/and_b0_22  (\sel0_b7/B22 , n57[7], n160);
  and \sel0_b7/and_b0_23  (\sel0_b7/B23 , n57[7], n159);
  and \sel0_b7/and_b0_24  (\sel0_b7/B24 , n57[7], n158);
  and \sel0_b7/and_b0_25  (\sel0_b7/B25 , n57[7], n157);
  and \sel0_b7/and_b0_26  (\sel0_b7/B26 , n57[7], n156);
  and \sel0_b7/and_b0_27  (\sel0_b7/B27 , n57[7], n155);
  and \sel0_b7/and_b0_28  (\sel0_b7/B28 , n57[7], n154);
  and \sel0_b7/and_b0_29  (\sel0_b7/B29 , n57[7], n153);
  and \sel0_b7/and_b0_3  (\sel0_b7/B3 , n70[7], n179);
  and \sel0_b7/and_b0_30  (\sel0_b7/B30 , n57[7], n152);
  and \sel0_b7/and_b0_31  (\sel0_b7/B31 , n57[7], n151);
  and \sel0_b7/and_b0_32  (\sel0_b7/B32 , n57[7], n150);
  and \sel0_b7/and_b0_33  (\sel0_b7/B33 , n57[7], n149);
  and \sel0_b7/and_b0_34  (\sel0_b7/B34 , n70[7], n148);
  and \sel0_b7/and_b0_35  (\sel0_b7/B35 , n57[7], n147);
  and \sel0_b7/and_b0_36  (\sel0_b7/B36 , n35[7], n146);
  and \sel0_b7/and_b0_4  (\sel0_b7/B4 , n57[7], n178);
  and \sel0_b7/and_b0_5  (\sel0_b7/B5 , n57[7], n177);
  and \sel0_b7/and_b0_6  (\sel0_b7/B6 , n57[7], n176);
  and \sel0_b7/and_b0_7  (\sel0_b7/B7 , n57[7], n175);
  and \sel0_b7/and_b0_8  (\sel0_b7/B8 , n57[7], n174);
  and \sel0_b7/and_b0_9  (\sel0_b7/B9 , n57[7], n173);
  or \sel0_b7/or_B0_B1  (\sel0_b7/or_B0_B1_o , \sel0_b7/B0 , \sel0_b7/B1 );
  or \sel0_b7/or_B11_B12  (\sel0_b7/or_B11_B12_o , \sel0_b7/B11 , \sel0_b7/B12 );
  or \sel0_b7/or_B13_B14  (\sel0_b7/or_B13_B14_o , \sel0_b7/B13 , \sel0_b7/B14 );
  or \sel0_b7/or_B15_or_B16_B17_o  (\sel0_b7/or_B15_or_B16_B17_o_o , \sel0_b7/B15 , \sel0_b7/or_B16_B17_o );
  or \sel0_b7/or_B16_B17  (\sel0_b7/or_B16_B17_o , \sel0_b7/B16 , \sel0_b7/B17 );
  or \sel0_b7/or_B18_B19  (\sel0_b7/or_B18_B19_o , \sel0_b7/B18 , \sel0_b7/B19 );
  or \sel0_b7/or_B20_B21  (\sel0_b7/or_B20_B21_o , \sel0_b7/B20 , \sel0_b7/B21 );
  or \sel0_b7/or_B22_B23  (\sel0_b7/or_B22_B23_o , \sel0_b7/B22 , \sel0_b7/B23 );
  or \sel0_b7/or_B24_or_B25_B26_o  (\sel0_b7/or_B24_or_B25_B26_o_o , \sel0_b7/B24 , \sel0_b7/or_B25_B26_o );
  or \sel0_b7/or_B25_B26  (\sel0_b7/or_B25_B26_o , \sel0_b7/B25 , \sel0_b7/B26 );
  or \sel0_b7/or_B27_B28  (\sel0_b7/or_B27_B28_o , \sel0_b7/B27 , \sel0_b7/B28 );
  or \sel0_b7/or_B29_or_B30_B31_o  (\sel0_b7/or_B29_or_B30_B31_o_o , \sel0_b7/B29 , \sel0_b7/or_B30_B31_o );
  or \sel0_b7/or_B2_B3  (\sel0_b7/or_B2_B3_o , \sel0_b7/B2 , \sel0_b7/B3 );
  or \sel0_b7/or_B30_B31  (\sel0_b7/or_B30_B31_o , \sel0_b7/B30 , \sel0_b7/B31 );
  or \sel0_b7/or_B32_B33  (\sel0_b7/or_B32_B33_o , \sel0_b7/B32 , \sel0_b7/B33 );
  or \sel0_b7/or_B34_or_B35_B36_o  (\sel0_b7/or_B34_or_B35_B36_o_o , \sel0_b7/B34 , \sel0_b7/or_B35_B36_o );
  or \sel0_b7/or_B35_B36  (\sel0_b7/or_B35_B36_o , \sel0_b7/B35 , \sel0_b7/B36 );
  or \sel0_b7/or_B4_B5  (\sel0_b7/or_B4_B5_o , \sel0_b7/B4 , \sel0_b7/B5 );
  or \sel0_b7/or_B6_or_B7_B8_o  (\sel0_b7/or_B6_or_B7_B8_o_o , \sel0_b7/B6 , \sel0_b7/or_B7_B8_o );
  or \sel0_b7/or_B7_B8  (\sel0_b7/or_B7_B8_o , \sel0_b7/B7 , \sel0_b7/B8 );
  or \sel0_b7/or_B9_B10  (\sel0_b7/or_B9_B10_o , \sel0_b7/B9 , \sel0_b7/B10 );
  or \sel0_b7/or_or_B0_B1_o_or_B2_  (\sel0_b7/or_or_B0_B1_o_or_B2__o , \sel0_b7/or_B0_B1_o , \sel0_b7/or_B2_B3_o );
  or \sel0_b7/or_or_B13_B14_o_or_B  (\sel0_b7/or_or_B13_B14_o_or_B_o , \sel0_b7/or_B13_B14_o , \sel0_b7/or_B15_or_B16_B17_o_o );
  or \sel0_b7/or_or_B18_B19_o_or_B  (\sel0_b7/or_or_B18_B19_o_or_B_o , \sel0_b7/or_B18_B19_o , \sel0_b7/or_B20_B21_o );
  or \sel0_b7/or_or_B22_B23_o_or_B  (\sel0_b7/or_or_B22_B23_o_or_B_o , \sel0_b7/or_B22_B23_o , \sel0_b7/or_B24_or_B25_B26_o_o );
  or \sel0_b7/or_or_B27_B28_o_or_B  (\sel0_b7/or_or_B27_B28_o_or_B_o , \sel0_b7/or_B27_B28_o , \sel0_b7/or_B29_or_B30_B31_o_o );
  or \sel0_b7/or_or_B32_B33_o_or_B  (\sel0_b7/or_or_B32_B33_o_or_B_o , \sel0_b7/or_B32_B33_o , \sel0_b7/or_B34_or_B35_B36_o_o );
  or \sel0_b7/or_or_B4_B5_o_or_B6_  (\sel0_b7/or_or_B4_B5_o_or_B6__o , \sel0_b7/or_B4_B5_o , \sel0_b7/or_B6_or_B7_B8_o_o );
  or \sel0_b7/or_or_B9_B10_o_or_B1  (\sel0_b7/or_or_B9_B10_o_or_B1_o , \sel0_b7/or_B9_B10_o , \sel0_b7/or_B11_B12_o );
  or \sel0_b7/or_or_or_B0_B1_o_or_  (\sel0_b7/or_or_or_B0_B1_o_or__o , \sel0_b7/or_or_B0_B1_o_or_B2__o , \sel0_b7/or_or_B4_B5_o_or_B6__o );
  or \sel0_b7/or_or_or_B18_B19_o_o  (\sel0_b7/or_or_or_B18_B19_o_o_o , \sel0_b7/or_or_B18_B19_o_or_B_o , \sel0_b7/or_or_B22_B23_o_or_B_o );
  or \sel0_b7/or_or_or_B27_B28_o_o  (\sel0_b7/or_or_or_B27_B28_o_o_o , \sel0_b7/or_or_B27_B28_o_or_B_o , \sel0_b7/or_or_B32_B33_o_or_B_o );
  or \sel0_b7/or_or_or_B9_B10_o_or  (\sel0_b7/or_or_or_B9_B10_o_or_o , \sel0_b7/or_or_B9_B10_o_or_B1_o , \sel0_b7/or_or_B13_B14_o_or_B_o );
  or \sel0_b7/or_or_or_or_B0_B1_o_  (\sel0_b7/or_or_or_or_B0_B1_o__o , \sel0_b7/or_or_or_B0_B1_o_or__o , \sel0_b7/or_or_or_B9_B10_o_or_o );
  or \sel0_b7/or_or_or_or_B18_B19_  (\sel0_b7/or_or_or_or_B18_B19__o , \sel0_b7/or_or_or_B18_B19_o_o_o , \sel0_b7/or_or_or_B27_B28_o_o_o );
  or \sel0_b7/or_or_or_or_or_B0_B1  (n99[7], \sel0_b7/or_or_or_or_B0_B1_o__o , \sel0_b7/or_or_or_or_B18_B19__o );
  and \sel1/and_b0_0  (\sel1/B0 , sda, n181);
  and \sel1/and_b0_1  (\sel1/B1 , n145, n180);
  and \sel1/and_b0_10  (\sel1/B10 , n136, n171);
  and \sel1/and_b0_11  (\sel1/B11 , n135, n170);
  and \sel1/and_b0_12  (\sel1/B12 , n134, n169);
  and \sel1/and_b0_13  (\sel1/B13 , n106, n168);
  and \sel1/and_b0_14  (\sel1/B14 , n106, n167);
  and \sel1/and_b0_15  (\sel1/B15 , n133, n166);
  and \sel1/and_b0_16  (\sel1/B16 , n132, n165);
  and \sel1/and_b0_17  (\sel1/B17 , n131, n164);
  and \sel1/and_b0_18  (\sel1/B18 , n130, n163);
  and \sel1/and_b0_19  (\sel1/B19 , n129, n162);
  and \sel1/and_b0_2  (\sel1/B2 , n112, n179);
  and \sel1/and_b0_20  (\sel1/B20 , n128, n161);
  and \sel1/and_b0_21  (\sel1/B21 , n127, n160);
  and \sel1/and_b0_22  (\sel1/B22 , n126, n159);
  and \sel1/and_b0_23  (\sel1/B23 , n106, n158);
  and \sel1/and_b0_24  (\sel1/B24 , n106, n157);
  and \sel1/and_b0_25  (\sel1/B25 , n123, n156);
  and \sel1/and_b0_26  (\sel1/B26 , n122, n155);
  and \sel1/and_b0_27  (\sel1/B27 , n121, n154);
  and \sel1/and_b0_28  (\sel1/B28 , n120, n153);
  and \sel1/and_b0_29  (\sel1/B29 , n119, n152);
  and \sel1/and_b0_3  (\sel1/B3 , n106, n178);
  and \sel1/and_b0_30  (\sel1/B30 , n118, n151);
  and \sel1/and_b0_31  (\sel1/B31 , n117, n150);
  and \sel1/and_b0_32  (\sel1/B32 , n116, n149);
  and \sel1/and_b0_33  (\sel1/B33 , n112, n148);
  and \sel1/and_b0_34  (\sel1/B34 , n106, n147);
  and \sel1/and_b0_4  (\sel1/B4 , n106, n177);
  and \sel1/and_b0_5  (\sel1/B5 , n141, n176);
  and \sel1/and_b0_6  (\sel1/B6 , n140, n175);
  and \sel1/and_b0_7  (\sel1/B7 , n139, n174);
  and \sel1/and_b0_8  (\sel1/B8 , n138, n173);
  and \sel1/and_b0_9  (\sel1/B9 , n137, n172);
  or \sel1/or_B0_B1  (\sel1/or_B0_B1_o , \sel1/B0 , \sel1/B1 );
  or \sel1/or_B11_B12  (\sel1/or_B11_B12_o , \sel1/B11 , \sel1/B12 );
  or \sel1/or_B13_B14  (\sel1/or_B13_B14_o , \sel1/B13 , \sel1/B14 );
  or \sel1/or_B15_or_B16_B17_o  (\sel1/or_B15_or_B16_B17_o_o , \sel1/B15 , \sel1/or_B16_B17_o );
  or \sel1/or_B16_B17  (\sel1/or_B16_B17_o , \sel1/B16 , \sel1/B17 );
  or \sel1/or_B18_B19  (\sel1/or_B18_B19_o , \sel1/B18 , \sel1/B19 );
  or \sel1/or_B20_B21  (\sel1/or_B20_B21_o , \sel1/B20 , \sel1/B21 );
  or \sel1/or_B22_B23  (\sel1/or_B22_B23_o , \sel1/B22 , \sel1/B23 );
  or \sel1/or_B24_or_B25_B26_o  (\sel1/or_B24_or_B25_B26_o_o , \sel1/B24 , \sel1/or_B25_B26_o );
  or \sel1/or_B25_B26  (\sel1/or_B25_B26_o , \sel1/B25 , \sel1/B26 );
  or \sel1/or_B27_B28  (\sel1/or_B27_B28_o , \sel1/B27 , \sel1/B28 );
  or \sel1/or_B29_B30  (\sel1/or_B29_B30_o , \sel1/B29 , \sel1/B30 );
  or \sel1/or_B2_B3  (\sel1/or_B2_B3_o , \sel1/B2 , \sel1/B3 );
  or \sel1/or_B31_B32  (\sel1/or_B31_B32_o , \sel1/B31 , \sel1/B32 );
  or \sel1/or_B33_or_B34_B35_o  (\sel1/or_B33_or_B34_B35_o_o , \sel1/B33 , \sel1/or_B34_B35_o );
  or \sel1/or_B34_B35  (\sel1/or_B34_B35_o , \sel1/B34 , n183);
  or \sel1/or_B4_B5  (\sel1/or_B4_B5_o , \sel1/B4 , \sel1/B5 );
  or \sel1/or_B6_or_B7_B8_o  (\sel1/or_B6_or_B7_B8_o_o , \sel1/B6 , \sel1/or_B7_B8_o );
  or \sel1/or_B7_B8  (\sel1/or_B7_B8_o , \sel1/B7 , \sel1/B8 );
  or \sel1/or_B9_B10  (\sel1/or_B9_B10_o , \sel1/B9 , \sel1/B10 );
  or \sel1/or_or_B0_B1_o_or_B2_  (\sel1/or_or_B0_B1_o_or_B2__o , \sel1/or_B0_B1_o , \sel1/or_B2_B3_o );
  or \sel1/or_or_B13_B14_o_or_B  (\sel1/or_or_B13_B14_o_or_B_o , \sel1/or_B13_B14_o , \sel1/or_B15_or_B16_B17_o_o );
  or \sel1/or_or_B18_B19_o_or_B  (\sel1/or_or_B18_B19_o_or_B_o , \sel1/or_B18_B19_o , \sel1/or_B20_B21_o );
  or \sel1/or_or_B22_B23_o_or_B  (\sel1/or_or_B22_B23_o_or_B_o , \sel1/or_B22_B23_o , \sel1/or_B24_or_B25_B26_o_o );
  or \sel1/or_or_B27_B28_o_or_B  (\sel1/or_or_B27_B28_o_or_B_o , \sel1/or_B27_B28_o , \sel1/or_B29_B30_o );
  or \sel1/or_or_B31_B32_o_or_B  (\sel1/or_or_B31_B32_o_or_B_o , \sel1/or_B31_B32_o , \sel1/or_B33_or_B34_B35_o_o );
  or \sel1/or_or_B4_B5_o_or_B6_  (\sel1/or_or_B4_B5_o_or_B6__o , \sel1/or_B4_B5_o , \sel1/or_B6_or_B7_B8_o_o );
  or \sel1/or_or_B9_B10_o_or_B1  (\sel1/or_or_B9_B10_o_or_B1_o , \sel1/or_B9_B10_o , \sel1/or_B11_B12_o );
  or \sel1/or_or_or_B0_B1_o_or_  (\sel1/or_or_or_B0_B1_o_or__o , \sel1/or_or_B0_B1_o_or_B2__o , \sel1/or_or_B4_B5_o_or_B6__o );
  or \sel1/or_or_or_B18_B19_o_o  (\sel1/or_or_or_B18_B19_o_o_o , \sel1/or_or_B18_B19_o_or_B_o , \sel1/or_or_B22_B23_o_or_B_o );
  or \sel1/or_or_or_B27_B28_o_o  (\sel1/or_or_or_B27_B28_o_o_o , \sel1/or_or_B27_B28_o_or_B_o , \sel1/or_or_B31_B32_o_or_B_o );
  or \sel1/or_or_or_B9_B10_o_or  (\sel1/or_or_or_B9_B10_o_or_o , \sel1/or_or_B9_B10_o_or_B1_o , \sel1/or_or_B13_B14_o_or_B_o );
  or \sel1/or_or_or_or_B0_B1_o_  (\sel1/or_or_or_or_B0_B1_o__o , \sel1/or_or_or_B0_B1_o_or__o , \sel1/or_or_or_B9_B10_o_or_o );
  or \sel1/or_or_or_or_B18_B19_  (\sel1/or_or_or_or_B18_B19__o , \sel1/or_or_or_B18_B19_o_o_o , \sel1/or_or_or_B27_B28_o_o_o );
  or \sel1/or_or_or_or_or_B0_B1  (n184, \sel1/or_or_or_or_B0_B1_o__o , \sel1/or_or_or_or_B18_B19__o );
  and \sel2/and_b0_0  (\sel2/B0 , sda_oe, n181);
  and \sel2/and_b0_1  (\sel2/B1 , n105, n180);
  and \sel2/and_b0_10  (\sel2/B10 , n105, n171);
  and \sel2/and_b0_11  (\sel2/B11 , n105, n170);
  and \sel2/and_b0_12  (\sel2/B12 , n105, n169);
  and \sel2/and_b0_13  (\sel2/B13 , n105, n168);
  and \sel2/and_b0_14  (\sel2/B14 , n124, n167);
  and \sel2/and_b0_15  (\sel2/B15 , n105, n166);
  and \sel2/and_b0_16  (\sel2/B16 , n105, n165);
  and \sel2/and_b0_17  (\sel2/B17 , n105, n164);
  and \sel2/and_b0_18  (\sel2/B18 , n105, n163);
  and \sel2/and_b0_19  (\sel2/B19 , n105, n162);
  and \sel2/and_b0_2  (\sel2/B2 , n111, n179);
  and \sel2/and_b0_20  (\sel2/B20 , n105, n161);
  and \sel2/and_b0_21  (\sel2/B21 , n105, n160);
  and \sel2/and_b0_22  (\sel2/B22 , n105, n159);
  and \sel2/and_b0_23  (\sel2/B23 , n105, n158);
  and \sel2/and_b0_24  (\sel2/B24 , n124, n157);
  and \sel2/and_b0_25  (\sel2/B25 , n105, n156);
  and \sel2/and_b0_26  (\sel2/B26 , n105, n155);
  and \sel2/and_b0_27  (\sel2/B27 , n105, n154);
  and \sel2/and_b0_28  (\sel2/B28 , n105, n153);
  and \sel2/and_b0_29  (\sel2/B29 , n105, n152);
  and \sel2/and_b0_3  (\sel2/B3 , n105, n178);
  and \sel2/and_b0_30  (\sel2/B30 , n105, n151);
  and \sel2/and_b0_31  (\sel2/B31 , n105, n150);
  and \sel2/and_b0_32  (\sel2/B32 , n105, n149);
  and \sel2/and_b0_33  (\sel2/B33 , n111, n148);
  and \sel2/and_b0_34  (\sel2/B34 , n105, n147);
  and \sel2/and_b0_4  (\sel2/B4 , n124, n177);
  and \sel2/and_b0_5  (\sel2/B5 , n105, n176);
  and \sel2/and_b0_6  (\sel2/B6 , n105, n175);
  and \sel2/and_b0_7  (\sel2/B7 , n105, n174);
  and \sel2/and_b0_8  (\sel2/B8 , n105, n173);
  and \sel2/and_b0_9  (\sel2/B9 , n105, n172);
  or \sel2/or_B0_B1  (\sel2/or_B0_B1_o , \sel2/B0 , \sel2/B1 );
  or \sel2/or_B11_B12  (\sel2/or_B11_B12_o , \sel2/B11 , \sel2/B12 );
  or \sel2/or_B13_B14  (\sel2/or_B13_B14_o , \sel2/B13 , \sel2/B14 );
  or \sel2/or_B15_or_B16_B17_o  (\sel2/or_B15_or_B16_B17_o_o , \sel2/B15 , \sel2/or_B16_B17_o );
  or \sel2/or_B16_B17  (\sel2/or_B16_B17_o , \sel2/B16 , \sel2/B17 );
  or \sel2/or_B18_B19  (\sel2/or_B18_B19_o , \sel2/B18 , \sel2/B19 );
  or \sel2/or_B20_B21  (\sel2/or_B20_B21_o , \sel2/B20 , \sel2/B21 );
  or \sel2/or_B22_B23  (\sel2/or_B22_B23_o , \sel2/B22 , \sel2/B23 );
  or \sel2/or_B24_or_B25_B26_o  (\sel2/or_B24_or_B25_B26_o_o , \sel2/B24 , \sel2/or_B25_B26_o );
  or \sel2/or_B25_B26  (\sel2/or_B25_B26_o , \sel2/B25 , \sel2/B26 );
  or \sel2/or_B27_B28  (\sel2/or_B27_B28_o , \sel2/B27 , \sel2/B28 );
  or \sel2/or_B29_B30  (\sel2/or_B29_B30_o , \sel2/B29 , \sel2/B30 );
  or \sel2/or_B2_B3  (\sel2/or_B2_B3_o , \sel2/B2 , \sel2/B3 );
  or \sel2/or_B31_B32  (\sel2/or_B31_B32_o , \sel2/B31 , \sel2/B32 );
  or \sel2/or_B33_or_B34_B35_o  (\sel2/or_B33_or_B34_B35_o_o , \sel2/B33 , \sel2/or_B34_B35_o );
  or \sel2/or_B34_B35  (\sel2/or_B34_B35_o , \sel2/B34 , n183);
  or \sel2/or_B4_B5  (\sel2/or_B4_B5_o , \sel2/B4 , \sel2/B5 );
  or \sel2/or_B6_or_B7_B8_o  (\sel2/or_B6_or_B7_B8_o_o , \sel2/B6 , \sel2/or_B7_B8_o );
  or \sel2/or_B7_B8  (\sel2/or_B7_B8_o , \sel2/B7 , \sel2/B8 );
  or \sel2/or_B9_B10  (\sel2/or_B9_B10_o , \sel2/B9 , \sel2/B10 );
  or \sel2/or_or_B0_B1_o_or_B2_  (\sel2/or_or_B0_B1_o_or_B2__o , \sel2/or_B0_B1_o , \sel2/or_B2_B3_o );
  or \sel2/or_or_B13_B14_o_or_B  (\sel2/or_or_B13_B14_o_or_B_o , \sel2/or_B13_B14_o , \sel2/or_B15_or_B16_B17_o_o );
  or \sel2/or_or_B18_B19_o_or_B  (\sel2/or_or_B18_B19_o_or_B_o , \sel2/or_B18_B19_o , \sel2/or_B20_B21_o );
  or \sel2/or_or_B22_B23_o_or_B  (\sel2/or_or_B22_B23_o_or_B_o , \sel2/or_B22_B23_o , \sel2/or_B24_or_B25_B26_o_o );
  or \sel2/or_or_B27_B28_o_or_B  (\sel2/or_or_B27_B28_o_or_B_o , \sel2/or_B27_B28_o , \sel2/or_B29_B30_o );
  or \sel2/or_or_B31_B32_o_or_B  (\sel2/or_or_B31_B32_o_or_B_o , \sel2/or_B31_B32_o , \sel2/or_B33_or_B34_B35_o_o );
  or \sel2/or_or_B4_B5_o_or_B6_  (\sel2/or_or_B4_B5_o_or_B6__o , \sel2/or_B4_B5_o , \sel2/or_B6_or_B7_B8_o_o );
  or \sel2/or_or_B9_B10_o_or_B1  (\sel2/or_or_B9_B10_o_or_B1_o , \sel2/or_B9_B10_o , \sel2/or_B11_B12_o );
  or \sel2/or_or_or_B0_B1_o_or_  (\sel2/or_or_or_B0_B1_o_or__o , \sel2/or_or_B0_B1_o_or_B2__o , \sel2/or_or_B4_B5_o_or_B6__o );
  or \sel2/or_or_or_B18_B19_o_o  (\sel2/or_or_or_B18_B19_o_o_o , \sel2/or_or_B18_B19_o_or_B_o , \sel2/or_or_B22_B23_o_or_B_o );
  or \sel2/or_or_or_B27_B28_o_o  (\sel2/or_or_or_B27_B28_o_o_o , \sel2/or_or_B27_B28_o_or_B_o , \sel2/or_or_B31_B32_o_or_B_o );
  or \sel2/or_or_or_B9_B10_o_or  (\sel2/or_or_or_B9_B10_o_or_o , \sel2/or_or_B9_B10_o_or_B1_o , \sel2/or_or_B13_B14_o_or_B_o );
  or \sel2/or_or_or_or_B0_B1_o_  (\sel2/or_or_or_or_B0_B1_o__o , \sel2/or_or_or_B0_B1_o_or__o , \sel2/or_or_or_B9_B10_o_or_o );
  or \sel2/or_or_or_or_B18_B19_  (\sel2/or_or_or_or_B18_B19__o , \sel2/or_or_or_B18_B19_o_o_o , \sel2/or_or_or_B27_B28_o_o_o );
  or \sel2/or_or_or_or_or_B0_B1  (n186, \sel2/or_or_or_or_B0_B1_o__o , \sel2/or_or_or_or_B18_B19__o );
  and \sel3/and_b0_0  (\sel3/B0 , scl_output_enable, n181);
  and \sel3/and_b0_1  (\sel3/B1 , n104, n180);
  and \sel3/and_b0_10  (\sel3/B10 , n115, n171);
  and \sel3/and_b0_11  (\sel3/B11 , n115, n170);
  and \sel3/and_b0_12  (\sel3/B12 , n115, n169);
  and \sel3/and_b0_13  (\sel3/B13 , n104, n168);
  and \sel3/and_b0_14  (\sel3/B14 , n115, n167);
  and \sel3/and_b0_15  (\sel3/B15 , n115, n166);
  and \sel3/and_b0_16  (\sel3/B16 , n115, n165);
  and \sel3/and_b0_17  (\sel3/B17 , n115, n164);
  and \sel3/and_b0_18  (\sel3/B18 , n115, n163);
  and \sel3/and_b0_19  (\sel3/B19 , n115, n162);
  and \sel3/and_b0_2  (\sel3/B2 , n110, n179);
  and \sel3/and_b0_20  (\sel3/B20 , n115, n161);
  and \sel3/and_b0_21  (\sel3/B21 , n115, n160);
  and \sel3/and_b0_22  (\sel3/B22 , n115, n159);
  and \sel3/and_b0_23  (\sel3/B23 , n104, n158);
  and \sel3/and_b0_24  (\sel3/B24 , n115, n157);
  and \sel3/and_b0_25  (\sel3/B25 , n115, n156);
  and \sel3/and_b0_26  (\sel3/B26 , n115, n155);
  and \sel3/and_b0_27  (\sel3/B27 , n115, n154);
  and \sel3/and_b0_28  (\sel3/B28 , n115, n153);
  and \sel3/and_b0_29  (\sel3/B29 , n115, n152);
  and \sel3/and_b0_3  (\sel3/B3 , n142, n178);
  and \sel3/and_b0_30  (\sel3/B30 , n115, n151);
  and \sel3/and_b0_31  (\sel3/B31 , n115, n150);
  and \sel3/and_b0_32  (\sel3/B32 , n115, n149);
  and \sel3/and_b0_33  (\sel3/B33 , n110, n148);
  and \sel3/and_b0_34  (\sel3/B34 , n104, n147);
  and \sel3/and_b0_4  (\sel3/B4 , n115, n177);
  and \sel3/and_b0_5  (\sel3/B5 , n115, n176);
  and \sel3/and_b0_6  (\sel3/B6 , n115, n175);
  and \sel3/and_b0_7  (\sel3/B7 , n115, n174);
  and \sel3/and_b0_8  (\sel3/B8 , n115, n173);
  and \sel3/and_b0_9  (\sel3/B9 , n115, n172);
  or \sel3/or_B0_B1  (\sel3/or_B0_B1_o , \sel3/B0 , \sel3/B1 );
  or \sel3/or_B11_B12  (\sel3/or_B11_B12_o , \sel3/B11 , \sel3/B12 );
  or \sel3/or_B13_B14  (\sel3/or_B13_B14_o , \sel3/B13 , \sel3/B14 );
  or \sel3/or_B15_or_B16_B17_o  (\sel3/or_B15_or_B16_B17_o_o , \sel3/B15 , \sel3/or_B16_B17_o );
  or \sel3/or_B16_B17  (\sel3/or_B16_B17_o , \sel3/B16 , \sel3/B17 );
  or \sel3/or_B18_B19  (\sel3/or_B18_B19_o , \sel3/B18 , \sel3/B19 );
  or \sel3/or_B20_B21  (\sel3/or_B20_B21_o , \sel3/B20 , \sel3/B21 );
  or \sel3/or_B22_B23  (\sel3/or_B22_B23_o , \sel3/B22 , \sel3/B23 );
  or \sel3/or_B24_or_B25_B26_o  (\sel3/or_B24_or_B25_B26_o_o , \sel3/B24 , \sel3/or_B25_B26_o );
  or \sel3/or_B25_B26  (\sel3/or_B25_B26_o , \sel3/B25 , \sel3/B26 );
  or \sel3/or_B27_B28  (\sel3/or_B27_B28_o , \sel3/B27 , \sel3/B28 );
  or \sel3/or_B29_B30  (\sel3/or_B29_B30_o , \sel3/B29 , \sel3/B30 );
  or \sel3/or_B2_B3  (\sel3/or_B2_B3_o , \sel3/B2 , \sel3/B3 );
  or \sel3/or_B31_B32  (\sel3/or_B31_B32_o , \sel3/B31 , \sel3/B32 );
  or \sel3/or_B33_or_B34_B35_o  (\sel3/or_B33_or_B34_B35_o_o , \sel3/B33 , \sel3/B34 );
  or \sel3/or_B4_B5  (\sel3/or_B4_B5_o , \sel3/B4 , \sel3/B5 );
  or \sel3/or_B6_or_B7_B8_o  (\sel3/or_B6_or_B7_B8_o_o , \sel3/B6 , \sel3/or_B7_B8_o );
  or \sel3/or_B7_B8  (\sel3/or_B7_B8_o , \sel3/B7 , \sel3/B8 );
  or \sel3/or_B9_B10  (\sel3/or_B9_B10_o , \sel3/B9 , \sel3/B10 );
  or \sel3/or_or_B0_B1_o_or_B2_  (\sel3/or_or_B0_B1_o_or_B2__o , \sel3/or_B0_B1_o , \sel3/or_B2_B3_o );
  or \sel3/or_or_B13_B14_o_or_B  (\sel3/or_or_B13_B14_o_or_B_o , \sel3/or_B13_B14_o , \sel3/or_B15_or_B16_B17_o_o );
  or \sel3/or_or_B18_B19_o_or_B  (\sel3/or_or_B18_B19_o_or_B_o , \sel3/or_B18_B19_o , \sel3/or_B20_B21_o );
  or \sel3/or_or_B22_B23_o_or_B  (\sel3/or_or_B22_B23_o_or_B_o , \sel3/or_B22_B23_o , \sel3/or_B24_or_B25_B26_o_o );
  or \sel3/or_or_B27_B28_o_or_B  (\sel3/or_or_B27_B28_o_or_B_o , \sel3/or_B27_B28_o , \sel3/or_B29_B30_o );
  or \sel3/or_or_B31_B32_o_or_B  (\sel3/or_or_B31_B32_o_or_B_o , \sel3/or_B31_B32_o , \sel3/or_B33_or_B34_B35_o_o );
  or \sel3/or_or_B4_B5_o_or_B6_  (\sel3/or_or_B4_B5_o_or_B6__o , \sel3/or_B4_B5_o , \sel3/or_B6_or_B7_B8_o_o );
  or \sel3/or_or_B9_B10_o_or_B1  (\sel3/or_or_B9_B10_o_or_B1_o , \sel3/or_B9_B10_o , \sel3/or_B11_B12_o );
  or \sel3/or_or_or_B0_B1_o_or_  (\sel3/or_or_or_B0_B1_o_or__o , \sel3/or_or_B0_B1_o_or_B2__o , \sel3/or_or_B4_B5_o_or_B6__o );
  or \sel3/or_or_or_B18_B19_o_o  (\sel3/or_or_or_B18_B19_o_o_o , \sel3/or_or_B18_B19_o_or_B_o , \sel3/or_or_B22_B23_o_or_B_o );
  or \sel3/or_or_or_B27_B28_o_o  (\sel3/or_or_or_B27_B28_o_o_o , \sel3/or_or_B27_B28_o_or_B_o , \sel3/or_or_B31_B32_o_or_B_o );
  or \sel3/or_or_or_B9_B10_o_or  (\sel3/or_or_or_B9_B10_o_or_o , \sel3/or_or_B9_B10_o_or_B1_o , \sel3/or_or_B13_B14_o_or_B_o );
  or \sel3/or_or_or_or_B0_B1_o_  (\sel3/or_or_or_or_B0_B1_o__o , \sel3/or_or_or_B0_B1_o_or__o , \sel3/or_or_or_B9_B10_o_or_o );
  or \sel3/or_or_or_or_B18_B19_  (\sel3/or_or_or_or_B18_B19__o , \sel3/or_or_or_B18_B19_o_o_o , \sel3/or_or_or_B27_B28_o_o_o );
  or \sel3/or_or_or_or_or_B0_B1  (n188, \sel3/or_or_or_or_B0_B1_o__o , \sel3/or_or_or_or_B18_B19__o );
  and \sel4/and_b0_0  (\sel4/B0 , ready, n181);
  and \sel4/and_b0_1  (\sel4/B1 , n107, n180);
  and \sel4/and_b0_10  (\sel4/B10 , n107, n171);
  and \sel4/and_b0_11  (\sel4/B11 , n107, n170);
  and \sel4/and_b0_12  (\sel4/B12 , n107, n169);
  and \sel4/and_b0_13  (\sel4/B13 , n107, n168);
  and \sel4/and_b0_14  (\sel4/B14 , n107, n167);
  and \sel4/and_b0_15  (\sel4/B15 , n107, n166);
  and \sel4/and_b0_16  (\sel4/B16 , n107, n165);
  and \sel4/and_b0_17  (\sel4/B17 , n107, n164);
  and \sel4/and_b0_18  (\sel4/B18 , n107, n163);
  and \sel4/and_b0_19  (\sel4/B19 , n107, n162);
  and \sel4/and_b0_2  (\sel4/B2 , n113, n179);
  and \sel4/and_b0_20  (\sel4/B20 , n107, n161);
  and \sel4/and_b0_21  (\sel4/B21 , n107, n160);
  and \sel4/and_b0_22  (\sel4/B22 , n107, n159);
  and \sel4/and_b0_23  (\sel4/B23 , n107, n158);
  and \sel4/and_b0_24  (\sel4/B24 , n107, n157);
  and \sel4/and_b0_25  (\sel4/B25 , n107, n156);
  and \sel4/and_b0_26  (\sel4/B26 , n107, n155);
  and \sel4/and_b0_27  (\sel4/B27 , n107, n154);
  and \sel4/and_b0_28  (\sel4/B28 , n107, n153);
  and \sel4/and_b0_29  (\sel4/B29 , n107, n152);
  and \sel4/and_b0_3  (\sel4/B3 , n107, n178);
  and \sel4/and_b0_30  (\sel4/B30 , n107, n151);
  and \sel4/and_b0_31  (\sel4/B31 , n107, n150);
  and \sel4/and_b0_32  (\sel4/B32 , n107, n149);
  and \sel4/and_b0_33  (\sel4/B33 , n113, n148);
  and \sel4/and_b0_34  (\sel4/B34 , n107, n147);
  and \sel4/and_b0_4  (\sel4/B4 , n107, n177);
  and \sel4/and_b0_5  (\sel4/B5 , n107, n176);
  and \sel4/and_b0_6  (\sel4/B6 , n107, n175);
  and \sel4/and_b0_7  (\sel4/B7 , n107, n174);
  and \sel4/and_b0_8  (\sel4/B8 , n107, n173);
  and \sel4/and_b0_9  (\sel4/B9 , n107, n172);
  or \sel4/or_B0_B1  (\sel4/or_B0_B1_o , \sel4/B0 , \sel4/B1 );
  or \sel4/or_B11_B12  (\sel4/or_B11_B12_o , \sel4/B11 , \sel4/B12 );
  or \sel4/or_B13_B14  (\sel4/or_B13_B14_o , \sel4/B13 , \sel4/B14 );
  or \sel4/or_B15_or_B16_B17_o  (\sel4/or_B15_or_B16_B17_o_o , \sel4/B15 , \sel4/or_B16_B17_o );
  or \sel4/or_B16_B17  (\sel4/or_B16_B17_o , \sel4/B16 , \sel4/B17 );
  or \sel4/or_B18_B19  (\sel4/or_B18_B19_o , \sel4/B18 , \sel4/B19 );
  or \sel4/or_B20_B21  (\sel4/or_B20_B21_o , \sel4/B20 , \sel4/B21 );
  or \sel4/or_B22_B23  (\sel4/or_B22_B23_o , \sel4/B22 , \sel4/B23 );
  or \sel4/or_B24_or_B25_B26_o  (\sel4/or_B24_or_B25_B26_o_o , \sel4/B24 , \sel4/or_B25_B26_o );
  or \sel4/or_B25_B26  (\sel4/or_B25_B26_o , \sel4/B25 , \sel4/B26 );
  or \sel4/or_B27_B28  (\sel4/or_B27_B28_o , \sel4/B27 , \sel4/B28 );
  or \sel4/or_B29_B30  (\sel4/or_B29_B30_o , \sel4/B29 , \sel4/B30 );
  or \sel4/or_B2_B3  (\sel4/or_B2_B3_o , \sel4/B2 , \sel4/B3 );
  or \sel4/or_B31_B32  (\sel4/or_B31_B32_o , \sel4/B31 , \sel4/B32 );
  or \sel4/or_B33_or_B34_B35_o  (\sel4/or_B33_or_B34_B35_o_o , \sel4/B33 , \sel4/or_B34_B35_o );
  or \sel4/or_B34_B35  (\sel4/or_B34_B35_o , \sel4/B34 , n183);
  or \sel4/or_B4_B5  (\sel4/or_B4_B5_o , \sel4/B4 , \sel4/B5 );
  or \sel4/or_B6_or_B7_B8_o  (\sel4/or_B6_or_B7_B8_o_o , \sel4/B6 , \sel4/or_B7_B8_o );
  or \sel4/or_B7_B8  (\sel4/or_B7_B8_o , \sel4/B7 , \sel4/B8 );
  or \sel4/or_B9_B10  (\sel4/or_B9_B10_o , \sel4/B9 , \sel4/B10 );
  or \sel4/or_or_B0_B1_o_or_B2_  (\sel4/or_or_B0_B1_o_or_B2__o , \sel4/or_B0_B1_o , \sel4/or_B2_B3_o );
  or \sel4/or_or_B13_B14_o_or_B  (\sel4/or_or_B13_B14_o_or_B_o , \sel4/or_B13_B14_o , \sel4/or_B15_or_B16_B17_o_o );
  or \sel4/or_or_B18_B19_o_or_B  (\sel4/or_or_B18_B19_o_or_B_o , \sel4/or_B18_B19_o , \sel4/or_B20_B21_o );
  or \sel4/or_or_B22_B23_o_or_B  (\sel4/or_or_B22_B23_o_or_B_o , \sel4/or_B22_B23_o , \sel4/or_B24_or_B25_B26_o_o );
  or \sel4/or_or_B27_B28_o_or_B  (\sel4/or_or_B27_B28_o_or_B_o , \sel4/or_B27_B28_o , \sel4/or_B29_B30_o );
  or \sel4/or_or_B31_B32_o_or_B  (\sel4/or_or_B31_B32_o_or_B_o , \sel4/or_B31_B32_o , \sel4/or_B33_or_B34_B35_o_o );
  or \sel4/or_or_B4_B5_o_or_B6_  (\sel4/or_or_B4_B5_o_or_B6__o , \sel4/or_B4_B5_o , \sel4/or_B6_or_B7_B8_o_o );
  or \sel4/or_or_B9_B10_o_or_B1  (\sel4/or_or_B9_B10_o_or_B1_o , \sel4/or_B9_B10_o , \sel4/or_B11_B12_o );
  or \sel4/or_or_or_B0_B1_o_or_  (\sel4/or_or_or_B0_B1_o_or__o , \sel4/or_or_B0_B1_o_or_B2__o , \sel4/or_or_B4_B5_o_or_B6__o );
  or \sel4/or_or_or_B18_B19_o_o  (\sel4/or_or_or_B18_B19_o_o_o , \sel4/or_or_B18_B19_o_or_B_o , \sel4/or_or_B22_B23_o_or_B_o );
  or \sel4/or_or_or_B27_B28_o_o  (\sel4/or_or_or_B27_B28_o_o_o , \sel4/or_or_B27_B28_o_or_B_o , \sel4/or_or_B31_B32_o_or_B_o );
  or \sel4/or_or_or_B9_B10_o_or  (\sel4/or_or_or_B9_B10_o_or_o , \sel4/or_or_B9_B10_o_or_B1_o , \sel4/or_or_B13_B14_o_or_B_o );
  or \sel4/or_or_or_or_B0_B1_o_  (\sel4/or_or_or_or_B0_B1_o__o , \sel4/or_or_or_B0_B1_o_or__o , \sel4/or_or_or_B9_B10_o_or_o );
  or \sel4/or_or_or_or_B18_B19_  (\sel4/or_or_or_or_B18_B19__o , \sel4/or_or_or_B18_B19_o_o_o , \sel4/or_or_or_B27_B28_o_o_o );
  or \sel4/or_or_or_or_or_B0_B1  (n190, \sel4/or_or_or_or_B0_B1_o__o , \sel4/or_or_or_or_B18_B19__o );
  and \sel5/and_b0_0  (\sel5/B0 , success, n181);
  and \sel5/and_b0_1  (\sel5/B1 , n108, n180);
  and \sel5/and_b0_10  (\sel5/B10 , n108, n171);
  and \sel5/and_b0_11  (\sel5/B11 , n108, n170);
  and \sel5/and_b0_12  (\sel5/B12 , n108, n169);
  and \sel5/and_b0_13  (\sel5/B13 , n108, n168);
  and \sel5/and_b0_14  (\sel5/B14 , n108, n167);
  and \sel5/and_b0_15  (\sel5/B15 , n108, n166);
  and \sel5/and_b0_16  (\sel5/B16 , n108, n165);
  and \sel5/and_b0_17  (\sel5/B17 , n108, n164);
  and \sel5/and_b0_18  (\sel5/B18 , n108, n163);
  and \sel5/and_b0_19  (\sel5/B19 , n108, n162);
  and \sel5/and_b0_2  (\sel5/B2 , n114, n179);
  and \sel5/and_b0_20  (\sel5/B20 , n108, n161);
  and \sel5/and_b0_21  (\sel5/B21 , n108, n160);
  and \sel5/and_b0_22  (\sel5/B22 , n108, n159);
  and \sel5/and_b0_23  (\sel5/B23 , n108, n158);
  and \sel5/and_b0_24  (\sel5/B24 , n108, n157);
  and \sel5/and_b0_25  (\sel5/B25 , n108, n156);
  and \sel5/and_b0_26  (\sel5/B26 , n108, n155);
  and \sel5/and_b0_27  (\sel5/B27 , n108, n154);
  and \sel5/and_b0_28  (\sel5/B28 , n108, n153);
  and \sel5/and_b0_29  (\sel5/B29 , n108, n152);
  and \sel5/and_b0_3  (\sel5/B3 , n143, n178);
  and \sel5/and_b0_30  (\sel5/B30 , n108, n151);
  and \sel5/and_b0_31  (\sel5/B31 , n108, n150);
  and \sel5/and_b0_32  (\sel5/B32 , n108, n149);
  and \sel5/and_b0_33  (\sel5/B33 , n114, n148);
  and \sel5/and_b0_34  (\sel5/B34 , n108, n147);
  and \sel5/and_b0_4  (\sel5/B4 , n108, n177);
  and \sel5/and_b0_5  (\sel5/B5 , n108, n176);
  and \sel5/and_b0_6  (\sel5/B6 , n108, n175);
  and \sel5/and_b0_7  (\sel5/B7 , n108, n174);
  and \sel5/and_b0_8  (\sel5/B8 , n108, n173);
  and \sel5/and_b0_9  (\sel5/B9 , n108, n172);
  or \sel5/or_B0_B1  (\sel5/or_B0_B1_o , \sel5/B0 , \sel5/B1 );
  or \sel5/or_B11_B12  (\sel5/or_B11_B12_o , \sel5/B11 , \sel5/B12 );
  or \sel5/or_B13_B14  (\sel5/or_B13_B14_o , \sel5/B13 , \sel5/B14 );
  or \sel5/or_B15_or_B16_B17_o  (\sel5/or_B15_or_B16_B17_o_o , \sel5/B15 , \sel5/or_B16_B17_o );
  or \sel5/or_B16_B17  (\sel5/or_B16_B17_o , \sel5/B16 , \sel5/B17 );
  or \sel5/or_B18_B19  (\sel5/or_B18_B19_o , \sel5/B18 , \sel5/B19 );
  or \sel5/or_B20_B21  (\sel5/or_B20_B21_o , \sel5/B20 , \sel5/B21 );
  or \sel5/or_B22_B23  (\sel5/or_B22_B23_o , \sel5/B22 , \sel5/B23 );
  or \sel5/or_B24_or_B25_B26_o  (\sel5/or_B24_or_B25_B26_o_o , \sel5/B24 , \sel5/or_B25_B26_o );
  or \sel5/or_B25_B26  (\sel5/or_B25_B26_o , \sel5/B25 , \sel5/B26 );
  or \sel5/or_B27_B28  (\sel5/or_B27_B28_o , \sel5/B27 , \sel5/B28 );
  or \sel5/or_B29_B30  (\sel5/or_B29_B30_o , \sel5/B29 , \sel5/B30 );
  or \sel5/or_B2_B3  (\sel5/or_B2_B3_o , \sel5/B2 , \sel5/B3 );
  or \sel5/or_B31_B32  (\sel5/or_B31_B32_o , \sel5/B31 , \sel5/B32 );
  or \sel5/or_B33_or_B34_B35_o  (\sel5/or_B33_or_B34_B35_o_o , \sel5/B33 , \sel5/B34 );
  or \sel5/or_B4_B5  (\sel5/or_B4_B5_o , \sel5/B4 , \sel5/B5 );
  or \sel5/or_B6_or_B7_B8_o  (\sel5/or_B6_or_B7_B8_o_o , \sel5/B6 , \sel5/or_B7_B8_o );
  or \sel5/or_B7_B8  (\sel5/or_B7_B8_o , \sel5/B7 , \sel5/B8 );
  or \sel5/or_B9_B10  (\sel5/or_B9_B10_o , \sel5/B9 , \sel5/B10 );
  or \sel5/or_or_B0_B1_o_or_B2_  (\sel5/or_or_B0_B1_o_or_B2__o , \sel5/or_B0_B1_o , \sel5/or_B2_B3_o );
  or \sel5/or_or_B13_B14_o_or_B  (\sel5/or_or_B13_B14_o_or_B_o , \sel5/or_B13_B14_o , \sel5/or_B15_or_B16_B17_o_o );
  or \sel5/or_or_B18_B19_o_or_B  (\sel5/or_or_B18_B19_o_or_B_o , \sel5/or_B18_B19_o , \sel5/or_B20_B21_o );
  or \sel5/or_or_B22_B23_o_or_B  (\sel5/or_or_B22_B23_o_or_B_o , \sel5/or_B22_B23_o , \sel5/or_B24_or_B25_B26_o_o );
  or \sel5/or_or_B27_B28_o_or_B  (\sel5/or_or_B27_B28_o_or_B_o , \sel5/or_B27_B28_o , \sel5/or_B29_B30_o );
  or \sel5/or_or_B31_B32_o_or_B  (\sel5/or_or_B31_B32_o_or_B_o , \sel5/or_B31_B32_o , \sel5/or_B33_or_B34_B35_o_o );
  or \sel5/or_or_B4_B5_o_or_B6_  (\sel5/or_or_B4_B5_o_or_B6__o , \sel5/or_B4_B5_o , \sel5/or_B6_or_B7_B8_o_o );
  or \sel5/or_or_B9_B10_o_or_B1  (\sel5/or_or_B9_B10_o_or_B1_o , \sel5/or_B9_B10_o , \sel5/or_B11_B12_o );
  or \sel5/or_or_or_B0_B1_o_or_  (\sel5/or_or_or_B0_B1_o_or__o , \sel5/or_or_B0_B1_o_or_B2__o , \sel5/or_or_B4_B5_o_or_B6__o );
  or \sel5/or_or_or_B18_B19_o_o  (\sel5/or_or_or_B18_B19_o_o_o , \sel5/or_or_B18_B19_o_or_B_o , \sel5/or_or_B22_B23_o_or_B_o );
  or \sel5/or_or_or_B27_B28_o_o  (\sel5/or_or_or_B27_B28_o_o_o , \sel5/or_or_B27_B28_o_or_B_o , \sel5/or_or_B31_B32_o_or_B_o );
  or \sel5/or_or_or_B9_B10_o_or  (\sel5/or_or_or_B9_B10_o_or_o , \sel5/or_or_B9_B10_o_or_B1_o , \sel5/or_or_B13_B14_o_or_B_o );
  or \sel5/or_or_or_or_B0_B1_o_  (\sel5/or_or_or_or_B0_B1_o__o , \sel5/or_or_or_B0_B1_o_or__o , \sel5/or_or_or_B9_B10_o_or_o );
  or \sel5/or_or_or_or_B18_B19_  (\sel5/or_or_or_or_B18_B19__o , \sel5/or_or_or_B18_B19_o_o_o , \sel5/or_or_or_B27_B28_o_o_o );
  or \sel5/or_or_or_or_or_B0_B1  (n192, \sel5/or_or_or_or_B0_B1_o__o , \sel5/or_or_or_or_B18_B19__o );
  and \sel6/and_b0_0  (\sel6/B0 , scl_output_zero, n181);
  and \sel6/and_b0_1  (\sel6/B1 , n103, n180);
  and \sel6/and_b0_10  (\sel6/B10 , n103, n171);
  and \sel6/and_b0_11  (\sel6/B11 , n103, n170);
  and \sel6/and_b0_12  (\sel6/B12 , n103, n169);
  and \sel6/and_b0_13  (\sel6/B13 , n125, n168);
  and \sel6/and_b0_14  (\sel6/B14 , n103, n167);
  and \sel6/and_b0_15  (\sel6/B15 , n103, n166);
  and \sel6/and_b0_16  (\sel6/B16 , n103, n165);
  and \sel6/and_b0_17  (\sel6/B17 , n103, n164);
  and \sel6/and_b0_18  (\sel6/B18 , n103, n163);
  and \sel6/and_b0_19  (\sel6/B19 , n103, n162);
  and \sel6/and_b0_2  (\sel6/B2 , n144, n179);
  and \sel6/and_b0_20  (\sel6/B20 , n103, n161);
  and \sel6/and_b0_21  (\sel6/B21 , n103, n160);
  and \sel6/and_b0_22  (\sel6/B22 , n103, n159);
  and \sel6/and_b0_23  (\sel6/B23 , n125, n158);
  and \sel6/and_b0_24  (\sel6/B24 , n103, n157);
  and \sel6/and_b0_25  (\sel6/B25 , n103, n156);
  and \sel6/and_b0_26  (\sel6/B26 , n103, n155);
  and \sel6/and_b0_27  (\sel6/B27 , n103, n154);
  and \sel6/and_b0_28  (\sel6/B28 , n103, n153);
  and \sel6/and_b0_29  (\sel6/B29 , n103, n152);
  and \sel6/and_b0_3  (\sel6/B3 , n125, n178);
  and \sel6/and_b0_30  (\sel6/B30 , n103, n151);
  and \sel6/and_b0_31  (\sel6/B31 , n103, n150);
  and \sel6/and_b0_32  (\sel6/B32 , n103, n149);
  and \sel6/and_b0_33  (\sel6/B33 , n109, n148);
  and \sel6/and_b0_34  (\sel6/B34 , n103, n147);
  and \sel6/and_b0_4  (\sel6/B4 , n103, n177);
  and \sel6/and_b0_5  (\sel6/B5 , n103, n176);
  and \sel6/and_b0_6  (\sel6/B6 , n103, n175);
  and \sel6/and_b0_7  (\sel6/B7 , n103, n174);
  and \sel6/and_b0_8  (\sel6/B8 , n103, n173);
  and \sel6/and_b0_9  (\sel6/B9 , n103, n172);
  or \sel6/or_B0_B1  (\sel6/or_B0_B1_o , \sel6/B0 , \sel6/B1 );
  or \sel6/or_B11_B12  (\sel6/or_B11_B12_o , \sel6/B11 , \sel6/B12 );
  or \sel6/or_B13_B14  (\sel6/or_B13_B14_o , \sel6/B13 , \sel6/B14 );
  or \sel6/or_B15_or_B16_B17_o  (\sel6/or_B15_or_B16_B17_o_o , \sel6/B15 , \sel6/or_B16_B17_o );
  or \sel6/or_B16_B17  (\sel6/or_B16_B17_o , \sel6/B16 , \sel6/B17 );
  or \sel6/or_B18_B19  (\sel6/or_B18_B19_o , \sel6/B18 , \sel6/B19 );
  or \sel6/or_B20_B21  (\sel6/or_B20_B21_o , \sel6/B20 , \sel6/B21 );
  or \sel6/or_B22_B23  (\sel6/or_B22_B23_o , \sel6/B22 , \sel6/B23 );
  or \sel6/or_B24_or_B25_B26_o  (\sel6/or_B24_or_B25_B26_o_o , \sel6/B24 , \sel6/or_B25_B26_o );
  or \sel6/or_B25_B26  (\sel6/or_B25_B26_o , \sel6/B25 , \sel6/B26 );
  or \sel6/or_B27_B28  (\sel6/or_B27_B28_o , \sel6/B27 , \sel6/B28 );
  or \sel6/or_B29_B30  (\sel6/or_B29_B30_o , \sel6/B29 , \sel6/B30 );
  or \sel6/or_B2_B3  (\sel6/or_B2_B3_o , \sel6/B2 , \sel6/B3 );
  or \sel6/or_B31_B32  (\sel6/or_B31_B32_o , \sel6/B31 , \sel6/B32 );
  or \sel6/or_B33_or_B34_B35_o  (\sel6/or_B33_or_B34_B35_o_o , \sel6/B33 , \sel6/B34 );
  or \sel6/or_B4_B5  (\sel6/or_B4_B5_o , \sel6/B4 , \sel6/B5 );
  or \sel6/or_B6_or_B7_B8_o  (\sel6/or_B6_or_B7_B8_o_o , \sel6/B6 , \sel6/or_B7_B8_o );
  or \sel6/or_B7_B8  (\sel6/or_B7_B8_o , \sel6/B7 , \sel6/B8 );
  or \sel6/or_B9_B10  (\sel6/or_B9_B10_o , \sel6/B9 , \sel6/B10 );
  or \sel6/or_or_B0_B1_o_or_B2_  (\sel6/or_or_B0_B1_o_or_B2__o , \sel6/or_B0_B1_o , \sel6/or_B2_B3_o );
  or \sel6/or_or_B13_B14_o_or_B  (\sel6/or_or_B13_B14_o_or_B_o , \sel6/or_B13_B14_o , \sel6/or_B15_or_B16_B17_o_o );
  or \sel6/or_or_B18_B19_o_or_B  (\sel6/or_or_B18_B19_o_or_B_o , \sel6/or_B18_B19_o , \sel6/or_B20_B21_o );
  or \sel6/or_or_B22_B23_o_or_B  (\sel6/or_or_B22_B23_o_or_B_o , \sel6/or_B22_B23_o , \sel6/or_B24_or_B25_B26_o_o );
  or \sel6/or_or_B27_B28_o_or_B  (\sel6/or_or_B27_B28_o_or_B_o , \sel6/or_B27_B28_o , \sel6/or_B29_B30_o );
  or \sel6/or_or_B31_B32_o_or_B  (\sel6/or_or_B31_B32_o_or_B_o , \sel6/or_B31_B32_o , \sel6/or_B33_or_B34_B35_o_o );
  or \sel6/or_or_B4_B5_o_or_B6_  (\sel6/or_or_B4_B5_o_or_B6__o , \sel6/or_B4_B5_o , \sel6/or_B6_or_B7_B8_o_o );
  or \sel6/or_or_B9_B10_o_or_B1  (\sel6/or_or_B9_B10_o_or_B1_o , \sel6/or_B9_B10_o , \sel6/or_B11_B12_o );
  or \sel6/or_or_or_B0_B1_o_or_  (\sel6/or_or_or_B0_B1_o_or__o , \sel6/or_or_B0_B1_o_or_B2__o , \sel6/or_or_B4_B5_o_or_B6__o );
  or \sel6/or_or_or_B18_B19_o_o  (\sel6/or_or_or_B18_B19_o_o_o , \sel6/or_or_B18_B19_o_or_B_o , \sel6/or_or_B22_B23_o_or_B_o );
  or \sel6/or_or_or_B27_B28_o_o  (\sel6/or_or_or_B27_B28_o_o_o , \sel6/or_or_B27_B28_o_or_B_o , \sel6/or_or_B31_B32_o_or_B_o );
  or \sel6/or_or_or_B9_B10_o_or  (\sel6/or_or_or_B9_B10_o_or_o , \sel6/or_or_B9_B10_o_or_B1_o , \sel6/or_or_B13_B14_o_or_B_o );
  or \sel6/or_or_or_or_B0_B1_o_  (\sel6/or_or_or_or_B0_B1_o__o , \sel6/or_or_or_B0_B1_o_or__o , \sel6/or_or_or_B9_B10_o_or_o );
  or \sel6/or_or_or_or_B18_B19_  (\sel6/or_or_or_or_B18_B19__o , \sel6/or_or_or_B18_B19_o_o_o , \sel6/or_or_or_B27_B28_o_o_o );
  or \sel6/or_or_or_or_or_B0_B1  (n194, \sel6/or_or_or_or_B0_B1_o__o , \sel6/or_or_or_or_B18_B19__o );
  reg_ar_as_w1 success_out_reg (
    .clk(~divider2[7]),
    .d(n33),
    .en(n28),
    .reset(1'b0),
    .set(1'b0),
    .q(success_out));  // sources/rtl/i2c_module.v(167)
  reg_sr_as_w1 success_reg (
    .clk(~divider2[7]),
    .d(n192),
    .en(1'b1),
    .reset(~reset_n),
    .set(1'b0),
    .q(success));  // sources/rtl/i2c_module.v(1066)
  and u10 (n29, n27, n28);  // sources/rtl/i2c_module.v(147)
  and u12 (n31, n179, success);  // sources/rtl/i2c_module.v(160)
  AL_MUX u13 (
    .i0(success_out),
    .i1(1'b0),
    .sel(n147),
    .o(n32));  // sources/rtl/i2c_module.v(164)
  AL_MUX u14 (
    .i0(n32),
    .i1(1'b1),
    .sel(n31),
    .o(n33));  // sources/rtl/i2c_module.v(164)
  or u16 (n98, n181, n180);  // sources/rtl/i2c_module.v(1064)
  or u17 (n189, n177, n176);  // sources/rtl/i2c_module.v(1064)
  or u18 (n187, n174, n173);  // sources/rtl/i2c_module.v(1064)
  or u19 (n185, n175, n187);  // sources/rtl/i2c_module.v(1064)
  not u2 (n0, clk_div);  // sources/rtl/i2c_module.v(75)
  or u20 (n97, n189, n185);  // sources/rtl/i2c_module.v(1064)
  or u21 (n96, n191, n97);  // sources/rtl/i2c_module.v(1064)
  or u22 (n30, n172, n171);  // sources/rtl/i2c_module.v(1064)
  or u23 (n24, n170, n169);  // sources/rtl/i2c_module.v(1064)
  or u24 (n95, n30, n24);  // sources/rtl/i2c_module.v(1064)
  or u25 (n94, n168, n167);  // sources/rtl/i2c_module.v(1064)
  not u26 (n58[0], ack_ok);  // sources/rtl/i2c_module.v(381)
  or u27 (n93, n165, n164);  // sources/rtl/i2c_module.v(1064)
  or u28 (n92, n166, n93);  // sources/rtl/i2c_module.v(1064)
  or u29 (n91, n94, n92);  // sources/rtl/i2c_module.v(1064)
  or u30 (n90, n95, n91);  // sources/rtl/i2c_module.v(1064)
  or u31 (n89, n96, n90);  // sources/rtl/i2c_module.v(1064)
  or u32 (n88, n163, n162);  // sources/rtl/i2c_module.v(1064)
  or u33 (n87, n161, n160);  // sources/rtl/i2c_module.v(1064)
  or u34 (n22, n88, n87);  // sources/rtl/i2c_module.v(1064)
  or u35 (n86, n159, n158);  // sources/rtl/i2c_module.v(1064)
  or u36 (n85, n156, n155);  // sources/rtl/i2c_module.v(1064)
  or u37 (n84, n157, n85);  // sources/rtl/i2c_module.v(1064)
  or u38 (n83, n86, n84);  // sources/rtl/i2c_module.v(1064)
  or u39 (n82, n22, n83);  // sources/rtl/i2c_module.v(1064)
  not u4 (n18, scl_out);  // sources/rtl/i2c_module.v(127)
  or u40 (n81, n154, n153);  // sources/rtl/i2c_module.v(1064)
  or u41 (n80, n152, n151);  // sources/rtl/i2c_module.v(1064)
  or u42 (n79, n81, n80);  // sources/rtl/i2c_module.v(1064)
  or u43 (n78, n150, n149);  // sources/rtl/i2c_module.v(1064)
  or u44 (n21, n147, n146);  // sources/rtl/i2c_module.v(1064)
  or u45 (n77, n148, n21);  // sources/rtl/i2c_module.v(1064)
  or u46 (n76, n78, n77);  // sources/rtl/i2c_module.v(1064)
  or u47 (n75, n79, n76);  // sources/rtl/i2c_module.v(1064)
  or u48 (n193, n179, n178);  // sources/rtl/i2c_module.v(1064)
  or u49 (n74, n82, n75);  // sources/rtl/i2c_module.v(1064)
  AL_MUX u5 (
    .i0(n19),
    .i1(n18),
    .sel(n17),
    .o(n20));  // sources/rtl/i2c_module.v(135)
  or u50 (n191, n98, n193);  // sources/rtl/i2c_module.v(1064)
  not u51 (n102, reset_n);  // sources/rtl/i2c_module.v(514)
  AL_MUX u52 (
    .i0(scl_output_zero),
    .i1(1'b0),
    .sel(n36),
    .o(n103));  // sources/rtl/i2c_module.v(545)
  AL_MUX u53 (
    .i0(scl_output_enable),
    .i1(1'b0),
    .sel(n36),
    .o(n104));  // sources/rtl/i2c_module.v(545)
  AL_MUX u54 (
    .i0(sda_oe),
    .i1(1'b1),
    .sel(n36),
    .o(n105));  // sources/rtl/i2c_module.v(545)
  AL_MUX u55 (
    .i0(sda),
    .i1(1'b0),
    .sel(n36),
    .o(n106));  // sources/rtl/i2c_module.v(545)
  AL_MUX u56 (
    .i0(ready),
    .i1(1'b0),
    .sel(n36),
    .o(n107));  // sources/rtl/i2c_module.v(545)
  AL_MUX u57 (
    .i0(success),
    .i1(1'b0),
    .sel(n36),
    .o(n108));  // sources/rtl/i2c_module.v(545)
  AL_MUX u58 (
    .i0(scl_output_zero),
    .i1(1'b1),
    .sel(n28),
    .o(n109));  // sources/rtl/i2c_module.v(558)
  AL_MUX u59 (
    .i0(scl_output_enable),
    .i1(1'b0),
    .sel(n28),
    .o(n110));  // sources/rtl/i2c_module.v(558)
  or u6 (n23, n158, n168);  // sources/rtl/i2c_module.v(147)
  AL_MUX u60 (
    .i0(sda_oe),
    .i1(1'b1),
    .sel(n28),
    .o(n111));  // sources/rtl/i2c_module.v(558)
  AL_MUX u61 (
    .i0(sda),
    .i1(1'b0),
    .sel(n28),
    .o(n112));  // sources/rtl/i2c_module.v(558)
  AL_MUX u62 (
    .i0(ready),
    .i1(1'b0),
    .sel(n28),
    .o(n113));  // sources/rtl/i2c_module.v(558)
  AL_MUX u63 (
    .i0(success),
    .i1(1'b0),
    .sel(n28),
    .o(n114));  // sources/rtl/i2c_module.v(558)
  AL_MUX u64 (
    .i0(scl_output_enable),
    .i1(1'b1),
    .sel(n36),
    .o(n115));  // sources/rtl/i2c_module.v(571)
  AL_MUX u65 (
    .i0(sda),
    .i1(slave_address[7]),
    .sel(n36),
    .o(n116));  // sources/rtl/i2c_module.v(571)
  AL_MUX u66 (
    .i0(sda),
    .i1(slave_address[6]),
    .sel(n36),
    .o(n117));  // sources/rtl/i2c_module.v(584)
  AL_MUX u67 (
    .i0(sda),
    .i1(slave_address[5]),
    .sel(n36),
    .o(n118));  // sources/rtl/i2c_module.v(597)
  AL_MUX u68 (
    .i0(sda),
    .i1(slave_address[4]),
    .sel(n36),
    .o(n119));  // sources/rtl/i2c_module.v(610)
  AL_MUX u69 (
    .i0(sda),
    .i1(slave_address[3]),
    .sel(n36),
    .o(n120));  // sources/rtl/i2c_module.v(623)
  or u7 (n25, n23, n178);  // sources/rtl/i2c_module.v(147)
  AL_MUX u70 (
    .i0(sda),
    .i1(slave_address[2]),
    .sel(n36),
    .o(n121));  // sources/rtl/i2c_module.v(636)
  AL_MUX u71 (
    .i0(sda),
    .i1(slave_address[1]),
    .sel(n36),
    .o(n122));  // sources/rtl/i2c_module.v(649)
  AL_MUX u72 (
    .i0(sda),
    .i1(slave_address[0]),
    .sel(n36),
    .o(n123));  // sources/rtl/i2c_module.v(662)
  AL_MUX u73 (
    .i0(sda_oe),
    .i1(1'b0),
    .sel(n36),
    .o(n124));  // sources/rtl/i2c_module.v(675)
  AL_MUX u74 (
    .i0(scl_output_zero),
    .i1(1'b1),
    .sel(n36),
    .o(n125));  // sources/rtl/i2c_module.v(700)
  AL_MUX u75 (
    .i0(sda),
    .i1(slave_reg_address[7]),
    .sel(n36),
    .o(n126));  // sources/rtl/i2c_module.v(727)
  AL_MUX u76 (
    .i0(sda),
    .i1(slave_reg_address[6]),
    .sel(n36),
    .o(n127));  // sources/rtl/i2c_module.v(740)
  AL_MUX u77 (
    .i0(sda),
    .i1(slave_reg_address[5]),
    .sel(n36),
    .o(n128));  // sources/rtl/i2c_module.v(753)
  AL_MUX u78 (
    .i0(sda),
    .i1(slave_reg_address[4]),
    .sel(n36),
    .o(n129));  // sources/rtl/i2c_module.v(766)
  AL_MUX u79 (
    .i0(sda),
    .i1(slave_reg_address[3]),
    .sel(n36),
    .o(n130));  // sources/rtl/i2c_module.v(779)
  not u8 (n26, sda_in);  // sources/rtl/i2c_module.v(147)
  AL_MUX u80 (
    .i0(sda),
    .i1(slave_reg_address[2]),
    .sel(n36),
    .o(n131));  // sources/rtl/i2c_module.v(792)
  AL_MUX u81 (
    .i0(sda),
    .i1(slave_reg_address[1]),
    .sel(n36),
    .o(n132));  // sources/rtl/i2c_module.v(805)
  AL_MUX u82 (
    .i0(sda),
    .i1(slave_reg_address[0]),
    .sel(n36),
    .o(n133));  // sources/rtl/i2c_module.v(818)
  AL_MUX u83 (
    .i0(sda),
    .i1(slave_data_1[7]),
    .sel(n36),
    .o(n134));  // sources/rtl/i2c_module.v(878)
  AL_MUX u84 (
    .i0(sda),
    .i1(slave_data_1[6]),
    .sel(n36),
    .o(n135));  // sources/rtl/i2c_module.v(891)
  AL_MUX u85 (
    .i0(sda),
    .i1(slave_data_1[5]),
    .sel(n36),
    .o(n136));  // sources/rtl/i2c_module.v(904)
  AL_MUX u86 (
    .i0(sda),
    .i1(slave_data_1[4]),
    .sel(n36),
    .o(n137));  // sources/rtl/i2c_module.v(917)
  AL_MUX u87 (
    .i0(sda),
    .i1(slave_data_1[3]),
    .sel(n36),
    .o(n138));  // sources/rtl/i2c_module.v(930)
  AL_MUX u88 (
    .i0(sda),
    .i1(slave_data_1[2]),
    .sel(n36),
    .o(n139));  // sources/rtl/i2c_module.v(943)
  AL_MUX u89 (
    .i0(sda),
    .i1(slave_data_1[1]),
    .sel(n36),
    .o(n140));  // sources/rtl/i2c_module.v(956)
  and u9 (n27, n25, n26);  // sources/rtl/i2c_module.v(147)
  AL_MUX u90 (
    .i0(sda),
    .i1(slave_data_1[0]),
    .sel(n36),
    .o(n141));  // sources/rtl/i2c_module.v(969)
  AL_MUX u91 (
    .i0(scl_output_enable),
    .i1(ack_ok),
    .sel(n36),
    .o(n142));  // sources/rtl/i2c_module.v(1008)
  AL_MUX u92 (
    .i0(success),
    .i1(ack_ok),
    .sel(n36),
    .o(n143));  // sources/rtl/i2c_module.v(1008)
  AL_MUX u93 (
    .i0(scl_output_zero),
    .i1(1'b0),
    .sel(n28),
    .o(n144));  // sources/rtl/i2c_module.v(1030)
  AL_MUX u94 (
    .i0(sda),
    .i1(1'b1),
    .sel(n36),
    .o(n145));  // sources/rtl/i2c_module.v(1043)
  or u95 (n183, n146, n182);  // sources/rtl/i2c_module.v(1064)
  not u96 (n182, n73);  // sources/rtl/i2c_module.v(1064)
  or u97 (n73, n89, n74);  // sources/rtl/i2c_module.v(1064)

endmodule 

module add_pu11_pu11_o11
  (
  i0,
  i1,
  o
  );

  input [10:0] i0;
  input [10:0] i1;
  output [10:0] o;

  wire net_a0;
  wire net_a1;
  wire net_a10;
  wire net_a2;
  wire net_a3;
  wire net_a4;
  wire net_a5;
  wire net_a6;
  wire net_a7;
  wire net_a8;
  wire net_a9;
  wire net_b0;
  wire net_b1;
  wire net_b10;
  wire net_b2;
  wire net_b3;
  wire net_b4;
  wire net_b5;
  wire net_b6;
  wire net_b7;
  wire net_b8;
  wire net_b9;
  wire net_cout0;
  wire net_cout1;
  wire net_cout10;
  wire net_cout2;
  wire net_cout3;
  wire net_cout4;
  wire net_cout5;
  wire net_cout6;
  wire net_cout7;
  wire net_cout8;
  wire net_cout9;
  wire net_sum0;
  wire net_sum1;
  wire net_sum10;
  wire net_sum2;
  wire net_sum3;
  wire net_sum4;
  wire net_sum5;
  wire net_sum6;
  wire net_sum7;
  wire net_sum8;
  wire net_sum9;

  assign net_a10 = i0[10];
  assign net_a9 = i0[9];
  assign net_a8 = i0[8];
  assign net_a7 = i0[7];
  assign net_a6 = i0[6];
  assign net_a5 = i0[5];
  assign net_a4 = i0[4];
  assign net_a3 = i0[3];
  assign net_a2 = i0[2];
  assign net_a1 = i0[1];
  assign net_a0 = i0[0];
  assign net_b10 = i1[10];
  assign net_b9 = i1[9];
  assign net_b8 = i1[8];
  assign net_b7 = i1[7];
  assign net_b6 = i1[6];
  assign net_b5 = i1[5];
  assign net_b4 = i1[4];
  assign net_b3 = i1[3];
  assign net_b2 = i1[2];
  assign net_b1 = i1[1];
  assign net_b0 = i1[0];
  assign o[10] = net_sum10;
  assign o[9] = net_sum9;
  assign o[8] = net_sum8;
  assign o[7] = net_sum7;
  assign o[6] = net_sum6;
  assign o[5] = net_sum5;
  assign o[4] = net_sum4;
  assign o[3] = net_sum3;
  assign o[2] = net_sum2;
  assign o[1] = net_sum1;
  assign o[0] = net_sum0;
  AL_FADD comp_0 (
    .a(net_a0),
    .b(net_b0),
    .c(1'b0),
    .cout(net_cout0),
    .sum(net_sum0));
  AL_FADD comp_1 (
    .a(net_a1),
    .b(net_b1),
    .c(net_cout0),
    .cout(net_cout1),
    .sum(net_sum1));
  AL_FADD comp_10 (
    .a(net_a10),
    .b(net_b10),
    .c(net_cout9),
    .cout(net_cout10),
    .sum(net_sum10));
  AL_FADD comp_2 (
    .a(net_a2),
    .b(net_b2),
    .c(net_cout1),
    .cout(net_cout2),
    .sum(net_sum2));
  AL_FADD comp_3 (
    .a(net_a3),
    .b(net_b3),
    .c(net_cout2),
    .cout(net_cout3),
    .sum(net_sum3));
  AL_FADD comp_4 (
    .a(net_a4),
    .b(net_b4),
    .c(net_cout3),
    .cout(net_cout4),
    .sum(net_sum4));
  AL_FADD comp_5 (
    .a(net_a5),
    .b(net_b5),
    .c(net_cout4),
    .cout(net_cout5),
    .sum(net_sum5));
  AL_FADD comp_6 (
    .a(net_a6),
    .b(net_b6),
    .c(net_cout5),
    .cout(net_cout6),
    .sum(net_sum6));
  AL_FADD comp_7 (
    .a(net_a7),
    .b(net_b7),
    .c(net_cout6),
    .cout(net_cout7),
    .sum(net_sum7));
  AL_FADD comp_8 (
    .a(net_a8),
    .b(net_b8),
    .c(net_cout7),
    .cout(net_cout8),
    .sum(net_sum8));
  AL_FADD comp_9 (
    .a(net_a9),
    .b(net_b9),
    .c(net_cout8),
    .cout(net_cout9),
    .sum(net_sum9));

endmodule 

module eq_w11
  (
  i0,
  i1,
  o
  );

  input [10:0] i0;
  input [10:0] i1;
  output o;

  wire \or_or_or_xor_i0[0]_i_o ;
  wire \or_or_xor_i0[0]_i1[0_o ;
  wire \or_or_xor_i0[5]_i1[5_o ;
  wire \or_xor_i0[0]_i1[0]_o_o ;
  wire \or_xor_i0[2]_i1[2]_o_o ;
  wire \or_xor_i0[3]_i1[3]_o_o ;
  wire \or_xor_i0[5]_i1[5]_o_o ;
  wire \or_xor_i0[6]_i1[6]_o_o ;
  wire \or_xor_i0[8]_i1[8]_o_o ;
  wire \or_xor_i0[9]_i1[9]_o_o ;
  wire \xor_i0[0]_i1[0]_o ;
  wire \xor_i0[10]_i1[10]_o ;
  wire \xor_i0[1]_i1[1]_o ;
  wire \xor_i0[2]_i1[2]_o ;
  wire \xor_i0[3]_i1[3]_o ;
  wire \xor_i0[4]_i1[4]_o ;
  wire \xor_i0[5]_i1[5]_o ;
  wire \xor_i0[6]_i1[6]_o ;
  wire \xor_i0[7]_i1[7]_o ;
  wire \xor_i0[8]_i1[8]_o ;
  wire \xor_i0[9]_i1[9]_o ;

  not none_diff (o, \or_or_or_xor_i0[0]_i_o );
  or \or_or_or_xor_i0[0]_i  (\or_or_or_xor_i0[0]_i_o , \or_or_xor_i0[0]_i1[0_o , \or_or_xor_i0[5]_i1[5_o );
  or \or_or_xor_i0[0]_i1[0  (\or_or_xor_i0[0]_i1[0_o , \or_xor_i0[0]_i1[0]_o_o , \or_xor_i0[2]_i1[2]_o_o );
  or \or_or_xor_i0[5]_i1[5  (\or_or_xor_i0[5]_i1[5_o , \or_xor_i0[5]_i1[5]_o_o , \or_xor_i0[8]_i1[8]_o_o );
  or \or_xor_i0[0]_i1[0]_o  (\or_xor_i0[0]_i1[0]_o_o , \xor_i0[0]_i1[0]_o , \xor_i0[1]_i1[1]_o );
  or \or_xor_i0[2]_i1[2]_o  (\or_xor_i0[2]_i1[2]_o_o , \xor_i0[2]_i1[2]_o , \or_xor_i0[3]_i1[3]_o_o );
  or \or_xor_i0[3]_i1[3]_o  (\or_xor_i0[3]_i1[3]_o_o , \xor_i0[3]_i1[3]_o , \xor_i0[4]_i1[4]_o );
  or \or_xor_i0[5]_i1[5]_o  (\or_xor_i0[5]_i1[5]_o_o , \xor_i0[5]_i1[5]_o , \or_xor_i0[6]_i1[6]_o_o );
  or \or_xor_i0[6]_i1[6]_o  (\or_xor_i0[6]_i1[6]_o_o , \xor_i0[6]_i1[6]_o , \xor_i0[7]_i1[7]_o );
  or \or_xor_i0[8]_i1[8]_o  (\or_xor_i0[8]_i1[8]_o_o , \xor_i0[8]_i1[8]_o , \or_xor_i0[9]_i1[9]_o_o );
  or \or_xor_i0[9]_i1[9]_o  (\or_xor_i0[9]_i1[9]_o_o , \xor_i0[9]_i1[9]_o , \xor_i0[10]_i1[10]_o );
  xor \xor_i0[0]_i1[0]  (\xor_i0[0]_i1[0]_o , i0[0], i1[0]);
  xor \xor_i0[10]_i1[10]  (\xor_i0[10]_i1[10]_o , i0[10], i1[10]);
  xor \xor_i0[1]_i1[1]  (\xor_i0[1]_i1[1]_o , i0[1], i1[1]);
  xor \xor_i0[2]_i1[2]  (\xor_i0[2]_i1[2]_o , i0[2], i1[2]);
  xor \xor_i0[3]_i1[3]  (\xor_i0[3]_i1[3]_o , i0[3], i1[3]);
  xor \xor_i0[4]_i1[4]  (\xor_i0[4]_i1[4]_o , i0[4], i1[4]);
  xor \xor_i0[5]_i1[5]  (\xor_i0[5]_i1[5]_o , i0[5], i1[5]);
  xor \xor_i0[6]_i1[6]  (\xor_i0[6]_i1[6]_o , i0[6], i1[6]);
  xor \xor_i0[7]_i1[7]  (\xor_i0[7]_i1[7]_o , i0[7], i1[7]);
  xor \xor_i0[8]_i1[8]  (\xor_i0[8]_i1[8]_o , i0[8], i1[8]);
  xor \xor_i0[9]_i1[9]  (\xor_i0[9]_i1[9]_o , i0[9], i1[9]);

endmodule 

module lt_u11_u11
  (
  ci,
  i0,
  i1,
  o
  );

  input ci;
  input [10:0] i0;
  input [10:0] i1;
  output o;

  wire [10:0] diff;
  wire diff_6_10;
  wire less_6_10;
  wire \less_6_10_inst/diff_0 ;
  wire \less_6_10_inst/diff_1 ;
  wire \less_6_10_inst/diff_2 ;
  wire \less_6_10_inst/diff_3 ;
  wire \less_6_10_inst/diff_4 ;
  wire \less_6_10_inst/o_0 ;
  wire \less_6_10_inst/o_1 ;
  wire \less_6_10_inst/o_2 ;
  wire \less_6_10_inst/o_3 ;
  wire o_0;
  wire o_1;
  wire o_2;
  wire o_3;
  wire o_4;
  wire o_5;

  or any_diff_6_10 (diff_6_10, diff[6], diff[7], diff[8], diff[9], diff[10]);
  xor diff_0 (diff[0], i0[0], i1[0]);
  xor diff_1 (diff[1], i0[1], i1[1]);
  xor diff_10 (diff[10], i0[10], i1[10]);
  xor diff_2 (diff[2], i0[2], i1[2]);
  xor diff_3 (diff[3], i0[3], i1[3]);
  xor diff_4 (diff[4], i0[4], i1[4]);
  xor diff_5 (diff[5], i0[5], i1[5]);
  xor diff_6 (diff[6], i0[6], i1[6]);
  xor diff_7 (diff[7], i0[7], i1[7]);
  xor diff_8 (diff[8], i0[8], i1[8]);
  xor diff_9 (diff[9], i0[9], i1[9]);
  AL_MUX \less_6_10_inst/mux_0  (
    .i0(1'b0),
    .i1(i1[6]),
    .sel(\less_6_10_inst/diff_0 ),
    .o(\less_6_10_inst/o_0 ));
  AL_MUX \less_6_10_inst/mux_1  (
    .i0(\less_6_10_inst/o_0 ),
    .i1(i1[7]),
    .sel(\less_6_10_inst/diff_1 ),
    .o(\less_6_10_inst/o_1 ));
  AL_MUX \less_6_10_inst/mux_2  (
    .i0(\less_6_10_inst/o_1 ),
    .i1(i1[8]),
    .sel(\less_6_10_inst/diff_2 ),
    .o(\less_6_10_inst/o_2 ));
  AL_MUX \less_6_10_inst/mux_3  (
    .i0(\less_6_10_inst/o_2 ),
    .i1(i1[9]),
    .sel(\less_6_10_inst/diff_3 ),
    .o(\less_6_10_inst/o_3 ));
  AL_MUX \less_6_10_inst/mux_4  (
    .i0(\less_6_10_inst/o_3 ),
    .i1(i1[10]),
    .sel(\less_6_10_inst/diff_4 ),
    .o(less_6_10));
  xor \less_6_10_inst/xor_0  (\less_6_10_inst/diff_0 , i0[6], i1[6]);
  xor \less_6_10_inst/xor_1  (\less_6_10_inst/diff_1 , i0[7], i1[7]);
  xor \less_6_10_inst/xor_2  (\less_6_10_inst/diff_2 , i0[8], i1[8]);
  xor \less_6_10_inst/xor_3  (\less_6_10_inst/diff_3 , i0[9], i1[9]);
  xor \less_6_10_inst/xor_4  (\less_6_10_inst/diff_4 , i0[10], i1[10]);
  AL_MUX mux_0 (
    .i0(ci),
    .i1(i1[0]),
    .sel(diff[0]),
    .o(o_0));
  AL_MUX mux_1 (
    .i0(o_0),
    .i1(i1[1]),
    .sel(diff[1]),
    .o(o_1));
  AL_MUX mux_2 (
    .i0(o_1),
    .i1(i1[2]),
    .sel(diff[2]),
    .o(o_2));
  AL_MUX mux_3 (
    .i0(o_2),
    .i1(i1[3]),
    .sel(diff[3]),
    .o(o_3));
  AL_MUX mux_4 (
    .i0(o_3),
    .i1(i1[4]),
    .sel(diff[4]),
    .o(o_4));
  AL_MUX mux_5 (
    .i0(o_4),
    .i1(i1[5]),
    .sel(diff[5]),
    .o(o_5));
  AL_MUX mux_6 (
    .i0(o_5),
    .i1(less_6_10),
    .sel(diff_6_10),
    .o(o));

endmodule 

module lt_u12_u12
  (
  ci,
  i0,
  i1,
  o
  );

  input ci;
  input [11:0] i0;
  input [11:0] i1;
  output o;

  wire [11:0] diff;
  wire diff_6_11;
  wire less_6_11;
  wire \less_6_11_inst/diff_0 ;
  wire \less_6_11_inst/diff_1 ;
  wire \less_6_11_inst/diff_2 ;
  wire \less_6_11_inst/diff_3 ;
  wire \less_6_11_inst/diff_4 ;
  wire \less_6_11_inst/diff_5 ;
  wire \less_6_11_inst/o_0 ;
  wire \less_6_11_inst/o_1 ;
  wire \less_6_11_inst/o_2 ;
  wire \less_6_11_inst/o_3 ;
  wire \less_6_11_inst/o_4 ;
  wire o_0;
  wire o_1;
  wire o_2;
  wire o_3;
  wire o_4;
  wire o_5;

  or any_diff_6_11 (diff_6_11, diff[6], diff[7], diff[8], diff[9], diff[10], diff[11]);
  xor diff_0 (diff[0], i0[0], i1[0]);
  xor diff_1 (diff[1], i0[1], i1[1]);
  xor diff_10 (diff[10], i0[10], i1[10]);
  xor diff_11 (diff[11], i0[11], i1[11]);
  xor diff_2 (diff[2], i0[2], i1[2]);
  xor diff_3 (diff[3], i0[3], i1[3]);
  xor diff_4 (diff[4], i0[4], i1[4]);
  xor diff_5 (diff[5], i0[5], i1[5]);
  xor diff_6 (diff[6], i0[6], i1[6]);
  xor diff_7 (diff[7], i0[7], i1[7]);
  xor diff_8 (diff[8], i0[8], i1[8]);
  xor diff_9 (diff[9], i0[9], i1[9]);
  AL_MUX \less_6_11_inst/mux_0  (
    .i0(1'b0),
    .i1(i1[6]),
    .sel(\less_6_11_inst/diff_0 ),
    .o(\less_6_11_inst/o_0 ));
  AL_MUX \less_6_11_inst/mux_1  (
    .i0(\less_6_11_inst/o_0 ),
    .i1(i1[7]),
    .sel(\less_6_11_inst/diff_1 ),
    .o(\less_6_11_inst/o_1 ));
  AL_MUX \less_6_11_inst/mux_2  (
    .i0(\less_6_11_inst/o_1 ),
    .i1(i1[8]),
    .sel(\less_6_11_inst/diff_2 ),
    .o(\less_6_11_inst/o_2 ));
  AL_MUX \less_6_11_inst/mux_3  (
    .i0(\less_6_11_inst/o_2 ),
    .i1(i1[9]),
    .sel(\less_6_11_inst/diff_3 ),
    .o(\less_6_11_inst/o_3 ));
  AL_MUX \less_6_11_inst/mux_4  (
    .i0(\less_6_11_inst/o_3 ),
    .i1(i1[10]),
    .sel(\less_6_11_inst/diff_4 ),
    .o(\less_6_11_inst/o_4 ));
  AL_MUX \less_6_11_inst/mux_5  (
    .i0(\less_6_11_inst/o_4 ),
    .i1(i1[11]),
    .sel(\less_6_11_inst/diff_5 ),
    .o(less_6_11));
  xor \less_6_11_inst/xor_0  (\less_6_11_inst/diff_0 , i0[6], i1[6]);
  xor \less_6_11_inst/xor_1  (\less_6_11_inst/diff_1 , i0[7], i1[7]);
  xor \less_6_11_inst/xor_2  (\less_6_11_inst/diff_2 , i0[8], i1[8]);
  xor \less_6_11_inst/xor_3  (\less_6_11_inst/diff_3 , i0[9], i1[9]);
  xor \less_6_11_inst/xor_4  (\less_6_11_inst/diff_4 , i0[10], i1[10]);
  xor \less_6_11_inst/xor_5  (\less_6_11_inst/diff_5 , i0[11], i1[11]);
  AL_MUX mux_0 (
    .i0(ci),
    .i1(i1[0]),
    .sel(diff[0]),
    .o(o_0));
  AL_MUX mux_1 (
    .i0(o_0),
    .i1(i1[1]),
    .sel(diff[1]),
    .o(o_1));
  AL_MUX mux_2 (
    .i0(o_1),
    .i1(i1[2]),
    .sel(diff[2]),
    .o(o_2));
  AL_MUX mux_3 (
    .i0(o_2),
    .i1(i1[3]),
    .sel(diff[3]),
    .o(o_3));
  AL_MUX mux_4 (
    .i0(o_3),
    .i1(i1[4]),
    .sel(diff[4]),
    .o(o_4));
  AL_MUX mux_5 (
    .i0(o_4),
    .i1(i1[5]),
    .sel(diff[5]),
    .o(o_5));
  AL_MUX mux_6 (
    .i0(o_5),
    .i1(less_6_11),
    .sel(diff_6_11),
    .o(o));

endmodule 

module mult_u13_u5_o13
  (
  i0,
  i1,
  o
  );

  input [12:0] i0;
  input [4:0] i1;
  output [12:0] o;

  wire a0;
  wire a1;
  wire a10;
  wire a11;
  wire a12;
  wire a2;
  wire a3;
  wire a4;
  wire a5;
  wire a6;
  wire a7;
  wire a8;
  wire a9;
  wire b0;
  wire b1;
  wire b2;
  wire b3;
  wire b4;
  wire net_and_a0_b0;
  wire net_and_a0_b1;
  wire net_and_a0_b2;
  wire net_and_a0_b3;
  wire net_and_a0_b4;
  wire net_and_a10_b0;
  wire net_and_a10_b1;
  wire net_and_a10_b2;
  wire net_and_a11_b0;
  wire net_and_a11_b1;
  wire net_and_a12_b0;
  wire net_and_a1_b0;
  wire net_and_a1_b1;
  wire net_and_a1_b2;
  wire net_and_a1_b3;
  wire net_and_a1_b4;
  wire net_and_a2_b0;
  wire net_and_a2_b1;
  wire net_and_a2_b2;
  wire net_and_a2_b3;
  wire net_and_a2_b4;
  wire net_and_a3_b0;
  wire net_and_a3_b1;
  wire net_and_a3_b2;
  wire net_and_a3_b3;
  wire net_and_a3_b4;
  wire net_and_a4_b0;
  wire net_and_a4_b1;
  wire net_and_a4_b2;
  wire net_and_a4_b3;
  wire net_and_a4_b4;
  wire net_and_a5_b0;
  wire net_and_a5_b1;
  wire net_and_a5_b2;
  wire net_and_a5_b3;
  wire net_and_a5_b4;
  wire net_and_a6_b0;
  wire net_and_a6_b1;
  wire net_and_a6_b2;
  wire net_and_a6_b3;
  wire net_and_a6_b4;
  wire net_and_a7_b0;
  wire net_and_a7_b1;
  wire net_and_a7_b2;
  wire net_and_a7_b3;
  wire net_and_a7_b4;
  wire net_and_a8_b0;
  wire net_and_a8_b1;
  wire net_and_a8_b2;
  wire net_and_a8_b3;
  wire net_and_a8_b4;
  wire net_and_a9_b0;
  wire net_and_a9_b1;
  wire net_and_a9_b2;
  wire net_and_a9_b3;
  wire o_0;
  wire o_1;
  wire o_10;
  wire o_11;
  wire o_12;
  wire o_2;
  wire o_3;
  wire o_4;
  wire o_5;
  wire o_6;
  wire o_7;
  wire o_8;
  wire o_9;

  assign a12 = i0[12];
  assign a11 = i0[11];
  assign a10 = i0[10];
  assign a9 = i0[9];
  assign a8 = i0[8];
  assign a7 = i0[7];
  assign a6 = i0[6];
  assign a5 = i0[5];
  assign a4 = i0[4];
  assign a3 = i0[3];
  assign a2 = i0[2];
  assign a1 = i0[1];
  assign a0 = i0[0];
  assign b4 = i1[4];
  assign b3 = i1[3];
  assign b2 = i1[2];
  assign b1 = i1[1];
  assign b0 = i1[0];
  assign o[12] = o_12;
  assign o[11] = o_11;
  assign o[10] = o_10;
  assign o[9] = o_9;
  assign o[8] = o_8;
  assign o[7] = o_7;
  assign o[6] = o_6;
  assign o[5] = o_5;
  assign o[4] = o_4;
  assign o[3] = o_3;
  assign o[2] = o_2;
  assign o[1] = o_1;
  assign o[0] = o_0;
  and and_a0_b0 (net_and_a0_b0, a0, b0);
  and and_a0_b1 (net_and_a0_b1, a0, b1);
  and and_a0_b2 (net_and_a0_b2, a0, b2);
  and and_a0_b3 (net_and_a0_b3, a0, b3);
  and and_a0_b4 (net_and_a0_b4, a0, b4);
  and and_a10_b0 (net_and_a10_b0, a10, b0);
  and and_a10_b1 (net_and_a10_b1, a10, b1);
  and and_a10_b2 (net_and_a10_b2, a10, b2);
  and and_a11_b0 (net_and_a11_b0, a11, b0);
  and and_a11_b1 (net_and_a11_b1, a11, b1);
  and and_a12_b0 (net_and_a12_b0, a12, b0);
  and and_a1_b0 (net_and_a1_b0, a1, b0);
  and and_a1_b1 (net_and_a1_b1, a1, b1);
  and and_a1_b2 (net_and_a1_b2, a1, b2);
  and and_a1_b3 (net_and_a1_b3, a1, b3);
  and and_a1_b4 (net_and_a1_b4, a1, b4);
  and and_a2_b0 (net_and_a2_b0, a2, b0);
  and and_a2_b1 (net_and_a2_b1, a2, b1);
  and and_a2_b2 (net_and_a2_b2, a2, b2);
  and and_a2_b3 (net_and_a2_b3, a2, b3);
  and and_a2_b4 (net_and_a2_b4, a2, b4);
  and and_a3_b0 (net_and_a3_b0, a3, b0);
  and and_a3_b1 (net_and_a3_b1, a3, b1);
  and and_a3_b2 (net_and_a3_b2, a3, b2);
  and and_a3_b3 (net_and_a3_b3, a3, b3);
  and and_a3_b4 (net_and_a3_b4, a3, b4);
  and and_a4_b0 (net_and_a4_b0, a4, b0);
  and and_a4_b1 (net_and_a4_b1, a4, b1);
  and and_a4_b2 (net_and_a4_b2, a4, b2);
  and and_a4_b3 (net_and_a4_b3, a4, b3);
  and and_a4_b4 (net_and_a4_b4, a4, b4);
  and and_a5_b0 (net_and_a5_b0, a5, b0);
  and and_a5_b1 (net_and_a5_b1, a5, b1);
  and and_a5_b2 (net_and_a5_b2, a5, b2);
  and and_a5_b3 (net_and_a5_b3, a5, b3);
  and and_a5_b4 (net_and_a5_b4, a5, b4);
  and and_a6_b0 (net_and_a6_b0, a6, b0);
  and and_a6_b1 (net_and_a6_b1, a6, b1);
  and and_a6_b2 (net_and_a6_b2, a6, b2);
  and and_a6_b3 (net_and_a6_b3, a6, b3);
  and and_a6_b4 (net_and_a6_b4, a6, b4);
  and and_a7_b0 (net_and_a7_b0, a7, b0);
  and and_a7_b1 (net_and_a7_b1, a7, b1);
  and and_a7_b2 (net_and_a7_b2, a7, b2);
  and and_a7_b3 (net_and_a7_b3, a7, b3);
  and and_a7_b4 (net_and_a7_b4, a7, b4);
  and and_a8_b0 (net_and_a8_b0, a8, b0);
  and and_a8_b1 (net_and_a8_b1, a8, b1);
  and and_a8_b2 (net_and_a8_b2, a8, b2);
  and and_a8_b3 (net_and_a8_b3, a8, b3);
  and and_a8_b4 (net_and_a8_b4, a8, b4);
  and and_a9_b0 (net_and_a9_b0, a9, b0);
  and and_a9_b1 (net_and_a9_b1, a9, b1);
  and and_a9_b2 (net_and_a9_b2, a9, b2);
  and and_a9_b3 (net_and_a9_b3, a9, b3);
  add_pu13_pu13_pu13_pu13_pu13_o13 sum (
    .i0({net_and_a12_b0,net_and_a11_b0,net_and_a10_b0,net_and_a9_b0,net_and_a8_b0,net_and_a7_b0,net_and_a6_b0,net_and_a5_b0,net_and_a4_b0,net_and_a3_b0,net_and_a2_b0,net_and_a1_b0,net_and_a0_b0}),
    .i1({net_and_a11_b1,net_and_a10_b1,net_and_a9_b1,net_and_a8_b1,net_and_a7_b1,net_and_a6_b1,net_and_a5_b1,net_and_a4_b1,net_and_a3_b1,net_and_a2_b1,net_and_a1_b1,net_and_a0_b1,1'b0}),
    .i2({net_and_a10_b2,net_and_a9_b2,net_and_a8_b2,net_and_a7_b2,net_and_a6_b2,net_and_a5_b2,net_and_a4_b2,net_and_a3_b2,net_and_a2_b2,net_and_a1_b2,net_and_a0_b2,2'b00}),
    .i3({net_and_a9_b3,net_and_a8_b3,net_and_a7_b3,net_and_a6_b3,net_and_a5_b3,net_and_a4_b3,net_and_a3_b3,net_and_a2_b3,net_and_a1_b3,net_and_a0_b3,3'b000}),
    .i4({net_and_a8_b4,net_and_a7_b4,net_and_a6_b4,net_and_a5_b4,net_and_a4_b4,net_and_a3_b4,net_and_a2_b4,net_and_a1_b4,net_and_a0_b4,4'b0000}),
    .o({o_12,o_11,o_10,o_9,o_8,o_7,o_6,o_5,o_4,o_3,o_2,o_1,o_0}));

endmodule 

module ne_w11
  (
  i0,
  i1,
  o
  );

  input [10:0] i0;
  input [10:0] i1;
  output o;

  wire [10:0] diff;

  or any_diff (o, diff[0], diff[1], diff[2], diff[3], diff[4], diff[5], diff[6], diff[7], diff[8], diff[9], diff[10]);
  xor diff_0 (diff[0], i0[0], i1[0]);
  xor diff_1 (diff[1], i0[1], i1[1]);
  xor diff_10 (diff[10], i0[10], i1[10]);
  xor diff_2 (diff[2], i0[2], i1[2]);
  xor diff_3 (diff[3], i0[3], i1[3]);
  xor diff_4 (diff[4], i0[4], i1[4]);
  xor diff_5 (diff[5], i0[5], i1[5]);
  xor diff_6 (diff[6], i0[6], i1[6]);
  xor diff_7 (diff[7], i0[7], i1[7]);
  xor diff_8 (diff[8], i0[8], i1[8]);
  xor diff_9 (diff[9], i0[9], i1[9]);

endmodule 

module add_pu11_mu11_o12
  (
  i0,
  i1,
  o
  );

  input [10:0] i0;
  input [10:0] i1;
  output [11:0] o;

  wire net_a0;
  wire net_a1;
  wire net_a10;
  wire net_a2;
  wire net_a3;
  wire net_a4;
  wire net_a5;
  wire net_a6;
  wire net_a7;
  wire net_a8;
  wire net_a9;
  wire net_b0;
  wire net_b1;
  wire net_b10;
  wire net_b2;
  wire net_b3;
  wire net_b4;
  wire net_b5;
  wire net_b6;
  wire net_b7;
  wire net_b8;
  wire net_b9;
  wire net_cout0;
  wire net_cout1;
  wire net_cout10;
  wire net_cout2;
  wire net_cout3;
  wire net_cout4;
  wire net_cout5;
  wire net_cout6;
  wire net_cout7;
  wire net_cout8;
  wire net_cout9;
  wire net_nb0;
  wire net_nb1;
  wire net_nb10;
  wire net_nb2;
  wire net_nb3;
  wire net_nb4;
  wire net_nb5;
  wire net_nb6;
  wire net_nb7;
  wire net_nb8;
  wire net_nb9;
  wire net_ncout;
  wire net_sum0;
  wire net_sum1;
  wire net_sum10;
  wire net_sum2;
  wire net_sum3;
  wire net_sum4;
  wire net_sum5;
  wire net_sum6;
  wire net_sum7;
  wire net_sum8;
  wire net_sum9;

  assign net_a10 = i0[10];
  assign net_a9 = i0[9];
  assign net_a8 = i0[8];
  assign net_a7 = i0[7];
  assign net_a6 = i0[6];
  assign net_a5 = i0[5];
  assign net_a4 = i0[4];
  assign net_a3 = i0[3];
  assign net_a2 = i0[2];
  assign net_a1 = i0[1];
  assign net_a0 = i0[0];
  assign net_b10 = i1[10];
  assign net_b9 = i1[9];
  assign net_b8 = i1[8];
  assign net_b7 = i1[7];
  assign net_b6 = i1[6];
  assign net_b5 = i1[5];
  assign net_b4 = i1[4];
  assign net_b3 = i1[3];
  assign net_b2 = i1[2];
  assign net_b1 = i1[1];
  assign net_b0 = i1[0];
  assign o[11] = net_ncout;
  assign o[10] = net_sum10;
  assign o[9] = net_sum9;
  assign o[8] = net_sum8;
  assign o[7] = net_sum7;
  assign o[6] = net_sum6;
  assign o[5] = net_sum5;
  assign o[4] = net_sum4;
  assign o[3] = net_sum3;
  assign o[2] = net_sum2;
  assign o[1] = net_sum1;
  assign o[0] = net_sum0;
  AL_FADD comp_0 (
    .a(net_a0),
    .b(net_nb0),
    .c(1'b1),
    .cout(net_cout0),
    .sum(net_sum0));
  AL_FADD comp_1 (
    .a(net_a1),
    .b(net_nb1),
    .c(net_cout0),
    .cout(net_cout1),
    .sum(net_sum1));
  AL_FADD comp_10 (
    .a(net_a10),
    .b(net_nb10),
    .c(net_cout9),
    .cout(net_cout10),
    .sum(net_sum10));
  AL_FADD comp_2 (
    .a(net_a2),
    .b(net_nb2),
    .c(net_cout1),
    .cout(net_cout2),
    .sum(net_sum2));
  AL_FADD comp_3 (
    .a(net_a3),
    .b(net_nb3),
    .c(net_cout2),
    .cout(net_cout3),
    .sum(net_sum3));
  AL_FADD comp_4 (
    .a(net_a4),
    .b(net_nb4),
    .c(net_cout3),
    .cout(net_cout4),
    .sum(net_sum4));
  AL_FADD comp_5 (
    .a(net_a5),
    .b(net_nb5),
    .c(net_cout4),
    .cout(net_cout5),
    .sum(net_sum5));
  AL_FADD comp_6 (
    .a(net_a6),
    .b(net_nb6),
    .c(net_cout5),
    .cout(net_cout6),
    .sum(net_sum6));
  AL_FADD comp_7 (
    .a(net_a7),
    .b(net_nb7),
    .c(net_cout6),
    .cout(net_cout7),
    .sum(net_sum7));
  AL_FADD comp_8 (
    .a(net_a8),
    .b(net_nb8),
    .c(net_cout7),
    .cout(net_cout8),
    .sum(net_sum8));
  AL_FADD comp_9 (
    .a(net_a9),
    .b(net_nb9),
    .c(net_cout8),
    .cout(net_cout9),
    .sum(net_sum9));
  not inv_b0 (net_nb0, net_b0);
  not inv_b1 (net_nb1, net_b1);
  not inv_b10 (net_nb10, net_b10);
  not inv_b2 (net_nb2, net_b2);
  not inv_b3 (net_nb3, net_b3);
  not inv_b4 (net_nb4, net_b4);
  not inv_b5 (net_nb5, net_b5);
  not inv_b6 (net_nb6, net_b6);
  not inv_b7 (net_nb7, net_b7);
  not inv_b8 (net_nb8, net_b8);
  not inv_b9 (net_nb9, net_b9);
  not inv_cout (net_ncout, net_cout10);

endmodule 

module add_pu16_mu16_o16
  (
  i0,
  i1,
  o
  );

  input [15:0] i0;
  input [15:0] i1;
  output [15:0] o;

  wire net_a0;
  wire net_a1;
  wire net_a10;
  wire net_a11;
  wire net_a12;
  wire net_a13;
  wire net_a14;
  wire net_a15;
  wire net_a2;
  wire net_a3;
  wire net_a4;
  wire net_a5;
  wire net_a6;
  wire net_a7;
  wire net_a8;
  wire net_a9;
  wire net_b0;
  wire net_b1;
  wire net_b10;
  wire net_b11;
  wire net_b12;
  wire net_b13;
  wire net_b14;
  wire net_b15;
  wire net_b2;
  wire net_b3;
  wire net_b4;
  wire net_b5;
  wire net_b6;
  wire net_b7;
  wire net_b8;
  wire net_b9;
  wire net_cout0;
  wire net_cout1;
  wire net_cout10;
  wire net_cout11;
  wire net_cout12;
  wire net_cout13;
  wire net_cout14;
  wire net_cout15;
  wire net_cout2;
  wire net_cout3;
  wire net_cout4;
  wire net_cout5;
  wire net_cout6;
  wire net_cout7;
  wire net_cout8;
  wire net_cout9;
  wire net_nb0;
  wire net_nb1;
  wire net_nb10;
  wire net_nb11;
  wire net_nb12;
  wire net_nb13;
  wire net_nb14;
  wire net_nb15;
  wire net_nb2;
  wire net_nb3;
  wire net_nb4;
  wire net_nb5;
  wire net_nb6;
  wire net_nb7;
  wire net_nb8;
  wire net_nb9;
  wire net_sum0;
  wire net_sum1;
  wire net_sum10;
  wire net_sum11;
  wire net_sum12;
  wire net_sum13;
  wire net_sum14;
  wire net_sum15;
  wire net_sum2;
  wire net_sum3;
  wire net_sum4;
  wire net_sum5;
  wire net_sum6;
  wire net_sum7;
  wire net_sum8;
  wire net_sum9;

  assign net_a15 = i0[15];
  assign net_a14 = i0[14];
  assign net_a13 = i0[13];
  assign net_a12 = i0[12];
  assign net_a11 = i0[11];
  assign net_a10 = i0[10];
  assign net_a9 = i0[9];
  assign net_a8 = i0[8];
  assign net_a7 = i0[7];
  assign net_a6 = i0[6];
  assign net_a5 = i0[5];
  assign net_a4 = i0[4];
  assign net_a3 = i0[3];
  assign net_a2 = i0[2];
  assign net_a1 = i0[1];
  assign net_a0 = i0[0];
  assign net_b15 = i1[15];
  assign net_b14 = i1[14];
  assign net_b13 = i1[13];
  assign net_b12 = i1[12];
  assign net_b11 = i1[11];
  assign net_b10 = i1[10];
  assign net_b9 = i1[9];
  assign net_b8 = i1[8];
  assign net_b7 = i1[7];
  assign net_b6 = i1[6];
  assign net_b5 = i1[5];
  assign net_b4 = i1[4];
  assign net_b3 = i1[3];
  assign net_b2 = i1[2];
  assign net_b1 = i1[1];
  assign net_b0 = i1[0];
  assign o[15] = net_sum15;
  assign o[14] = net_sum14;
  assign o[13] = net_sum13;
  assign o[12] = net_sum12;
  assign o[11] = net_sum11;
  assign o[10] = net_sum10;
  assign o[9] = net_sum9;
  assign o[8] = net_sum8;
  assign o[7] = net_sum7;
  assign o[6] = net_sum6;
  assign o[5] = net_sum5;
  assign o[4] = net_sum4;
  assign o[3] = net_sum3;
  assign o[2] = net_sum2;
  assign o[1] = net_sum1;
  assign o[0] = net_sum0;
  AL_FADD comp_0 (
    .a(net_a0),
    .b(net_nb0),
    .c(1'b1),
    .cout(net_cout0),
    .sum(net_sum0));
  AL_FADD comp_1 (
    .a(net_a1),
    .b(net_nb1),
    .c(net_cout0),
    .cout(net_cout1),
    .sum(net_sum1));
  AL_FADD comp_10 (
    .a(net_a10),
    .b(net_nb10),
    .c(net_cout9),
    .cout(net_cout10),
    .sum(net_sum10));
  AL_FADD comp_11 (
    .a(net_a11),
    .b(net_nb11),
    .c(net_cout10),
    .cout(net_cout11),
    .sum(net_sum11));
  AL_FADD comp_12 (
    .a(net_a12),
    .b(net_nb12),
    .c(net_cout11),
    .cout(net_cout12),
    .sum(net_sum12));
  AL_FADD comp_13 (
    .a(net_a13),
    .b(net_nb13),
    .c(net_cout12),
    .cout(net_cout13),
    .sum(net_sum13));
  AL_FADD comp_14 (
    .a(net_a14),
    .b(net_nb14),
    .c(net_cout13),
    .cout(net_cout14),
    .sum(net_sum14));
  AL_FADD comp_15 (
    .a(net_a15),
    .b(net_nb15),
    .c(net_cout14),
    .cout(net_cout15),
    .sum(net_sum15));
  AL_FADD comp_2 (
    .a(net_a2),
    .b(net_nb2),
    .c(net_cout1),
    .cout(net_cout2),
    .sum(net_sum2));
  AL_FADD comp_3 (
    .a(net_a3),
    .b(net_nb3),
    .c(net_cout2),
    .cout(net_cout3),
    .sum(net_sum3));
  AL_FADD comp_4 (
    .a(net_a4),
    .b(net_nb4),
    .c(net_cout3),
    .cout(net_cout4),
    .sum(net_sum4));
  AL_FADD comp_5 (
    .a(net_a5),
    .b(net_nb5),
    .c(net_cout4),
    .cout(net_cout5),
    .sum(net_sum5));
  AL_FADD comp_6 (
    .a(net_a6),
    .b(net_nb6),
    .c(net_cout5),
    .cout(net_cout6),
    .sum(net_sum6));
  AL_FADD comp_7 (
    .a(net_a7),
    .b(net_nb7),
    .c(net_cout6),
    .cout(net_cout7),
    .sum(net_sum7));
  AL_FADD comp_8 (
    .a(net_a8),
    .b(net_nb8),
    .c(net_cout7),
    .cout(net_cout8),
    .sum(net_sum8));
  AL_FADD comp_9 (
    .a(net_a9),
    .b(net_nb9),
    .c(net_cout8),
    .cout(net_cout9),
    .sum(net_sum9));
  not inv_b0 (net_nb0, net_b0);
  not inv_b1 (net_nb1, net_b1);
  not inv_b10 (net_nb10, net_b10);
  not inv_b11 (net_nb11, net_b11);
  not inv_b12 (net_nb12, net_b12);
  not inv_b13 (net_nb13, net_b13);
  not inv_b14 (net_nb14, net_b14);
  not inv_b15 (net_nb15, net_b15);
  not inv_b2 (net_nb2, net_b2);
  not inv_b3 (net_nb3, net_b3);
  not inv_b4 (net_nb4, net_b4);
  not inv_b5 (net_nb5, net_b5);
  not inv_b6 (net_nb6, net_b6);
  not inv_b7 (net_nb7, net_b7);
  not inv_b8 (net_nb8, net_b8);
  not inv_b9 (net_nb9, net_b9);

endmodule 

module add_pu13_mu13_o13
  (
  i0,
  i1,
  o
  );

  input [12:0] i0;
  input [12:0] i1;
  output [12:0] o;

  wire net_a0;
  wire net_a1;
  wire net_a10;
  wire net_a11;
  wire net_a12;
  wire net_a2;
  wire net_a3;
  wire net_a4;
  wire net_a5;
  wire net_a6;
  wire net_a7;
  wire net_a8;
  wire net_a9;
  wire net_b0;
  wire net_b1;
  wire net_b10;
  wire net_b11;
  wire net_b12;
  wire net_b2;
  wire net_b3;
  wire net_b4;
  wire net_b5;
  wire net_b6;
  wire net_b7;
  wire net_b8;
  wire net_b9;
  wire net_cout0;
  wire net_cout1;
  wire net_cout10;
  wire net_cout11;
  wire net_cout12;
  wire net_cout2;
  wire net_cout3;
  wire net_cout4;
  wire net_cout5;
  wire net_cout6;
  wire net_cout7;
  wire net_cout8;
  wire net_cout9;
  wire net_nb0;
  wire net_nb1;
  wire net_nb10;
  wire net_nb11;
  wire net_nb12;
  wire net_nb2;
  wire net_nb3;
  wire net_nb4;
  wire net_nb5;
  wire net_nb6;
  wire net_nb7;
  wire net_nb8;
  wire net_nb9;
  wire net_sum0;
  wire net_sum1;
  wire net_sum10;
  wire net_sum11;
  wire net_sum12;
  wire net_sum2;
  wire net_sum3;
  wire net_sum4;
  wire net_sum5;
  wire net_sum6;
  wire net_sum7;
  wire net_sum8;
  wire net_sum9;

  assign net_a12 = i0[12];
  assign net_a11 = i0[11];
  assign net_a10 = i0[10];
  assign net_a9 = i0[9];
  assign net_a8 = i0[8];
  assign net_a7 = i0[7];
  assign net_a6 = i0[6];
  assign net_a5 = i0[5];
  assign net_a4 = i0[4];
  assign net_a3 = i0[3];
  assign net_a2 = i0[2];
  assign net_a1 = i0[1];
  assign net_a0 = i0[0];
  assign net_b12 = i1[12];
  assign net_b11 = i1[11];
  assign net_b10 = i1[10];
  assign net_b9 = i1[9];
  assign net_b8 = i1[8];
  assign net_b7 = i1[7];
  assign net_b6 = i1[6];
  assign net_b5 = i1[5];
  assign net_b4 = i1[4];
  assign net_b3 = i1[3];
  assign net_b2 = i1[2];
  assign net_b1 = i1[1];
  assign net_b0 = i1[0];
  assign o[12] = net_sum12;
  assign o[11] = net_sum11;
  assign o[10] = net_sum10;
  assign o[9] = net_sum9;
  assign o[8] = net_sum8;
  assign o[7] = net_sum7;
  assign o[6] = net_sum6;
  assign o[5] = net_sum5;
  assign o[4] = net_sum4;
  assign o[3] = net_sum3;
  assign o[2] = net_sum2;
  assign o[1] = net_sum1;
  assign o[0] = net_sum0;
  AL_FADD comp_0 (
    .a(net_a0),
    .b(net_nb0),
    .c(1'b1),
    .cout(net_cout0),
    .sum(net_sum0));
  AL_FADD comp_1 (
    .a(net_a1),
    .b(net_nb1),
    .c(net_cout0),
    .cout(net_cout1),
    .sum(net_sum1));
  AL_FADD comp_10 (
    .a(net_a10),
    .b(net_nb10),
    .c(net_cout9),
    .cout(net_cout10),
    .sum(net_sum10));
  AL_FADD comp_11 (
    .a(net_a11),
    .b(net_nb11),
    .c(net_cout10),
    .cout(net_cout11),
    .sum(net_sum11));
  AL_FADD comp_12 (
    .a(net_a12),
    .b(net_nb12),
    .c(net_cout11),
    .cout(net_cout12),
    .sum(net_sum12));
  AL_FADD comp_2 (
    .a(net_a2),
    .b(net_nb2),
    .c(net_cout1),
    .cout(net_cout2),
    .sum(net_sum2));
  AL_FADD comp_3 (
    .a(net_a3),
    .b(net_nb3),
    .c(net_cout2),
    .cout(net_cout3),
    .sum(net_sum3));
  AL_FADD comp_4 (
    .a(net_a4),
    .b(net_nb4),
    .c(net_cout3),
    .cout(net_cout4),
    .sum(net_sum4));
  AL_FADD comp_5 (
    .a(net_a5),
    .b(net_nb5),
    .c(net_cout4),
    .cout(net_cout5),
    .sum(net_sum5));
  AL_FADD comp_6 (
    .a(net_a6),
    .b(net_nb6),
    .c(net_cout5),
    .cout(net_cout6),
    .sum(net_sum6));
  AL_FADD comp_7 (
    .a(net_a7),
    .b(net_nb7),
    .c(net_cout6),
    .cout(net_cout7),
    .sum(net_sum7));
  AL_FADD comp_8 (
    .a(net_a8),
    .b(net_nb8),
    .c(net_cout7),
    .cout(net_cout8),
    .sum(net_sum8));
  AL_FADD comp_9 (
    .a(net_a9),
    .b(net_nb9),
    .c(net_cout8),
    .cout(net_cout9),
    .sum(net_sum9));
  not inv_b0 (net_nb0, net_b0);
  not inv_b1 (net_nb1, net_b1);
  not inv_b10 (net_nb10, net_b10);
  not inv_b11 (net_nb11, net_b11);
  not inv_b12 (net_nb12, net_b12);
  not inv_b2 (net_nb2, net_b2);
  not inv_b3 (net_nb3, net_b3);
  not inv_b4 (net_nb4, net_b4);
  not inv_b5 (net_nb5, net_b5);
  not inv_b6 (net_nb6, net_b6);
  not inv_b7 (net_nb7, net_b7);
  not inv_b8 (net_nb8, net_b8);
  not inv_b9 (net_nb9, net_b9);

endmodule 

module ne_w8
  (
  i0,
  i1,
  o
  );

  input [7:0] i0;
  input [7:0] i1;
  output o;

  wire [7:0] diff;

  or any_diff (o, diff[0], diff[1], diff[2], diff[3], diff[4], diff[5], diff[6], diff[7]);
  xor diff_0 (diff[0], i0[0], i1[0]);
  xor diff_1 (diff[1], i0[1], i1[1]);
  xor diff_2 (diff[2], i0[2], i1[2]);
  xor diff_3 (diff[3], i0[3], i1[3]);
  xor diff_4 (diff[4], i0[4], i1[4]);
  xor diff_5 (diff[5], i0[5], i1[5]);
  xor diff_6 (diff[6], i0[6], i1[6]);
  xor diff_7 (diff[7], i0[7], i1[7]);

endmodule 

module reg_sr_as_w1
  (
  clk,
  d,
  en,
  reset,
  set,
  q
  );

  input clk;
  input d;
  input en;
  input reset;
  input set;
  output q;

  parameter REGSET = "RESET";
  wire enout;
  wire resetout;

  AL_MUX u_en0 (
    .i0(q),
    .i1(d),
    .sel(en),
    .o(enout));
  AL_MUX u_reset0 (
    .i0(enout),
    .i1(1'b0),
    .sel(reset),
    .o(resetout));
  AL_DFF #(
    .INI((REGSET == "SET") ? 1'b1 : 1'b0))
    u_seq0 (
    .clk(clk),
    .d(resetout),
    .reset(1'b0),
    .set(set),
    .q(q));

endmodule 

module add_pu13_pu13_pu13_pu13_pu13_o13
  (
  i0,
  i1,
  i2,
  i3,
  i4,
  o
  );

  input [12:0] i0;
  input [12:0] i1;
  input [12:0] i2;
  input [12:0] i3;
  input [12:0] i4;
  output [12:0] o;

  wire net_a0_0;
  wire net_a0_1;
  wire net_a0_10;
  wire net_a0_11;
  wire net_a0_12;
  wire net_a0_2;
  wire net_a0_3;
  wire net_a0_4;
  wire net_a0_5;
  wire net_a0_6;
  wire net_a0_7;
  wire net_a0_8;
  wire net_a0_9;
  wire net_a1_0;
  wire net_a1_1;
  wire net_a1_10;
  wire net_a1_11;
  wire net_a1_12;
  wire net_a1_2;
  wire net_a1_3;
  wire net_a1_4;
  wire net_a1_5;
  wire net_a1_6;
  wire net_a1_7;
  wire net_a1_8;
  wire net_a1_9;
  wire net_a2_0;
  wire net_a2_1;
  wire net_a2_10;
  wire net_a2_11;
  wire net_a2_12;
  wire net_a2_2;
  wire net_a2_3;
  wire net_a2_4;
  wire net_a2_5;
  wire net_a2_6;
  wire net_a2_7;
  wire net_a2_8;
  wire net_a2_9;
  wire net_a3_0;
  wire net_a3_1;
  wire net_a3_10;
  wire net_a3_11;
  wire net_a3_12;
  wire net_a3_2;
  wire net_a3_3;
  wire net_a3_4;
  wire net_a3_5;
  wire net_a3_6;
  wire net_a3_7;
  wire net_a3_8;
  wire net_a3_9;
  wire net_a4_0;
  wire net_a4_1;
  wire net_a4_10;
  wire net_a4_11;
  wire net_a4_12;
  wire net_a4_2;
  wire net_a4_3;
  wire net_a4_4;
  wire net_a4_5;
  wire net_a4_6;
  wire net_a4_7;
  wire net_a4_8;
  wire net_a4_9;
  wire net_cout1_0;
  wire net_cout1_1;
  wire net_cout1_10;
  wire net_cout1_11;
  wire net_cout1_12;
  wire net_cout1_2;
  wire net_cout1_3;
  wire net_cout1_4;
  wire net_cout1_5;
  wire net_cout1_6;
  wire net_cout1_7;
  wire net_cout1_8;
  wire net_cout1_9;
  wire net_cout2_0;
  wire net_cout2_1;
  wire net_cout2_10;
  wire net_cout2_11;
  wire net_cout2_12;
  wire net_cout2_2;
  wire net_cout2_3;
  wire net_cout2_4;
  wire net_cout2_5;
  wire net_cout2_6;
  wire net_cout2_7;
  wire net_cout2_8;
  wire net_cout2_9;
  wire net_cout3_0;
  wire net_cout3_1;
  wire net_cout3_10;
  wire net_cout3_11;
  wire net_cout3_12;
  wire net_cout3_2;
  wire net_cout3_3;
  wire net_cout3_4;
  wire net_cout3_5;
  wire net_cout3_6;
  wire net_cout3_7;
  wire net_cout3_8;
  wire net_cout3_9;
  wire net_cout4_0;
  wire net_cout4_1;
  wire net_cout4_10;
  wire net_cout4_11;
  wire net_cout4_12;
  wire net_cout4_2;
  wire net_cout4_3;
  wire net_cout4_4;
  wire net_cout4_5;
  wire net_cout4_6;
  wire net_cout4_7;
  wire net_cout4_8;
  wire net_cout4_9;
  wire net_sum1_0;
  wire net_sum1_1;
  wire net_sum1_10;
  wire net_sum1_11;
  wire net_sum1_12;
  wire net_sum1_2;
  wire net_sum1_3;
  wire net_sum1_4;
  wire net_sum1_5;
  wire net_sum1_6;
  wire net_sum1_7;
  wire net_sum1_8;
  wire net_sum1_9;
  wire net_sum2_0;
  wire net_sum2_1;
  wire net_sum2_10;
  wire net_sum2_11;
  wire net_sum2_12;
  wire net_sum2_2;
  wire net_sum2_3;
  wire net_sum2_4;
  wire net_sum2_5;
  wire net_sum2_6;
  wire net_sum2_7;
  wire net_sum2_8;
  wire net_sum2_9;
  wire net_sum3_0;
  wire net_sum3_1;
  wire net_sum3_10;
  wire net_sum3_11;
  wire net_sum3_12;
  wire net_sum3_2;
  wire net_sum3_3;
  wire net_sum3_4;
  wire net_sum3_5;
  wire net_sum3_6;
  wire net_sum3_7;
  wire net_sum3_8;
  wire net_sum3_9;
  wire net_sum4_0;
  wire net_sum4_1;
  wire net_sum4_10;
  wire net_sum4_11;
  wire net_sum4_12;
  wire net_sum4_2;
  wire net_sum4_3;
  wire net_sum4_4;
  wire net_sum4_5;
  wire net_sum4_6;
  wire net_sum4_7;
  wire net_sum4_8;
  wire net_sum4_9;

  assign net_a0_12 = i0[12];
  assign net_a0_11 = i0[11];
  assign net_a0_10 = i0[10];
  assign net_a0_9 = i0[9];
  assign net_a0_8 = i0[8];
  assign net_a0_7 = i0[7];
  assign net_a0_6 = i0[6];
  assign net_a0_5 = i0[5];
  assign net_a0_4 = i0[4];
  assign net_a0_3 = i0[3];
  assign net_a0_2 = i0[2];
  assign net_a0_1 = i0[1];
  assign net_a0_0 = i0[0];
  assign net_a1_12 = i1[12];
  assign net_a1_11 = i1[11];
  assign net_a1_10 = i1[10];
  assign net_a1_9 = i1[9];
  assign net_a1_8 = i1[8];
  assign net_a1_7 = i1[7];
  assign net_a1_6 = i1[6];
  assign net_a1_5 = i1[5];
  assign net_a1_4 = i1[4];
  assign net_a1_3 = i1[3];
  assign net_a1_2 = i1[2];
  assign net_a1_1 = i1[1];
  assign net_a1_0 = i1[0];
  assign net_a2_12 = i2[12];
  assign net_a2_11 = i2[11];
  assign net_a2_10 = i2[10];
  assign net_a2_9 = i2[9];
  assign net_a2_8 = i2[8];
  assign net_a2_7 = i2[7];
  assign net_a2_6 = i2[6];
  assign net_a2_5 = i2[5];
  assign net_a2_4 = i2[4];
  assign net_a2_3 = i2[3];
  assign net_a2_2 = i2[2];
  assign net_a2_1 = i2[1];
  assign net_a2_0 = i2[0];
  assign net_a3_12 = i3[12];
  assign net_a3_11 = i3[11];
  assign net_a3_10 = i3[10];
  assign net_a3_9 = i3[9];
  assign net_a3_8 = i3[8];
  assign net_a3_7 = i3[7];
  assign net_a3_6 = i3[6];
  assign net_a3_5 = i3[5];
  assign net_a3_4 = i3[4];
  assign net_a3_3 = i3[3];
  assign net_a3_2 = i3[2];
  assign net_a3_1 = i3[1];
  assign net_a3_0 = i3[0];
  assign net_a4_12 = i4[12];
  assign net_a4_11 = i4[11];
  assign net_a4_10 = i4[10];
  assign net_a4_9 = i4[9];
  assign net_a4_8 = i4[8];
  assign net_a4_7 = i4[7];
  assign net_a4_6 = i4[6];
  assign net_a4_5 = i4[5];
  assign net_a4_4 = i4[4];
  assign net_a4_3 = i4[3];
  assign net_a4_2 = i4[2];
  assign net_a4_1 = i4[1];
  assign net_a4_0 = i4[0];
  assign o[12] = net_sum4_12;
  assign o[11] = net_sum4_11;
  assign o[10] = net_sum4_10;
  assign o[9] = net_sum4_9;
  assign o[8] = net_sum4_8;
  assign o[7] = net_sum4_7;
  assign o[6] = net_sum4_6;
  assign o[5] = net_sum4_5;
  assign o[4] = net_sum4_4;
  assign o[3] = net_sum4_3;
  assign o[2] = net_sum4_2;
  assign o[1] = net_sum4_1;
  assign o[0] = net_sum4_0;
  AL_FADD comp1_0 (
    .a(net_a1_0),
    .b(net_a0_0),
    .c(1'b0),
    .cout(net_cout1_0),
    .sum(net_sum1_0));
  AL_FADD comp1_1 (
    .a(net_a1_1),
    .b(net_a0_1),
    .c(net_cout1_0),
    .cout(net_cout1_1),
    .sum(net_sum1_1));
  AL_FADD comp1_10 (
    .a(net_a1_10),
    .b(net_a0_10),
    .c(net_cout1_9),
    .cout(net_cout1_10),
    .sum(net_sum1_10));
  AL_FADD comp1_11 (
    .a(net_a1_11),
    .b(net_a0_11),
    .c(net_cout1_10),
    .cout(net_cout1_11),
    .sum(net_sum1_11));
  AL_FADD comp1_12 (
    .a(net_a1_12),
    .b(net_a0_12),
    .c(net_cout1_11),
    .cout(net_cout1_12),
    .sum(net_sum1_12));
  AL_FADD comp1_2 (
    .a(net_a1_2),
    .b(net_a0_2),
    .c(net_cout1_1),
    .cout(net_cout1_2),
    .sum(net_sum1_2));
  AL_FADD comp1_3 (
    .a(net_a1_3),
    .b(net_a0_3),
    .c(net_cout1_2),
    .cout(net_cout1_3),
    .sum(net_sum1_3));
  AL_FADD comp1_4 (
    .a(net_a1_4),
    .b(net_a0_4),
    .c(net_cout1_3),
    .cout(net_cout1_4),
    .sum(net_sum1_4));
  AL_FADD comp1_5 (
    .a(net_a1_5),
    .b(net_a0_5),
    .c(net_cout1_4),
    .cout(net_cout1_5),
    .sum(net_sum1_5));
  AL_FADD comp1_6 (
    .a(net_a1_6),
    .b(net_a0_6),
    .c(net_cout1_5),
    .cout(net_cout1_6),
    .sum(net_sum1_6));
  AL_FADD comp1_7 (
    .a(net_a1_7),
    .b(net_a0_7),
    .c(net_cout1_6),
    .cout(net_cout1_7),
    .sum(net_sum1_7));
  AL_FADD comp1_8 (
    .a(net_a1_8),
    .b(net_a0_8),
    .c(net_cout1_7),
    .cout(net_cout1_8),
    .sum(net_sum1_8));
  AL_FADD comp1_9 (
    .a(net_a1_9),
    .b(net_a0_9),
    .c(net_cout1_8),
    .cout(net_cout1_9),
    .sum(net_sum1_9));
  AL_FADD comp2_0 (
    .a(net_a2_0),
    .b(net_sum1_0),
    .c(1'b0),
    .cout(net_cout2_0),
    .sum(net_sum2_0));
  AL_FADD comp2_1 (
    .a(net_a2_1),
    .b(net_sum1_1),
    .c(net_cout2_0),
    .cout(net_cout2_1),
    .sum(net_sum2_1));
  AL_FADD comp2_10 (
    .a(net_a2_10),
    .b(net_sum1_10),
    .c(net_cout2_9),
    .cout(net_cout2_10),
    .sum(net_sum2_10));
  AL_FADD comp2_11 (
    .a(net_a2_11),
    .b(net_sum1_11),
    .c(net_cout2_10),
    .cout(net_cout2_11),
    .sum(net_sum2_11));
  AL_FADD comp2_12 (
    .a(net_a2_12),
    .b(net_sum1_12),
    .c(net_cout2_11),
    .cout(net_cout2_12),
    .sum(net_sum2_12));
  AL_FADD comp2_2 (
    .a(net_a2_2),
    .b(net_sum1_2),
    .c(net_cout2_1),
    .cout(net_cout2_2),
    .sum(net_sum2_2));
  AL_FADD comp2_3 (
    .a(net_a2_3),
    .b(net_sum1_3),
    .c(net_cout2_2),
    .cout(net_cout2_3),
    .sum(net_sum2_3));
  AL_FADD comp2_4 (
    .a(net_a2_4),
    .b(net_sum1_4),
    .c(net_cout2_3),
    .cout(net_cout2_4),
    .sum(net_sum2_4));
  AL_FADD comp2_5 (
    .a(net_a2_5),
    .b(net_sum1_5),
    .c(net_cout2_4),
    .cout(net_cout2_5),
    .sum(net_sum2_5));
  AL_FADD comp2_6 (
    .a(net_a2_6),
    .b(net_sum1_6),
    .c(net_cout2_5),
    .cout(net_cout2_6),
    .sum(net_sum2_6));
  AL_FADD comp2_7 (
    .a(net_a2_7),
    .b(net_sum1_7),
    .c(net_cout2_6),
    .cout(net_cout2_7),
    .sum(net_sum2_7));
  AL_FADD comp2_8 (
    .a(net_a2_8),
    .b(net_sum1_8),
    .c(net_cout2_7),
    .cout(net_cout2_8),
    .sum(net_sum2_8));
  AL_FADD comp2_9 (
    .a(net_a2_9),
    .b(net_sum1_9),
    .c(net_cout2_8),
    .cout(net_cout2_9),
    .sum(net_sum2_9));
  AL_FADD comp3_0 (
    .a(net_a3_0),
    .b(net_sum2_0),
    .c(1'b0),
    .cout(net_cout3_0),
    .sum(net_sum3_0));
  AL_FADD comp3_1 (
    .a(net_a3_1),
    .b(net_sum2_1),
    .c(net_cout3_0),
    .cout(net_cout3_1),
    .sum(net_sum3_1));
  AL_FADD comp3_10 (
    .a(net_a3_10),
    .b(net_sum2_10),
    .c(net_cout3_9),
    .cout(net_cout3_10),
    .sum(net_sum3_10));
  AL_FADD comp3_11 (
    .a(net_a3_11),
    .b(net_sum2_11),
    .c(net_cout3_10),
    .cout(net_cout3_11),
    .sum(net_sum3_11));
  AL_FADD comp3_12 (
    .a(net_a3_12),
    .b(net_sum2_12),
    .c(net_cout3_11),
    .cout(net_cout3_12),
    .sum(net_sum3_12));
  AL_FADD comp3_2 (
    .a(net_a3_2),
    .b(net_sum2_2),
    .c(net_cout3_1),
    .cout(net_cout3_2),
    .sum(net_sum3_2));
  AL_FADD comp3_3 (
    .a(net_a3_3),
    .b(net_sum2_3),
    .c(net_cout3_2),
    .cout(net_cout3_3),
    .sum(net_sum3_3));
  AL_FADD comp3_4 (
    .a(net_a3_4),
    .b(net_sum2_4),
    .c(net_cout3_3),
    .cout(net_cout3_4),
    .sum(net_sum3_4));
  AL_FADD comp3_5 (
    .a(net_a3_5),
    .b(net_sum2_5),
    .c(net_cout3_4),
    .cout(net_cout3_5),
    .sum(net_sum3_5));
  AL_FADD comp3_6 (
    .a(net_a3_6),
    .b(net_sum2_6),
    .c(net_cout3_5),
    .cout(net_cout3_6),
    .sum(net_sum3_6));
  AL_FADD comp3_7 (
    .a(net_a3_7),
    .b(net_sum2_7),
    .c(net_cout3_6),
    .cout(net_cout3_7),
    .sum(net_sum3_7));
  AL_FADD comp3_8 (
    .a(net_a3_8),
    .b(net_sum2_8),
    .c(net_cout3_7),
    .cout(net_cout3_8),
    .sum(net_sum3_8));
  AL_FADD comp3_9 (
    .a(net_a3_9),
    .b(net_sum2_9),
    .c(net_cout3_8),
    .cout(net_cout3_9),
    .sum(net_sum3_9));
  AL_FADD comp4_0 (
    .a(net_a4_0),
    .b(net_sum3_0),
    .c(1'b0),
    .cout(net_cout4_0),
    .sum(net_sum4_0));
  AL_FADD comp4_1 (
    .a(net_a4_1),
    .b(net_sum3_1),
    .c(net_cout4_0),
    .cout(net_cout4_1),
    .sum(net_sum4_1));
  AL_FADD comp4_10 (
    .a(net_a4_10),
    .b(net_sum3_10),
    .c(net_cout4_9),
    .cout(net_cout4_10),
    .sum(net_sum4_10));
  AL_FADD comp4_11 (
    .a(net_a4_11),
    .b(net_sum3_11),
    .c(net_cout4_10),
    .cout(net_cout4_11),
    .sum(net_sum4_11));
  AL_FADD comp4_12 (
    .a(net_a4_12),
    .b(net_sum3_12),
    .c(net_cout4_11),
    .cout(net_cout4_12),
    .sum(net_sum4_12));
  AL_FADD comp4_2 (
    .a(net_a4_2),
    .b(net_sum3_2),
    .c(net_cout4_1),
    .cout(net_cout4_2),
    .sum(net_sum4_2));
  AL_FADD comp4_3 (
    .a(net_a4_3),
    .b(net_sum3_3),
    .c(net_cout4_2),
    .cout(net_cout4_3),
    .sum(net_sum4_3));
  AL_FADD comp4_4 (
    .a(net_a4_4),
    .b(net_sum3_4),
    .c(net_cout4_3),
    .cout(net_cout4_4),
    .sum(net_sum4_4));
  AL_FADD comp4_5 (
    .a(net_a4_5),
    .b(net_sum3_5),
    .c(net_cout4_4),
    .cout(net_cout4_5),
    .sum(net_sum4_5));
  AL_FADD comp4_6 (
    .a(net_a4_6),
    .b(net_sum3_6),
    .c(net_cout4_5),
    .cout(net_cout4_6),
    .sum(net_sum4_6));
  AL_FADD comp4_7 (
    .a(net_a4_7),
    .b(net_sum3_7),
    .c(net_cout4_6),
    .cout(net_cout4_7),
    .sum(net_sum4_7));
  AL_FADD comp4_8 (
    .a(net_a4_8),
    .b(net_sum3_8),
    .c(net_cout4_7),
    .cout(net_cout4_8),
    .sum(net_sum4_8));
  AL_FADD comp4_9 (
    .a(net_a4_9),
    .b(net_sum3_9),
    .c(net_cout4_8),
    .cout(net_cout4_9),
    .sum(net_sum4_9));

endmodule 

module AL_MUX
  (
  input i0,
  input i1,
  input sel,
  output o
  );

  wire not_sel, sel_i0, sel_i1;
  not u0 (not_sel, sel);
  and u1 (sel_i1, sel, i1);
  and u2 (sel_i0, not_sel, i0);
  or u3 (o, sel_i1, sel_i0);

endmodule

module AL_FADD
  (
  input a,
  input b,
  input c,
  output sum,
  output cout
  );

  wire prop;
  wire not_prop;
  wire sel_i0;
  wire sel_i1;

  xor u0 (prop, a, b);
  xor u1 (sum, prop, c);
  not u2 (not_prop, prop);
  and u3 (sel_i1, prop, c);
  and u4 (sel_i0, not_prop, a);
  or  u5 (cout, sel_i0, sel_i1);

endmodule

module AL_DFF
  (
  input reset,
  input set,
  input clk,
  input d,
  output reg q
  );

  parameter INI = 1'b0;

  always @(posedge reset or posedge set or posedge clk)
  begin
    if (reset)
      q <= 1'b0;
    else if (set)
      q <= 1'b1;
    else
      q <= d;
  end

endmodule

